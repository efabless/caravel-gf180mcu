VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_power_routing
  CLASS BLOCK ;
  FOREIGN caravel_power_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.400 BY 25.350 ;
  OBS
      LAYER Metal2 ;
        RECT 1896.360 4698.600 1905.860 4720.000 ;
        RECT 1908.760 4698.600 1919.010 4720.000 ;
        RECT 1920.610 4698.600 1930.860 4720.000 ;
        RECT 1934.140 4698.600 1944.390 4720.000 ;
        RECT 1945.990 4698.600 1956.240 4720.000 ;
        RECT 1959.140 4698.600 1968.640 4720.000 ;
        RECT 2996.360 4698.600 3005.860 4720.000 ;
        RECT 3008.760 4698.600 3019.010 4720.000 ;
        RECT 3020.610 4698.600 3030.860 4720.000 ;
        RECT 3034.140 4698.600 3044.390 4720.000 ;
        RECT 3045.990 4698.600 3056.240 4720.000 ;
        RECT 3059.140 4698.600 3068.640 4720.000 ;
        RECT 350.000 4384.140 352.440 4393.640 ;
        RECT 350.000 4370.990 352.440 4381.240 ;
        RECT 3527.560 4379.140 3530.000 4388.640 ;
        RECT 350.000 4359.140 352.440 4369.390 ;
        RECT 3527.560 4365.990 3530.000 4376.240 ;
        RECT 350.000 4345.610 352.440 4355.860 ;
        RECT 3527.560 4354.140 3530.000 4364.390 ;
        RECT 350.000 4333.760 352.440 4344.010 ;
        RECT 3527.560 4340.610 3530.000 4350.860 ;
        RECT 350.000 4321.360 352.440 4330.860 ;
        RECT 3527.560 4328.760 3530.000 4339.010 ;
        RECT 3527.560 4316.360 3530.000 4325.860 ;
        RECT 350.000 4179.140 352.440 4188.640 ;
        RECT 350.000 4165.990 352.440 4176.240 ;
        RECT 350.000 4154.140 352.440 4164.390 ;
        RECT 350.000 4140.610 352.440 4150.860 ;
        RECT 350.000 4128.760 352.440 4139.010 ;
        RECT 350.000 4116.360 352.440 4125.860 ;
        RECT 350.000 3974.140 352.440 3983.640 ;
        RECT 350.000 3960.990 352.440 3971.240 ;
        RECT 350.000 3949.140 352.440 3959.390 ;
        RECT 3527.560 3949.140 3530.000 3958.640 ;
        RECT 350.000 3935.610 352.440 3945.860 ;
        RECT 3527.560 3935.990 3530.000 3946.240 ;
        RECT 350.000 3923.760 352.440 3934.010 ;
        RECT 3527.560 3924.140 3530.000 3934.390 ;
        RECT 350.000 3911.360 352.440 3920.860 ;
        RECT 3527.560 3910.610 3530.000 3920.860 ;
        RECT 3527.560 3898.760 3530.000 3909.010 ;
        RECT 3527.560 3886.360 3530.000 3895.860 ;
        RECT 3527.560 2444.140 3530.000 2453.640 ;
        RECT 3527.560 2430.990 3530.000 2441.240 ;
        RECT 3527.560 2419.140 3530.000 2429.390 ;
        RECT 3527.560 2405.610 3530.000 2415.860 ;
        RECT 3527.560 2393.760 3530.000 2404.010 ;
        RECT 3527.560 2381.360 3530.000 2390.860 ;
        RECT 350.000 2334.140 352.440 2343.640 ;
        RECT 350.000 2320.990 352.440 2331.240 ;
        RECT 350.000 2309.140 352.440 2319.390 ;
        RECT 350.000 2295.610 352.440 2305.860 ;
        RECT 350.000 2283.760 352.440 2294.010 ;
        RECT 350.000 2271.360 352.440 2280.860 ;
        RECT 3527.560 2229.140 3530.000 2238.640 ;
        RECT 3527.560 2215.990 3530.000 2226.240 ;
        RECT 3527.560 2204.140 3530.000 2214.390 ;
        RECT 3527.560 2190.610 3530.000 2200.860 ;
        RECT 3527.560 2178.760 3530.000 2189.010 ;
        RECT 3527.560 2166.360 3530.000 2175.860 ;
        RECT 350.000 2129.140 352.440 2138.640 ;
        RECT 350.000 2115.990 352.440 2126.240 ;
        RECT 350.000 2104.140 352.440 2114.390 ;
        RECT 350.000 2090.610 352.440 2100.860 ;
        RECT 350.000 2078.760 352.440 2089.010 ;
        RECT 350.000 2066.360 352.440 2075.860 ;
        RECT 3527.560 2014.140 3530.000 2023.640 ;
        RECT 3527.560 2000.990 3530.000 2011.240 ;
        RECT 3527.560 1989.140 3530.000 1999.390 ;
        RECT 3527.560 1975.610 3530.000 1985.860 ;
        RECT 3527.560 1963.760 3530.000 1974.010 ;
        RECT 3527.560 1951.360 3530.000 1960.860 ;
        RECT 350.000 694.140 352.440 703.640 ;
        RECT 350.000 680.990 352.440 691.240 ;
        RECT 350.000 669.140 352.440 679.390 ;
        RECT 350.000 655.610 352.440 665.860 ;
        RECT 350.000 643.760 352.440 654.010 ;
        RECT 350.000 631.360 352.440 640.860 ;
        RECT 350.000 489.140 352.440 498.640 ;
        RECT 350.000 475.990 352.440 486.240 ;
        RECT 350.000 464.140 352.440 474.390 ;
        RECT 350.000 450.610 352.440 460.860 ;
        RECT 350.000 438.760 352.440 449.010 ;
        RECT 350.000 426.360 352.440 435.860 ;
        RECT 526.360 350.000 535.860 370.440 ;
        RECT 538.760 350.000 549.010 370.440 ;
        RECT 550.610 350.000 560.860 370.440 ;
        RECT 564.140 350.000 574.390 370.440 ;
        RECT 575.990 350.000 586.240 370.440 ;
        RECT 589.140 350.000 598.640 370.440 ;
        RECT 1351.360 350.000 1360.860 370.440 ;
        RECT 1363.760 350.000 1374.010 370.440 ;
        RECT 1375.610 350.000 1385.860 370.440 ;
        RECT 1389.140 350.000 1399.390 370.440 ;
        RECT 1400.990 350.000 1411.240 370.440 ;
        RECT 1414.140 350.000 1423.640 370.440 ;
        RECT 3001.360 350.000 3010.860 370.440 ;
        RECT 3013.760 350.000 3024.010 370.440 ;
        RECT 3025.610 350.000 3035.860 370.440 ;
        RECT 3039.140 350.000 3049.390 370.440 ;
        RECT 3050.990 350.000 3061.240 370.440 ;
        RECT 3064.140 350.000 3073.640 370.440 ;
        RECT 3276.360 350.000 3285.860 380.440 ;
        RECT 3288.760 350.000 3299.010 380.440 ;
        RECT 3300.610 350.000 3310.860 380.440 ;
        RECT 3314.140 350.000 3324.390 380.440 ;
        RECT 3325.990 350.000 3336.240 380.440 ;
        RECT 3339.140 350.000 3348.640 380.440 ;
      LAYER Via2 ;
        RECT 1896.630 4707.995 1896.910 4708.275 ;
        RECT 1897.250 4707.995 1897.530 4708.275 ;
        RECT 1897.870 4707.995 1898.150 4708.275 ;
        RECT 1898.490 4707.995 1898.770 4708.275 ;
        RECT 1899.110 4707.995 1899.390 4708.275 ;
        RECT 1899.730 4707.995 1900.010 4708.275 ;
        RECT 1896.630 4707.375 1896.910 4707.655 ;
        RECT 1897.250 4707.375 1897.530 4707.655 ;
        RECT 1897.870 4707.375 1898.150 4707.655 ;
        RECT 1898.490 4707.375 1898.770 4707.655 ;
        RECT 1899.110 4707.375 1899.390 4707.655 ;
        RECT 1899.730 4707.375 1900.010 4707.655 ;
        RECT 1896.630 4706.755 1896.910 4707.035 ;
        RECT 1897.250 4706.755 1897.530 4707.035 ;
        RECT 1897.870 4706.755 1898.150 4707.035 ;
        RECT 1898.490 4706.755 1898.770 4707.035 ;
        RECT 1899.110 4706.755 1899.390 4707.035 ;
        RECT 1899.730 4706.755 1900.010 4707.035 ;
        RECT 1896.630 4706.135 1896.910 4706.415 ;
        RECT 1897.250 4706.135 1897.530 4706.415 ;
        RECT 1897.870 4706.135 1898.150 4706.415 ;
        RECT 1898.490 4706.135 1898.770 4706.415 ;
        RECT 1899.110 4706.135 1899.390 4706.415 ;
        RECT 1899.730 4706.135 1900.010 4706.415 ;
        RECT 1896.630 4705.515 1896.910 4705.795 ;
        RECT 1897.250 4705.515 1897.530 4705.795 ;
        RECT 1897.870 4705.515 1898.150 4705.795 ;
        RECT 1898.490 4705.515 1898.770 4705.795 ;
        RECT 1899.110 4705.515 1899.390 4705.795 ;
        RECT 1899.730 4705.515 1900.010 4705.795 ;
        RECT 1896.630 4704.895 1896.910 4705.175 ;
        RECT 1897.250 4704.895 1897.530 4705.175 ;
        RECT 1897.870 4704.895 1898.150 4705.175 ;
        RECT 1898.490 4704.895 1898.770 4705.175 ;
        RECT 1899.110 4704.895 1899.390 4705.175 ;
        RECT 1899.730 4704.895 1900.010 4705.175 ;
        RECT 1896.630 4704.275 1896.910 4704.555 ;
        RECT 1897.250 4704.275 1897.530 4704.555 ;
        RECT 1897.870 4704.275 1898.150 4704.555 ;
        RECT 1898.490 4704.275 1898.770 4704.555 ;
        RECT 1899.110 4704.275 1899.390 4704.555 ;
        RECT 1899.730 4704.275 1900.010 4704.555 ;
        RECT 1896.630 4703.655 1896.910 4703.935 ;
        RECT 1897.250 4703.655 1897.530 4703.935 ;
        RECT 1897.870 4703.655 1898.150 4703.935 ;
        RECT 1898.490 4703.655 1898.770 4703.935 ;
        RECT 1899.110 4703.655 1899.390 4703.935 ;
        RECT 1899.730 4703.655 1900.010 4703.935 ;
        RECT 1896.630 4703.035 1896.910 4703.315 ;
        RECT 1897.250 4703.035 1897.530 4703.315 ;
        RECT 1897.870 4703.035 1898.150 4703.315 ;
        RECT 1898.490 4703.035 1898.770 4703.315 ;
        RECT 1899.110 4703.035 1899.390 4703.315 ;
        RECT 1899.730 4703.035 1900.010 4703.315 ;
        RECT 1896.630 4702.415 1896.910 4702.695 ;
        RECT 1897.250 4702.415 1897.530 4702.695 ;
        RECT 1897.870 4702.415 1898.150 4702.695 ;
        RECT 1898.490 4702.415 1898.770 4702.695 ;
        RECT 1899.110 4702.415 1899.390 4702.695 ;
        RECT 1899.730 4702.415 1900.010 4702.695 ;
        RECT 1896.630 4701.795 1896.910 4702.075 ;
        RECT 1897.250 4701.795 1897.530 4702.075 ;
        RECT 1897.870 4701.795 1898.150 4702.075 ;
        RECT 1898.490 4701.795 1898.770 4702.075 ;
        RECT 1899.110 4701.795 1899.390 4702.075 ;
        RECT 1899.730 4701.795 1900.010 4702.075 ;
        RECT 1896.630 4701.175 1896.910 4701.455 ;
        RECT 1897.250 4701.175 1897.530 4701.455 ;
        RECT 1897.870 4701.175 1898.150 4701.455 ;
        RECT 1898.490 4701.175 1898.770 4701.455 ;
        RECT 1899.110 4701.175 1899.390 4701.455 ;
        RECT 1899.730 4701.175 1900.010 4701.455 ;
        RECT 1896.630 4700.555 1896.910 4700.835 ;
        RECT 1897.250 4700.555 1897.530 4700.835 ;
        RECT 1897.870 4700.555 1898.150 4700.835 ;
        RECT 1898.490 4700.555 1898.770 4700.835 ;
        RECT 1899.110 4700.555 1899.390 4700.835 ;
        RECT 1899.730 4700.555 1900.010 4700.835 ;
        RECT 1896.630 4699.935 1896.910 4700.215 ;
        RECT 1897.250 4699.935 1897.530 4700.215 ;
        RECT 1897.870 4699.935 1898.150 4700.215 ;
        RECT 1898.490 4699.935 1898.770 4700.215 ;
        RECT 1899.110 4699.935 1899.390 4700.215 ;
        RECT 1899.730 4699.935 1900.010 4700.215 ;
        RECT 1896.630 4699.315 1896.910 4699.595 ;
        RECT 1897.250 4699.315 1897.530 4699.595 ;
        RECT 1897.870 4699.315 1898.150 4699.595 ;
        RECT 1898.490 4699.315 1898.770 4699.595 ;
        RECT 1899.110 4699.315 1899.390 4699.595 ;
        RECT 1899.730 4699.315 1900.010 4699.595 ;
        RECT 1909.160 4707.995 1909.440 4708.275 ;
        RECT 1909.780 4707.995 1910.060 4708.275 ;
        RECT 1910.400 4707.995 1910.680 4708.275 ;
        RECT 1911.020 4707.995 1911.300 4708.275 ;
        RECT 1911.640 4707.995 1911.920 4708.275 ;
        RECT 1912.260 4707.995 1912.540 4708.275 ;
        RECT 1912.880 4707.995 1913.160 4708.275 ;
        RECT 1913.500 4707.995 1913.780 4708.275 ;
        RECT 1914.120 4707.995 1914.400 4708.275 ;
        RECT 1914.740 4707.995 1915.020 4708.275 ;
        RECT 1915.360 4707.995 1915.640 4708.275 ;
        RECT 1915.980 4707.995 1916.260 4708.275 ;
        RECT 1916.600 4707.995 1916.880 4708.275 ;
        RECT 1917.220 4707.995 1917.500 4708.275 ;
        RECT 1917.840 4707.995 1918.120 4708.275 ;
        RECT 1918.460 4707.995 1918.740 4708.275 ;
        RECT 1909.160 4707.375 1909.440 4707.655 ;
        RECT 1909.780 4707.375 1910.060 4707.655 ;
        RECT 1910.400 4707.375 1910.680 4707.655 ;
        RECT 1911.020 4707.375 1911.300 4707.655 ;
        RECT 1911.640 4707.375 1911.920 4707.655 ;
        RECT 1912.260 4707.375 1912.540 4707.655 ;
        RECT 1912.880 4707.375 1913.160 4707.655 ;
        RECT 1913.500 4707.375 1913.780 4707.655 ;
        RECT 1914.120 4707.375 1914.400 4707.655 ;
        RECT 1914.740 4707.375 1915.020 4707.655 ;
        RECT 1915.360 4707.375 1915.640 4707.655 ;
        RECT 1915.980 4707.375 1916.260 4707.655 ;
        RECT 1916.600 4707.375 1916.880 4707.655 ;
        RECT 1917.220 4707.375 1917.500 4707.655 ;
        RECT 1917.840 4707.375 1918.120 4707.655 ;
        RECT 1918.460 4707.375 1918.740 4707.655 ;
        RECT 1909.160 4706.755 1909.440 4707.035 ;
        RECT 1909.780 4706.755 1910.060 4707.035 ;
        RECT 1910.400 4706.755 1910.680 4707.035 ;
        RECT 1911.020 4706.755 1911.300 4707.035 ;
        RECT 1911.640 4706.755 1911.920 4707.035 ;
        RECT 1912.260 4706.755 1912.540 4707.035 ;
        RECT 1912.880 4706.755 1913.160 4707.035 ;
        RECT 1913.500 4706.755 1913.780 4707.035 ;
        RECT 1914.120 4706.755 1914.400 4707.035 ;
        RECT 1914.740 4706.755 1915.020 4707.035 ;
        RECT 1915.360 4706.755 1915.640 4707.035 ;
        RECT 1915.980 4706.755 1916.260 4707.035 ;
        RECT 1916.600 4706.755 1916.880 4707.035 ;
        RECT 1917.220 4706.755 1917.500 4707.035 ;
        RECT 1917.840 4706.755 1918.120 4707.035 ;
        RECT 1918.460 4706.755 1918.740 4707.035 ;
        RECT 1909.160 4706.135 1909.440 4706.415 ;
        RECT 1909.780 4706.135 1910.060 4706.415 ;
        RECT 1910.400 4706.135 1910.680 4706.415 ;
        RECT 1911.020 4706.135 1911.300 4706.415 ;
        RECT 1911.640 4706.135 1911.920 4706.415 ;
        RECT 1912.260 4706.135 1912.540 4706.415 ;
        RECT 1912.880 4706.135 1913.160 4706.415 ;
        RECT 1913.500 4706.135 1913.780 4706.415 ;
        RECT 1914.120 4706.135 1914.400 4706.415 ;
        RECT 1914.740 4706.135 1915.020 4706.415 ;
        RECT 1915.360 4706.135 1915.640 4706.415 ;
        RECT 1915.980 4706.135 1916.260 4706.415 ;
        RECT 1916.600 4706.135 1916.880 4706.415 ;
        RECT 1917.220 4706.135 1917.500 4706.415 ;
        RECT 1917.840 4706.135 1918.120 4706.415 ;
        RECT 1918.460 4706.135 1918.740 4706.415 ;
        RECT 1909.160 4705.515 1909.440 4705.795 ;
        RECT 1909.780 4705.515 1910.060 4705.795 ;
        RECT 1910.400 4705.515 1910.680 4705.795 ;
        RECT 1911.020 4705.515 1911.300 4705.795 ;
        RECT 1911.640 4705.515 1911.920 4705.795 ;
        RECT 1912.260 4705.515 1912.540 4705.795 ;
        RECT 1912.880 4705.515 1913.160 4705.795 ;
        RECT 1913.500 4705.515 1913.780 4705.795 ;
        RECT 1914.120 4705.515 1914.400 4705.795 ;
        RECT 1914.740 4705.515 1915.020 4705.795 ;
        RECT 1915.360 4705.515 1915.640 4705.795 ;
        RECT 1915.980 4705.515 1916.260 4705.795 ;
        RECT 1916.600 4705.515 1916.880 4705.795 ;
        RECT 1917.220 4705.515 1917.500 4705.795 ;
        RECT 1917.840 4705.515 1918.120 4705.795 ;
        RECT 1918.460 4705.515 1918.740 4705.795 ;
        RECT 1909.160 4704.895 1909.440 4705.175 ;
        RECT 1909.780 4704.895 1910.060 4705.175 ;
        RECT 1910.400 4704.895 1910.680 4705.175 ;
        RECT 1911.020 4704.895 1911.300 4705.175 ;
        RECT 1911.640 4704.895 1911.920 4705.175 ;
        RECT 1912.260 4704.895 1912.540 4705.175 ;
        RECT 1912.880 4704.895 1913.160 4705.175 ;
        RECT 1913.500 4704.895 1913.780 4705.175 ;
        RECT 1914.120 4704.895 1914.400 4705.175 ;
        RECT 1914.740 4704.895 1915.020 4705.175 ;
        RECT 1915.360 4704.895 1915.640 4705.175 ;
        RECT 1915.980 4704.895 1916.260 4705.175 ;
        RECT 1916.600 4704.895 1916.880 4705.175 ;
        RECT 1917.220 4704.895 1917.500 4705.175 ;
        RECT 1917.840 4704.895 1918.120 4705.175 ;
        RECT 1918.460 4704.895 1918.740 4705.175 ;
        RECT 1909.160 4704.275 1909.440 4704.555 ;
        RECT 1909.780 4704.275 1910.060 4704.555 ;
        RECT 1910.400 4704.275 1910.680 4704.555 ;
        RECT 1911.020 4704.275 1911.300 4704.555 ;
        RECT 1911.640 4704.275 1911.920 4704.555 ;
        RECT 1912.260 4704.275 1912.540 4704.555 ;
        RECT 1912.880 4704.275 1913.160 4704.555 ;
        RECT 1913.500 4704.275 1913.780 4704.555 ;
        RECT 1914.120 4704.275 1914.400 4704.555 ;
        RECT 1914.740 4704.275 1915.020 4704.555 ;
        RECT 1915.360 4704.275 1915.640 4704.555 ;
        RECT 1915.980 4704.275 1916.260 4704.555 ;
        RECT 1916.600 4704.275 1916.880 4704.555 ;
        RECT 1917.220 4704.275 1917.500 4704.555 ;
        RECT 1917.840 4704.275 1918.120 4704.555 ;
        RECT 1918.460 4704.275 1918.740 4704.555 ;
        RECT 1909.160 4703.655 1909.440 4703.935 ;
        RECT 1909.780 4703.655 1910.060 4703.935 ;
        RECT 1910.400 4703.655 1910.680 4703.935 ;
        RECT 1911.020 4703.655 1911.300 4703.935 ;
        RECT 1911.640 4703.655 1911.920 4703.935 ;
        RECT 1912.260 4703.655 1912.540 4703.935 ;
        RECT 1912.880 4703.655 1913.160 4703.935 ;
        RECT 1913.500 4703.655 1913.780 4703.935 ;
        RECT 1914.120 4703.655 1914.400 4703.935 ;
        RECT 1914.740 4703.655 1915.020 4703.935 ;
        RECT 1915.360 4703.655 1915.640 4703.935 ;
        RECT 1915.980 4703.655 1916.260 4703.935 ;
        RECT 1916.600 4703.655 1916.880 4703.935 ;
        RECT 1917.220 4703.655 1917.500 4703.935 ;
        RECT 1917.840 4703.655 1918.120 4703.935 ;
        RECT 1918.460 4703.655 1918.740 4703.935 ;
        RECT 1909.160 4703.035 1909.440 4703.315 ;
        RECT 1909.780 4703.035 1910.060 4703.315 ;
        RECT 1910.400 4703.035 1910.680 4703.315 ;
        RECT 1911.020 4703.035 1911.300 4703.315 ;
        RECT 1911.640 4703.035 1911.920 4703.315 ;
        RECT 1912.260 4703.035 1912.540 4703.315 ;
        RECT 1912.880 4703.035 1913.160 4703.315 ;
        RECT 1913.500 4703.035 1913.780 4703.315 ;
        RECT 1914.120 4703.035 1914.400 4703.315 ;
        RECT 1914.740 4703.035 1915.020 4703.315 ;
        RECT 1915.360 4703.035 1915.640 4703.315 ;
        RECT 1915.980 4703.035 1916.260 4703.315 ;
        RECT 1916.600 4703.035 1916.880 4703.315 ;
        RECT 1917.220 4703.035 1917.500 4703.315 ;
        RECT 1917.840 4703.035 1918.120 4703.315 ;
        RECT 1918.460 4703.035 1918.740 4703.315 ;
        RECT 1909.160 4702.415 1909.440 4702.695 ;
        RECT 1909.780 4702.415 1910.060 4702.695 ;
        RECT 1910.400 4702.415 1910.680 4702.695 ;
        RECT 1911.020 4702.415 1911.300 4702.695 ;
        RECT 1911.640 4702.415 1911.920 4702.695 ;
        RECT 1912.260 4702.415 1912.540 4702.695 ;
        RECT 1912.880 4702.415 1913.160 4702.695 ;
        RECT 1913.500 4702.415 1913.780 4702.695 ;
        RECT 1914.120 4702.415 1914.400 4702.695 ;
        RECT 1914.740 4702.415 1915.020 4702.695 ;
        RECT 1915.360 4702.415 1915.640 4702.695 ;
        RECT 1915.980 4702.415 1916.260 4702.695 ;
        RECT 1916.600 4702.415 1916.880 4702.695 ;
        RECT 1917.220 4702.415 1917.500 4702.695 ;
        RECT 1917.840 4702.415 1918.120 4702.695 ;
        RECT 1918.460 4702.415 1918.740 4702.695 ;
        RECT 1909.160 4701.795 1909.440 4702.075 ;
        RECT 1909.780 4701.795 1910.060 4702.075 ;
        RECT 1910.400 4701.795 1910.680 4702.075 ;
        RECT 1911.020 4701.795 1911.300 4702.075 ;
        RECT 1911.640 4701.795 1911.920 4702.075 ;
        RECT 1912.260 4701.795 1912.540 4702.075 ;
        RECT 1912.880 4701.795 1913.160 4702.075 ;
        RECT 1913.500 4701.795 1913.780 4702.075 ;
        RECT 1914.120 4701.795 1914.400 4702.075 ;
        RECT 1914.740 4701.795 1915.020 4702.075 ;
        RECT 1915.360 4701.795 1915.640 4702.075 ;
        RECT 1915.980 4701.795 1916.260 4702.075 ;
        RECT 1916.600 4701.795 1916.880 4702.075 ;
        RECT 1917.220 4701.795 1917.500 4702.075 ;
        RECT 1917.840 4701.795 1918.120 4702.075 ;
        RECT 1918.460 4701.795 1918.740 4702.075 ;
        RECT 1909.160 4701.175 1909.440 4701.455 ;
        RECT 1909.780 4701.175 1910.060 4701.455 ;
        RECT 1910.400 4701.175 1910.680 4701.455 ;
        RECT 1911.020 4701.175 1911.300 4701.455 ;
        RECT 1911.640 4701.175 1911.920 4701.455 ;
        RECT 1912.260 4701.175 1912.540 4701.455 ;
        RECT 1912.880 4701.175 1913.160 4701.455 ;
        RECT 1913.500 4701.175 1913.780 4701.455 ;
        RECT 1914.120 4701.175 1914.400 4701.455 ;
        RECT 1914.740 4701.175 1915.020 4701.455 ;
        RECT 1915.360 4701.175 1915.640 4701.455 ;
        RECT 1915.980 4701.175 1916.260 4701.455 ;
        RECT 1916.600 4701.175 1916.880 4701.455 ;
        RECT 1917.220 4701.175 1917.500 4701.455 ;
        RECT 1917.840 4701.175 1918.120 4701.455 ;
        RECT 1918.460 4701.175 1918.740 4701.455 ;
        RECT 1909.160 4700.555 1909.440 4700.835 ;
        RECT 1909.780 4700.555 1910.060 4700.835 ;
        RECT 1910.400 4700.555 1910.680 4700.835 ;
        RECT 1911.020 4700.555 1911.300 4700.835 ;
        RECT 1911.640 4700.555 1911.920 4700.835 ;
        RECT 1912.260 4700.555 1912.540 4700.835 ;
        RECT 1912.880 4700.555 1913.160 4700.835 ;
        RECT 1913.500 4700.555 1913.780 4700.835 ;
        RECT 1914.120 4700.555 1914.400 4700.835 ;
        RECT 1914.740 4700.555 1915.020 4700.835 ;
        RECT 1915.360 4700.555 1915.640 4700.835 ;
        RECT 1915.980 4700.555 1916.260 4700.835 ;
        RECT 1916.600 4700.555 1916.880 4700.835 ;
        RECT 1917.220 4700.555 1917.500 4700.835 ;
        RECT 1917.840 4700.555 1918.120 4700.835 ;
        RECT 1918.460 4700.555 1918.740 4700.835 ;
        RECT 1909.160 4699.935 1909.440 4700.215 ;
        RECT 1909.780 4699.935 1910.060 4700.215 ;
        RECT 1910.400 4699.935 1910.680 4700.215 ;
        RECT 1911.020 4699.935 1911.300 4700.215 ;
        RECT 1911.640 4699.935 1911.920 4700.215 ;
        RECT 1912.260 4699.935 1912.540 4700.215 ;
        RECT 1912.880 4699.935 1913.160 4700.215 ;
        RECT 1913.500 4699.935 1913.780 4700.215 ;
        RECT 1914.120 4699.935 1914.400 4700.215 ;
        RECT 1914.740 4699.935 1915.020 4700.215 ;
        RECT 1915.360 4699.935 1915.640 4700.215 ;
        RECT 1915.980 4699.935 1916.260 4700.215 ;
        RECT 1916.600 4699.935 1916.880 4700.215 ;
        RECT 1917.220 4699.935 1917.500 4700.215 ;
        RECT 1917.840 4699.935 1918.120 4700.215 ;
        RECT 1918.460 4699.935 1918.740 4700.215 ;
        RECT 1909.160 4699.315 1909.440 4699.595 ;
        RECT 1909.780 4699.315 1910.060 4699.595 ;
        RECT 1910.400 4699.315 1910.680 4699.595 ;
        RECT 1911.020 4699.315 1911.300 4699.595 ;
        RECT 1911.640 4699.315 1911.920 4699.595 ;
        RECT 1912.260 4699.315 1912.540 4699.595 ;
        RECT 1912.880 4699.315 1913.160 4699.595 ;
        RECT 1913.500 4699.315 1913.780 4699.595 ;
        RECT 1914.120 4699.315 1914.400 4699.595 ;
        RECT 1914.740 4699.315 1915.020 4699.595 ;
        RECT 1915.360 4699.315 1915.640 4699.595 ;
        RECT 1915.980 4699.315 1916.260 4699.595 ;
        RECT 1916.600 4699.315 1916.880 4699.595 ;
        RECT 1917.220 4699.315 1917.500 4699.595 ;
        RECT 1917.840 4699.315 1918.120 4699.595 ;
        RECT 1918.460 4699.315 1918.740 4699.595 ;
        RECT 1921.010 4707.995 1921.290 4708.275 ;
        RECT 1921.630 4707.995 1921.910 4708.275 ;
        RECT 1922.250 4707.995 1922.530 4708.275 ;
        RECT 1922.870 4707.995 1923.150 4708.275 ;
        RECT 1923.490 4707.995 1923.770 4708.275 ;
        RECT 1924.110 4707.995 1924.390 4708.275 ;
        RECT 1924.730 4707.995 1925.010 4708.275 ;
        RECT 1925.350 4707.995 1925.630 4708.275 ;
        RECT 1925.970 4707.995 1926.250 4708.275 ;
        RECT 1926.590 4707.995 1926.870 4708.275 ;
        RECT 1927.210 4707.995 1927.490 4708.275 ;
        RECT 1927.830 4707.995 1928.110 4708.275 ;
        RECT 1928.450 4707.995 1928.730 4708.275 ;
        RECT 1929.070 4707.995 1929.350 4708.275 ;
        RECT 1929.690 4707.995 1929.970 4708.275 ;
        RECT 1930.310 4707.995 1930.590 4708.275 ;
        RECT 1921.010 4707.375 1921.290 4707.655 ;
        RECT 1921.630 4707.375 1921.910 4707.655 ;
        RECT 1922.250 4707.375 1922.530 4707.655 ;
        RECT 1922.870 4707.375 1923.150 4707.655 ;
        RECT 1923.490 4707.375 1923.770 4707.655 ;
        RECT 1924.110 4707.375 1924.390 4707.655 ;
        RECT 1924.730 4707.375 1925.010 4707.655 ;
        RECT 1925.350 4707.375 1925.630 4707.655 ;
        RECT 1925.970 4707.375 1926.250 4707.655 ;
        RECT 1926.590 4707.375 1926.870 4707.655 ;
        RECT 1927.210 4707.375 1927.490 4707.655 ;
        RECT 1927.830 4707.375 1928.110 4707.655 ;
        RECT 1928.450 4707.375 1928.730 4707.655 ;
        RECT 1929.070 4707.375 1929.350 4707.655 ;
        RECT 1929.690 4707.375 1929.970 4707.655 ;
        RECT 1930.310 4707.375 1930.590 4707.655 ;
        RECT 1921.010 4706.755 1921.290 4707.035 ;
        RECT 1921.630 4706.755 1921.910 4707.035 ;
        RECT 1922.250 4706.755 1922.530 4707.035 ;
        RECT 1922.870 4706.755 1923.150 4707.035 ;
        RECT 1923.490 4706.755 1923.770 4707.035 ;
        RECT 1924.110 4706.755 1924.390 4707.035 ;
        RECT 1924.730 4706.755 1925.010 4707.035 ;
        RECT 1925.350 4706.755 1925.630 4707.035 ;
        RECT 1925.970 4706.755 1926.250 4707.035 ;
        RECT 1926.590 4706.755 1926.870 4707.035 ;
        RECT 1927.210 4706.755 1927.490 4707.035 ;
        RECT 1927.830 4706.755 1928.110 4707.035 ;
        RECT 1928.450 4706.755 1928.730 4707.035 ;
        RECT 1929.070 4706.755 1929.350 4707.035 ;
        RECT 1929.690 4706.755 1929.970 4707.035 ;
        RECT 1930.310 4706.755 1930.590 4707.035 ;
        RECT 1921.010 4706.135 1921.290 4706.415 ;
        RECT 1921.630 4706.135 1921.910 4706.415 ;
        RECT 1922.250 4706.135 1922.530 4706.415 ;
        RECT 1922.870 4706.135 1923.150 4706.415 ;
        RECT 1923.490 4706.135 1923.770 4706.415 ;
        RECT 1924.110 4706.135 1924.390 4706.415 ;
        RECT 1924.730 4706.135 1925.010 4706.415 ;
        RECT 1925.350 4706.135 1925.630 4706.415 ;
        RECT 1925.970 4706.135 1926.250 4706.415 ;
        RECT 1926.590 4706.135 1926.870 4706.415 ;
        RECT 1927.210 4706.135 1927.490 4706.415 ;
        RECT 1927.830 4706.135 1928.110 4706.415 ;
        RECT 1928.450 4706.135 1928.730 4706.415 ;
        RECT 1929.070 4706.135 1929.350 4706.415 ;
        RECT 1929.690 4706.135 1929.970 4706.415 ;
        RECT 1930.310 4706.135 1930.590 4706.415 ;
        RECT 1921.010 4705.515 1921.290 4705.795 ;
        RECT 1921.630 4705.515 1921.910 4705.795 ;
        RECT 1922.250 4705.515 1922.530 4705.795 ;
        RECT 1922.870 4705.515 1923.150 4705.795 ;
        RECT 1923.490 4705.515 1923.770 4705.795 ;
        RECT 1924.110 4705.515 1924.390 4705.795 ;
        RECT 1924.730 4705.515 1925.010 4705.795 ;
        RECT 1925.350 4705.515 1925.630 4705.795 ;
        RECT 1925.970 4705.515 1926.250 4705.795 ;
        RECT 1926.590 4705.515 1926.870 4705.795 ;
        RECT 1927.210 4705.515 1927.490 4705.795 ;
        RECT 1927.830 4705.515 1928.110 4705.795 ;
        RECT 1928.450 4705.515 1928.730 4705.795 ;
        RECT 1929.070 4705.515 1929.350 4705.795 ;
        RECT 1929.690 4705.515 1929.970 4705.795 ;
        RECT 1930.310 4705.515 1930.590 4705.795 ;
        RECT 1921.010 4704.895 1921.290 4705.175 ;
        RECT 1921.630 4704.895 1921.910 4705.175 ;
        RECT 1922.250 4704.895 1922.530 4705.175 ;
        RECT 1922.870 4704.895 1923.150 4705.175 ;
        RECT 1923.490 4704.895 1923.770 4705.175 ;
        RECT 1924.110 4704.895 1924.390 4705.175 ;
        RECT 1924.730 4704.895 1925.010 4705.175 ;
        RECT 1925.350 4704.895 1925.630 4705.175 ;
        RECT 1925.970 4704.895 1926.250 4705.175 ;
        RECT 1926.590 4704.895 1926.870 4705.175 ;
        RECT 1927.210 4704.895 1927.490 4705.175 ;
        RECT 1927.830 4704.895 1928.110 4705.175 ;
        RECT 1928.450 4704.895 1928.730 4705.175 ;
        RECT 1929.070 4704.895 1929.350 4705.175 ;
        RECT 1929.690 4704.895 1929.970 4705.175 ;
        RECT 1930.310 4704.895 1930.590 4705.175 ;
        RECT 1921.010 4704.275 1921.290 4704.555 ;
        RECT 1921.630 4704.275 1921.910 4704.555 ;
        RECT 1922.250 4704.275 1922.530 4704.555 ;
        RECT 1922.870 4704.275 1923.150 4704.555 ;
        RECT 1923.490 4704.275 1923.770 4704.555 ;
        RECT 1924.110 4704.275 1924.390 4704.555 ;
        RECT 1924.730 4704.275 1925.010 4704.555 ;
        RECT 1925.350 4704.275 1925.630 4704.555 ;
        RECT 1925.970 4704.275 1926.250 4704.555 ;
        RECT 1926.590 4704.275 1926.870 4704.555 ;
        RECT 1927.210 4704.275 1927.490 4704.555 ;
        RECT 1927.830 4704.275 1928.110 4704.555 ;
        RECT 1928.450 4704.275 1928.730 4704.555 ;
        RECT 1929.070 4704.275 1929.350 4704.555 ;
        RECT 1929.690 4704.275 1929.970 4704.555 ;
        RECT 1930.310 4704.275 1930.590 4704.555 ;
        RECT 1921.010 4703.655 1921.290 4703.935 ;
        RECT 1921.630 4703.655 1921.910 4703.935 ;
        RECT 1922.250 4703.655 1922.530 4703.935 ;
        RECT 1922.870 4703.655 1923.150 4703.935 ;
        RECT 1923.490 4703.655 1923.770 4703.935 ;
        RECT 1924.110 4703.655 1924.390 4703.935 ;
        RECT 1924.730 4703.655 1925.010 4703.935 ;
        RECT 1925.350 4703.655 1925.630 4703.935 ;
        RECT 1925.970 4703.655 1926.250 4703.935 ;
        RECT 1926.590 4703.655 1926.870 4703.935 ;
        RECT 1927.210 4703.655 1927.490 4703.935 ;
        RECT 1927.830 4703.655 1928.110 4703.935 ;
        RECT 1928.450 4703.655 1928.730 4703.935 ;
        RECT 1929.070 4703.655 1929.350 4703.935 ;
        RECT 1929.690 4703.655 1929.970 4703.935 ;
        RECT 1930.310 4703.655 1930.590 4703.935 ;
        RECT 1921.010 4703.035 1921.290 4703.315 ;
        RECT 1921.630 4703.035 1921.910 4703.315 ;
        RECT 1922.250 4703.035 1922.530 4703.315 ;
        RECT 1922.870 4703.035 1923.150 4703.315 ;
        RECT 1923.490 4703.035 1923.770 4703.315 ;
        RECT 1924.110 4703.035 1924.390 4703.315 ;
        RECT 1924.730 4703.035 1925.010 4703.315 ;
        RECT 1925.350 4703.035 1925.630 4703.315 ;
        RECT 1925.970 4703.035 1926.250 4703.315 ;
        RECT 1926.590 4703.035 1926.870 4703.315 ;
        RECT 1927.210 4703.035 1927.490 4703.315 ;
        RECT 1927.830 4703.035 1928.110 4703.315 ;
        RECT 1928.450 4703.035 1928.730 4703.315 ;
        RECT 1929.070 4703.035 1929.350 4703.315 ;
        RECT 1929.690 4703.035 1929.970 4703.315 ;
        RECT 1930.310 4703.035 1930.590 4703.315 ;
        RECT 1921.010 4702.415 1921.290 4702.695 ;
        RECT 1921.630 4702.415 1921.910 4702.695 ;
        RECT 1922.250 4702.415 1922.530 4702.695 ;
        RECT 1922.870 4702.415 1923.150 4702.695 ;
        RECT 1923.490 4702.415 1923.770 4702.695 ;
        RECT 1924.110 4702.415 1924.390 4702.695 ;
        RECT 1924.730 4702.415 1925.010 4702.695 ;
        RECT 1925.350 4702.415 1925.630 4702.695 ;
        RECT 1925.970 4702.415 1926.250 4702.695 ;
        RECT 1926.590 4702.415 1926.870 4702.695 ;
        RECT 1927.210 4702.415 1927.490 4702.695 ;
        RECT 1927.830 4702.415 1928.110 4702.695 ;
        RECT 1928.450 4702.415 1928.730 4702.695 ;
        RECT 1929.070 4702.415 1929.350 4702.695 ;
        RECT 1929.690 4702.415 1929.970 4702.695 ;
        RECT 1930.310 4702.415 1930.590 4702.695 ;
        RECT 1921.010 4701.795 1921.290 4702.075 ;
        RECT 1921.630 4701.795 1921.910 4702.075 ;
        RECT 1922.250 4701.795 1922.530 4702.075 ;
        RECT 1922.870 4701.795 1923.150 4702.075 ;
        RECT 1923.490 4701.795 1923.770 4702.075 ;
        RECT 1924.110 4701.795 1924.390 4702.075 ;
        RECT 1924.730 4701.795 1925.010 4702.075 ;
        RECT 1925.350 4701.795 1925.630 4702.075 ;
        RECT 1925.970 4701.795 1926.250 4702.075 ;
        RECT 1926.590 4701.795 1926.870 4702.075 ;
        RECT 1927.210 4701.795 1927.490 4702.075 ;
        RECT 1927.830 4701.795 1928.110 4702.075 ;
        RECT 1928.450 4701.795 1928.730 4702.075 ;
        RECT 1929.070 4701.795 1929.350 4702.075 ;
        RECT 1929.690 4701.795 1929.970 4702.075 ;
        RECT 1930.310 4701.795 1930.590 4702.075 ;
        RECT 1921.010 4701.175 1921.290 4701.455 ;
        RECT 1921.630 4701.175 1921.910 4701.455 ;
        RECT 1922.250 4701.175 1922.530 4701.455 ;
        RECT 1922.870 4701.175 1923.150 4701.455 ;
        RECT 1923.490 4701.175 1923.770 4701.455 ;
        RECT 1924.110 4701.175 1924.390 4701.455 ;
        RECT 1924.730 4701.175 1925.010 4701.455 ;
        RECT 1925.350 4701.175 1925.630 4701.455 ;
        RECT 1925.970 4701.175 1926.250 4701.455 ;
        RECT 1926.590 4701.175 1926.870 4701.455 ;
        RECT 1927.210 4701.175 1927.490 4701.455 ;
        RECT 1927.830 4701.175 1928.110 4701.455 ;
        RECT 1928.450 4701.175 1928.730 4701.455 ;
        RECT 1929.070 4701.175 1929.350 4701.455 ;
        RECT 1929.690 4701.175 1929.970 4701.455 ;
        RECT 1930.310 4701.175 1930.590 4701.455 ;
        RECT 1921.010 4700.555 1921.290 4700.835 ;
        RECT 1921.630 4700.555 1921.910 4700.835 ;
        RECT 1922.250 4700.555 1922.530 4700.835 ;
        RECT 1922.870 4700.555 1923.150 4700.835 ;
        RECT 1923.490 4700.555 1923.770 4700.835 ;
        RECT 1924.110 4700.555 1924.390 4700.835 ;
        RECT 1924.730 4700.555 1925.010 4700.835 ;
        RECT 1925.350 4700.555 1925.630 4700.835 ;
        RECT 1925.970 4700.555 1926.250 4700.835 ;
        RECT 1926.590 4700.555 1926.870 4700.835 ;
        RECT 1927.210 4700.555 1927.490 4700.835 ;
        RECT 1927.830 4700.555 1928.110 4700.835 ;
        RECT 1928.450 4700.555 1928.730 4700.835 ;
        RECT 1929.070 4700.555 1929.350 4700.835 ;
        RECT 1929.690 4700.555 1929.970 4700.835 ;
        RECT 1930.310 4700.555 1930.590 4700.835 ;
        RECT 1921.010 4699.935 1921.290 4700.215 ;
        RECT 1921.630 4699.935 1921.910 4700.215 ;
        RECT 1922.250 4699.935 1922.530 4700.215 ;
        RECT 1922.870 4699.935 1923.150 4700.215 ;
        RECT 1923.490 4699.935 1923.770 4700.215 ;
        RECT 1924.110 4699.935 1924.390 4700.215 ;
        RECT 1924.730 4699.935 1925.010 4700.215 ;
        RECT 1925.350 4699.935 1925.630 4700.215 ;
        RECT 1925.970 4699.935 1926.250 4700.215 ;
        RECT 1926.590 4699.935 1926.870 4700.215 ;
        RECT 1927.210 4699.935 1927.490 4700.215 ;
        RECT 1927.830 4699.935 1928.110 4700.215 ;
        RECT 1928.450 4699.935 1928.730 4700.215 ;
        RECT 1929.070 4699.935 1929.350 4700.215 ;
        RECT 1929.690 4699.935 1929.970 4700.215 ;
        RECT 1930.310 4699.935 1930.590 4700.215 ;
        RECT 1921.010 4699.315 1921.290 4699.595 ;
        RECT 1921.630 4699.315 1921.910 4699.595 ;
        RECT 1922.250 4699.315 1922.530 4699.595 ;
        RECT 1922.870 4699.315 1923.150 4699.595 ;
        RECT 1923.490 4699.315 1923.770 4699.595 ;
        RECT 1924.110 4699.315 1924.390 4699.595 ;
        RECT 1924.730 4699.315 1925.010 4699.595 ;
        RECT 1925.350 4699.315 1925.630 4699.595 ;
        RECT 1925.970 4699.315 1926.250 4699.595 ;
        RECT 1926.590 4699.315 1926.870 4699.595 ;
        RECT 1927.210 4699.315 1927.490 4699.595 ;
        RECT 1927.830 4699.315 1928.110 4699.595 ;
        RECT 1928.450 4699.315 1928.730 4699.595 ;
        RECT 1929.070 4699.315 1929.350 4699.595 ;
        RECT 1929.690 4699.315 1929.970 4699.595 ;
        RECT 1930.310 4699.315 1930.590 4699.595 ;
        RECT 1934.540 4707.995 1934.820 4708.275 ;
        RECT 1935.160 4707.995 1935.440 4708.275 ;
        RECT 1935.780 4707.995 1936.060 4708.275 ;
        RECT 1936.400 4707.995 1936.680 4708.275 ;
        RECT 1937.020 4707.995 1937.300 4708.275 ;
        RECT 1937.640 4707.995 1937.920 4708.275 ;
        RECT 1938.260 4707.995 1938.540 4708.275 ;
        RECT 1938.880 4707.995 1939.160 4708.275 ;
        RECT 1939.500 4707.995 1939.780 4708.275 ;
        RECT 1940.120 4707.995 1940.400 4708.275 ;
        RECT 1940.740 4707.995 1941.020 4708.275 ;
        RECT 1941.360 4707.995 1941.640 4708.275 ;
        RECT 1941.980 4707.995 1942.260 4708.275 ;
        RECT 1942.600 4707.995 1942.880 4708.275 ;
        RECT 1943.220 4707.995 1943.500 4708.275 ;
        RECT 1943.840 4707.995 1944.120 4708.275 ;
        RECT 1934.540 4707.375 1934.820 4707.655 ;
        RECT 1935.160 4707.375 1935.440 4707.655 ;
        RECT 1935.780 4707.375 1936.060 4707.655 ;
        RECT 1936.400 4707.375 1936.680 4707.655 ;
        RECT 1937.020 4707.375 1937.300 4707.655 ;
        RECT 1937.640 4707.375 1937.920 4707.655 ;
        RECT 1938.260 4707.375 1938.540 4707.655 ;
        RECT 1938.880 4707.375 1939.160 4707.655 ;
        RECT 1939.500 4707.375 1939.780 4707.655 ;
        RECT 1940.120 4707.375 1940.400 4707.655 ;
        RECT 1940.740 4707.375 1941.020 4707.655 ;
        RECT 1941.360 4707.375 1941.640 4707.655 ;
        RECT 1941.980 4707.375 1942.260 4707.655 ;
        RECT 1942.600 4707.375 1942.880 4707.655 ;
        RECT 1943.220 4707.375 1943.500 4707.655 ;
        RECT 1943.840 4707.375 1944.120 4707.655 ;
        RECT 1934.540 4706.755 1934.820 4707.035 ;
        RECT 1935.160 4706.755 1935.440 4707.035 ;
        RECT 1935.780 4706.755 1936.060 4707.035 ;
        RECT 1936.400 4706.755 1936.680 4707.035 ;
        RECT 1937.020 4706.755 1937.300 4707.035 ;
        RECT 1937.640 4706.755 1937.920 4707.035 ;
        RECT 1938.260 4706.755 1938.540 4707.035 ;
        RECT 1938.880 4706.755 1939.160 4707.035 ;
        RECT 1939.500 4706.755 1939.780 4707.035 ;
        RECT 1940.120 4706.755 1940.400 4707.035 ;
        RECT 1940.740 4706.755 1941.020 4707.035 ;
        RECT 1941.360 4706.755 1941.640 4707.035 ;
        RECT 1941.980 4706.755 1942.260 4707.035 ;
        RECT 1942.600 4706.755 1942.880 4707.035 ;
        RECT 1943.220 4706.755 1943.500 4707.035 ;
        RECT 1943.840 4706.755 1944.120 4707.035 ;
        RECT 1934.540 4706.135 1934.820 4706.415 ;
        RECT 1935.160 4706.135 1935.440 4706.415 ;
        RECT 1935.780 4706.135 1936.060 4706.415 ;
        RECT 1936.400 4706.135 1936.680 4706.415 ;
        RECT 1937.020 4706.135 1937.300 4706.415 ;
        RECT 1937.640 4706.135 1937.920 4706.415 ;
        RECT 1938.260 4706.135 1938.540 4706.415 ;
        RECT 1938.880 4706.135 1939.160 4706.415 ;
        RECT 1939.500 4706.135 1939.780 4706.415 ;
        RECT 1940.120 4706.135 1940.400 4706.415 ;
        RECT 1940.740 4706.135 1941.020 4706.415 ;
        RECT 1941.360 4706.135 1941.640 4706.415 ;
        RECT 1941.980 4706.135 1942.260 4706.415 ;
        RECT 1942.600 4706.135 1942.880 4706.415 ;
        RECT 1943.220 4706.135 1943.500 4706.415 ;
        RECT 1943.840 4706.135 1944.120 4706.415 ;
        RECT 1934.540 4705.515 1934.820 4705.795 ;
        RECT 1935.160 4705.515 1935.440 4705.795 ;
        RECT 1935.780 4705.515 1936.060 4705.795 ;
        RECT 1936.400 4705.515 1936.680 4705.795 ;
        RECT 1937.020 4705.515 1937.300 4705.795 ;
        RECT 1937.640 4705.515 1937.920 4705.795 ;
        RECT 1938.260 4705.515 1938.540 4705.795 ;
        RECT 1938.880 4705.515 1939.160 4705.795 ;
        RECT 1939.500 4705.515 1939.780 4705.795 ;
        RECT 1940.120 4705.515 1940.400 4705.795 ;
        RECT 1940.740 4705.515 1941.020 4705.795 ;
        RECT 1941.360 4705.515 1941.640 4705.795 ;
        RECT 1941.980 4705.515 1942.260 4705.795 ;
        RECT 1942.600 4705.515 1942.880 4705.795 ;
        RECT 1943.220 4705.515 1943.500 4705.795 ;
        RECT 1943.840 4705.515 1944.120 4705.795 ;
        RECT 1934.540 4704.895 1934.820 4705.175 ;
        RECT 1935.160 4704.895 1935.440 4705.175 ;
        RECT 1935.780 4704.895 1936.060 4705.175 ;
        RECT 1936.400 4704.895 1936.680 4705.175 ;
        RECT 1937.020 4704.895 1937.300 4705.175 ;
        RECT 1937.640 4704.895 1937.920 4705.175 ;
        RECT 1938.260 4704.895 1938.540 4705.175 ;
        RECT 1938.880 4704.895 1939.160 4705.175 ;
        RECT 1939.500 4704.895 1939.780 4705.175 ;
        RECT 1940.120 4704.895 1940.400 4705.175 ;
        RECT 1940.740 4704.895 1941.020 4705.175 ;
        RECT 1941.360 4704.895 1941.640 4705.175 ;
        RECT 1941.980 4704.895 1942.260 4705.175 ;
        RECT 1942.600 4704.895 1942.880 4705.175 ;
        RECT 1943.220 4704.895 1943.500 4705.175 ;
        RECT 1943.840 4704.895 1944.120 4705.175 ;
        RECT 1934.540 4704.275 1934.820 4704.555 ;
        RECT 1935.160 4704.275 1935.440 4704.555 ;
        RECT 1935.780 4704.275 1936.060 4704.555 ;
        RECT 1936.400 4704.275 1936.680 4704.555 ;
        RECT 1937.020 4704.275 1937.300 4704.555 ;
        RECT 1937.640 4704.275 1937.920 4704.555 ;
        RECT 1938.260 4704.275 1938.540 4704.555 ;
        RECT 1938.880 4704.275 1939.160 4704.555 ;
        RECT 1939.500 4704.275 1939.780 4704.555 ;
        RECT 1940.120 4704.275 1940.400 4704.555 ;
        RECT 1940.740 4704.275 1941.020 4704.555 ;
        RECT 1941.360 4704.275 1941.640 4704.555 ;
        RECT 1941.980 4704.275 1942.260 4704.555 ;
        RECT 1942.600 4704.275 1942.880 4704.555 ;
        RECT 1943.220 4704.275 1943.500 4704.555 ;
        RECT 1943.840 4704.275 1944.120 4704.555 ;
        RECT 1934.540 4703.655 1934.820 4703.935 ;
        RECT 1935.160 4703.655 1935.440 4703.935 ;
        RECT 1935.780 4703.655 1936.060 4703.935 ;
        RECT 1936.400 4703.655 1936.680 4703.935 ;
        RECT 1937.020 4703.655 1937.300 4703.935 ;
        RECT 1937.640 4703.655 1937.920 4703.935 ;
        RECT 1938.260 4703.655 1938.540 4703.935 ;
        RECT 1938.880 4703.655 1939.160 4703.935 ;
        RECT 1939.500 4703.655 1939.780 4703.935 ;
        RECT 1940.120 4703.655 1940.400 4703.935 ;
        RECT 1940.740 4703.655 1941.020 4703.935 ;
        RECT 1941.360 4703.655 1941.640 4703.935 ;
        RECT 1941.980 4703.655 1942.260 4703.935 ;
        RECT 1942.600 4703.655 1942.880 4703.935 ;
        RECT 1943.220 4703.655 1943.500 4703.935 ;
        RECT 1943.840 4703.655 1944.120 4703.935 ;
        RECT 1934.540 4703.035 1934.820 4703.315 ;
        RECT 1935.160 4703.035 1935.440 4703.315 ;
        RECT 1935.780 4703.035 1936.060 4703.315 ;
        RECT 1936.400 4703.035 1936.680 4703.315 ;
        RECT 1937.020 4703.035 1937.300 4703.315 ;
        RECT 1937.640 4703.035 1937.920 4703.315 ;
        RECT 1938.260 4703.035 1938.540 4703.315 ;
        RECT 1938.880 4703.035 1939.160 4703.315 ;
        RECT 1939.500 4703.035 1939.780 4703.315 ;
        RECT 1940.120 4703.035 1940.400 4703.315 ;
        RECT 1940.740 4703.035 1941.020 4703.315 ;
        RECT 1941.360 4703.035 1941.640 4703.315 ;
        RECT 1941.980 4703.035 1942.260 4703.315 ;
        RECT 1942.600 4703.035 1942.880 4703.315 ;
        RECT 1943.220 4703.035 1943.500 4703.315 ;
        RECT 1943.840 4703.035 1944.120 4703.315 ;
        RECT 1934.540 4702.415 1934.820 4702.695 ;
        RECT 1935.160 4702.415 1935.440 4702.695 ;
        RECT 1935.780 4702.415 1936.060 4702.695 ;
        RECT 1936.400 4702.415 1936.680 4702.695 ;
        RECT 1937.020 4702.415 1937.300 4702.695 ;
        RECT 1937.640 4702.415 1937.920 4702.695 ;
        RECT 1938.260 4702.415 1938.540 4702.695 ;
        RECT 1938.880 4702.415 1939.160 4702.695 ;
        RECT 1939.500 4702.415 1939.780 4702.695 ;
        RECT 1940.120 4702.415 1940.400 4702.695 ;
        RECT 1940.740 4702.415 1941.020 4702.695 ;
        RECT 1941.360 4702.415 1941.640 4702.695 ;
        RECT 1941.980 4702.415 1942.260 4702.695 ;
        RECT 1942.600 4702.415 1942.880 4702.695 ;
        RECT 1943.220 4702.415 1943.500 4702.695 ;
        RECT 1943.840 4702.415 1944.120 4702.695 ;
        RECT 1934.540 4701.795 1934.820 4702.075 ;
        RECT 1935.160 4701.795 1935.440 4702.075 ;
        RECT 1935.780 4701.795 1936.060 4702.075 ;
        RECT 1936.400 4701.795 1936.680 4702.075 ;
        RECT 1937.020 4701.795 1937.300 4702.075 ;
        RECT 1937.640 4701.795 1937.920 4702.075 ;
        RECT 1938.260 4701.795 1938.540 4702.075 ;
        RECT 1938.880 4701.795 1939.160 4702.075 ;
        RECT 1939.500 4701.795 1939.780 4702.075 ;
        RECT 1940.120 4701.795 1940.400 4702.075 ;
        RECT 1940.740 4701.795 1941.020 4702.075 ;
        RECT 1941.360 4701.795 1941.640 4702.075 ;
        RECT 1941.980 4701.795 1942.260 4702.075 ;
        RECT 1942.600 4701.795 1942.880 4702.075 ;
        RECT 1943.220 4701.795 1943.500 4702.075 ;
        RECT 1943.840 4701.795 1944.120 4702.075 ;
        RECT 1934.540 4701.175 1934.820 4701.455 ;
        RECT 1935.160 4701.175 1935.440 4701.455 ;
        RECT 1935.780 4701.175 1936.060 4701.455 ;
        RECT 1936.400 4701.175 1936.680 4701.455 ;
        RECT 1937.020 4701.175 1937.300 4701.455 ;
        RECT 1937.640 4701.175 1937.920 4701.455 ;
        RECT 1938.260 4701.175 1938.540 4701.455 ;
        RECT 1938.880 4701.175 1939.160 4701.455 ;
        RECT 1939.500 4701.175 1939.780 4701.455 ;
        RECT 1940.120 4701.175 1940.400 4701.455 ;
        RECT 1940.740 4701.175 1941.020 4701.455 ;
        RECT 1941.360 4701.175 1941.640 4701.455 ;
        RECT 1941.980 4701.175 1942.260 4701.455 ;
        RECT 1942.600 4701.175 1942.880 4701.455 ;
        RECT 1943.220 4701.175 1943.500 4701.455 ;
        RECT 1943.840 4701.175 1944.120 4701.455 ;
        RECT 1934.540 4700.555 1934.820 4700.835 ;
        RECT 1935.160 4700.555 1935.440 4700.835 ;
        RECT 1935.780 4700.555 1936.060 4700.835 ;
        RECT 1936.400 4700.555 1936.680 4700.835 ;
        RECT 1937.020 4700.555 1937.300 4700.835 ;
        RECT 1937.640 4700.555 1937.920 4700.835 ;
        RECT 1938.260 4700.555 1938.540 4700.835 ;
        RECT 1938.880 4700.555 1939.160 4700.835 ;
        RECT 1939.500 4700.555 1939.780 4700.835 ;
        RECT 1940.120 4700.555 1940.400 4700.835 ;
        RECT 1940.740 4700.555 1941.020 4700.835 ;
        RECT 1941.360 4700.555 1941.640 4700.835 ;
        RECT 1941.980 4700.555 1942.260 4700.835 ;
        RECT 1942.600 4700.555 1942.880 4700.835 ;
        RECT 1943.220 4700.555 1943.500 4700.835 ;
        RECT 1943.840 4700.555 1944.120 4700.835 ;
        RECT 1934.540 4699.935 1934.820 4700.215 ;
        RECT 1935.160 4699.935 1935.440 4700.215 ;
        RECT 1935.780 4699.935 1936.060 4700.215 ;
        RECT 1936.400 4699.935 1936.680 4700.215 ;
        RECT 1937.020 4699.935 1937.300 4700.215 ;
        RECT 1937.640 4699.935 1937.920 4700.215 ;
        RECT 1938.260 4699.935 1938.540 4700.215 ;
        RECT 1938.880 4699.935 1939.160 4700.215 ;
        RECT 1939.500 4699.935 1939.780 4700.215 ;
        RECT 1940.120 4699.935 1940.400 4700.215 ;
        RECT 1940.740 4699.935 1941.020 4700.215 ;
        RECT 1941.360 4699.935 1941.640 4700.215 ;
        RECT 1941.980 4699.935 1942.260 4700.215 ;
        RECT 1942.600 4699.935 1942.880 4700.215 ;
        RECT 1943.220 4699.935 1943.500 4700.215 ;
        RECT 1943.840 4699.935 1944.120 4700.215 ;
        RECT 1934.540 4699.315 1934.820 4699.595 ;
        RECT 1935.160 4699.315 1935.440 4699.595 ;
        RECT 1935.780 4699.315 1936.060 4699.595 ;
        RECT 1936.400 4699.315 1936.680 4699.595 ;
        RECT 1937.020 4699.315 1937.300 4699.595 ;
        RECT 1937.640 4699.315 1937.920 4699.595 ;
        RECT 1938.260 4699.315 1938.540 4699.595 ;
        RECT 1938.880 4699.315 1939.160 4699.595 ;
        RECT 1939.500 4699.315 1939.780 4699.595 ;
        RECT 1940.120 4699.315 1940.400 4699.595 ;
        RECT 1940.740 4699.315 1941.020 4699.595 ;
        RECT 1941.360 4699.315 1941.640 4699.595 ;
        RECT 1941.980 4699.315 1942.260 4699.595 ;
        RECT 1942.600 4699.315 1942.880 4699.595 ;
        RECT 1943.220 4699.315 1943.500 4699.595 ;
        RECT 1943.840 4699.315 1944.120 4699.595 ;
        RECT 1946.390 4707.995 1946.670 4708.275 ;
        RECT 1947.010 4707.995 1947.290 4708.275 ;
        RECT 1947.630 4707.995 1947.910 4708.275 ;
        RECT 1948.250 4707.995 1948.530 4708.275 ;
        RECT 1948.870 4707.995 1949.150 4708.275 ;
        RECT 1949.490 4707.995 1949.770 4708.275 ;
        RECT 1950.110 4707.995 1950.390 4708.275 ;
        RECT 1950.730 4707.995 1951.010 4708.275 ;
        RECT 1951.350 4707.995 1951.630 4708.275 ;
        RECT 1951.970 4707.995 1952.250 4708.275 ;
        RECT 1952.590 4707.995 1952.870 4708.275 ;
        RECT 1953.210 4707.995 1953.490 4708.275 ;
        RECT 1953.830 4707.995 1954.110 4708.275 ;
        RECT 1954.450 4707.995 1954.730 4708.275 ;
        RECT 1955.070 4707.995 1955.350 4708.275 ;
        RECT 1955.690 4707.995 1955.970 4708.275 ;
        RECT 1946.390 4707.375 1946.670 4707.655 ;
        RECT 1947.010 4707.375 1947.290 4707.655 ;
        RECT 1947.630 4707.375 1947.910 4707.655 ;
        RECT 1948.250 4707.375 1948.530 4707.655 ;
        RECT 1948.870 4707.375 1949.150 4707.655 ;
        RECT 1949.490 4707.375 1949.770 4707.655 ;
        RECT 1950.110 4707.375 1950.390 4707.655 ;
        RECT 1950.730 4707.375 1951.010 4707.655 ;
        RECT 1951.350 4707.375 1951.630 4707.655 ;
        RECT 1951.970 4707.375 1952.250 4707.655 ;
        RECT 1952.590 4707.375 1952.870 4707.655 ;
        RECT 1953.210 4707.375 1953.490 4707.655 ;
        RECT 1953.830 4707.375 1954.110 4707.655 ;
        RECT 1954.450 4707.375 1954.730 4707.655 ;
        RECT 1955.070 4707.375 1955.350 4707.655 ;
        RECT 1955.690 4707.375 1955.970 4707.655 ;
        RECT 1946.390 4706.755 1946.670 4707.035 ;
        RECT 1947.010 4706.755 1947.290 4707.035 ;
        RECT 1947.630 4706.755 1947.910 4707.035 ;
        RECT 1948.250 4706.755 1948.530 4707.035 ;
        RECT 1948.870 4706.755 1949.150 4707.035 ;
        RECT 1949.490 4706.755 1949.770 4707.035 ;
        RECT 1950.110 4706.755 1950.390 4707.035 ;
        RECT 1950.730 4706.755 1951.010 4707.035 ;
        RECT 1951.350 4706.755 1951.630 4707.035 ;
        RECT 1951.970 4706.755 1952.250 4707.035 ;
        RECT 1952.590 4706.755 1952.870 4707.035 ;
        RECT 1953.210 4706.755 1953.490 4707.035 ;
        RECT 1953.830 4706.755 1954.110 4707.035 ;
        RECT 1954.450 4706.755 1954.730 4707.035 ;
        RECT 1955.070 4706.755 1955.350 4707.035 ;
        RECT 1955.690 4706.755 1955.970 4707.035 ;
        RECT 1946.390 4706.135 1946.670 4706.415 ;
        RECT 1947.010 4706.135 1947.290 4706.415 ;
        RECT 1947.630 4706.135 1947.910 4706.415 ;
        RECT 1948.250 4706.135 1948.530 4706.415 ;
        RECT 1948.870 4706.135 1949.150 4706.415 ;
        RECT 1949.490 4706.135 1949.770 4706.415 ;
        RECT 1950.110 4706.135 1950.390 4706.415 ;
        RECT 1950.730 4706.135 1951.010 4706.415 ;
        RECT 1951.350 4706.135 1951.630 4706.415 ;
        RECT 1951.970 4706.135 1952.250 4706.415 ;
        RECT 1952.590 4706.135 1952.870 4706.415 ;
        RECT 1953.210 4706.135 1953.490 4706.415 ;
        RECT 1953.830 4706.135 1954.110 4706.415 ;
        RECT 1954.450 4706.135 1954.730 4706.415 ;
        RECT 1955.070 4706.135 1955.350 4706.415 ;
        RECT 1955.690 4706.135 1955.970 4706.415 ;
        RECT 1946.390 4705.515 1946.670 4705.795 ;
        RECT 1947.010 4705.515 1947.290 4705.795 ;
        RECT 1947.630 4705.515 1947.910 4705.795 ;
        RECT 1948.250 4705.515 1948.530 4705.795 ;
        RECT 1948.870 4705.515 1949.150 4705.795 ;
        RECT 1949.490 4705.515 1949.770 4705.795 ;
        RECT 1950.110 4705.515 1950.390 4705.795 ;
        RECT 1950.730 4705.515 1951.010 4705.795 ;
        RECT 1951.350 4705.515 1951.630 4705.795 ;
        RECT 1951.970 4705.515 1952.250 4705.795 ;
        RECT 1952.590 4705.515 1952.870 4705.795 ;
        RECT 1953.210 4705.515 1953.490 4705.795 ;
        RECT 1953.830 4705.515 1954.110 4705.795 ;
        RECT 1954.450 4705.515 1954.730 4705.795 ;
        RECT 1955.070 4705.515 1955.350 4705.795 ;
        RECT 1955.690 4705.515 1955.970 4705.795 ;
        RECT 1946.390 4704.895 1946.670 4705.175 ;
        RECT 1947.010 4704.895 1947.290 4705.175 ;
        RECT 1947.630 4704.895 1947.910 4705.175 ;
        RECT 1948.250 4704.895 1948.530 4705.175 ;
        RECT 1948.870 4704.895 1949.150 4705.175 ;
        RECT 1949.490 4704.895 1949.770 4705.175 ;
        RECT 1950.110 4704.895 1950.390 4705.175 ;
        RECT 1950.730 4704.895 1951.010 4705.175 ;
        RECT 1951.350 4704.895 1951.630 4705.175 ;
        RECT 1951.970 4704.895 1952.250 4705.175 ;
        RECT 1952.590 4704.895 1952.870 4705.175 ;
        RECT 1953.210 4704.895 1953.490 4705.175 ;
        RECT 1953.830 4704.895 1954.110 4705.175 ;
        RECT 1954.450 4704.895 1954.730 4705.175 ;
        RECT 1955.070 4704.895 1955.350 4705.175 ;
        RECT 1955.690 4704.895 1955.970 4705.175 ;
        RECT 1946.390 4704.275 1946.670 4704.555 ;
        RECT 1947.010 4704.275 1947.290 4704.555 ;
        RECT 1947.630 4704.275 1947.910 4704.555 ;
        RECT 1948.250 4704.275 1948.530 4704.555 ;
        RECT 1948.870 4704.275 1949.150 4704.555 ;
        RECT 1949.490 4704.275 1949.770 4704.555 ;
        RECT 1950.110 4704.275 1950.390 4704.555 ;
        RECT 1950.730 4704.275 1951.010 4704.555 ;
        RECT 1951.350 4704.275 1951.630 4704.555 ;
        RECT 1951.970 4704.275 1952.250 4704.555 ;
        RECT 1952.590 4704.275 1952.870 4704.555 ;
        RECT 1953.210 4704.275 1953.490 4704.555 ;
        RECT 1953.830 4704.275 1954.110 4704.555 ;
        RECT 1954.450 4704.275 1954.730 4704.555 ;
        RECT 1955.070 4704.275 1955.350 4704.555 ;
        RECT 1955.690 4704.275 1955.970 4704.555 ;
        RECT 1946.390 4703.655 1946.670 4703.935 ;
        RECT 1947.010 4703.655 1947.290 4703.935 ;
        RECT 1947.630 4703.655 1947.910 4703.935 ;
        RECT 1948.250 4703.655 1948.530 4703.935 ;
        RECT 1948.870 4703.655 1949.150 4703.935 ;
        RECT 1949.490 4703.655 1949.770 4703.935 ;
        RECT 1950.110 4703.655 1950.390 4703.935 ;
        RECT 1950.730 4703.655 1951.010 4703.935 ;
        RECT 1951.350 4703.655 1951.630 4703.935 ;
        RECT 1951.970 4703.655 1952.250 4703.935 ;
        RECT 1952.590 4703.655 1952.870 4703.935 ;
        RECT 1953.210 4703.655 1953.490 4703.935 ;
        RECT 1953.830 4703.655 1954.110 4703.935 ;
        RECT 1954.450 4703.655 1954.730 4703.935 ;
        RECT 1955.070 4703.655 1955.350 4703.935 ;
        RECT 1955.690 4703.655 1955.970 4703.935 ;
        RECT 1946.390 4703.035 1946.670 4703.315 ;
        RECT 1947.010 4703.035 1947.290 4703.315 ;
        RECT 1947.630 4703.035 1947.910 4703.315 ;
        RECT 1948.250 4703.035 1948.530 4703.315 ;
        RECT 1948.870 4703.035 1949.150 4703.315 ;
        RECT 1949.490 4703.035 1949.770 4703.315 ;
        RECT 1950.110 4703.035 1950.390 4703.315 ;
        RECT 1950.730 4703.035 1951.010 4703.315 ;
        RECT 1951.350 4703.035 1951.630 4703.315 ;
        RECT 1951.970 4703.035 1952.250 4703.315 ;
        RECT 1952.590 4703.035 1952.870 4703.315 ;
        RECT 1953.210 4703.035 1953.490 4703.315 ;
        RECT 1953.830 4703.035 1954.110 4703.315 ;
        RECT 1954.450 4703.035 1954.730 4703.315 ;
        RECT 1955.070 4703.035 1955.350 4703.315 ;
        RECT 1955.690 4703.035 1955.970 4703.315 ;
        RECT 1946.390 4702.415 1946.670 4702.695 ;
        RECT 1947.010 4702.415 1947.290 4702.695 ;
        RECT 1947.630 4702.415 1947.910 4702.695 ;
        RECT 1948.250 4702.415 1948.530 4702.695 ;
        RECT 1948.870 4702.415 1949.150 4702.695 ;
        RECT 1949.490 4702.415 1949.770 4702.695 ;
        RECT 1950.110 4702.415 1950.390 4702.695 ;
        RECT 1950.730 4702.415 1951.010 4702.695 ;
        RECT 1951.350 4702.415 1951.630 4702.695 ;
        RECT 1951.970 4702.415 1952.250 4702.695 ;
        RECT 1952.590 4702.415 1952.870 4702.695 ;
        RECT 1953.210 4702.415 1953.490 4702.695 ;
        RECT 1953.830 4702.415 1954.110 4702.695 ;
        RECT 1954.450 4702.415 1954.730 4702.695 ;
        RECT 1955.070 4702.415 1955.350 4702.695 ;
        RECT 1955.690 4702.415 1955.970 4702.695 ;
        RECT 1946.390 4701.795 1946.670 4702.075 ;
        RECT 1947.010 4701.795 1947.290 4702.075 ;
        RECT 1947.630 4701.795 1947.910 4702.075 ;
        RECT 1948.250 4701.795 1948.530 4702.075 ;
        RECT 1948.870 4701.795 1949.150 4702.075 ;
        RECT 1949.490 4701.795 1949.770 4702.075 ;
        RECT 1950.110 4701.795 1950.390 4702.075 ;
        RECT 1950.730 4701.795 1951.010 4702.075 ;
        RECT 1951.350 4701.795 1951.630 4702.075 ;
        RECT 1951.970 4701.795 1952.250 4702.075 ;
        RECT 1952.590 4701.795 1952.870 4702.075 ;
        RECT 1953.210 4701.795 1953.490 4702.075 ;
        RECT 1953.830 4701.795 1954.110 4702.075 ;
        RECT 1954.450 4701.795 1954.730 4702.075 ;
        RECT 1955.070 4701.795 1955.350 4702.075 ;
        RECT 1955.690 4701.795 1955.970 4702.075 ;
        RECT 1946.390 4701.175 1946.670 4701.455 ;
        RECT 1947.010 4701.175 1947.290 4701.455 ;
        RECT 1947.630 4701.175 1947.910 4701.455 ;
        RECT 1948.250 4701.175 1948.530 4701.455 ;
        RECT 1948.870 4701.175 1949.150 4701.455 ;
        RECT 1949.490 4701.175 1949.770 4701.455 ;
        RECT 1950.110 4701.175 1950.390 4701.455 ;
        RECT 1950.730 4701.175 1951.010 4701.455 ;
        RECT 1951.350 4701.175 1951.630 4701.455 ;
        RECT 1951.970 4701.175 1952.250 4701.455 ;
        RECT 1952.590 4701.175 1952.870 4701.455 ;
        RECT 1953.210 4701.175 1953.490 4701.455 ;
        RECT 1953.830 4701.175 1954.110 4701.455 ;
        RECT 1954.450 4701.175 1954.730 4701.455 ;
        RECT 1955.070 4701.175 1955.350 4701.455 ;
        RECT 1955.690 4701.175 1955.970 4701.455 ;
        RECT 1946.390 4700.555 1946.670 4700.835 ;
        RECT 1947.010 4700.555 1947.290 4700.835 ;
        RECT 1947.630 4700.555 1947.910 4700.835 ;
        RECT 1948.250 4700.555 1948.530 4700.835 ;
        RECT 1948.870 4700.555 1949.150 4700.835 ;
        RECT 1949.490 4700.555 1949.770 4700.835 ;
        RECT 1950.110 4700.555 1950.390 4700.835 ;
        RECT 1950.730 4700.555 1951.010 4700.835 ;
        RECT 1951.350 4700.555 1951.630 4700.835 ;
        RECT 1951.970 4700.555 1952.250 4700.835 ;
        RECT 1952.590 4700.555 1952.870 4700.835 ;
        RECT 1953.210 4700.555 1953.490 4700.835 ;
        RECT 1953.830 4700.555 1954.110 4700.835 ;
        RECT 1954.450 4700.555 1954.730 4700.835 ;
        RECT 1955.070 4700.555 1955.350 4700.835 ;
        RECT 1955.690 4700.555 1955.970 4700.835 ;
        RECT 1946.390 4699.935 1946.670 4700.215 ;
        RECT 1947.010 4699.935 1947.290 4700.215 ;
        RECT 1947.630 4699.935 1947.910 4700.215 ;
        RECT 1948.250 4699.935 1948.530 4700.215 ;
        RECT 1948.870 4699.935 1949.150 4700.215 ;
        RECT 1949.490 4699.935 1949.770 4700.215 ;
        RECT 1950.110 4699.935 1950.390 4700.215 ;
        RECT 1950.730 4699.935 1951.010 4700.215 ;
        RECT 1951.350 4699.935 1951.630 4700.215 ;
        RECT 1951.970 4699.935 1952.250 4700.215 ;
        RECT 1952.590 4699.935 1952.870 4700.215 ;
        RECT 1953.210 4699.935 1953.490 4700.215 ;
        RECT 1953.830 4699.935 1954.110 4700.215 ;
        RECT 1954.450 4699.935 1954.730 4700.215 ;
        RECT 1955.070 4699.935 1955.350 4700.215 ;
        RECT 1955.690 4699.935 1955.970 4700.215 ;
        RECT 1946.390 4699.315 1946.670 4699.595 ;
        RECT 1947.010 4699.315 1947.290 4699.595 ;
        RECT 1947.630 4699.315 1947.910 4699.595 ;
        RECT 1948.250 4699.315 1948.530 4699.595 ;
        RECT 1948.870 4699.315 1949.150 4699.595 ;
        RECT 1949.490 4699.315 1949.770 4699.595 ;
        RECT 1950.110 4699.315 1950.390 4699.595 ;
        RECT 1950.730 4699.315 1951.010 4699.595 ;
        RECT 1951.350 4699.315 1951.630 4699.595 ;
        RECT 1951.970 4699.315 1952.250 4699.595 ;
        RECT 1952.590 4699.315 1952.870 4699.595 ;
        RECT 1953.210 4699.315 1953.490 4699.595 ;
        RECT 1953.830 4699.315 1954.110 4699.595 ;
        RECT 1954.450 4699.315 1954.730 4699.595 ;
        RECT 1955.070 4699.315 1955.350 4699.595 ;
        RECT 1955.690 4699.315 1955.970 4699.595 ;
        RECT 1959.410 4707.995 1959.690 4708.275 ;
        RECT 1960.030 4707.995 1960.310 4708.275 ;
        RECT 1960.650 4707.995 1960.930 4708.275 ;
        RECT 1961.270 4707.995 1961.550 4708.275 ;
        RECT 1961.890 4707.995 1962.170 4708.275 ;
        RECT 1962.510 4707.995 1962.790 4708.275 ;
        RECT 1963.130 4707.995 1963.410 4708.275 ;
        RECT 1963.750 4707.995 1964.030 4708.275 ;
        RECT 1964.370 4707.995 1964.650 4708.275 ;
        RECT 1964.990 4707.995 1965.270 4708.275 ;
        RECT 1965.610 4707.995 1965.890 4708.275 ;
        RECT 1966.230 4707.995 1966.510 4708.275 ;
        RECT 1966.850 4707.995 1967.130 4708.275 ;
        RECT 1967.470 4707.995 1967.750 4708.275 ;
        RECT 1968.090 4707.995 1968.370 4708.275 ;
        RECT 1959.410 4707.375 1959.690 4707.655 ;
        RECT 1960.030 4707.375 1960.310 4707.655 ;
        RECT 1960.650 4707.375 1960.930 4707.655 ;
        RECT 1961.270 4707.375 1961.550 4707.655 ;
        RECT 1961.890 4707.375 1962.170 4707.655 ;
        RECT 1962.510 4707.375 1962.790 4707.655 ;
        RECT 1963.130 4707.375 1963.410 4707.655 ;
        RECT 1963.750 4707.375 1964.030 4707.655 ;
        RECT 1964.370 4707.375 1964.650 4707.655 ;
        RECT 1964.990 4707.375 1965.270 4707.655 ;
        RECT 1965.610 4707.375 1965.890 4707.655 ;
        RECT 1966.230 4707.375 1966.510 4707.655 ;
        RECT 1966.850 4707.375 1967.130 4707.655 ;
        RECT 1967.470 4707.375 1967.750 4707.655 ;
        RECT 1968.090 4707.375 1968.370 4707.655 ;
        RECT 1959.410 4706.755 1959.690 4707.035 ;
        RECT 1960.030 4706.755 1960.310 4707.035 ;
        RECT 1960.650 4706.755 1960.930 4707.035 ;
        RECT 1961.270 4706.755 1961.550 4707.035 ;
        RECT 1961.890 4706.755 1962.170 4707.035 ;
        RECT 1962.510 4706.755 1962.790 4707.035 ;
        RECT 1963.130 4706.755 1963.410 4707.035 ;
        RECT 1963.750 4706.755 1964.030 4707.035 ;
        RECT 1964.370 4706.755 1964.650 4707.035 ;
        RECT 1964.990 4706.755 1965.270 4707.035 ;
        RECT 1965.610 4706.755 1965.890 4707.035 ;
        RECT 1966.230 4706.755 1966.510 4707.035 ;
        RECT 1966.850 4706.755 1967.130 4707.035 ;
        RECT 1967.470 4706.755 1967.750 4707.035 ;
        RECT 1968.090 4706.755 1968.370 4707.035 ;
        RECT 1959.410 4706.135 1959.690 4706.415 ;
        RECT 1960.030 4706.135 1960.310 4706.415 ;
        RECT 1960.650 4706.135 1960.930 4706.415 ;
        RECT 1961.270 4706.135 1961.550 4706.415 ;
        RECT 1961.890 4706.135 1962.170 4706.415 ;
        RECT 1962.510 4706.135 1962.790 4706.415 ;
        RECT 1963.130 4706.135 1963.410 4706.415 ;
        RECT 1963.750 4706.135 1964.030 4706.415 ;
        RECT 1964.370 4706.135 1964.650 4706.415 ;
        RECT 1964.990 4706.135 1965.270 4706.415 ;
        RECT 1965.610 4706.135 1965.890 4706.415 ;
        RECT 1966.230 4706.135 1966.510 4706.415 ;
        RECT 1966.850 4706.135 1967.130 4706.415 ;
        RECT 1967.470 4706.135 1967.750 4706.415 ;
        RECT 1968.090 4706.135 1968.370 4706.415 ;
        RECT 1959.410 4705.515 1959.690 4705.795 ;
        RECT 1960.030 4705.515 1960.310 4705.795 ;
        RECT 1960.650 4705.515 1960.930 4705.795 ;
        RECT 1961.270 4705.515 1961.550 4705.795 ;
        RECT 1961.890 4705.515 1962.170 4705.795 ;
        RECT 1962.510 4705.515 1962.790 4705.795 ;
        RECT 1963.130 4705.515 1963.410 4705.795 ;
        RECT 1963.750 4705.515 1964.030 4705.795 ;
        RECT 1964.370 4705.515 1964.650 4705.795 ;
        RECT 1964.990 4705.515 1965.270 4705.795 ;
        RECT 1965.610 4705.515 1965.890 4705.795 ;
        RECT 1966.230 4705.515 1966.510 4705.795 ;
        RECT 1966.850 4705.515 1967.130 4705.795 ;
        RECT 1967.470 4705.515 1967.750 4705.795 ;
        RECT 1968.090 4705.515 1968.370 4705.795 ;
        RECT 1959.410 4704.895 1959.690 4705.175 ;
        RECT 1960.030 4704.895 1960.310 4705.175 ;
        RECT 1960.650 4704.895 1960.930 4705.175 ;
        RECT 1961.270 4704.895 1961.550 4705.175 ;
        RECT 1961.890 4704.895 1962.170 4705.175 ;
        RECT 1962.510 4704.895 1962.790 4705.175 ;
        RECT 1963.130 4704.895 1963.410 4705.175 ;
        RECT 1963.750 4704.895 1964.030 4705.175 ;
        RECT 1964.370 4704.895 1964.650 4705.175 ;
        RECT 1964.990 4704.895 1965.270 4705.175 ;
        RECT 1965.610 4704.895 1965.890 4705.175 ;
        RECT 1966.230 4704.895 1966.510 4705.175 ;
        RECT 1966.850 4704.895 1967.130 4705.175 ;
        RECT 1967.470 4704.895 1967.750 4705.175 ;
        RECT 1968.090 4704.895 1968.370 4705.175 ;
        RECT 1959.410 4704.275 1959.690 4704.555 ;
        RECT 1960.030 4704.275 1960.310 4704.555 ;
        RECT 1960.650 4704.275 1960.930 4704.555 ;
        RECT 1961.270 4704.275 1961.550 4704.555 ;
        RECT 1961.890 4704.275 1962.170 4704.555 ;
        RECT 1962.510 4704.275 1962.790 4704.555 ;
        RECT 1963.130 4704.275 1963.410 4704.555 ;
        RECT 1963.750 4704.275 1964.030 4704.555 ;
        RECT 1964.370 4704.275 1964.650 4704.555 ;
        RECT 1964.990 4704.275 1965.270 4704.555 ;
        RECT 1965.610 4704.275 1965.890 4704.555 ;
        RECT 1966.230 4704.275 1966.510 4704.555 ;
        RECT 1966.850 4704.275 1967.130 4704.555 ;
        RECT 1967.470 4704.275 1967.750 4704.555 ;
        RECT 1968.090 4704.275 1968.370 4704.555 ;
        RECT 1959.410 4703.655 1959.690 4703.935 ;
        RECT 1960.030 4703.655 1960.310 4703.935 ;
        RECT 1960.650 4703.655 1960.930 4703.935 ;
        RECT 1961.270 4703.655 1961.550 4703.935 ;
        RECT 1961.890 4703.655 1962.170 4703.935 ;
        RECT 1962.510 4703.655 1962.790 4703.935 ;
        RECT 1963.130 4703.655 1963.410 4703.935 ;
        RECT 1963.750 4703.655 1964.030 4703.935 ;
        RECT 1964.370 4703.655 1964.650 4703.935 ;
        RECT 1964.990 4703.655 1965.270 4703.935 ;
        RECT 1965.610 4703.655 1965.890 4703.935 ;
        RECT 1966.230 4703.655 1966.510 4703.935 ;
        RECT 1966.850 4703.655 1967.130 4703.935 ;
        RECT 1967.470 4703.655 1967.750 4703.935 ;
        RECT 1968.090 4703.655 1968.370 4703.935 ;
        RECT 1959.410 4703.035 1959.690 4703.315 ;
        RECT 1960.030 4703.035 1960.310 4703.315 ;
        RECT 1960.650 4703.035 1960.930 4703.315 ;
        RECT 1961.270 4703.035 1961.550 4703.315 ;
        RECT 1961.890 4703.035 1962.170 4703.315 ;
        RECT 1962.510 4703.035 1962.790 4703.315 ;
        RECT 1963.130 4703.035 1963.410 4703.315 ;
        RECT 1963.750 4703.035 1964.030 4703.315 ;
        RECT 1964.370 4703.035 1964.650 4703.315 ;
        RECT 1964.990 4703.035 1965.270 4703.315 ;
        RECT 1965.610 4703.035 1965.890 4703.315 ;
        RECT 1966.230 4703.035 1966.510 4703.315 ;
        RECT 1966.850 4703.035 1967.130 4703.315 ;
        RECT 1967.470 4703.035 1967.750 4703.315 ;
        RECT 1968.090 4703.035 1968.370 4703.315 ;
        RECT 1959.410 4702.415 1959.690 4702.695 ;
        RECT 1960.030 4702.415 1960.310 4702.695 ;
        RECT 1960.650 4702.415 1960.930 4702.695 ;
        RECT 1961.270 4702.415 1961.550 4702.695 ;
        RECT 1961.890 4702.415 1962.170 4702.695 ;
        RECT 1962.510 4702.415 1962.790 4702.695 ;
        RECT 1963.130 4702.415 1963.410 4702.695 ;
        RECT 1963.750 4702.415 1964.030 4702.695 ;
        RECT 1964.370 4702.415 1964.650 4702.695 ;
        RECT 1964.990 4702.415 1965.270 4702.695 ;
        RECT 1965.610 4702.415 1965.890 4702.695 ;
        RECT 1966.230 4702.415 1966.510 4702.695 ;
        RECT 1966.850 4702.415 1967.130 4702.695 ;
        RECT 1967.470 4702.415 1967.750 4702.695 ;
        RECT 1968.090 4702.415 1968.370 4702.695 ;
        RECT 1959.410 4701.795 1959.690 4702.075 ;
        RECT 1960.030 4701.795 1960.310 4702.075 ;
        RECT 1960.650 4701.795 1960.930 4702.075 ;
        RECT 1961.270 4701.795 1961.550 4702.075 ;
        RECT 1961.890 4701.795 1962.170 4702.075 ;
        RECT 1962.510 4701.795 1962.790 4702.075 ;
        RECT 1963.130 4701.795 1963.410 4702.075 ;
        RECT 1963.750 4701.795 1964.030 4702.075 ;
        RECT 1964.370 4701.795 1964.650 4702.075 ;
        RECT 1964.990 4701.795 1965.270 4702.075 ;
        RECT 1965.610 4701.795 1965.890 4702.075 ;
        RECT 1966.230 4701.795 1966.510 4702.075 ;
        RECT 1966.850 4701.795 1967.130 4702.075 ;
        RECT 1967.470 4701.795 1967.750 4702.075 ;
        RECT 1968.090 4701.795 1968.370 4702.075 ;
        RECT 1959.410 4701.175 1959.690 4701.455 ;
        RECT 1960.030 4701.175 1960.310 4701.455 ;
        RECT 1960.650 4701.175 1960.930 4701.455 ;
        RECT 1961.270 4701.175 1961.550 4701.455 ;
        RECT 1961.890 4701.175 1962.170 4701.455 ;
        RECT 1962.510 4701.175 1962.790 4701.455 ;
        RECT 1963.130 4701.175 1963.410 4701.455 ;
        RECT 1963.750 4701.175 1964.030 4701.455 ;
        RECT 1964.370 4701.175 1964.650 4701.455 ;
        RECT 1964.990 4701.175 1965.270 4701.455 ;
        RECT 1965.610 4701.175 1965.890 4701.455 ;
        RECT 1966.230 4701.175 1966.510 4701.455 ;
        RECT 1966.850 4701.175 1967.130 4701.455 ;
        RECT 1967.470 4701.175 1967.750 4701.455 ;
        RECT 1968.090 4701.175 1968.370 4701.455 ;
        RECT 1959.410 4700.555 1959.690 4700.835 ;
        RECT 1960.030 4700.555 1960.310 4700.835 ;
        RECT 1960.650 4700.555 1960.930 4700.835 ;
        RECT 1961.270 4700.555 1961.550 4700.835 ;
        RECT 1961.890 4700.555 1962.170 4700.835 ;
        RECT 1962.510 4700.555 1962.790 4700.835 ;
        RECT 1963.130 4700.555 1963.410 4700.835 ;
        RECT 1963.750 4700.555 1964.030 4700.835 ;
        RECT 1964.370 4700.555 1964.650 4700.835 ;
        RECT 1964.990 4700.555 1965.270 4700.835 ;
        RECT 1965.610 4700.555 1965.890 4700.835 ;
        RECT 1966.230 4700.555 1966.510 4700.835 ;
        RECT 1966.850 4700.555 1967.130 4700.835 ;
        RECT 1967.470 4700.555 1967.750 4700.835 ;
        RECT 1968.090 4700.555 1968.370 4700.835 ;
        RECT 1959.410 4699.935 1959.690 4700.215 ;
        RECT 1960.030 4699.935 1960.310 4700.215 ;
        RECT 1960.650 4699.935 1960.930 4700.215 ;
        RECT 1961.270 4699.935 1961.550 4700.215 ;
        RECT 1961.890 4699.935 1962.170 4700.215 ;
        RECT 1962.510 4699.935 1962.790 4700.215 ;
        RECT 1963.130 4699.935 1963.410 4700.215 ;
        RECT 1963.750 4699.935 1964.030 4700.215 ;
        RECT 1964.370 4699.935 1964.650 4700.215 ;
        RECT 1964.990 4699.935 1965.270 4700.215 ;
        RECT 1965.610 4699.935 1965.890 4700.215 ;
        RECT 1966.230 4699.935 1966.510 4700.215 ;
        RECT 1966.850 4699.935 1967.130 4700.215 ;
        RECT 1967.470 4699.935 1967.750 4700.215 ;
        RECT 1968.090 4699.935 1968.370 4700.215 ;
        RECT 1959.410 4699.315 1959.690 4699.595 ;
        RECT 1960.030 4699.315 1960.310 4699.595 ;
        RECT 1960.650 4699.315 1960.930 4699.595 ;
        RECT 1961.270 4699.315 1961.550 4699.595 ;
        RECT 1961.890 4699.315 1962.170 4699.595 ;
        RECT 1962.510 4699.315 1962.790 4699.595 ;
        RECT 1963.130 4699.315 1963.410 4699.595 ;
        RECT 1963.750 4699.315 1964.030 4699.595 ;
        RECT 1964.370 4699.315 1964.650 4699.595 ;
        RECT 1964.990 4699.315 1965.270 4699.595 ;
        RECT 1965.610 4699.315 1965.890 4699.595 ;
        RECT 1966.230 4699.315 1966.510 4699.595 ;
        RECT 1966.850 4699.315 1967.130 4699.595 ;
        RECT 1967.470 4699.315 1967.750 4699.595 ;
        RECT 1968.090 4699.315 1968.370 4699.595 ;
        RECT 2996.630 4707.995 2996.910 4708.275 ;
        RECT 2997.250 4707.995 2997.530 4708.275 ;
        RECT 2997.870 4707.995 2998.150 4708.275 ;
        RECT 2998.490 4707.995 2998.770 4708.275 ;
        RECT 2999.110 4707.995 2999.390 4708.275 ;
        RECT 2999.730 4707.995 3000.010 4708.275 ;
        RECT 3000.350 4707.995 3000.630 4708.275 ;
        RECT 3000.970 4707.995 3001.250 4708.275 ;
        RECT 3001.590 4707.995 3001.870 4708.275 ;
        RECT 3002.210 4707.995 3002.490 4708.275 ;
        RECT 3002.830 4707.995 3003.110 4708.275 ;
        RECT 3003.450 4707.995 3003.730 4708.275 ;
        RECT 3004.070 4707.995 3004.350 4708.275 ;
        RECT 3004.690 4707.995 3004.970 4708.275 ;
        RECT 3005.310 4707.995 3005.590 4708.275 ;
        RECT 2996.630 4707.375 2996.910 4707.655 ;
        RECT 2997.250 4707.375 2997.530 4707.655 ;
        RECT 2997.870 4707.375 2998.150 4707.655 ;
        RECT 2998.490 4707.375 2998.770 4707.655 ;
        RECT 2999.110 4707.375 2999.390 4707.655 ;
        RECT 2999.730 4707.375 3000.010 4707.655 ;
        RECT 3000.350 4707.375 3000.630 4707.655 ;
        RECT 3000.970 4707.375 3001.250 4707.655 ;
        RECT 3001.590 4707.375 3001.870 4707.655 ;
        RECT 3002.210 4707.375 3002.490 4707.655 ;
        RECT 3002.830 4707.375 3003.110 4707.655 ;
        RECT 3003.450 4707.375 3003.730 4707.655 ;
        RECT 3004.070 4707.375 3004.350 4707.655 ;
        RECT 3004.690 4707.375 3004.970 4707.655 ;
        RECT 3005.310 4707.375 3005.590 4707.655 ;
        RECT 2996.630 4706.755 2996.910 4707.035 ;
        RECT 2997.250 4706.755 2997.530 4707.035 ;
        RECT 2997.870 4706.755 2998.150 4707.035 ;
        RECT 2998.490 4706.755 2998.770 4707.035 ;
        RECT 2999.110 4706.755 2999.390 4707.035 ;
        RECT 2999.730 4706.755 3000.010 4707.035 ;
        RECT 3000.350 4706.755 3000.630 4707.035 ;
        RECT 3000.970 4706.755 3001.250 4707.035 ;
        RECT 3001.590 4706.755 3001.870 4707.035 ;
        RECT 3002.210 4706.755 3002.490 4707.035 ;
        RECT 3002.830 4706.755 3003.110 4707.035 ;
        RECT 3003.450 4706.755 3003.730 4707.035 ;
        RECT 3004.070 4706.755 3004.350 4707.035 ;
        RECT 3004.690 4706.755 3004.970 4707.035 ;
        RECT 3005.310 4706.755 3005.590 4707.035 ;
        RECT 2996.630 4706.135 2996.910 4706.415 ;
        RECT 2997.250 4706.135 2997.530 4706.415 ;
        RECT 2997.870 4706.135 2998.150 4706.415 ;
        RECT 2998.490 4706.135 2998.770 4706.415 ;
        RECT 2999.110 4706.135 2999.390 4706.415 ;
        RECT 2999.730 4706.135 3000.010 4706.415 ;
        RECT 3000.350 4706.135 3000.630 4706.415 ;
        RECT 3000.970 4706.135 3001.250 4706.415 ;
        RECT 3001.590 4706.135 3001.870 4706.415 ;
        RECT 3002.210 4706.135 3002.490 4706.415 ;
        RECT 3002.830 4706.135 3003.110 4706.415 ;
        RECT 3003.450 4706.135 3003.730 4706.415 ;
        RECT 3004.070 4706.135 3004.350 4706.415 ;
        RECT 3004.690 4706.135 3004.970 4706.415 ;
        RECT 3005.310 4706.135 3005.590 4706.415 ;
        RECT 2996.630 4705.515 2996.910 4705.795 ;
        RECT 2997.250 4705.515 2997.530 4705.795 ;
        RECT 2997.870 4705.515 2998.150 4705.795 ;
        RECT 2998.490 4705.515 2998.770 4705.795 ;
        RECT 2999.110 4705.515 2999.390 4705.795 ;
        RECT 2999.730 4705.515 3000.010 4705.795 ;
        RECT 3000.350 4705.515 3000.630 4705.795 ;
        RECT 3000.970 4705.515 3001.250 4705.795 ;
        RECT 3001.590 4705.515 3001.870 4705.795 ;
        RECT 3002.210 4705.515 3002.490 4705.795 ;
        RECT 3002.830 4705.515 3003.110 4705.795 ;
        RECT 3003.450 4705.515 3003.730 4705.795 ;
        RECT 3004.070 4705.515 3004.350 4705.795 ;
        RECT 3004.690 4705.515 3004.970 4705.795 ;
        RECT 3005.310 4705.515 3005.590 4705.795 ;
        RECT 2996.630 4704.895 2996.910 4705.175 ;
        RECT 2997.250 4704.895 2997.530 4705.175 ;
        RECT 2997.870 4704.895 2998.150 4705.175 ;
        RECT 2998.490 4704.895 2998.770 4705.175 ;
        RECT 2999.110 4704.895 2999.390 4705.175 ;
        RECT 2999.730 4704.895 3000.010 4705.175 ;
        RECT 3000.350 4704.895 3000.630 4705.175 ;
        RECT 3000.970 4704.895 3001.250 4705.175 ;
        RECT 3001.590 4704.895 3001.870 4705.175 ;
        RECT 3002.210 4704.895 3002.490 4705.175 ;
        RECT 3002.830 4704.895 3003.110 4705.175 ;
        RECT 3003.450 4704.895 3003.730 4705.175 ;
        RECT 3004.070 4704.895 3004.350 4705.175 ;
        RECT 3004.690 4704.895 3004.970 4705.175 ;
        RECT 3005.310 4704.895 3005.590 4705.175 ;
        RECT 2996.630 4704.275 2996.910 4704.555 ;
        RECT 2997.250 4704.275 2997.530 4704.555 ;
        RECT 2997.870 4704.275 2998.150 4704.555 ;
        RECT 2998.490 4704.275 2998.770 4704.555 ;
        RECT 2999.110 4704.275 2999.390 4704.555 ;
        RECT 2999.730 4704.275 3000.010 4704.555 ;
        RECT 3000.350 4704.275 3000.630 4704.555 ;
        RECT 3000.970 4704.275 3001.250 4704.555 ;
        RECT 3001.590 4704.275 3001.870 4704.555 ;
        RECT 3002.210 4704.275 3002.490 4704.555 ;
        RECT 3002.830 4704.275 3003.110 4704.555 ;
        RECT 3003.450 4704.275 3003.730 4704.555 ;
        RECT 3004.070 4704.275 3004.350 4704.555 ;
        RECT 3004.690 4704.275 3004.970 4704.555 ;
        RECT 3005.310 4704.275 3005.590 4704.555 ;
        RECT 2996.630 4703.655 2996.910 4703.935 ;
        RECT 2997.250 4703.655 2997.530 4703.935 ;
        RECT 2997.870 4703.655 2998.150 4703.935 ;
        RECT 2998.490 4703.655 2998.770 4703.935 ;
        RECT 2999.110 4703.655 2999.390 4703.935 ;
        RECT 2999.730 4703.655 3000.010 4703.935 ;
        RECT 3000.350 4703.655 3000.630 4703.935 ;
        RECT 3000.970 4703.655 3001.250 4703.935 ;
        RECT 3001.590 4703.655 3001.870 4703.935 ;
        RECT 3002.210 4703.655 3002.490 4703.935 ;
        RECT 3002.830 4703.655 3003.110 4703.935 ;
        RECT 3003.450 4703.655 3003.730 4703.935 ;
        RECT 3004.070 4703.655 3004.350 4703.935 ;
        RECT 3004.690 4703.655 3004.970 4703.935 ;
        RECT 3005.310 4703.655 3005.590 4703.935 ;
        RECT 2996.630 4703.035 2996.910 4703.315 ;
        RECT 2997.250 4703.035 2997.530 4703.315 ;
        RECT 2997.870 4703.035 2998.150 4703.315 ;
        RECT 2998.490 4703.035 2998.770 4703.315 ;
        RECT 2999.110 4703.035 2999.390 4703.315 ;
        RECT 2999.730 4703.035 3000.010 4703.315 ;
        RECT 3000.350 4703.035 3000.630 4703.315 ;
        RECT 3000.970 4703.035 3001.250 4703.315 ;
        RECT 3001.590 4703.035 3001.870 4703.315 ;
        RECT 3002.210 4703.035 3002.490 4703.315 ;
        RECT 3002.830 4703.035 3003.110 4703.315 ;
        RECT 3003.450 4703.035 3003.730 4703.315 ;
        RECT 3004.070 4703.035 3004.350 4703.315 ;
        RECT 3004.690 4703.035 3004.970 4703.315 ;
        RECT 3005.310 4703.035 3005.590 4703.315 ;
        RECT 2996.630 4702.415 2996.910 4702.695 ;
        RECT 2997.250 4702.415 2997.530 4702.695 ;
        RECT 2997.870 4702.415 2998.150 4702.695 ;
        RECT 2998.490 4702.415 2998.770 4702.695 ;
        RECT 2999.110 4702.415 2999.390 4702.695 ;
        RECT 2999.730 4702.415 3000.010 4702.695 ;
        RECT 3000.350 4702.415 3000.630 4702.695 ;
        RECT 3000.970 4702.415 3001.250 4702.695 ;
        RECT 3001.590 4702.415 3001.870 4702.695 ;
        RECT 3002.210 4702.415 3002.490 4702.695 ;
        RECT 3002.830 4702.415 3003.110 4702.695 ;
        RECT 3003.450 4702.415 3003.730 4702.695 ;
        RECT 3004.070 4702.415 3004.350 4702.695 ;
        RECT 3004.690 4702.415 3004.970 4702.695 ;
        RECT 3005.310 4702.415 3005.590 4702.695 ;
        RECT 2996.630 4701.795 2996.910 4702.075 ;
        RECT 2997.250 4701.795 2997.530 4702.075 ;
        RECT 2997.870 4701.795 2998.150 4702.075 ;
        RECT 2998.490 4701.795 2998.770 4702.075 ;
        RECT 2999.110 4701.795 2999.390 4702.075 ;
        RECT 2999.730 4701.795 3000.010 4702.075 ;
        RECT 3000.350 4701.795 3000.630 4702.075 ;
        RECT 3000.970 4701.795 3001.250 4702.075 ;
        RECT 3001.590 4701.795 3001.870 4702.075 ;
        RECT 3002.210 4701.795 3002.490 4702.075 ;
        RECT 3002.830 4701.795 3003.110 4702.075 ;
        RECT 3003.450 4701.795 3003.730 4702.075 ;
        RECT 3004.070 4701.795 3004.350 4702.075 ;
        RECT 3004.690 4701.795 3004.970 4702.075 ;
        RECT 3005.310 4701.795 3005.590 4702.075 ;
        RECT 2996.630 4701.175 2996.910 4701.455 ;
        RECT 2997.250 4701.175 2997.530 4701.455 ;
        RECT 2997.870 4701.175 2998.150 4701.455 ;
        RECT 2998.490 4701.175 2998.770 4701.455 ;
        RECT 2999.110 4701.175 2999.390 4701.455 ;
        RECT 2999.730 4701.175 3000.010 4701.455 ;
        RECT 3000.350 4701.175 3000.630 4701.455 ;
        RECT 3000.970 4701.175 3001.250 4701.455 ;
        RECT 3001.590 4701.175 3001.870 4701.455 ;
        RECT 3002.210 4701.175 3002.490 4701.455 ;
        RECT 3002.830 4701.175 3003.110 4701.455 ;
        RECT 3003.450 4701.175 3003.730 4701.455 ;
        RECT 3004.070 4701.175 3004.350 4701.455 ;
        RECT 3004.690 4701.175 3004.970 4701.455 ;
        RECT 3005.310 4701.175 3005.590 4701.455 ;
        RECT 2996.630 4700.555 2996.910 4700.835 ;
        RECT 2997.250 4700.555 2997.530 4700.835 ;
        RECT 2997.870 4700.555 2998.150 4700.835 ;
        RECT 2998.490 4700.555 2998.770 4700.835 ;
        RECT 2999.110 4700.555 2999.390 4700.835 ;
        RECT 2999.730 4700.555 3000.010 4700.835 ;
        RECT 3000.350 4700.555 3000.630 4700.835 ;
        RECT 3000.970 4700.555 3001.250 4700.835 ;
        RECT 3001.590 4700.555 3001.870 4700.835 ;
        RECT 3002.210 4700.555 3002.490 4700.835 ;
        RECT 3002.830 4700.555 3003.110 4700.835 ;
        RECT 3003.450 4700.555 3003.730 4700.835 ;
        RECT 3004.070 4700.555 3004.350 4700.835 ;
        RECT 3004.690 4700.555 3004.970 4700.835 ;
        RECT 3005.310 4700.555 3005.590 4700.835 ;
        RECT 2996.630 4699.935 2996.910 4700.215 ;
        RECT 2997.250 4699.935 2997.530 4700.215 ;
        RECT 2997.870 4699.935 2998.150 4700.215 ;
        RECT 2998.490 4699.935 2998.770 4700.215 ;
        RECT 2999.110 4699.935 2999.390 4700.215 ;
        RECT 2999.730 4699.935 3000.010 4700.215 ;
        RECT 3000.350 4699.935 3000.630 4700.215 ;
        RECT 3000.970 4699.935 3001.250 4700.215 ;
        RECT 3001.590 4699.935 3001.870 4700.215 ;
        RECT 3002.210 4699.935 3002.490 4700.215 ;
        RECT 3002.830 4699.935 3003.110 4700.215 ;
        RECT 3003.450 4699.935 3003.730 4700.215 ;
        RECT 3004.070 4699.935 3004.350 4700.215 ;
        RECT 3004.690 4699.935 3004.970 4700.215 ;
        RECT 3005.310 4699.935 3005.590 4700.215 ;
        RECT 2996.630 4699.315 2996.910 4699.595 ;
        RECT 2997.250 4699.315 2997.530 4699.595 ;
        RECT 2997.870 4699.315 2998.150 4699.595 ;
        RECT 2998.490 4699.315 2998.770 4699.595 ;
        RECT 2999.110 4699.315 2999.390 4699.595 ;
        RECT 2999.730 4699.315 3000.010 4699.595 ;
        RECT 3000.350 4699.315 3000.630 4699.595 ;
        RECT 3000.970 4699.315 3001.250 4699.595 ;
        RECT 3001.590 4699.315 3001.870 4699.595 ;
        RECT 3002.210 4699.315 3002.490 4699.595 ;
        RECT 3002.830 4699.315 3003.110 4699.595 ;
        RECT 3003.450 4699.315 3003.730 4699.595 ;
        RECT 3004.070 4699.315 3004.350 4699.595 ;
        RECT 3004.690 4699.315 3004.970 4699.595 ;
        RECT 3005.310 4699.315 3005.590 4699.595 ;
        RECT 3009.160 4707.995 3009.440 4708.275 ;
        RECT 3009.780 4707.995 3010.060 4708.275 ;
        RECT 3010.400 4707.995 3010.680 4708.275 ;
        RECT 3011.020 4707.995 3011.300 4708.275 ;
        RECT 3011.640 4707.995 3011.920 4708.275 ;
        RECT 3012.260 4707.995 3012.540 4708.275 ;
        RECT 3012.880 4707.995 3013.160 4708.275 ;
        RECT 3013.500 4707.995 3013.780 4708.275 ;
        RECT 3014.120 4707.995 3014.400 4708.275 ;
        RECT 3014.740 4707.995 3015.020 4708.275 ;
        RECT 3015.360 4707.995 3015.640 4708.275 ;
        RECT 3015.980 4707.995 3016.260 4708.275 ;
        RECT 3016.600 4707.995 3016.880 4708.275 ;
        RECT 3017.220 4707.995 3017.500 4708.275 ;
        RECT 3017.840 4707.995 3018.120 4708.275 ;
        RECT 3018.460 4707.995 3018.740 4708.275 ;
        RECT 3009.160 4707.375 3009.440 4707.655 ;
        RECT 3009.780 4707.375 3010.060 4707.655 ;
        RECT 3010.400 4707.375 3010.680 4707.655 ;
        RECT 3011.020 4707.375 3011.300 4707.655 ;
        RECT 3011.640 4707.375 3011.920 4707.655 ;
        RECT 3012.260 4707.375 3012.540 4707.655 ;
        RECT 3012.880 4707.375 3013.160 4707.655 ;
        RECT 3013.500 4707.375 3013.780 4707.655 ;
        RECT 3014.120 4707.375 3014.400 4707.655 ;
        RECT 3014.740 4707.375 3015.020 4707.655 ;
        RECT 3015.360 4707.375 3015.640 4707.655 ;
        RECT 3015.980 4707.375 3016.260 4707.655 ;
        RECT 3016.600 4707.375 3016.880 4707.655 ;
        RECT 3017.220 4707.375 3017.500 4707.655 ;
        RECT 3017.840 4707.375 3018.120 4707.655 ;
        RECT 3018.460 4707.375 3018.740 4707.655 ;
        RECT 3009.160 4706.755 3009.440 4707.035 ;
        RECT 3009.780 4706.755 3010.060 4707.035 ;
        RECT 3010.400 4706.755 3010.680 4707.035 ;
        RECT 3011.020 4706.755 3011.300 4707.035 ;
        RECT 3011.640 4706.755 3011.920 4707.035 ;
        RECT 3012.260 4706.755 3012.540 4707.035 ;
        RECT 3012.880 4706.755 3013.160 4707.035 ;
        RECT 3013.500 4706.755 3013.780 4707.035 ;
        RECT 3014.120 4706.755 3014.400 4707.035 ;
        RECT 3014.740 4706.755 3015.020 4707.035 ;
        RECT 3015.360 4706.755 3015.640 4707.035 ;
        RECT 3015.980 4706.755 3016.260 4707.035 ;
        RECT 3016.600 4706.755 3016.880 4707.035 ;
        RECT 3017.220 4706.755 3017.500 4707.035 ;
        RECT 3017.840 4706.755 3018.120 4707.035 ;
        RECT 3018.460 4706.755 3018.740 4707.035 ;
        RECT 3009.160 4706.135 3009.440 4706.415 ;
        RECT 3009.780 4706.135 3010.060 4706.415 ;
        RECT 3010.400 4706.135 3010.680 4706.415 ;
        RECT 3011.020 4706.135 3011.300 4706.415 ;
        RECT 3011.640 4706.135 3011.920 4706.415 ;
        RECT 3012.260 4706.135 3012.540 4706.415 ;
        RECT 3012.880 4706.135 3013.160 4706.415 ;
        RECT 3013.500 4706.135 3013.780 4706.415 ;
        RECT 3014.120 4706.135 3014.400 4706.415 ;
        RECT 3014.740 4706.135 3015.020 4706.415 ;
        RECT 3015.360 4706.135 3015.640 4706.415 ;
        RECT 3015.980 4706.135 3016.260 4706.415 ;
        RECT 3016.600 4706.135 3016.880 4706.415 ;
        RECT 3017.220 4706.135 3017.500 4706.415 ;
        RECT 3017.840 4706.135 3018.120 4706.415 ;
        RECT 3018.460 4706.135 3018.740 4706.415 ;
        RECT 3009.160 4705.515 3009.440 4705.795 ;
        RECT 3009.780 4705.515 3010.060 4705.795 ;
        RECT 3010.400 4705.515 3010.680 4705.795 ;
        RECT 3011.020 4705.515 3011.300 4705.795 ;
        RECT 3011.640 4705.515 3011.920 4705.795 ;
        RECT 3012.260 4705.515 3012.540 4705.795 ;
        RECT 3012.880 4705.515 3013.160 4705.795 ;
        RECT 3013.500 4705.515 3013.780 4705.795 ;
        RECT 3014.120 4705.515 3014.400 4705.795 ;
        RECT 3014.740 4705.515 3015.020 4705.795 ;
        RECT 3015.360 4705.515 3015.640 4705.795 ;
        RECT 3015.980 4705.515 3016.260 4705.795 ;
        RECT 3016.600 4705.515 3016.880 4705.795 ;
        RECT 3017.220 4705.515 3017.500 4705.795 ;
        RECT 3017.840 4705.515 3018.120 4705.795 ;
        RECT 3018.460 4705.515 3018.740 4705.795 ;
        RECT 3009.160 4704.895 3009.440 4705.175 ;
        RECT 3009.780 4704.895 3010.060 4705.175 ;
        RECT 3010.400 4704.895 3010.680 4705.175 ;
        RECT 3011.020 4704.895 3011.300 4705.175 ;
        RECT 3011.640 4704.895 3011.920 4705.175 ;
        RECT 3012.260 4704.895 3012.540 4705.175 ;
        RECT 3012.880 4704.895 3013.160 4705.175 ;
        RECT 3013.500 4704.895 3013.780 4705.175 ;
        RECT 3014.120 4704.895 3014.400 4705.175 ;
        RECT 3014.740 4704.895 3015.020 4705.175 ;
        RECT 3015.360 4704.895 3015.640 4705.175 ;
        RECT 3015.980 4704.895 3016.260 4705.175 ;
        RECT 3016.600 4704.895 3016.880 4705.175 ;
        RECT 3017.220 4704.895 3017.500 4705.175 ;
        RECT 3017.840 4704.895 3018.120 4705.175 ;
        RECT 3018.460 4704.895 3018.740 4705.175 ;
        RECT 3009.160 4704.275 3009.440 4704.555 ;
        RECT 3009.780 4704.275 3010.060 4704.555 ;
        RECT 3010.400 4704.275 3010.680 4704.555 ;
        RECT 3011.020 4704.275 3011.300 4704.555 ;
        RECT 3011.640 4704.275 3011.920 4704.555 ;
        RECT 3012.260 4704.275 3012.540 4704.555 ;
        RECT 3012.880 4704.275 3013.160 4704.555 ;
        RECT 3013.500 4704.275 3013.780 4704.555 ;
        RECT 3014.120 4704.275 3014.400 4704.555 ;
        RECT 3014.740 4704.275 3015.020 4704.555 ;
        RECT 3015.360 4704.275 3015.640 4704.555 ;
        RECT 3015.980 4704.275 3016.260 4704.555 ;
        RECT 3016.600 4704.275 3016.880 4704.555 ;
        RECT 3017.220 4704.275 3017.500 4704.555 ;
        RECT 3017.840 4704.275 3018.120 4704.555 ;
        RECT 3018.460 4704.275 3018.740 4704.555 ;
        RECT 3009.160 4703.655 3009.440 4703.935 ;
        RECT 3009.780 4703.655 3010.060 4703.935 ;
        RECT 3010.400 4703.655 3010.680 4703.935 ;
        RECT 3011.020 4703.655 3011.300 4703.935 ;
        RECT 3011.640 4703.655 3011.920 4703.935 ;
        RECT 3012.260 4703.655 3012.540 4703.935 ;
        RECT 3012.880 4703.655 3013.160 4703.935 ;
        RECT 3013.500 4703.655 3013.780 4703.935 ;
        RECT 3014.120 4703.655 3014.400 4703.935 ;
        RECT 3014.740 4703.655 3015.020 4703.935 ;
        RECT 3015.360 4703.655 3015.640 4703.935 ;
        RECT 3015.980 4703.655 3016.260 4703.935 ;
        RECT 3016.600 4703.655 3016.880 4703.935 ;
        RECT 3017.220 4703.655 3017.500 4703.935 ;
        RECT 3017.840 4703.655 3018.120 4703.935 ;
        RECT 3018.460 4703.655 3018.740 4703.935 ;
        RECT 3009.160 4703.035 3009.440 4703.315 ;
        RECT 3009.780 4703.035 3010.060 4703.315 ;
        RECT 3010.400 4703.035 3010.680 4703.315 ;
        RECT 3011.020 4703.035 3011.300 4703.315 ;
        RECT 3011.640 4703.035 3011.920 4703.315 ;
        RECT 3012.260 4703.035 3012.540 4703.315 ;
        RECT 3012.880 4703.035 3013.160 4703.315 ;
        RECT 3013.500 4703.035 3013.780 4703.315 ;
        RECT 3014.120 4703.035 3014.400 4703.315 ;
        RECT 3014.740 4703.035 3015.020 4703.315 ;
        RECT 3015.360 4703.035 3015.640 4703.315 ;
        RECT 3015.980 4703.035 3016.260 4703.315 ;
        RECT 3016.600 4703.035 3016.880 4703.315 ;
        RECT 3017.220 4703.035 3017.500 4703.315 ;
        RECT 3017.840 4703.035 3018.120 4703.315 ;
        RECT 3018.460 4703.035 3018.740 4703.315 ;
        RECT 3009.160 4702.415 3009.440 4702.695 ;
        RECT 3009.780 4702.415 3010.060 4702.695 ;
        RECT 3010.400 4702.415 3010.680 4702.695 ;
        RECT 3011.020 4702.415 3011.300 4702.695 ;
        RECT 3011.640 4702.415 3011.920 4702.695 ;
        RECT 3012.260 4702.415 3012.540 4702.695 ;
        RECT 3012.880 4702.415 3013.160 4702.695 ;
        RECT 3013.500 4702.415 3013.780 4702.695 ;
        RECT 3014.120 4702.415 3014.400 4702.695 ;
        RECT 3014.740 4702.415 3015.020 4702.695 ;
        RECT 3015.360 4702.415 3015.640 4702.695 ;
        RECT 3015.980 4702.415 3016.260 4702.695 ;
        RECT 3016.600 4702.415 3016.880 4702.695 ;
        RECT 3017.220 4702.415 3017.500 4702.695 ;
        RECT 3017.840 4702.415 3018.120 4702.695 ;
        RECT 3018.460 4702.415 3018.740 4702.695 ;
        RECT 3009.160 4701.795 3009.440 4702.075 ;
        RECT 3009.780 4701.795 3010.060 4702.075 ;
        RECT 3010.400 4701.795 3010.680 4702.075 ;
        RECT 3011.020 4701.795 3011.300 4702.075 ;
        RECT 3011.640 4701.795 3011.920 4702.075 ;
        RECT 3012.260 4701.795 3012.540 4702.075 ;
        RECT 3012.880 4701.795 3013.160 4702.075 ;
        RECT 3013.500 4701.795 3013.780 4702.075 ;
        RECT 3014.120 4701.795 3014.400 4702.075 ;
        RECT 3014.740 4701.795 3015.020 4702.075 ;
        RECT 3015.360 4701.795 3015.640 4702.075 ;
        RECT 3015.980 4701.795 3016.260 4702.075 ;
        RECT 3016.600 4701.795 3016.880 4702.075 ;
        RECT 3017.220 4701.795 3017.500 4702.075 ;
        RECT 3017.840 4701.795 3018.120 4702.075 ;
        RECT 3018.460 4701.795 3018.740 4702.075 ;
        RECT 3009.160 4701.175 3009.440 4701.455 ;
        RECT 3009.780 4701.175 3010.060 4701.455 ;
        RECT 3010.400 4701.175 3010.680 4701.455 ;
        RECT 3011.020 4701.175 3011.300 4701.455 ;
        RECT 3011.640 4701.175 3011.920 4701.455 ;
        RECT 3012.260 4701.175 3012.540 4701.455 ;
        RECT 3012.880 4701.175 3013.160 4701.455 ;
        RECT 3013.500 4701.175 3013.780 4701.455 ;
        RECT 3014.120 4701.175 3014.400 4701.455 ;
        RECT 3014.740 4701.175 3015.020 4701.455 ;
        RECT 3015.360 4701.175 3015.640 4701.455 ;
        RECT 3015.980 4701.175 3016.260 4701.455 ;
        RECT 3016.600 4701.175 3016.880 4701.455 ;
        RECT 3017.220 4701.175 3017.500 4701.455 ;
        RECT 3017.840 4701.175 3018.120 4701.455 ;
        RECT 3018.460 4701.175 3018.740 4701.455 ;
        RECT 3009.160 4700.555 3009.440 4700.835 ;
        RECT 3009.780 4700.555 3010.060 4700.835 ;
        RECT 3010.400 4700.555 3010.680 4700.835 ;
        RECT 3011.020 4700.555 3011.300 4700.835 ;
        RECT 3011.640 4700.555 3011.920 4700.835 ;
        RECT 3012.260 4700.555 3012.540 4700.835 ;
        RECT 3012.880 4700.555 3013.160 4700.835 ;
        RECT 3013.500 4700.555 3013.780 4700.835 ;
        RECT 3014.120 4700.555 3014.400 4700.835 ;
        RECT 3014.740 4700.555 3015.020 4700.835 ;
        RECT 3015.360 4700.555 3015.640 4700.835 ;
        RECT 3015.980 4700.555 3016.260 4700.835 ;
        RECT 3016.600 4700.555 3016.880 4700.835 ;
        RECT 3017.220 4700.555 3017.500 4700.835 ;
        RECT 3017.840 4700.555 3018.120 4700.835 ;
        RECT 3018.460 4700.555 3018.740 4700.835 ;
        RECT 3009.160 4699.935 3009.440 4700.215 ;
        RECT 3009.780 4699.935 3010.060 4700.215 ;
        RECT 3010.400 4699.935 3010.680 4700.215 ;
        RECT 3011.020 4699.935 3011.300 4700.215 ;
        RECT 3011.640 4699.935 3011.920 4700.215 ;
        RECT 3012.260 4699.935 3012.540 4700.215 ;
        RECT 3012.880 4699.935 3013.160 4700.215 ;
        RECT 3013.500 4699.935 3013.780 4700.215 ;
        RECT 3014.120 4699.935 3014.400 4700.215 ;
        RECT 3014.740 4699.935 3015.020 4700.215 ;
        RECT 3015.360 4699.935 3015.640 4700.215 ;
        RECT 3015.980 4699.935 3016.260 4700.215 ;
        RECT 3016.600 4699.935 3016.880 4700.215 ;
        RECT 3017.220 4699.935 3017.500 4700.215 ;
        RECT 3017.840 4699.935 3018.120 4700.215 ;
        RECT 3018.460 4699.935 3018.740 4700.215 ;
        RECT 3009.160 4699.315 3009.440 4699.595 ;
        RECT 3009.780 4699.315 3010.060 4699.595 ;
        RECT 3010.400 4699.315 3010.680 4699.595 ;
        RECT 3011.020 4699.315 3011.300 4699.595 ;
        RECT 3011.640 4699.315 3011.920 4699.595 ;
        RECT 3012.260 4699.315 3012.540 4699.595 ;
        RECT 3012.880 4699.315 3013.160 4699.595 ;
        RECT 3013.500 4699.315 3013.780 4699.595 ;
        RECT 3014.120 4699.315 3014.400 4699.595 ;
        RECT 3014.740 4699.315 3015.020 4699.595 ;
        RECT 3015.360 4699.315 3015.640 4699.595 ;
        RECT 3015.980 4699.315 3016.260 4699.595 ;
        RECT 3016.600 4699.315 3016.880 4699.595 ;
        RECT 3017.220 4699.315 3017.500 4699.595 ;
        RECT 3017.840 4699.315 3018.120 4699.595 ;
        RECT 3018.460 4699.315 3018.740 4699.595 ;
        RECT 3025.350 4707.995 3025.630 4708.275 ;
        RECT 3025.970 4707.995 3026.250 4708.275 ;
        RECT 3026.590 4707.995 3026.870 4708.275 ;
        RECT 3027.210 4707.995 3027.490 4708.275 ;
        RECT 3027.830 4707.995 3028.110 4708.275 ;
        RECT 3028.450 4707.995 3028.730 4708.275 ;
        RECT 3029.070 4707.995 3029.350 4708.275 ;
        RECT 3029.690 4707.995 3029.970 4708.275 ;
        RECT 3030.310 4707.995 3030.590 4708.275 ;
        RECT 3025.350 4707.375 3025.630 4707.655 ;
        RECT 3025.970 4707.375 3026.250 4707.655 ;
        RECT 3026.590 4707.375 3026.870 4707.655 ;
        RECT 3027.210 4707.375 3027.490 4707.655 ;
        RECT 3027.830 4707.375 3028.110 4707.655 ;
        RECT 3028.450 4707.375 3028.730 4707.655 ;
        RECT 3029.070 4707.375 3029.350 4707.655 ;
        RECT 3029.690 4707.375 3029.970 4707.655 ;
        RECT 3030.310 4707.375 3030.590 4707.655 ;
        RECT 3025.350 4706.755 3025.630 4707.035 ;
        RECT 3025.970 4706.755 3026.250 4707.035 ;
        RECT 3026.590 4706.755 3026.870 4707.035 ;
        RECT 3027.210 4706.755 3027.490 4707.035 ;
        RECT 3027.830 4706.755 3028.110 4707.035 ;
        RECT 3028.450 4706.755 3028.730 4707.035 ;
        RECT 3029.070 4706.755 3029.350 4707.035 ;
        RECT 3029.690 4706.755 3029.970 4707.035 ;
        RECT 3030.310 4706.755 3030.590 4707.035 ;
        RECT 3025.350 4706.135 3025.630 4706.415 ;
        RECT 3025.970 4706.135 3026.250 4706.415 ;
        RECT 3026.590 4706.135 3026.870 4706.415 ;
        RECT 3027.210 4706.135 3027.490 4706.415 ;
        RECT 3027.830 4706.135 3028.110 4706.415 ;
        RECT 3028.450 4706.135 3028.730 4706.415 ;
        RECT 3029.070 4706.135 3029.350 4706.415 ;
        RECT 3029.690 4706.135 3029.970 4706.415 ;
        RECT 3030.310 4706.135 3030.590 4706.415 ;
        RECT 3025.350 4705.515 3025.630 4705.795 ;
        RECT 3025.970 4705.515 3026.250 4705.795 ;
        RECT 3026.590 4705.515 3026.870 4705.795 ;
        RECT 3027.210 4705.515 3027.490 4705.795 ;
        RECT 3027.830 4705.515 3028.110 4705.795 ;
        RECT 3028.450 4705.515 3028.730 4705.795 ;
        RECT 3029.070 4705.515 3029.350 4705.795 ;
        RECT 3029.690 4705.515 3029.970 4705.795 ;
        RECT 3030.310 4705.515 3030.590 4705.795 ;
        RECT 3025.350 4704.895 3025.630 4705.175 ;
        RECT 3025.970 4704.895 3026.250 4705.175 ;
        RECT 3026.590 4704.895 3026.870 4705.175 ;
        RECT 3027.210 4704.895 3027.490 4705.175 ;
        RECT 3027.830 4704.895 3028.110 4705.175 ;
        RECT 3028.450 4704.895 3028.730 4705.175 ;
        RECT 3029.070 4704.895 3029.350 4705.175 ;
        RECT 3029.690 4704.895 3029.970 4705.175 ;
        RECT 3030.310 4704.895 3030.590 4705.175 ;
        RECT 3025.350 4704.275 3025.630 4704.555 ;
        RECT 3025.970 4704.275 3026.250 4704.555 ;
        RECT 3026.590 4704.275 3026.870 4704.555 ;
        RECT 3027.210 4704.275 3027.490 4704.555 ;
        RECT 3027.830 4704.275 3028.110 4704.555 ;
        RECT 3028.450 4704.275 3028.730 4704.555 ;
        RECT 3029.070 4704.275 3029.350 4704.555 ;
        RECT 3029.690 4704.275 3029.970 4704.555 ;
        RECT 3030.310 4704.275 3030.590 4704.555 ;
        RECT 3025.350 4703.655 3025.630 4703.935 ;
        RECT 3025.970 4703.655 3026.250 4703.935 ;
        RECT 3026.590 4703.655 3026.870 4703.935 ;
        RECT 3027.210 4703.655 3027.490 4703.935 ;
        RECT 3027.830 4703.655 3028.110 4703.935 ;
        RECT 3028.450 4703.655 3028.730 4703.935 ;
        RECT 3029.070 4703.655 3029.350 4703.935 ;
        RECT 3029.690 4703.655 3029.970 4703.935 ;
        RECT 3030.310 4703.655 3030.590 4703.935 ;
        RECT 3025.350 4703.035 3025.630 4703.315 ;
        RECT 3025.970 4703.035 3026.250 4703.315 ;
        RECT 3026.590 4703.035 3026.870 4703.315 ;
        RECT 3027.210 4703.035 3027.490 4703.315 ;
        RECT 3027.830 4703.035 3028.110 4703.315 ;
        RECT 3028.450 4703.035 3028.730 4703.315 ;
        RECT 3029.070 4703.035 3029.350 4703.315 ;
        RECT 3029.690 4703.035 3029.970 4703.315 ;
        RECT 3030.310 4703.035 3030.590 4703.315 ;
        RECT 3025.350 4702.415 3025.630 4702.695 ;
        RECT 3025.970 4702.415 3026.250 4702.695 ;
        RECT 3026.590 4702.415 3026.870 4702.695 ;
        RECT 3027.210 4702.415 3027.490 4702.695 ;
        RECT 3027.830 4702.415 3028.110 4702.695 ;
        RECT 3028.450 4702.415 3028.730 4702.695 ;
        RECT 3029.070 4702.415 3029.350 4702.695 ;
        RECT 3029.690 4702.415 3029.970 4702.695 ;
        RECT 3030.310 4702.415 3030.590 4702.695 ;
        RECT 3025.350 4701.795 3025.630 4702.075 ;
        RECT 3025.970 4701.795 3026.250 4702.075 ;
        RECT 3026.590 4701.795 3026.870 4702.075 ;
        RECT 3027.210 4701.795 3027.490 4702.075 ;
        RECT 3027.830 4701.795 3028.110 4702.075 ;
        RECT 3028.450 4701.795 3028.730 4702.075 ;
        RECT 3029.070 4701.795 3029.350 4702.075 ;
        RECT 3029.690 4701.795 3029.970 4702.075 ;
        RECT 3030.310 4701.795 3030.590 4702.075 ;
        RECT 3025.350 4701.175 3025.630 4701.455 ;
        RECT 3025.970 4701.175 3026.250 4701.455 ;
        RECT 3026.590 4701.175 3026.870 4701.455 ;
        RECT 3027.210 4701.175 3027.490 4701.455 ;
        RECT 3027.830 4701.175 3028.110 4701.455 ;
        RECT 3028.450 4701.175 3028.730 4701.455 ;
        RECT 3029.070 4701.175 3029.350 4701.455 ;
        RECT 3029.690 4701.175 3029.970 4701.455 ;
        RECT 3030.310 4701.175 3030.590 4701.455 ;
        RECT 3025.350 4700.555 3025.630 4700.835 ;
        RECT 3025.970 4700.555 3026.250 4700.835 ;
        RECT 3026.590 4700.555 3026.870 4700.835 ;
        RECT 3027.210 4700.555 3027.490 4700.835 ;
        RECT 3027.830 4700.555 3028.110 4700.835 ;
        RECT 3028.450 4700.555 3028.730 4700.835 ;
        RECT 3029.070 4700.555 3029.350 4700.835 ;
        RECT 3029.690 4700.555 3029.970 4700.835 ;
        RECT 3030.310 4700.555 3030.590 4700.835 ;
        RECT 3025.350 4699.935 3025.630 4700.215 ;
        RECT 3025.970 4699.935 3026.250 4700.215 ;
        RECT 3026.590 4699.935 3026.870 4700.215 ;
        RECT 3027.210 4699.935 3027.490 4700.215 ;
        RECT 3027.830 4699.935 3028.110 4700.215 ;
        RECT 3028.450 4699.935 3028.730 4700.215 ;
        RECT 3029.070 4699.935 3029.350 4700.215 ;
        RECT 3029.690 4699.935 3029.970 4700.215 ;
        RECT 3030.310 4699.935 3030.590 4700.215 ;
        RECT 3025.350 4699.315 3025.630 4699.595 ;
        RECT 3025.970 4699.315 3026.250 4699.595 ;
        RECT 3026.590 4699.315 3026.870 4699.595 ;
        RECT 3027.210 4699.315 3027.490 4699.595 ;
        RECT 3027.830 4699.315 3028.110 4699.595 ;
        RECT 3028.450 4699.315 3028.730 4699.595 ;
        RECT 3029.070 4699.315 3029.350 4699.595 ;
        RECT 3029.690 4699.315 3029.970 4699.595 ;
        RECT 3030.310 4699.315 3030.590 4699.595 ;
        RECT 3034.540 4707.995 3034.820 4708.275 ;
        RECT 3035.160 4707.995 3035.440 4708.275 ;
        RECT 3035.780 4707.995 3036.060 4708.275 ;
        RECT 3036.400 4707.995 3036.680 4708.275 ;
        RECT 3037.020 4707.995 3037.300 4708.275 ;
        RECT 3037.640 4707.995 3037.920 4708.275 ;
        RECT 3038.260 4707.995 3038.540 4708.275 ;
        RECT 3038.880 4707.995 3039.160 4708.275 ;
        RECT 3039.500 4707.995 3039.780 4708.275 ;
        RECT 3040.120 4707.995 3040.400 4708.275 ;
        RECT 3040.740 4707.995 3041.020 4708.275 ;
        RECT 3041.360 4707.995 3041.640 4708.275 ;
        RECT 3041.980 4707.995 3042.260 4708.275 ;
        RECT 3042.600 4707.995 3042.880 4708.275 ;
        RECT 3043.220 4707.995 3043.500 4708.275 ;
        RECT 3043.840 4707.995 3044.120 4708.275 ;
        RECT 3034.540 4707.375 3034.820 4707.655 ;
        RECT 3035.160 4707.375 3035.440 4707.655 ;
        RECT 3035.780 4707.375 3036.060 4707.655 ;
        RECT 3036.400 4707.375 3036.680 4707.655 ;
        RECT 3037.020 4707.375 3037.300 4707.655 ;
        RECT 3037.640 4707.375 3037.920 4707.655 ;
        RECT 3038.260 4707.375 3038.540 4707.655 ;
        RECT 3038.880 4707.375 3039.160 4707.655 ;
        RECT 3039.500 4707.375 3039.780 4707.655 ;
        RECT 3040.120 4707.375 3040.400 4707.655 ;
        RECT 3040.740 4707.375 3041.020 4707.655 ;
        RECT 3041.360 4707.375 3041.640 4707.655 ;
        RECT 3041.980 4707.375 3042.260 4707.655 ;
        RECT 3042.600 4707.375 3042.880 4707.655 ;
        RECT 3043.220 4707.375 3043.500 4707.655 ;
        RECT 3043.840 4707.375 3044.120 4707.655 ;
        RECT 3034.540 4706.755 3034.820 4707.035 ;
        RECT 3035.160 4706.755 3035.440 4707.035 ;
        RECT 3035.780 4706.755 3036.060 4707.035 ;
        RECT 3036.400 4706.755 3036.680 4707.035 ;
        RECT 3037.020 4706.755 3037.300 4707.035 ;
        RECT 3037.640 4706.755 3037.920 4707.035 ;
        RECT 3038.260 4706.755 3038.540 4707.035 ;
        RECT 3038.880 4706.755 3039.160 4707.035 ;
        RECT 3039.500 4706.755 3039.780 4707.035 ;
        RECT 3040.120 4706.755 3040.400 4707.035 ;
        RECT 3040.740 4706.755 3041.020 4707.035 ;
        RECT 3041.360 4706.755 3041.640 4707.035 ;
        RECT 3041.980 4706.755 3042.260 4707.035 ;
        RECT 3042.600 4706.755 3042.880 4707.035 ;
        RECT 3043.220 4706.755 3043.500 4707.035 ;
        RECT 3043.840 4706.755 3044.120 4707.035 ;
        RECT 3034.540 4706.135 3034.820 4706.415 ;
        RECT 3035.160 4706.135 3035.440 4706.415 ;
        RECT 3035.780 4706.135 3036.060 4706.415 ;
        RECT 3036.400 4706.135 3036.680 4706.415 ;
        RECT 3037.020 4706.135 3037.300 4706.415 ;
        RECT 3037.640 4706.135 3037.920 4706.415 ;
        RECT 3038.260 4706.135 3038.540 4706.415 ;
        RECT 3038.880 4706.135 3039.160 4706.415 ;
        RECT 3039.500 4706.135 3039.780 4706.415 ;
        RECT 3040.120 4706.135 3040.400 4706.415 ;
        RECT 3040.740 4706.135 3041.020 4706.415 ;
        RECT 3041.360 4706.135 3041.640 4706.415 ;
        RECT 3041.980 4706.135 3042.260 4706.415 ;
        RECT 3042.600 4706.135 3042.880 4706.415 ;
        RECT 3043.220 4706.135 3043.500 4706.415 ;
        RECT 3043.840 4706.135 3044.120 4706.415 ;
        RECT 3034.540 4705.515 3034.820 4705.795 ;
        RECT 3035.160 4705.515 3035.440 4705.795 ;
        RECT 3035.780 4705.515 3036.060 4705.795 ;
        RECT 3036.400 4705.515 3036.680 4705.795 ;
        RECT 3037.020 4705.515 3037.300 4705.795 ;
        RECT 3037.640 4705.515 3037.920 4705.795 ;
        RECT 3038.260 4705.515 3038.540 4705.795 ;
        RECT 3038.880 4705.515 3039.160 4705.795 ;
        RECT 3039.500 4705.515 3039.780 4705.795 ;
        RECT 3040.120 4705.515 3040.400 4705.795 ;
        RECT 3040.740 4705.515 3041.020 4705.795 ;
        RECT 3041.360 4705.515 3041.640 4705.795 ;
        RECT 3041.980 4705.515 3042.260 4705.795 ;
        RECT 3042.600 4705.515 3042.880 4705.795 ;
        RECT 3043.220 4705.515 3043.500 4705.795 ;
        RECT 3043.840 4705.515 3044.120 4705.795 ;
        RECT 3034.540 4704.895 3034.820 4705.175 ;
        RECT 3035.160 4704.895 3035.440 4705.175 ;
        RECT 3035.780 4704.895 3036.060 4705.175 ;
        RECT 3036.400 4704.895 3036.680 4705.175 ;
        RECT 3037.020 4704.895 3037.300 4705.175 ;
        RECT 3037.640 4704.895 3037.920 4705.175 ;
        RECT 3038.260 4704.895 3038.540 4705.175 ;
        RECT 3038.880 4704.895 3039.160 4705.175 ;
        RECT 3039.500 4704.895 3039.780 4705.175 ;
        RECT 3040.120 4704.895 3040.400 4705.175 ;
        RECT 3040.740 4704.895 3041.020 4705.175 ;
        RECT 3041.360 4704.895 3041.640 4705.175 ;
        RECT 3041.980 4704.895 3042.260 4705.175 ;
        RECT 3042.600 4704.895 3042.880 4705.175 ;
        RECT 3043.220 4704.895 3043.500 4705.175 ;
        RECT 3043.840 4704.895 3044.120 4705.175 ;
        RECT 3034.540 4704.275 3034.820 4704.555 ;
        RECT 3035.160 4704.275 3035.440 4704.555 ;
        RECT 3035.780 4704.275 3036.060 4704.555 ;
        RECT 3036.400 4704.275 3036.680 4704.555 ;
        RECT 3037.020 4704.275 3037.300 4704.555 ;
        RECT 3037.640 4704.275 3037.920 4704.555 ;
        RECT 3038.260 4704.275 3038.540 4704.555 ;
        RECT 3038.880 4704.275 3039.160 4704.555 ;
        RECT 3039.500 4704.275 3039.780 4704.555 ;
        RECT 3040.120 4704.275 3040.400 4704.555 ;
        RECT 3040.740 4704.275 3041.020 4704.555 ;
        RECT 3041.360 4704.275 3041.640 4704.555 ;
        RECT 3041.980 4704.275 3042.260 4704.555 ;
        RECT 3042.600 4704.275 3042.880 4704.555 ;
        RECT 3043.220 4704.275 3043.500 4704.555 ;
        RECT 3043.840 4704.275 3044.120 4704.555 ;
        RECT 3034.540 4703.655 3034.820 4703.935 ;
        RECT 3035.160 4703.655 3035.440 4703.935 ;
        RECT 3035.780 4703.655 3036.060 4703.935 ;
        RECT 3036.400 4703.655 3036.680 4703.935 ;
        RECT 3037.020 4703.655 3037.300 4703.935 ;
        RECT 3037.640 4703.655 3037.920 4703.935 ;
        RECT 3038.260 4703.655 3038.540 4703.935 ;
        RECT 3038.880 4703.655 3039.160 4703.935 ;
        RECT 3039.500 4703.655 3039.780 4703.935 ;
        RECT 3040.120 4703.655 3040.400 4703.935 ;
        RECT 3040.740 4703.655 3041.020 4703.935 ;
        RECT 3041.360 4703.655 3041.640 4703.935 ;
        RECT 3041.980 4703.655 3042.260 4703.935 ;
        RECT 3042.600 4703.655 3042.880 4703.935 ;
        RECT 3043.220 4703.655 3043.500 4703.935 ;
        RECT 3043.840 4703.655 3044.120 4703.935 ;
        RECT 3034.540 4703.035 3034.820 4703.315 ;
        RECT 3035.160 4703.035 3035.440 4703.315 ;
        RECT 3035.780 4703.035 3036.060 4703.315 ;
        RECT 3036.400 4703.035 3036.680 4703.315 ;
        RECT 3037.020 4703.035 3037.300 4703.315 ;
        RECT 3037.640 4703.035 3037.920 4703.315 ;
        RECT 3038.260 4703.035 3038.540 4703.315 ;
        RECT 3038.880 4703.035 3039.160 4703.315 ;
        RECT 3039.500 4703.035 3039.780 4703.315 ;
        RECT 3040.120 4703.035 3040.400 4703.315 ;
        RECT 3040.740 4703.035 3041.020 4703.315 ;
        RECT 3041.360 4703.035 3041.640 4703.315 ;
        RECT 3041.980 4703.035 3042.260 4703.315 ;
        RECT 3042.600 4703.035 3042.880 4703.315 ;
        RECT 3043.220 4703.035 3043.500 4703.315 ;
        RECT 3043.840 4703.035 3044.120 4703.315 ;
        RECT 3034.540 4702.415 3034.820 4702.695 ;
        RECT 3035.160 4702.415 3035.440 4702.695 ;
        RECT 3035.780 4702.415 3036.060 4702.695 ;
        RECT 3036.400 4702.415 3036.680 4702.695 ;
        RECT 3037.020 4702.415 3037.300 4702.695 ;
        RECT 3037.640 4702.415 3037.920 4702.695 ;
        RECT 3038.260 4702.415 3038.540 4702.695 ;
        RECT 3038.880 4702.415 3039.160 4702.695 ;
        RECT 3039.500 4702.415 3039.780 4702.695 ;
        RECT 3040.120 4702.415 3040.400 4702.695 ;
        RECT 3040.740 4702.415 3041.020 4702.695 ;
        RECT 3041.360 4702.415 3041.640 4702.695 ;
        RECT 3041.980 4702.415 3042.260 4702.695 ;
        RECT 3042.600 4702.415 3042.880 4702.695 ;
        RECT 3043.220 4702.415 3043.500 4702.695 ;
        RECT 3043.840 4702.415 3044.120 4702.695 ;
        RECT 3034.540 4701.795 3034.820 4702.075 ;
        RECT 3035.160 4701.795 3035.440 4702.075 ;
        RECT 3035.780 4701.795 3036.060 4702.075 ;
        RECT 3036.400 4701.795 3036.680 4702.075 ;
        RECT 3037.020 4701.795 3037.300 4702.075 ;
        RECT 3037.640 4701.795 3037.920 4702.075 ;
        RECT 3038.260 4701.795 3038.540 4702.075 ;
        RECT 3038.880 4701.795 3039.160 4702.075 ;
        RECT 3039.500 4701.795 3039.780 4702.075 ;
        RECT 3040.120 4701.795 3040.400 4702.075 ;
        RECT 3040.740 4701.795 3041.020 4702.075 ;
        RECT 3041.360 4701.795 3041.640 4702.075 ;
        RECT 3041.980 4701.795 3042.260 4702.075 ;
        RECT 3042.600 4701.795 3042.880 4702.075 ;
        RECT 3043.220 4701.795 3043.500 4702.075 ;
        RECT 3043.840 4701.795 3044.120 4702.075 ;
        RECT 3034.540 4701.175 3034.820 4701.455 ;
        RECT 3035.160 4701.175 3035.440 4701.455 ;
        RECT 3035.780 4701.175 3036.060 4701.455 ;
        RECT 3036.400 4701.175 3036.680 4701.455 ;
        RECT 3037.020 4701.175 3037.300 4701.455 ;
        RECT 3037.640 4701.175 3037.920 4701.455 ;
        RECT 3038.260 4701.175 3038.540 4701.455 ;
        RECT 3038.880 4701.175 3039.160 4701.455 ;
        RECT 3039.500 4701.175 3039.780 4701.455 ;
        RECT 3040.120 4701.175 3040.400 4701.455 ;
        RECT 3040.740 4701.175 3041.020 4701.455 ;
        RECT 3041.360 4701.175 3041.640 4701.455 ;
        RECT 3041.980 4701.175 3042.260 4701.455 ;
        RECT 3042.600 4701.175 3042.880 4701.455 ;
        RECT 3043.220 4701.175 3043.500 4701.455 ;
        RECT 3043.840 4701.175 3044.120 4701.455 ;
        RECT 3034.540 4700.555 3034.820 4700.835 ;
        RECT 3035.160 4700.555 3035.440 4700.835 ;
        RECT 3035.780 4700.555 3036.060 4700.835 ;
        RECT 3036.400 4700.555 3036.680 4700.835 ;
        RECT 3037.020 4700.555 3037.300 4700.835 ;
        RECT 3037.640 4700.555 3037.920 4700.835 ;
        RECT 3038.260 4700.555 3038.540 4700.835 ;
        RECT 3038.880 4700.555 3039.160 4700.835 ;
        RECT 3039.500 4700.555 3039.780 4700.835 ;
        RECT 3040.120 4700.555 3040.400 4700.835 ;
        RECT 3040.740 4700.555 3041.020 4700.835 ;
        RECT 3041.360 4700.555 3041.640 4700.835 ;
        RECT 3041.980 4700.555 3042.260 4700.835 ;
        RECT 3042.600 4700.555 3042.880 4700.835 ;
        RECT 3043.220 4700.555 3043.500 4700.835 ;
        RECT 3043.840 4700.555 3044.120 4700.835 ;
        RECT 3034.540 4699.935 3034.820 4700.215 ;
        RECT 3035.160 4699.935 3035.440 4700.215 ;
        RECT 3035.780 4699.935 3036.060 4700.215 ;
        RECT 3036.400 4699.935 3036.680 4700.215 ;
        RECT 3037.020 4699.935 3037.300 4700.215 ;
        RECT 3037.640 4699.935 3037.920 4700.215 ;
        RECT 3038.260 4699.935 3038.540 4700.215 ;
        RECT 3038.880 4699.935 3039.160 4700.215 ;
        RECT 3039.500 4699.935 3039.780 4700.215 ;
        RECT 3040.120 4699.935 3040.400 4700.215 ;
        RECT 3040.740 4699.935 3041.020 4700.215 ;
        RECT 3041.360 4699.935 3041.640 4700.215 ;
        RECT 3041.980 4699.935 3042.260 4700.215 ;
        RECT 3042.600 4699.935 3042.880 4700.215 ;
        RECT 3043.220 4699.935 3043.500 4700.215 ;
        RECT 3043.840 4699.935 3044.120 4700.215 ;
        RECT 3034.540 4699.315 3034.820 4699.595 ;
        RECT 3035.160 4699.315 3035.440 4699.595 ;
        RECT 3035.780 4699.315 3036.060 4699.595 ;
        RECT 3036.400 4699.315 3036.680 4699.595 ;
        RECT 3037.020 4699.315 3037.300 4699.595 ;
        RECT 3037.640 4699.315 3037.920 4699.595 ;
        RECT 3038.260 4699.315 3038.540 4699.595 ;
        RECT 3038.880 4699.315 3039.160 4699.595 ;
        RECT 3039.500 4699.315 3039.780 4699.595 ;
        RECT 3040.120 4699.315 3040.400 4699.595 ;
        RECT 3040.740 4699.315 3041.020 4699.595 ;
        RECT 3041.360 4699.315 3041.640 4699.595 ;
        RECT 3041.980 4699.315 3042.260 4699.595 ;
        RECT 3042.600 4699.315 3042.880 4699.595 ;
        RECT 3043.220 4699.315 3043.500 4699.595 ;
        RECT 3043.840 4699.315 3044.120 4699.595 ;
        RECT 3046.390 4707.995 3046.670 4708.275 ;
        RECT 3047.010 4707.995 3047.290 4708.275 ;
        RECT 3047.630 4707.995 3047.910 4708.275 ;
        RECT 3048.250 4707.995 3048.530 4708.275 ;
        RECT 3048.870 4707.995 3049.150 4708.275 ;
        RECT 3049.490 4707.995 3049.770 4708.275 ;
        RECT 3050.110 4707.995 3050.390 4708.275 ;
        RECT 3050.730 4707.995 3051.010 4708.275 ;
        RECT 3051.350 4707.995 3051.630 4708.275 ;
        RECT 3051.970 4707.995 3052.250 4708.275 ;
        RECT 3052.590 4707.995 3052.870 4708.275 ;
        RECT 3053.210 4707.995 3053.490 4708.275 ;
        RECT 3053.830 4707.995 3054.110 4708.275 ;
        RECT 3054.450 4707.995 3054.730 4708.275 ;
        RECT 3055.070 4707.995 3055.350 4708.275 ;
        RECT 3055.690 4707.995 3055.970 4708.275 ;
        RECT 3046.390 4707.375 3046.670 4707.655 ;
        RECT 3047.010 4707.375 3047.290 4707.655 ;
        RECT 3047.630 4707.375 3047.910 4707.655 ;
        RECT 3048.250 4707.375 3048.530 4707.655 ;
        RECT 3048.870 4707.375 3049.150 4707.655 ;
        RECT 3049.490 4707.375 3049.770 4707.655 ;
        RECT 3050.110 4707.375 3050.390 4707.655 ;
        RECT 3050.730 4707.375 3051.010 4707.655 ;
        RECT 3051.350 4707.375 3051.630 4707.655 ;
        RECT 3051.970 4707.375 3052.250 4707.655 ;
        RECT 3052.590 4707.375 3052.870 4707.655 ;
        RECT 3053.210 4707.375 3053.490 4707.655 ;
        RECT 3053.830 4707.375 3054.110 4707.655 ;
        RECT 3054.450 4707.375 3054.730 4707.655 ;
        RECT 3055.070 4707.375 3055.350 4707.655 ;
        RECT 3055.690 4707.375 3055.970 4707.655 ;
        RECT 3046.390 4706.755 3046.670 4707.035 ;
        RECT 3047.010 4706.755 3047.290 4707.035 ;
        RECT 3047.630 4706.755 3047.910 4707.035 ;
        RECT 3048.250 4706.755 3048.530 4707.035 ;
        RECT 3048.870 4706.755 3049.150 4707.035 ;
        RECT 3049.490 4706.755 3049.770 4707.035 ;
        RECT 3050.110 4706.755 3050.390 4707.035 ;
        RECT 3050.730 4706.755 3051.010 4707.035 ;
        RECT 3051.350 4706.755 3051.630 4707.035 ;
        RECT 3051.970 4706.755 3052.250 4707.035 ;
        RECT 3052.590 4706.755 3052.870 4707.035 ;
        RECT 3053.210 4706.755 3053.490 4707.035 ;
        RECT 3053.830 4706.755 3054.110 4707.035 ;
        RECT 3054.450 4706.755 3054.730 4707.035 ;
        RECT 3055.070 4706.755 3055.350 4707.035 ;
        RECT 3055.690 4706.755 3055.970 4707.035 ;
        RECT 3046.390 4706.135 3046.670 4706.415 ;
        RECT 3047.010 4706.135 3047.290 4706.415 ;
        RECT 3047.630 4706.135 3047.910 4706.415 ;
        RECT 3048.250 4706.135 3048.530 4706.415 ;
        RECT 3048.870 4706.135 3049.150 4706.415 ;
        RECT 3049.490 4706.135 3049.770 4706.415 ;
        RECT 3050.110 4706.135 3050.390 4706.415 ;
        RECT 3050.730 4706.135 3051.010 4706.415 ;
        RECT 3051.350 4706.135 3051.630 4706.415 ;
        RECT 3051.970 4706.135 3052.250 4706.415 ;
        RECT 3052.590 4706.135 3052.870 4706.415 ;
        RECT 3053.210 4706.135 3053.490 4706.415 ;
        RECT 3053.830 4706.135 3054.110 4706.415 ;
        RECT 3054.450 4706.135 3054.730 4706.415 ;
        RECT 3055.070 4706.135 3055.350 4706.415 ;
        RECT 3055.690 4706.135 3055.970 4706.415 ;
        RECT 3046.390 4705.515 3046.670 4705.795 ;
        RECT 3047.010 4705.515 3047.290 4705.795 ;
        RECT 3047.630 4705.515 3047.910 4705.795 ;
        RECT 3048.250 4705.515 3048.530 4705.795 ;
        RECT 3048.870 4705.515 3049.150 4705.795 ;
        RECT 3049.490 4705.515 3049.770 4705.795 ;
        RECT 3050.110 4705.515 3050.390 4705.795 ;
        RECT 3050.730 4705.515 3051.010 4705.795 ;
        RECT 3051.350 4705.515 3051.630 4705.795 ;
        RECT 3051.970 4705.515 3052.250 4705.795 ;
        RECT 3052.590 4705.515 3052.870 4705.795 ;
        RECT 3053.210 4705.515 3053.490 4705.795 ;
        RECT 3053.830 4705.515 3054.110 4705.795 ;
        RECT 3054.450 4705.515 3054.730 4705.795 ;
        RECT 3055.070 4705.515 3055.350 4705.795 ;
        RECT 3055.690 4705.515 3055.970 4705.795 ;
        RECT 3046.390 4704.895 3046.670 4705.175 ;
        RECT 3047.010 4704.895 3047.290 4705.175 ;
        RECT 3047.630 4704.895 3047.910 4705.175 ;
        RECT 3048.250 4704.895 3048.530 4705.175 ;
        RECT 3048.870 4704.895 3049.150 4705.175 ;
        RECT 3049.490 4704.895 3049.770 4705.175 ;
        RECT 3050.110 4704.895 3050.390 4705.175 ;
        RECT 3050.730 4704.895 3051.010 4705.175 ;
        RECT 3051.350 4704.895 3051.630 4705.175 ;
        RECT 3051.970 4704.895 3052.250 4705.175 ;
        RECT 3052.590 4704.895 3052.870 4705.175 ;
        RECT 3053.210 4704.895 3053.490 4705.175 ;
        RECT 3053.830 4704.895 3054.110 4705.175 ;
        RECT 3054.450 4704.895 3054.730 4705.175 ;
        RECT 3055.070 4704.895 3055.350 4705.175 ;
        RECT 3055.690 4704.895 3055.970 4705.175 ;
        RECT 3046.390 4704.275 3046.670 4704.555 ;
        RECT 3047.010 4704.275 3047.290 4704.555 ;
        RECT 3047.630 4704.275 3047.910 4704.555 ;
        RECT 3048.250 4704.275 3048.530 4704.555 ;
        RECT 3048.870 4704.275 3049.150 4704.555 ;
        RECT 3049.490 4704.275 3049.770 4704.555 ;
        RECT 3050.110 4704.275 3050.390 4704.555 ;
        RECT 3050.730 4704.275 3051.010 4704.555 ;
        RECT 3051.350 4704.275 3051.630 4704.555 ;
        RECT 3051.970 4704.275 3052.250 4704.555 ;
        RECT 3052.590 4704.275 3052.870 4704.555 ;
        RECT 3053.210 4704.275 3053.490 4704.555 ;
        RECT 3053.830 4704.275 3054.110 4704.555 ;
        RECT 3054.450 4704.275 3054.730 4704.555 ;
        RECT 3055.070 4704.275 3055.350 4704.555 ;
        RECT 3055.690 4704.275 3055.970 4704.555 ;
        RECT 3046.390 4703.655 3046.670 4703.935 ;
        RECT 3047.010 4703.655 3047.290 4703.935 ;
        RECT 3047.630 4703.655 3047.910 4703.935 ;
        RECT 3048.250 4703.655 3048.530 4703.935 ;
        RECT 3048.870 4703.655 3049.150 4703.935 ;
        RECT 3049.490 4703.655 3049.770 4703.935 ;
        RECT 3050.110 4703.655 3050.390 4703.935 ;
        RECT 3050.730 4703.655 3051.010 4703.935 ;
        RECT 3051.350 4703.655 3051.630 4703.935 ;
        RECT 3051.970 4703.655 3052.250 4703.935 ;
        RECT 3052.590 4703.655 3052.870 4703.935 ;
        RECT 3053.210 4703.655 3053.490 4703.935 ;
        RECT 3053.830 4703.655 3054.110 4703.935 ;
        RECT 3054.450 4703.655 3054.730 4703.935 ;
        RECT 3055.070 4703.655 3055.350 4703.935 ;
        RECT 3055.690 4703.655 3055.970 4703.935 ;
        RECT 3046.390 4703.035 3046.670 4703.315 ;
        RECT 3047.010 4703.035 3047.290 4703.315 ;
        RECT 3047.630 4703.035 3047.910 4703.315 ;
        RECT 3048.250 4703.035 3048.530 4703.315 ;
        RECT 3048.870 4703.035 3049.150 4703.315 ;
        RECT 3049.490 4703.035 3049.770 4703.315 ;
        RECT 3050.110 4703.035 3050.390 4703.315 ;
        RECT 3050.730 4703.035 3051.010 4703.315 ;
        RECT 3051.350 4703.035 3051.630 4703.315 ;
        RECT 3051.970 4703.035 3052.250 4703.315 ;
        RECT 3052.590 4703.035 3052.870 4703.315 ;
        RECT 3053.210 4703.035 3053.490 4703.315 ;
        RECT 3053.830 4703.035 3054.110 4703.315 ;
        RECT 3054.450 4703.035 3054.730 4703.315 ;
        RECT 3055.070 4703.035 3055.350 4703.315 ;
        RECT 3055.690 4703.035 3055.970 4703.315 ;
        RECT 3046.390 4702.415 3046.670 4702.695 ;
        RECT 3047.010 4702.415 3047.290 4702.695 ;
        RECT 3047.630 4702.415 3047.910 4702.695 ;
        RECT 3048.250 4702.415 3048.530 4702.695 ;
        RECT 3048.870 4702.415 3049.150 4702.695 ;
        RECT 3049.490 4702.415 3049.770 4702.695 ;
        RECT 3050.110 4702.415 3050.390 4702.695 ;
        RECT 3050.730 4702.415 3051.010 4702.695 ;
        RECT 3051.350 4702.415 3051.630 4702.695 ;
        RECT 3051.970 4702.415 3052.250 4702.695 ;
        RECT 3052.590 4702.415 3052.870 4702.695 ;
        RECT 3053.210 4702.415 3053.490 4702.695 ;
        RECT 3053.830 4702.415 3054.110 4702.695 ;
        RECT 3054.450 4702.415 3054.730 4702.695 ;
        RECT 3055.070 4702.415 3055.350 4702.695 ;
        RECT 3055.690 4702.415 3055.970 4702.695 ;
        RECT 3046.390 4701.795 3046.670 4702.075 ;
        RECT 3047.010 4701.795 3047.290 4702.075 ;
        RECT 3047.630 4701.795 3047.910 4702.075 ;
        RECT 3048.250 4701.795 3048.530 4702.075 ;
        RECT 3048.870 4701.795 3049.150 4702.075 ;
        RECT 3049.490 4701.795 3049.770 4702.075 ;
        RECT 3050.110 4701.795 3050.390 4702.075 ;
        RECT 3050.730 4701.795 3051.010 4702.075 ;
        RECT 3051.350 4701.795 3051.630 4702.075 ;
        RECT 3051.970 4701.795 3052.250 4702.075 ;
        RECT 3052.590 4701.795 3052.870 4702.075 ;
        RECT 3053.210 4701.795 3053.490 4702.075 ;
        RECT 3053.830 4701.795 3054.110 4702.075 ;
        RECT 3054.450 4701.795 3054.730 4702.075 ;
        RECT 3055.070 4701.795 3055.350 4702.075 ;
        RECT 3055.690 4701.795 3055.970 4702.075 ;
        RECT 3046.390 4701.175 3046.670 4701.455 ;
        RECT 3047.010 4701.175 3047.290 4701.455 ;
        RECT 3047.630 4701.175 3047.910 4701.455 ;
        RECT 3048.250 4701.175 3048.530 4701.455 ;
        RECT 3048.870 4701.175 3049.150 4701.455 ;
        RECT 3049.490 4701.175 3049.770 4701.455 ;
        RECT 3050.110 4701.175 3050.390 4701.455 ;
        RECT 3050.730 4701.175 3051.010 4701.455 ;
        RECT 3051.350 4701.175 3051.630 4701.455 ;
        RECT 3051.970 4701.175 3052.250 4701.455 ;
        RECT 3052.590 4701.175 3052.870 4701.455 ;
        RECT 3053.210 4701.175 3053.490 4701.455 ;
        RECT 3053.830 4701.175 3054.110 4701.455 ;
        RECT 3054.450 4701.175 3054.730 4701.455 ;
        RECT 3055.070 4701.175 3055.350 4701.455 ;
        RECT 3055.690 4701.175 3055.970 4701.455 ;
        RECT 3046.390 4700.555 3046.670 4700.835 ;
        RECT 3047.010 4700.555 3047.290 4700.835 ;
        RECT 3047.630 4700.555 3047.910 4700.835 ;
        RECT 3048.250 4700.555 3048.530 4700.835 ;
        RECT 3048.870 4700.555 3049.150 4700.835 ;
        RECT 3049.490 4700.555 3049.770 4700.835 ;
        RECT 3050.110 4700.555 3050.390 4700.835 ;
        RECT 3050.730 4700.555 3051.010 4700.835 ;
        RECT 3051.350 4700.555 3051.630 4700.835 ;
        RECT 3051.970 4700.555 3052.250 4700.835 ;
        RECT 3052.590 4700.555 3052.870 4700.835 ;
        RECT 3053.210 4700.555 3053.490 4700.835 ;
        RECT 3053.830 4700.555 3054.110 4700.835 ;
        RECT 3054.450 4700.555 3054.730 4700.835 ;
        RECT 3055.070 4700.555 3055.350 4700.835 ;
        RECT 3055.690 4700.555 3055.970 4700.835 ;
        RECT 3046.390 4699.935 3046.670 4700.215 ;
        RECT 3047.010 4699.935 3047.290 4700.215 ;
        RECT 3047.630 4699.935 3047.910 4700.215 ;
        RECT 3048.250 4699.935 3048.530 4700.215 ;
        RECT 3048.870 4699.935 3049.150 4700.215 ;
        RECT 3049.490 4699.935 3049.770 4700.215 ;
        RECT 3050.110 4699.935 3050.390 4700.215 ;
        RECT 3050.730 4699.935 3051.010 4700.215 ;
        RECT 3051.350 4699.935 3051.630 4700.215 ;
        RECT 3051.970 4699.935 3052.250 4700.215 ;
        RECT 3052.590 4699.935 3052.870 4700.215 ;
        RECT 3053.210 4699.935 3053.490 4700.215 ;
        RECT 3053.830 4699.935 3054.110 4700.215 ;
        RECT 3054.450 4699.935 3054.730 4700.215 ;
        RECT 3055.070 4699.935 3055.350 4700.215 ;
        RECT 3055.690 4699.935 3055.970 4700.215 ;
        RECT 3046.390 4699.315 3046.670 4699.595 ;
        RECT 3047.010 4699.315 3047.290 4699.595 ;
        RECT 3047.630 4699.315 3047.910 4699.595 ;
        RECT 3048.250 4699.315 3048.530 4699.595 ;
        RECT 3048.870 4699.315 3049.150 4699.595 ;
        RECT 3049.490 4699.315 3049.770 4699.595 ;
        RECT 3050.110 4699.315 3050.390 4699.595 ;
        RECT 3050.730 4699.315 3051.010 4699.595 ;
        RECT 3051.350 4699.315 3051.630 4699.595 ;
        RECT 3051.970 4699.315 3052.250 4699.595 ;
        RECT 3052.590 4699.315 3052.870 4699.595 ;
        RECT 3053.210 4699.315 3053.490 4699.595 ;
        RECT 3053.830 4699.315 3054.110 4699.595 ;
        RECT 3054.450 4699.315 3054.730 4699.595 ;
        RECT 3055.070 4699.315 3055.350 4699.595 ;
        RECT 3055.690 4699.315 3055.970 4699.595 ;
        RECT 3059.410 4707.995 3059.690 4708.275 ;
        RECT 3060.030 4707.995 3060.310 4708.275 ;
        RECT 3060.650 4707.995 3060.930 4708.275 ;
        RECT 3061.270 4707.995 3061.550 4708.275 ;
        RECT 3061.890 4707.995 3062.170 4708.275 ;
        RECT 3062.510 4707.995 3062.790 4708.275 ;
        RECT 3063.130 4707.995 3063.410 4708.275 ;
        RECT 3063.750 4707.995 3064.030 4708.275 ;
        RECT 3064.370 4707.995 3064.650 4708.275 ;
        RECT 3064.990 4707.995 3065.270 4708.275 ;
        RECT 3065.610 4707.995 3065.890 4708.275 ;
        RECT 3066.230 4707.995 3066.510 4708.275 ;
        RECT 3066.850 4707.995 3067.130 4708.275 ;
        RECT 3067.470 4707.995 3067.750 4708.275 ;
        RECT 3068.090 4707.995 3068.370 4708.275 ;
        RECT 3059.410 4707.375 3059.690 4707.655 ;
        RECT 3060.030 4707.375 3060.310 4707.655 ;
        RECT 3060.650 4707.375 3060.930 4707.655 ;
        RECT 3061.270 4707.375 3061.550 4707.655 ;
        RECT 3061.890 4707.375 3062.170 4707.655 ;
        RECT 3062.510 4707.375 3062.790 4707.655 ;
        RECT 3063.130 4707.375 3063.410 4707.655 ;
        RECT 3063.750 4707.375 3064.030 4707.655 ;
        RECT 3064.370 4707.375 3064.650 4707.655 ;
        RECT 3064.990 4707.375 3065.270 4707.655 ;
        RECT 3065.610 4707.375 3065.890 4707.655 ;
        RECT 3066.230 4707.375 3066.510 4707.655 ;
        RECT 3066.850 4707.375 3067.130 4707.655 ;
        RECT 3067.470 4707.375 3067.750 4707.655 ;
        RECT 3068.090 4707.375 3068.370 4707.655 ;
        RECT 3059.410 4706.755 3059.690 4707.035 ;
        RECT 3060.030 4706.755 3060.310 4707.035 ;
        RECT 3060.650 4706.755 3060.930 4707.035 ;
        RECT 3061.270 4706.755 3061.550 4707.035 ;
        RECT 3061.890 4706.755 3062.170 4707.035 ;
        RECT 3062.510 4706.755 3062.790 4707.035 ;
        RECT 3063.130 4706.755 3063.410 4707.035 ;
        RECT 3063.750 4706.755 3064.030 4707.035 ;
        RECT 3064.370 4706.755 3064.650 4707.035 ;
        RECT 3064.990 4706.755 3065.270 4707.035 ;
        RECT 3065.610 4706.755 3065.890 4707.035 ;
        RECT 3066.230 4706.755 3066.510 4707.035 ;
        RECT 3066.850 4706.755 3067.130 4707.035 ;
        RECT 3067.470 4706.755 3067.750 4707.035 ;
        RECT 3068.090 4706.755 3068.370 4707.035 ;
        RECT 3059.410 4706.135 3059.690 4706.415 ;
        RECT 3060.030 4706.135 3060.310 4706.415 ;
        RECT 3060.650 4706.135 3060.930 4706.415 ;
        RECT 3061.270 4706.135 3061.550 4706.415 ;
        RECT 3061.890 4706.135 3062.170 4706.415 ;
        RECT 3062.510 4706.135 3062.790 4706.415 ;
        RECT 3063.130 4706.135 3063.410 4706.415 ;
        RECT 3063.750 4706.135 3064.030 4706.415 ;
        RECT 3064.370 4706.135 3064.650 4706.415 ;
        RECT 3064.990 4706.135 3065.270 4706.415 ;
        RECT 3065.610 4706.135 3065.890 4706.415 ;
        RECT 3066.230 4706.135 3066.510 4706.415 ;
        RECT 3066.850 4706.135 3067.130 4706.415 ;
        RECT 3067.470 4706.135 3067.750 4706.415 ;
        RECT 3068.090 4706.135 3068.370 4706.415 ;
        RECT 3059.410 4705.515 3059.690 4705.795 ;
        RECT 3060.030 4705.515 3060.310 4705.795 ;
        RECT 3060.650 4705.515 3060.930 4705.795 ;
        RECT 3061.270 4705.515 3061.550 4705.795 ;
        RECT 3061.890 4705.515 3062.170 4705.795 ;
        RECT 3062.510 4705.515 3062.790 4705.795 ;
        RECT 3063.130 4705.515 3063.410 4705.795 ;
        RECT 3063.750 4705.515 3064.030 4705.795 ;
        RECT 3064.370 4705.515 3064.650 4705.795 ;
        RECT 3064.990 4705.515 3065.270 4705.795 ;
        RECT 3065.610 4705.515 3065.890 4705.795 ;
        RECT 3066.230 4705.515 3066.510 4705.795 ;
        RECT 3066.850 4705.515 3067.130 4705.795 ;
        RECT 3067.470 4705.515 3067.750 4705.795 ;
        RECT 3068.090 4705.515 3068.370 4705.795 ;
        RECT 3059.410 4704.895 3059.690 4705.175 ;
        RECT 3060.030 4704.895 3060.310 4705.175 ;
        RECT 3060.650 4704.895 3060.930 4705.175 ;
        RECT 3061.270 4704.895 3061.550 4705.175 ;
        RECT 3061.890 4704.895 3062.170 4705.175 ;
        RECT 3062.510 4704.895 3062.790 4705.175 ;
        RECT 3063.130 4704.895 3063.410 4705.175 ;
        RECT 3063.750 4704.895 3064.030 4705.175 ;
        RECT 3064.370 4704.895 3064.650 4705.175 ;
        RECT 3064.990 4704.895 3065.270 4705.175 ;
        RECT 3065.610 4704.895 3065.890 4705.175 ;
        RECT 3066.230 4704.895 3066.510 4705.175 ;
        RECT 3066.850 4704.895 3067.130 4705.175 ;
        RECT 3067.470 4704.895 3067.750 4705.175 ;
        RECT 3068.090 4704.895 3068.370 4705.175 ;
        RECT 3059.410 4704.275 3059.690 4704.555 ;
        RECT 3060.030 4704.275 3060.310 4704.555 ;
        RECT 3060.650 4704.275 3060.930 4704.555 ;
        RECT 3061.270 4704.275 3061.550 4704.555 ;
        RECT 3061.890 4704.275 3062.170 4704.555 ;
        RECT 3062.510 4704.275 3062.790 4704.555 ;
        RECT 3063.130 4704.275 3063.410 4704.555 ;
        RECT 3063.750 4704.275 3064.030 4704.555 ;
        RECT 3064.370 4704.275 3064.650 4704.555 ;
        RECT 3064.990 4704.275 3065.270 4704.555 ;
        RECT 3065.610 4704.275 3065.890 4704.555 ;
        RECT 3066.230 4704.275 3066.510 4704.555 ;
        RECT 3066.850 4704.275 3067.130 4704.555 ;
        RECT 3067.470 4704.275 3067.750 4704.555 ;
        RECT 3068.090 4704.275 3068.370 4704.555 ;
        RECT 3059.410 4703.655 3059.690 4703.935 ;
        RECT 3060.030 4703.655 3060.310 4703.935 ;
        RECT 3060.650 4703.655 3060.930 4703.935 ;
        RECT 3061.270 4703.655 3061.550 4703.935 ;
        RECT 3061.890 4703.655 3062.170 4703.935 ;
        RECT 3062.510 4703.655 3062.790 4703.935 ;
        RECT 3063.130 4703.655 3063.410 4703.935 ;
        RECT 3063.750 4703.655 3064.030 4703.935 ;
        RECT 3064.370 4703.655 3064.650 4703.935 ;
        RECT 3064.990 4703.655 3065.270 4703.935 ;
        RECT 3065.610 4703.655 3065.890 4703.935 ;
        RECT 3066.230 4703.655 3066.510 4703.935 ;
        RECT 3066.850 4703.655 3067.130 4703.935 ;
        RECT 3067.470 4703.655 3067.750 4703.935 ;
        RECT 3068.090 4703.655 3068.370 4703.935 ;
        RECT 3059.410 4703.035 3059.690 4703.315 ;
        RECT 3060.030 4703.035 3060.310 4703.315 ;
        RECT 3060.650 4703.035 3060.930 4703.315 ;
        RECT 3061.270 4703.035 3061.550 4703.315 ;
        RECT 3061.890 4703.035 3062.170 4703.315 ;
        RECT 3062.510 4703.035 3062.790 4703.315 ;
        RECT 3063.130 4703.035 3063.410 4703.315 ;
        RECT 3063.750 4703.035 3064.030 4703.315 ;
        RECT 3064.370 4703.035 3064.650 4703.315 ;
        RECT 3064.990 4703.035 3065.270 4703.315 ;
        RECT 3065.610 4703.035 3065.890 4703.315 ;
        RECT 3066.230 4703.035 3066.510 4703.315 ;
        RECT 3066.850 4703.035 3067.130 4703.315 ;
        RECT 3067.470 4703.035 3067.750 4703.315 ;
        RECT 3068.090 4703.035 3068.370 4703.315 ;
        RECT 3059.410 4702.415 3059.690 4702.695 ;
        RECT 3060.030 4702.415 3060.310 4702.695 ;
        RECT 3060.650 4702.415 3060.930 4702.695 ;
        RECT 3061.270 4702.415 3061.550 4702.695 ;
        RECT 3061.890 4702.415 3062.170 4702.695 ;
        RECT 3062.510 4702.415 3062.790 4702.695 ;
        RECT 3063.130 4702.415 3063.410 4702.695 ;
        RECT 3063.750 4702.415 3064.030 4702.695 ;
        RECT 3064.370 4702.415 3064.650 4702.695 ;
        RECT 3064.990 4702.415 3065.270 4702.695 ;
        RECT 3065.610 4702.415 3065.890 4702.695 ;
        RECT 3066.230 4702.415 3066.510 4702.695 ;
        RECT 3066.850 4702.415 3067.130 4702.695 ;
        RECT 3067.470 4702.415 3067.750 4702.695 ;
        RECT 3068.090 4702.415 3068.370 4702.695 ;
        RECT 3059.410 4701.795 3059.690 4702.075 ;
        RECT 3060.030 4701.795 3060.310 4702.075 ;
        RECT 3060.650 4701.795 3060.930 4702.075 ;
        RECT 3061.270 4701.795 3061.550 4702.075 ;
        RECT 3061.890 4701.795 3062.170 4702.075 ;
        RECT 3062.510 4701.795 3062.790 4702.075 ;
        RECT 3063.130 4701.795 3063.410 4702.075 ;
        RECT 3063.750 4701.795 3064.030 4702.075 ;
        RECT 3064.370 4701.795 3064.650 4702.075 ;
        RECT 3064.990 4701.795 3065.270 4702.075 ;
        RECT 3065.610 4701.795 3065.890 4702.075 ;
        RECT 3066.230 4701.795 3066.510 4702.075 ;
        RECT 3066.850 4701.795 3067.130 4702.075 ;
        RECT 3067.470 4701.795 3067.750 4702.075 ;
        RECT 3068.090 4701.795 3068.370 4702.075 ;
        RECT 3059.410 4701.175 3059.690 4701.455 ;
        RECT 3060.030 4701.175 3060.310 4701.455 ;
        RECT 3060.650 4701.175 3060.930 4701.455 ;
        RECT 3061.270 4701.175 3061.550 4701.455 ;
        RECT 3061.890 4701.175 3062.170 4701.455 ;
        RECT 3062.510 4701.175 3062.790 4701.455 ;
        RECT 3063.130 4701.175 3063.410 4701.455 ;
        RECT 3063.750 4701.175 3064.030 4701.455 ;
        RECT 3064.370 4701.175 3064.650 4701.455 ;
        RECT 3064.990 4701.175 3065.270 4701.455 ;
        RECT 3065.610 4701.175 3065.890 4701.455 ;
        RECT 3066.230 4701.175 3066.510 4701.455 ;
        RECT 3066.850 4701.175 3067.130 4701.455 ;
        RECT 3067.470 4701.175 3067.750 4701.455 ;
        RECT 3068.090 4701.175 3068.370 4701.455 ;
        RECT 3059.410 4700.555 3059.690 4700.835 ;
        RECT 3060.030 4700.555 3060.310 4700.835 ;
        RECT 3060.650 4700.555 3060.930 4700.835 ;
        RECT 3061.270 4700.555 3061.550 4700.835 ;
        RECT 3061.890 4700.555 3062.170 4700.835 ;
        RECT 3062.510 4700.555 3062.790 4700.835 ;
        RECT 3063.130 4700.555 3063.410 4700.835 ;
        RECT 3063.750 4700.555 3064.030 4700.835 ;
        RECT 3064.370 4700.555 3064.650 4700.835 ;
        RECT 3064.990 4700.555 3065.270 4700.835 ;
        RECT 3065.610 4700.555 3065.890 4700.835 ;
        RECT 3066.230 4700.555 3066.510 4700.835 ;
        RECT 3066.850 4700.555 3067.130 4700.835 ;
        RECT 3067.470 4700.555 3067.750 4700.835 ;
        RECT 3068.090 4700.555 3068.370 4700.835 ;
        RECT 3059.410 4699.935 3059.690 4700.215 ;
        RECT 3060.030 4699.935 3060.310 4700.215 ;
        RECT 3060.650 4699.935 3060.930 4700.215 ;
        RECT 3061.270 4699.935 3061.550 4700.215 ;
        RECT 3061.890 4699.935 3062.170 4700.215 ;
        RECT 3062.510 4699.935 3062.790 4700.215 ;
        RECT 3063.130 4699.935 3063.410 4700.215 ;
        RECT 3063.750 4699.935 3064.030 4700.215 ;
        RECT 3064.370 4699.935 3064.650 4700.215 ;
        RECT 3064.990 4699.935 3065.270 4700.215 ;
        RECT 3065.610 4699.935 3065.890 4700.215 ;
        RECT 3066.230 4699.935 3066.510 4700.215 ;
        RECT 3066.850 4699.935 3067.130 4700.215 ;
        RECT 3067.470 4699.935 3067.750 4700.215 ;
        RECT 3068.090 4699.935 3068.370 4700.215 ;
        RECT 3059.410 4699.315 3059.690 4699.595 ;
        RECT 3060.030 4699.315 3060.310 4699.595 ;
        RECT 3060.650 4699.315 3060.930 4699.595 ;
        RECT 3061.270 4699.315 3061.550 4699.595 ;
        RECT 3061.890 4699.315 3062.170 4699.595 ;
        RECT 3062.510 4699.315 3062.790 4699.595 ;
        RECT 3063.130 4699.315 3063.410 4699.595 ;
        RECT 3063.750 4699.315 3064.030 4699.595 ;
        RECT 3064.370 4699.315 3064.650 4699.595 ;
        RECT 3064.990 4699.315 3065.270 4699.595 ;
        RECT 3065.610 4699.315 3065.890 4699.595 ;
        RECT 3066.230 4699.315 3066.510 4699.595 ;
        RECT 3066.850 4699.315 3067.130 4699.595 ;
        RECT 3067.470 4699.315 3067.750 4699.595 ;
        RECT 3068.090 4699.315 3068.370 4699.595 ;
        RECT 350.235 4393.025 350.515 4393.305 ;
        RECT 350.855 4393.025 351.135 4393.305 ;
        RECT 351.475 4393.025 351.755 4393.305 ;
        RECT 352.095 4393.025 352.375 4393.305 ;
        RECT 350.235 4392.405 350.515 4392.685 ;
        RECT 350.855 4392.405 351.135 4392.685 ;
        RECT 351.475 4392.405 351.755 4392.685 ;
        RECT 352.095 4392.405 352.375 4392.685 ;
        RECT 350.235 4391.785 350.515 4392.065 ;
        RECT 350.855 4391.785 351.135 4392.065 ;
        RECT 351.475 4391.785 351.755 4392.065 ;
        RECT 352.095 4391.785 352.375 4392.065 ;
        RECT 350.235 4391.165 350.515 4391.445 ;
        RECT 350.855 4391.165 351.135 4391.445 ;
        RECT 351.475 4391.165 351.755 4391.445 ;
        RECT 352.095 4391.165 352.375 4391.445 ;
        RECT 350.235 4390.545 350.515 4390.825 ;
        RECT 350.855 4390.545 351.135 4390.825 ;
        RECT 351.475 4390.545 351.755 4390.825 ;
        RECT 352.095 4390.545 352.375 4390.825 ;
        RECT 350.235 4389.925 350.515 4390.205 ;
        RECT 350.855 4389.925 351.135 4390.205 ;
        RECT 351.475 4389.925 351.755 4390.205 ;
        RECT 352.095 4389.925 352.375 4390.205 ;
        RECT 350.235 4389.305 350.515 4389.585 ;
        RECT 350.855 4389.305 351.135 4389.585 ;
        RECT 351.475 4389.305 351.755 4389.585 ;
        RECT 352.095 4389.305 352.375 4389.585 ;
        RECT 350.235 4388.685 350.515 4388.965 ;
        RECT 350.855 4388.685 351.135 4388.965 ;
        RECT 351.475 4388.685 351.755 4388.965 ;
        RECT 352.095 4388.685 352.375 4388.965 ;
        RECT 350.235 4388.065 350.515 4388.345 ;
        RECT 350.855 4388.065 351.135 4388.345 ;
        RECT 351.475 4388.065 351.755 4388.345 ;
        RECT 352.095 4388.065 352.375 4388.345 ;
        RECT 350.235 4387.445 350.515 4387.725 ;
        RECT 350.855 4387.445 351.135 4387.725 ;
        RECT 351.475 4387.445 351.755 4387.725 ;
        RECT 352.095 4387.445 352.375 4387.725 ;
        RECT 350.235 4386.825 350.515 4387.105 ;
        RECT 350.855 4386.825 351.135 4387.105 ;
        RECT 351.475 4386.825 351.755 4387.105 ;
        RECT 352.095 4386.825 352.375 4387.105 ;
        RECT 350.235 4386.205 350.515 4386.485 ;
        RECT 350.855 4386.205 351.135 4386.485 ;
        RECT 351.475 4386.205 351.755 4386.485 ;
        RECT 352.095 4386.205 352.375 4386.485 ;
        RECT 350.235 4385.585 350.515 4385.865 ;
        RECT 350.855 4385.585 351.135 4385.865 ;
        RECT 351.475 4385.585 351.755 4385.865 ;
        RECT 352.095 4385.585 352.375 4385.865 ;
        RECT 350.235 4384.965 350.515 4385.245 ;
        RECT 350.855 4384.965 351.135 4385.245 ;
        RECT 351.475 4384.965 351.755 4385.245 ;
        RECT 352.095 4384.965 352.375 4385.245 ;
        RECT 350.235 4384.345 350.515 4384.625 ;
        RECT 350.855 4384.345 351.135 4384.625 ;
        RECT 351.475 4384.345 351.755 4384.625 ;
        RECT 352.095 4384.345 352.375 4384.625 ;
        RECT 3527.625 4388.155 3527.905 4388.435 ;
        RECT 3528.245 4388.155 3528.525 4388.435 ;
        RECT 3528.865 4388.155 3529.145 4388.435 ;
        RECT 3529.485 4388.155 3529.765 4388.435 ;
        RECT 3527.625 4387.535 3527.905 4387.815 ;
        RECT 3528.245 4387.535 3528.525 4387.815 ;
        RECT 3528.865 4387.535 3529.145 4387.815 ;
        RECT 3529.485 4387.535 3529.765 4387.815 ;
        RECT 3527.625 4386.915 3527.905 4387.195 ;
        RECT 3528.245 4386.915 3528.525 4387.195 ;
        RECT 3528.865 4386.915 3529.145 4387.195 ;
        RECT 3529.485 4386.915 3529.765 4387.195 ;
        RECT 3527.625 4386.295 3527.905 4386.575 ;
        RECT 3528.245 4386.295 3528.525 4386.575 ;
        RECT 3528.865 4386.295 3529.145 4386.575 ;
        RECT 3529.485 4386.295 3529.765 4386.575 ;
        RECT 3527.625 4385.675 3527.905 4385.955 ;
        RECT 3528.245 4385.675 3528.525 4385.955 ;
        RECT 3528.865 4385.675 3529.145 4385.955 ;
        RECT 3529.485 4385.675 3529.765 4385.955 ;
        RECT 3527.625 4385.055 3527.905 4385.335 ;
        RECT 3528.245 4385.055 3528.525 4385.335 ;
        RECT 3528.865 4385.055 3529.145 4385.335 ;
        RECT 3529.485 4385.055 3529.765 4385.335 ;
        RECT 3527.625 4384.435 3527.905 4384.715 ;
        RECT 3528.245 4384.435 3528.525 4384.715 ;
        RECT 3528.865 4384.435 3529.145 4384.715 ;
        RECT 3529.485 4384.435 3529.765 4384.715 ;
        RECT 3527.625 4383.815 3527.905 4384.095 ;
        RECT 3528.245 4383.815 3528.525 4384.095 ;
        RECT 3528.865 4383.815 3529.145 4384.095 ;
        RECT 3529.485 4383.815 3529.765 4384.095 ;
        RECT 3527.625 4383.195 3527.905 4383.475 ;
        RECT 3528.245 4383.195 3528.525 4383.475 ;
        RECT 3528.865 4383.195 3529.145 4383.475 ;
        RECT 3529.485 4383.195 3529.765 4383.475 ;
        RECT 3527.625 4382.575 3527.905 4382.855 ;
        RECT 3528.245 4382.575 3528.525 4382.855 ;
        RECT 3528.865 4382.575 3529.145 4382.855 ;
        RECT 3529.485 4382.575 3529.765 4382.855 ;
        RECT 3527.625 4381.955 3527.905 4382.235 ;
        RECT 3528.245 4381.955 3528.525 4382.235 ;
        RECT 3528.865 4381.955 3529.145 4382.235 ;
        RECT 3529.485 4381.955 3529.765 4382.235 ;
        RECT 3527.625 4381.335 3527.905 4381.615 ;
        RECT 3528.245 4381.335 3528.525 4381.615 ;
        RECT 3528.865 4381.335 3529.145 4381.615 ;
        RECT 3529.485 4381.335 3529.765 4381.615 ;
        RECT 350.235 4380.625 350.515 4380.905 ;
        RECT 350.855 4380.625 351.135 4380.905 ;
        RECT 351.475 4380.625 351.755 4380.905 ;
        RECT 352.095 4380.625 352.375 4380.905 ;
        RECT 350.235 4380.005 350.515 4380.285 ;
        RECT 350.855 4380.005 351.135 4380.285 ;
        RECT 351.475 4380.005 351.755 4380.285 ;
        RECT 352.095 4380.005 352.375 4380.285 ;
        RECT 350.235 4379.385 350.515 4379.665 ;
        RECT 350.855 4379.385 351.135 4379.665 ;
        RECT 351.475 4379.385 351.755 4379.665 ;
        RECT 352.095 4379.385 352.375 4379.665 ;
        RECT 3527.625 4380.715 3527.905 4380.995 ;
        RECT 3528.245 4380.715 3528.525 4380.995 ;
        RECT 3528.865 4380.715 3529.145 4380.995 ;
        RECT 3529.485 4380.715 3529.765 4380.995 ;
        RECT 3527.625 4380.095 3527.905 4380.375 ;
        RECT 3528.245 4380.095 3528.525 4380.375 ;
        RECT 3528.865 4380.095 3529.145 4380.375 ;
        RECT 3529.485 4380.095 3529.765 4380.375 ;
        RECT 3527.625 4379.475 3527.905 4379.755 ;
        RECT 3528.245 4379.475 3528.525 4379.755 ;
        RECT 3528.865 4379.475 3529.145 4379.755 ;
        RECT 3529.485 4379.475 3529.765 4379.755 ;
        RECT 350.235 4378.765 350.515 4379.045 ;
        RECT 350.855 4378.765 351.135 4379.045 ;
        RECT 351.475 4378.765 351.755 4379.045 ;
        RECT 352.095 4378.765 352.375 4379.045 ;
        RECT 350.235 4378.145 350.515 4378.425 ;
        RECT 350.855 4378.145 351.135 4378.425 ;
        RECT 351.475 4378.145 351.755 4378.425 ;
        RECT 352.095 4378.145 352.375 4378.425 ;
        RECT 350.235 4377.525 350.515 4377.805 ;
        RECT 350.855 4377.525 351.135 4377.805 ;
        RECT 351.475 4377.525 351.755 4377.805 ;
        RECT 352.095 4377.525 352.375 4377.805 ;
        RECT 350.235 4376.905 350.515 4377.185 ;
        RECT 350.855 4376.905 351.135 4377.185 ;
        RECT 351.475 4376.905 351.755 4377.185 ;
        RECT 352.095 4376.905 352.375 4377.185 ;
        RECT 350.235 4376.285 350.515 4376.565 ;
        RECT 350.855 4376.285 351.135 4376.565 ;
        RECT 351.475 4376.285 351.755 4376.565 ;
        RECT 352.095 4376.285 352.375 4376.565 ;
        RECT 350.235 4375.665 350.515 4375.945 ;
        RECT 350.855 4375.665 351.135 4375.945 ;
        RECT 351.475 4375.665 351.755 4375.945 ;
        RECT 352.095 4375.665 352.375 4375.945 ;
        RECT 350.235 4375.045 350.515 4375.325 ;
        RECT 350.855 4375.045 351.135 4375.325 ;
        RECT 351.475 4375.045 351.755 4375.325 ;
        RECT 352.095 4375.045 352.375 4375.325 ;
        RECT 350.235 4374.425 350.515 4374.705 ;
        RECT 350.855 4374.425 351.135 4374.705 ;
        RECT 351.475 4374.425 351.755 4374.705 ;
        RECT 352.095 4374.425 352.375 4374.705 ;
        RECT 350.235 4373.805 350.515 4374.085 ;
        RECT 350.855 4373.805 351.135 4374.085 ;
        RECT 351.475 4373.805 351.755 4374.085 ;
        RECT 352.095 4373.805 352.375 4374.085 ;
        RECT 350.235 4373.185 350.515 4373.465 ;
        RECT 350.855 4373.185 351.135 4373.465 ;
        RECT 351.475 4373.185 351.755 4373.465 ;
        RECT 352.095 4373.185 352.375 4373.465 ;
        RECT 350.235 4372.565 350.515 4372.845 ;
        RECT 350.855 4372.565 351.135 4372.845 ;
        RECT 351.475 4372.565 351.755 4372.845 ;
        RECT 352.095 4372.565 352.375 4372.845 ;
        RECT 350.235 4371.945 350.515 4372.225 ;
        RECT 350.855 4371.945 351.135 4372.225 ;
        RECT 351.475 4371.945 351.755 4372.225 ;
        RECT 352.095 4371.945 352.375 4372.225 ;
        RECT 350.235 4371.325 350.515 4371.605 ;
        RECT 350.855 4371.325 351.135 4371.605 ;
        RECT 351.475 4371.325 351.755 4371.605 ;
        RECT 352.095 4371.325 352.375 4371.605 ;
        RECT 3527.625 4375.625 3527.905 4375.905 ;
        RECT 3528.245 4375.625 3528.525 4375.905 ;
        RECT 3528.865 4375.625 3529.145 4375.905 ;
        RECT 3529.485 4375.625 3529.765 4375.905 ;
        RECT 3527.625 4375.005 3527.905 4375.285 ;
        RECT 3528.245 4375.005 3528.525 4375.285 ;
        RECT 3528.865 4375.005 3529.145 4375.285 ;
        RECT 3529.485 4375.005 3529.765 4375.285 ;
        RECT 3527.625 4374.385 3527.905 4374.665 ;
        RECT 3528.245 4374.385 3528.525 4374.665 ;
        RECT 3528.865 4374.385 3529.145 4374.665 ;
        RECT 3529.485 4374.385 3529.765 4374.665 ;
        RECT 3527.625 4373.765 3527.905 4374.045 ;
        RECT 3528.245 4373.765 3528.525 4374.045 ;
        RECT 3528.865 4373.765 3529.145 4374.045 ;
        RECT 3529.485 4373.765 3529.765 4374.045 ;
        RECT 3527.625 4373.145 3527.905 4373.425 ;
        RECT 3528.245 4373.145 3528.525 4373.425 ;
        RECT 3528.865 4373.145 3529.145 4373.425 ;
        RECT 3529.485 4373.145 3529.765 4373.425 ;
        RECT 3527.625 4372.525 3527.905 4372.805 ;
        RECT 3528.245 4372.525 3528.525 4372.805 ;
        RECT 3528.865 4372.525 3529.145 4372.805 ;
        RECT 3529.485 4372.525 3529.765 4372.805 ;
        RECT 3527.625 4371.905 3527.905 4372.185 ;
        RECT 3528.245 4371.905 3528.525 4372.185 ;
        RECT 3528.865 4371.905 3529.145 4372.185 ;
        RECT 3529.485 4371.905 3529.765 4372.185 ;
        RECT 3527.625 4371.285 3527.905 4371.565 ;
        RECT 3528.245 4371.285 3528.525 4371.565 ;
        RECT 3528.865 4371.285 3529.145 4371.565 ;
        RECT 3529.485 4371.285 3529.765 4371.565 ;
        RECT 3527.625 4370.665 3527.905 4370.945 ;
        RECT 3528.245 4370.665 3528.525 4370.945 ;
        RECT 3528.865 4370.665 3529.145 4370.945 ;
        RECT 3529.485 4370.665 3529.765 4370.945 ;
        RECT 3527.625 4370.045 3527.905 4370.325 ;
        RECT 3528.245 4370.045 3528.525 4370.325 ;
        RECT 3528.865 4370.045 3529.145 4370.325 ;
        RECT 3529.485 4370.045 3529.765 4370.325 ;
        RECT 3527.625 4369.425 3527.905 4369.705 ;
        RECT 3528.245 4369.425 3528.525 4369.705 ;
        RECT 3528.865 4369.425 3529.145 4369.705 ;
        RECT 3529.485 4369.425 3529.765 4369.705 ;
        RECT 350.235 4368.775 350.515 4369.055 ;
        RECT 350.855 4368.775 351.135 4369.055 ;
        RECT 351.475 4368.775 351.755 4369.055 ;
        RECT 352.095 4368.775 352.375 4369.055 ;
        RECT 350.235 4368.155 350.515 4368.435 ;
        RECT 350.855 4368.155 351.135 4368.435 ;
        RECT 351.475 4368.155 351.755 4368.435 ;
        RECT 352.095 4368.155 352.375 4368.435 ;
        RECT 350.235 4367.535 350.515 4367.815 ;
        RECT 350.855 4367.535 351.135 4367.815 ;
        RECT 351.475 4367.535 351.755 4367.815 ;
        RECT 352.095 4367.535 352.375 4367.815 ;
        RECT 350.235 4366.915 350.515 4367.195 ;
        RECT 350.855 4366.915 351.135 4367.195 ;
        RECT 351.475 4366.915 351.755 4367.195 ;
        RECT 352.095 4366.915 352.375 4367.195 ;
        RECT 350.235 4366.295 350.515 4366.575 ;
        RECT 350.855 4366.295 351.135 4366.575 ;
        RECT 351.475 4366.295 351.755 4366.575 ;
        RECT 352.095 4366.295 352.375 4366.575 ;
        RECT 3527.625 4368.805 3527.905 4369.085 ;
        RECT 3528.245 4368.805 3528.525 4369.085 ;
        RECT 3528.865 4368.805 3529.145 4369.085 ;
        RECT 3529.485 4368.805 3529.765 4369.085 ;
        RECT 3527.625 4368.185 3527.905 4368.465 ;
        RECT 3528.245 4368.185 3528.525 4368.465 ;
        RECT 3528.865 4368.185 3529.145 4368.465 ;
        RECT 3529.485 4368.185 3529.765 4368.465 ;
        RECT 3527.625 4367.565 3527.905 4367.845 ;
        RECT 3528.245 4367.565 3528.525 4367.845 ;
        RECT 3528.865 4367.565 3529.145 4367.845 ;
        RECT 3529.485 4367.565 3529.765 4367.845 ;
        RECT 3527.625 4366.945 3527.905 4367.225 ;
        RECT 3528.245 4366.945 3528.525 4367.225 ;
        RECT 3528.865 4366.945 3529.145 4367.225 ;
        RECT 3529.485 4366.945 3529.765 4367.225 ;
        RECT 3527.625 4366.325 3527.905 4366.605 ;
        RECT 3528.245 4366.325 3528.525 4366.605 ;
        RECT 3528.865 4366.325 3529.145 4366.605 ;
        RECT 3529.485 4366.325 3529.765 4366.605 ;
        RECT 350.235 4365.675 350.515 4365.955 ;
        RECT 350.855 4365.675 351.135 4365.955 ;
        RECT 351.475 4365.675 351.755 4365.955 ;
        RECT 352.095 4365.675 352.375 4365.955 ;
        RECT 350.235 4365.055 350.515 4365.335 ;
        RECT 350.855 4365.055 351.135 4365.335 ;
        RECT 351.475 4365.055 351.755 4365.335 ;
        RECT 352.095 4365.055 352.375 4365.335 ;
        RECT 350.235 4364.435 350.515 4364.715 ;
        RECT 350.855 4364.435 351.135 4364.715 ;
        RECT 351.475 4364.435 351.755 4364.715 ;
        RECT 352.095 4364.435 352.375 4364.715 ;
        RECT 350.235 4363.815 350.515 4364.095 ;
        RECT 350.855 4363.815 351.135 4364.095 ;
        RECT 351.475 4363.815 351.755 4364.095 ;
        RECT 352.095 4363.815 352.375 4364.095 ;
        RECT 350.235 4363.195 350.515 4363.475 ;
        RECT 350.855 4363.195 351.135 4363.475 ;
        RECT 351.475 4363.195 351.755 4363.475 ;
        RECT 352.095 4363.195 352.375 4363.475 ;
        RECT 350.235 4362.575 350.515 4362.855 ;
        RECT 350.855 4362.575 351.135 4362.855 ;
        RECT 351.475 4362.575 351.755 4362.855 ;
        RECT 352.095 4362.575 352.375 4362.855 ;
        RECT 350.235 4361.955 350.515 4362.235 ;
        RECT 350.855 4361.955 351.135 4362.235 ;
        RECT 351.475 4361.955 351.755 4362.235 ;
        RECT 352.095 4361.955 352.375 4362.235 ;
        RECT 350.235 4361.335 350.515 4361.615 ;
        RECT 350.855 4361.335 351.135 4361.615 ;
        RECT 351.475 4361.335 351.755 4361.615 ;
        RECT 352.095 4361.335 352.375 4361.615 ;
        RECT 350.235 4360.715 350.515 4360.995 ;
        RECT 350.855 4360.715 351.135 4360.995 ;
        RECT 351.475 4360.715 351.755 4360.995 ;
        RECT 352.095 4360.715 352.375 4360.995 ;
        RECT 350.235 4360.095 350.515 4360.375 ;
        RECT 350.855 4360.095 351.135 4360.375 ;
        RECT 351.475 4360.095 351.755 4360.375 ;
        RECT 352.095 4360.095 352.375 4360.375 ;
        RECT 350.235 4359.475 350.515 4359.755 ;
        RECT 350.855 4359.475 351.135 4359.755 ;
        RECT 351.475 4359.475 351.755 4359.755 ;
        RECT 352.095 4359.475 352.375 4359.755 ;
        RECT 3527.625 4363.775 3527.905 4364.055 ;
        RECT 3528.245 4363.775 3528.525 4364.055 ;
        RECT 3528.865 4363.775 3529.145 4364.055 ;
        RECT 3529.485 4363.775 3529.765 4364.055 ;
        RECT 3527.625 4363.155 3527.905 4363.435 ;
        RECT 3528.245 4363.155 3528.525 4363.435 ;
        RECT 3528.865 4363.155 3529.145 4363.435 ;
        RECT 3529.485 4363.155 3529.765 4363.435 ;
        RECT 3527.625 4362.535 3527.905 4362.815 ;
        RECT 3528.245 4362.535 3528.525 4362.815 ;
        RECT 3528.865 4362.535 3529.145 4362.815 ;
        RECT 3529.485 4362.535 3529.765 4362.815 ;
        RECT 3527.625 4361.915 3527.905 4362.195 ;
        RECT 3528.245 4361.915 3528.525 4362.195 ;
        RECT 3528.865 4361.915 3529.145 4362.195 ;
        RECT 3529.485 4361.915 3529.765 4362.195 ;
        RECT 3527.625 4361.295 3527.905 4361.575 ;
        RECT 3528.245 4361.295 3528.525 4361.575 ;
        RECT 3528.865 4361.295 3529.145 4361.575 ;
        RECT 3529.485 4361.295 3529.765 4361.575 ;
        RECT 3527.625 4360.675 3527.905 4360.955 ;
        RECT 3528.245 4360.675 3528.525 4360.955 ;
        RECT 3528.865 4360.675 3529.145 4360.955 ;
        RECT 3529.485 4360.675 3529.765 4360.955 ;
        RECT 3527.625 4360.055 3527.905 4360.335 ;
        RECT 3528.245 4360.055 3528.525 4360.335 ;
        RECT 3528.865 4360.055 3529.145 4360.335 ;
        RECT 3529.485 4360.055 3529.765 4360.335 ;
        RECT 3527.625 4359.435 3527.905 4359.715 ;
        RECT 3528.245 4359.435 3528.525 4359.715 ;
        RECT 3528.865 4359.435 3529.145 4359.715 ;
        RECT 3529.485 4359.435 3529.765 4359.715 ;
        RECT 3527.625 4358.815 3527.905 4359.095 ;
        RECT 3528.245 4358.815 3528.525 4359.095 ;
        RECT 3528.865 4358.815 3529.145 4359.095 ;
        RECT 3529.485 4358.815 3529.765 4359.095 ;
        RECT 3527.625 4358.195 3527.905 4358.475 ;
        RECT 3528.245 4358.195 3528.525 4358.475 ;
        RECT 3528.865 4358.195 3529.145 4358.475 ;
        RECT 3529.485 4358.195 3529.765 4358.475 ;
        RECT 3527.625 4357.575 3527.905 4357.855 ;
        RECT 3528.245 4357.575 3528.525 4357.855 ;
        RECT 3528.865 4357.575 3529.145 4357.855 ;
        RECT 3529.485 4357.575 3529.765 4357.855 ;
        RECT 3527.625 4356.955 3527.905 4357.235 ;
        RECT 3528.245 4356.955 3528.525 4357.235 ;
        RECT 3528.865 4356.955 3529.145 4357.235 ;
        RECT 3529.485 4356.955 3529.765 4357.235 ;
        RECT 3527.625 4356.335 3527.905 4356.615 ;
        RECT 3528.245 4356.335 3528.525 4356.615 ;
        RECT 3528.865 4356.335 3529.145 4356.615 ;
        RECT 3529.485 4356.335 3529.765 4356.615 ;
        RECT 350.235 4355.245 350.515 4355.525 ;
        RECT 350.855 4355.245 351.135 4355.525 ;
        RECT 351.475 4355.245 351.755 4355.525 ;
        RECT 352.095 4355.245 352.375 4355.525 ;
        RECT 350.235 4354.625 350.515 4354.905 ;
        RECT 350.855 4354.625 351.135 4354.905 ;
        RECT 351.475 4354.625 351.755 4354.905 ;
        RECT 352.095 4354.625 352.375 4354.905 ;
        RECT 350.235 4354.005 350.515 4354.285 ;
        RECT 350.855 4354.005 351.135 4354.285 ;
        RECT 351.475 4354.005 351.755 4354.285 ;
        RECT 352.095 4354.005 352.375 4354.285 ;
        RECT 3527.625 4355.715 3527.905 4355.995 ;
        RECT 3528.245 4355.715 3528.525 4355.995 ;
        RECT 3528.865 4355.715 3529.145 4355.995 ;
        RECT 3529.485 4355.715 3529.765 4355.995 ;
        RECT 3527.625 4355.095 3527.905 4355.375 ;
        RECT 3528.245 4355.095 3528.525 4355.375 ;
        RECT 3528.865 4355.095 3529.145 4355.375 ;
        RECT 3529.485 4355.095 3529.765 4355.375 ;
        RECT 3527.625 4354.475 3527.905 4354.755 ;
        RECT 3528.245 4354.475 3528.525 4354.755 ;
        RECT 3528.865 4354.475 3529.145 4354.755 ;
        RECT 3529.485 4354.475 3529.765 4354.755 ;
        RECT 350.235 4353.385 350.515 4353.665 ;
        RECT 350.855 4353.385 351.135 4353.665 ;
        RECT 351.475 4353.385 351.755 4353.665 ;
        RECT 352.095 4353.385 352.375 4353.665 ;
        RECT 350.235 4352.765 350.515 4353.045 ;
        RECT 350.855 4352.765 351.135 4353.045 ;
        RECT 351.475 4352.765 351.755 4353.045 ;
        RECT 352.095 4352.765 352.375 4353.045 ;
        RECT 350.235 4352.145 350.515 4352.425 ;
        RECT 350.855 4352.145 351.135 4352.425 ;
        RECT 351.475 4352.145 351.755 4352.425 ;
        RECT 352.095 4352.145 352.375 4352.425 ;
        RECT 350.235 4351.525 350.515 4351.805 ;
        RECT 350.855 4351.525 351.135 4351.805 ;
        RECT 351.475 4351.525 351.755 4351.805 ;
        RECT 352.095 4351.525 352.375 4351.805 ;
        RECT 350.235 4350.905 350.515 4351.185 ;
        RECT 350.855 4350.905 351.135 4351.185 ;
        RECT 351.475 4350.905 351.755 4351.185 ;
        RECT 352.095 4350.905 352.375 4351.185 ;
        RECT 350.235 4350.285 350.515 4350.565 ;
        RECT 350.855 4350.285 351.135 4350.565 ;
        RECT 351.475 4350.285 351.755 4350.565 ;
        RECT 352.095 4350.285 352.375 4350.565 ;
        RECT 350.235 4349.665 350.515 4349.945 ;
        RECT 350.855 4349.665 351.135 4349.945 ;
        RECT 351.475 4349.665 351.755 4349.945 ;
        RECT 352.095 4349.665 352.375 4349.945 ;
        RECT 350.235 4349.045 350.515 4349.325 ;
        RECT 350.855 4349.045 351.135 4349.325 ;
        RECT 351.475 4349.045 351.755 4349.325 ;
        RECT 352.095 4349.045 352.375 4349.325 ;
        RECT 350.235 4348.425 350.515 4348.705 ;
        RECT 350.855 4348.425 351.135 4348.705 ;
        RECT 351.475 4348.425 351.755 4348.705 ;
        RECT 352.095 4348.425 352.375 4348.705 ;
        RECT 350.235 4347.805 350.515 4348.085 ;
        RECT 350.855 4347.805 351.135 4348.085 ;
        RECT 351.475 4347.805 351.755 4348.085 ;
        RECT 352.095 4347.805 352.375 4348.085 ;
        RECT 350.235 4347.185 350.515 4347.465 ;
        RECT 350.855 4347.185 351.135 4347.465 ;
        RECT 351.475 4347.185 351.755 4347.465 ;
        RECT 352.095 4347.185 352.375 4347.465 ;
        RECT 350.235 4346.565 350.515 4346.845 ;
        RECT 350.855 4346.565 351.135 4346.845 ;
        RECT 351.475 4346.565 351.755 4346.845 ;
        RECT 352.095 4346.565 352.375 4346.845 ;
        RECT 350.235 4345.945 350.515 4346.225 ;
        RECT 350.855 4345.945 351.135 4346.225 ;
        RECT 351.475 4345.945 351.755 4346.225 ;
        RECT 352.095 4345.945 352.375 4346.225 ;
        RECT 3527.625 4350.245 3527.905 4350.525 ;
        RECT 3528.245 4350.245 3528.525 4350.525 ;
        RECT 3528.865 4350.245 3529.145 4350.525 ;
        RECT 3529.485 4350.245 3529.765 4350.525 ;
        RECT 3527.625 4349.625 3527.905 4349.905 ;
        RECT 3528.245 4349.625 3528.525 4349.905 ;
        RECT 3528.865 4349.625 3529.145 4349.905 ;
        RECT 3529.485 4349.625 3529.765 4349.905 ;
        RECT 3527.625 4349.005 3527.905 4349.285 ;
        RECT 3528.245 4349.005 3528.525 4349.285 ;
        RECT 3528.865 4349.005 3529.145 4349.285 ;
        RECT 3529.485 4349.005 3529.765 4349.285 ;
        RECT 3527.625 4348.385 3527.905 4348.665 ;
        RECT 3528.245 4348.385 3528.525 4348.665 ;
        RECT 3528.865 4348.385 3529.145 4348.665 ;
        RECT 3529.485 4348.385 3529.765 4348.665 ;
        RECT 3527.625 4347.765 3527.905 4348.045 ;
        RECT 3528.245 4347.765 3528.525 4348.045 ;
        RECT 3528.865 4347.765 3529.145 4348.045 ;
        RECT 3529.485 4347.765 3529.765 4348.045 ;
        RECT 3527.625 4347.145 3527.905 4347.425 ;
        RECT 3528.245 4347.145 3528.525 4347.425 ;
        RECT 3528.865 4347.145 3529.145 4347.425 ;
        RECT 3529.485 4347.145 3529.765 4347.425 ;
        RECT 3527.625 4346.525 3527.905 4346.805 ;
        RECT 3528.245 4346.525 3528.525 4346.805 ;
        RECT 3528.865 4346.525 3529.145 4346.805 ;
        RECT 3529.485 4346.525 3529.765 4346.805 ;
        RECT 3527.625 4345.905 3527.905 4346.185 ;
        RECT 3528.245 4345.905 3528.525 4346.185 ;
        RECT 3528.865 4345.905 3529.145 4346.185 ;
        RECT 3529.485 4345.905 3529.765 4346.185 ;
        RECT 3527.625 4345.285 3527.905 4345.565 ;
        RECT 3528.245 4345.285 3528.525 4345.565 ;
        RECT 3528.865 4345.285 3529.145 4345.565 ;
        RECT 3529.485 4345.285 3529.765 4345.565 ;
        RECT 3527.625 4344.665 3527.905 4344.945 ;
        RECT 3528.245 4344.665 3528.525 4344.945 ;
        RECT 3528.865 4344.665 3529.145 4344.945 ;
        RECT 3529.485 4344.665 3529.765 4344.945 ;
        RECT 3527.625 4344.045 3527.905 4344.325 ;
        RECT 3528.245 4344.045 3528.525 4344.325 ;
        RECT 3528.865 4344.045 3529.145 4344.325 ;
        RECT 3529.485 4344.045 3529.765 4344.325 ;
        RECT 350.235 4343.395 350.515 4343.675 ;
        RECT 350.855 4343.395 351.135 4343.675 ;
        RECT 351.475 4343.395 351.755 4343.675 ;
        RECT 352.095 4343.395 352.375 4343.675 ;
        RECT 350.235 4342.775 350.515 4343.055 ;
        RECT 350.855 4342.775 351.135 4343.055 ;
        RECT 351.475 4342.775 351.755 4343.055 ;
        RECT 352.095 4342.775 352.375 4343.055 ;
        RECT 350.235 4342.155 350.515 4342.435 ;
        RECT 350.855 4342.155 351.135 4342.435 ;
        RECT 351.475 4342.155 351.755 4342.435 ;
        RECT 352.095 4342.155 352.375 4342.435 ;
        RECT 350.235 4341.535 350.515 4341.815 ;
        RECT 350.855 4341.535 351.135 4341.815 ;
        RECT 351.475 4341.535 351.755 4341.815 ;
        RECT 352.095 4341.535 352.375 4341.815 ;
        RECT 350.235 4340.915 350.515 4341.195 ;
        RECT 350.855 4340.915 351.135 4341.195 ;
        RECT 351.475 4340.915 351.755 4341.195 ;
        RECT 352.095 4340.915 352.375 4341.195 ;
        RECT 3527.625 4343.425 3527.905 4343.705 ;
        RECT 3528.245 4343.425 3528.525 4343.705 ;
        RECT 3528.865 4343.425 3529.145 4343.705 ;
        RECT 3529.485 4343.425 3529.765 4343.705 ;
        RECT 3527.625 4342.805 3527.905 4343.085 ;
        RECT 3528.245 4342.805 3528.525 4343.085 ;
        RECT 3528.865 4342.805 3529.145 4343.085 ;
        RECT 3529.485 4342.805 3529.765 4343.085 ;
        RECT 3527.625 4342.185 3527.905 4342.465 ;
        RECT 3528.245 4342.185 3528.525 4342.465 ;
        RECT 3528.865 4342.185 3529.145 4342.465 ;
        RECT 3529.485 4342.185 3529.765 4342.465 ;
        RECT 3527.625 4341.565 3527.905 4341.845 ;
        RECT 3528.245 4341.565 3528.525 4341.845 ;
        RECT 3528.865 4341.565 3529.145 4341.845 ;
        RECT 3529.485 4341.565 3529.765 4341.845 ;
        RECT 3527.625 4340.945 3527.905 4341.225 ;
        RECT 3528.245 4340.945 3528.525 4341.225 ;
        RECT 3528.865 4340.945 3529.145 4341.225 ;
        RECT 3529.485 4340.945 3529.765 4341.225 ;
        RECT 350.235 4340.295 350.515 4340.575 ;
        RECT 350.855 4340.295 351.135 4340.575 ;
        RECT 351.475 4340.295 351.755 4340.575 ;
        RECT 352.095 4340.295 352.375 4340.575 ;
        RECT 350.235 4339.675 350.515 4339.955 ;
        RECT 350.855 4339.675 351.135 4339.955 ;
        RECT 351.475 4339.675 351.755 4339.955 ;
        RECT 352.095 4339.675 352.375 4339.955 ;
        RECT 350.235 4339.055 350.515 4339.335 ;
        RECT 350.855 4339.055 351.135 4339.335 ;
        RECT 351.475 4339.055 351.755 4339.335 ;
        RECT 352.095 4339.055 352.375 4339.335 ;
        RECT 350.235 4338.435 350.515 4338.715 ;
        RECT 350.855 4338.435 351.135 4338.715 ;
        RECT 351.475 4338.435 351.755 4338.715 ;
        RECT 352.095 4338.435 352.375 4338.715 ;
        RECT 350.235 4337.815 350.515 4338.095 ;
        RECT 350.855 4337.815 351.135 4338.095 ;
        RECT 351.475 4337.815 351.755 4338.095 ;
        RECT 352.095 4337.815 352.375 4338.095 ;
        RECT 350.235 4337.195 350.515 4337.475 ;
        RECT 350.855 4337.195 351.135 4337.475 ;
        RECT 351.475 4337.195 351.755 4337.475 ;
        RECT 352.095 4337.195 352.375 4337.475 ;
        RECT 350.235 4336.575 350.515 4336.855 ;
        RECT 350.855 4336.575 351.135 4336.855 ;
        RECT 351.475 4336.575 351.755 4336.855 ;
        RECT 352.095 4336.575 352.375 4336.855 ;
        RECT 350.235 4335.955 350.515 4336.235 ;
        RECT 350.855 4335.955 351.135 4336.235 ;
        RECT 351.475 4335.955 351.755 4336.235 ;
        RECT 352.095 4335.955 352.375 4336.235 ;
        RECT 350.235 4335.335 350.515 4335.615 ;
        RECT 350.855 4335.335 351.135 4335.615 ;
        RECT 351.475 4335.335 351.755 4335.615 ;
        RECT 352.095 4335.335 352.375 4335.615 ;
        RECT 350.235 4334.715 350.515 4334.995 ;
        RECT 350.855 4334.715 351.135 4334.995 ;
        RECT 351.475 4334.715 351.755 4334.995 ;
        RECT 352.095 4334.715 352.375 4334.995 ;
        RECT 350.235 4334.095 350.515 4334.375 ;
        RECT 350.855 4334.095 351.135 4334.375 ;
        RECT 351.475 4334.095 351.755 4334.375 ;
        RECT 352.095 4334.095 352.375 4334.375 ;
        RECT 3527.625 4338.395 3527.905 4338.675 ;
        RECT 3528.245 4338.395 3528.525 4338.675 ;
        RECT 3528.865 4338.395 3529.145 4338.675 ;
        RECT 3529.485 4338.395 3529.765 4338.675 ;
        RECT 3527.625 4337.775 3527.905 4338.055 ;
        RECT 3528.245 4337.775 3528.525 4338.055 ;
        RECT 3528.865 4337.775 3529.145 4338.055 ;
        RECT 3529.485 4337.775 3529.765 4338.055 ;
        RECT 3527.625 4337.155 3527.905 4337.435 ;
        RECT 3528.245 4337.155 3528.525 4337.435 ;
        RECT 3528.865 4337.155 3529.145 4337.435 ;
        RECT 3529.485 4337.155 3529.765 4337.435 ;
        RECT 3527.625 4336.535 3527.905 4336.815 ;
        RECT 3528.245 4336.535 3528.525 4336.815 ;
        RECT 3528.865 4336.535 3529.145 4336.815 ;
        RECT 3529.485 4336.535 3529.765 4336.815 ;
        RECT 3527.625 4335.915 3527.905 4336.195 ;
        RECT 3528.245 4335.915 3528.525 4336.195 ;
        RECT 3528.865 4335.915 3529.145 4336.195 ;
        RECT 3529.485 4335.915 3529.765 4336.195 ;
        RECT 3527.625 4335.295 3527.905 4335.575 ;
        RECT 3528.245 4335.295 3528.525 4335.575 ;
        RECT 3528.865 4335.295 3529.145 4335.575 ;
        RECT 3529.485 4335.295 3529.765 4335.575 ;
        RECT 3527.625 4334.675 3527.905 4334.955 ;
        RECT 3528.245 4334.675 3528.525 4334.955 ;
        RECT 3528.865 4334.675 3529.145 4334.955 ;
        RECT 3529.485 4334.675 3529.765 4334.955 ;
        RECT 3527.625 4334.055 3527.905 4334.335 ;
        RECT 3528.245 4334.055 3528.525 4334.335 ;
        RECT 3528.865 4334.055 3529.145 4334.335 ;
        RECT 3529.485 4334.055 3529.765 4334.335 ;
        RECT 3527.625 4333.435 3527.905 4333.715 ;
        RECT 3528.245 4333.435 3528.525 4333.715 ;
        RECT 3528.865 4333.435 3529.145 4333.715 ;
        RECT 3529.485 4333.435 3529.765 4333.715 ;
        RECT 3527.625 4332.815 3527.905 4333.095 ;
        RECT 3528.245 4332.815 3528.525 4333.095 ;
        RECT 3528.865 4332.815 3529.145 4333.095 ;
        RECT 3529.485 4332.815 3529.765 4333.095 ;
        RECT 3527.625 4332.195 3527.905 4332.475 ;
        RECT 3528.245 4332.195 3528.525 4332.475 ;
        RECT 3528.865 4332.195 3529.145 4332.475 ;
        RECT 3529.485 4332.195 3529.765 4332.475 ;
        RECT 3527.625 4331.575 3527.905 4331.855 ;
        RECT 3528.245 4331.575 3528.525 4331.855 ;
        RECT 3528.865 4331.575 3529.145 4331.855 ;
        RECT 3529.485 4331.575 3529.765 4331.855 ;
        RECT 3527.625 4330.955 3527.905 4331.235 ;
        RECT 3528.245 4330.955 3528.525 4331.235 ;
        RECT 3528.865 4330.955 3529.145 4331.235 ;
        RECT 3529.485 4330.955 3529.765 4331.235 ;
        RECT 350.235 4330.245 350.515 4330.525 ;
        RECT 350.855 4330.245 351.135 4330.525 ;
        RECT 351.475 4330.245 351.755 4330.525 ;
        RECT 352.095 4330.245 352.375 4330.525 ;
        RECT 350.235 4329.625 350.515 4329.905 ;
        RECT 350.855 4329.625 351.135 4329.905 ;
        RECT 351.475 4329.625 351.755 4329.905 ;
        RECT 352.095 4329.625 352.375 4329.905 ;
        RECT 350.235 4329.005 350.515 4329.285 ;
        RECT 350.855 4329.005 351.135 4329.285 ;
        RECT 351.475 4329.005 351.755 4329.285 ;
        RECT 352.095 4329.005 352.375 4329.285 ;
        RECT 3527.625 4330.335 3527.905 4330.615 ;
        RECT 3528.245 4330.335 3528.525 4330.615 ;
        RECT 3528.865 4330.335 3529.145 4330.615 ;
        RECT 3529.485 4330.335 3529.765 4330.615 ;
        RECT 3527.625 4329.715 3527.905 4329.995 ;
        RECT 3528.245 4329.715 3528.525 4329.995 ;
        RECT 3528.865 4329.715 3529.145 4329.995 ;
        RECT 3529.485 4329.715 3529.765 4329.995 ;
        RECT 3527.625 4329.095 3527.905 4329.375 ;
        RECT 3528.245 4329.095 3528.525 4329.375 ;
        RECT 3528.865 4329.095 3529.145 4329.375 ;
        RECT 3529.485 4329.095 3529.765 4329.375 ;
        RECT 350.235 4328.385 350.515 4328.665 ;
        RECT 350.855 4328.385 351.135 4328.665 ;
        RECT 351.475 4328.385 351.755 4328.665 ;
        RECT 352.095 4328.385 352.375 4328.665 ;
        RECT 350.235 4327.765 350.515 4328.045 ;
        RECT 350.855 4327.765 351.135 4328.045 ;
        RECT 351.475 4327.765 351.755 4328.045 ;
        RECT 352.095 4327.765 352.375 4328.045 ;
        RECT 350.235 4327.145 350.515 4327.425 ;
        RECT 350.855 4327.145 351.135 4327.425 ;
        RECT 351.475 4327.145 351.755 4327.425 ;
        RECT 352.095 4327.145 352.375 4327.425 ;
        RECT 350.235 4326.525 350.515 4326.805 ;
        RECT 350.855 4326.525 351.135 4326.805 ;
        RECT 351.475 4326.525 351.755 4326.805 ;
        RECT 352.095 4326.525 352.375 4326.805 ;
        RECT 350.235 4325.905 350.515 4326.185 ;
        RECT 350.855 4325.905 351.135 4326.185 ;
        RECT 351.475 4325.905 351.755 4326.185 ;
        RECT 352.095 4325.905 352.375 4326.185 ;
        RECT 350.235 4325.285 350.515 4325.565 ;
        RECT 350.855 4325.285 351.135 4325.565 ;
        RECT 351.475 4325.285 351.755 4325.565 ;
        RECT 352.095 4325.285 352.375 4325.565 ;
        RECT 350.235 4324.665 350.515 4324.945 ;
        RECT 350.855 4324.665 351.135 4324.945 ;
        RECT 351.475 4324.665 351.755 4324.945 ;
        RECT 352.095 4324.665 352.375 4324.945 ;
        RECT 350.235 4324.045 350.515 4324.325 ;
        RECT 350.855 4324.045 351.135 4324.325 ;
        RECT 351.475 4324.045 351.755 4324.325 ;
        RECT 352.095 4324.045 352.375 4324.325 ;
        RECT 350.235 4323.425 350.515 4323.705 ;
        RECT 350.855 4323.425 351.135 4323.705 ;
        RECT 351.475 4323.425 351.755 4323.705 ;
        RECT 352.095 4323.425 352.375 4323.705 ;
        RECT 350.235 4322.805 350.515 4323.085 ;
        RECT 350.855 4322.805 351.135 4323.085 ;
        RECT 351.475 4322.805 351.755 4323.085 ;
        RECT 352.095 4322.805 352.375 4323.085 ;
        RECT 350.235 4322.185 350.515 4322.465 ;
        RECT 350.855 4322.185 351.135 4322.465 ;
        RECT 351.475 4322.185 351.755 4322.465 ;
        RECT 352.095 4322.185 352.375 4322.465 ;
        RECT 350.235 4321.565 350.515 4321.845 ;
        RECT 350.855 4321.565 351.135 4321.845 ;
        RECT 351.475 4321.565 351.755 4321.845 ;
        RECT 352.095 4321.565 352.375 4321.845 ;
        RECT 3527.625 4325.375 3527.905 4325.655 ;
        RECT 3528.245 4325.375 3528.525 4325.655 ;
        RECT 3528.865 4325.375 3529.145 4325.655 ;
        RECT 3529.485 4325.375 3529.765 4325.655 ;
        RECT 3527.625 4324.755 3527.905 4325.035 ;
        RECT 3528.245 4324.755 3528.525 4325.035 ;
        RECT 3528.865 4324.755 3529.145 4325.035 ;
        RECT 3529.485 4324.755 3529.765 4325.035 ;
        RECT 3527.625 4324.135 3527.905 4324.415 ;
        RECT 3528.245 4324.135 3528.525 4324.415 ;
        RECT 3528.865 4324.135 3529.145 4324.415 ;
        RECT 3529.485 4324.135 3529.765 4324.415 ;
        RECT 3527.625 4323.515 3527.905 4323.795 ;
        RECT 3528.245 4323.515 3528.525 4323.795 ;
        RECT 3528.865 4323.515 3529.145 4323.795 ;
        RECT 3529.485 4323.515 3529.765 4323.795 ;
        RECT 3527.625 4322.895 3527.905 4323.175 ;
        RECT 3528.245 4322.895 3528.525 4323.175 ;
        RECT 3528.865 4322.895 3529.145 4323.175 ;
        RECT 3529.485 4322.895 3529.765 4323.175 ;
        RECT 3527.625 4322.275 3527.905 4322.555 ;
        RECT 3528.245 4322.275 3528.525 4322.555 ;
        RECT 3528.865 4322.275 3529.145 4322.555 ;
        RECT 3529.485 4322.275 3529.765 4322.555 ;
        RECT 3527.625 4321.655 3527.905 4321.935 ;
        RECT 3528.245 4321.655 3528.525 4321.935 ;
        RECT 3528.865 4321.655 3529.145 4321.935 ;
        RECT 3529.485 4321.655 3529.765 4321.935 ;
        RECT 3527.625 4321.035 3527.905 4321.315 ;
        RECT 3528.245 4321.035 3528.525 4321.315 ;
        RECT 3528.865 4321.035 3529.145 4321.315 ;
        RECT 3529.485 4321.035 3529.765 4321.315 ;
        RECT 3527.625 4320.415 3527.905 4320.695 ;
        RECT 3528.245 4320.415 3528.525 4320.695 ;
        RECT 3528.865 4320.415 3529.145 4320.695 ;
        RECT 3529.485 4320.415 3529.765 4320.695 ;
        RECT 3527.625 4319.795 3527.905 4320.075 ;
        RECT 3528.245 4319.795 3528.525 4320.075 ;
        RECT 3528.865 4319.795 3529.145 4320.075 ;
        RECT 3529.485 4319.795 3529.765 4320.075 ;
        RECT 3527.625 4319.175 3527.905 4319.455 ;
        RECT 3528.245 4319.175 3528.525 4319.455 ;
        RECT 3528.865 4319.175 3529.145 4319.455 ;
        RECT 3529.485 4319.175 3529.765 4319.455 ;
        RECT 3527.625 4318.555 3527.905 4318.835 ;
        RECT 3528.245 4318.555 3528.525 4318.835 ;
        RECT 3528.865 4318.555 3529.145 4318.835 ;
        RECT 3529.485 4318.555 3529.765 4318.835 ;
        RECT 3527.625 4317.935 3527.905 4318.215 ;
        RECT 3528.245 4317.935 3528.525 4318.215 ;
        RECT 3528.865 4317.935 3529.145 4318.215 ;
        RECT 3529.485 4317.935 3529.765 4318.215 ;
        RECT 3527.625 4317.315 3527.905 4317.595 ;
        RECT 3528.245 4317.315 3528.525 4317.595 ;
        RECT 3528.865 4317.315 3529.145 4317.595 ;
        RECT 3529.485 4317.315 3529.765 4317.595 ;
        RECT 3527.625 4316.695 3527.905 4316.975 ;
        RECT 3528.245 4316.695 3528.525 4316.975 ;
        RECT 3528.865 4316.695 3529.145 4316.975 ;
        RECT 3529.485 4316.695 3529.765 4316.975 ;
        RECT 350.235 4188.025 350.515 4188.305 ;
        RECT 350.855 4188.025 351.135 4188.305 ;
        RECT 351.475 4188.025 351.755 4188.305 ;
        RECT 352.095 4188.025 352.375 4188.305 ;
        RECT 350.235 4187.405 350.515 4187.685 ;
        RECT 350.855 4187.405 351.135 4187.685 ;
        RECT 351.475 4187.405 351.755 4187.685 ;
        RECT 352.095 4187.405 352.375 4187.685 ;
        RECT 350.235 4186.785 350.515 4187.065 ;
        RECT 350.855 4186.785 351.135 4187.065 ;
        RECT 351.475 4186.785 351.755 4187.065 ;
        RECT 352.095 4186.785 352.375 4187.065 ;
        RECT 350.235 4186.165 350.515 4186.445 ;
        RECT 350.855 4186.165 351.135 4186.445 ;
        RECT 351.475 4186.165 351.755 4186.445 ;
        RECT 352.095 4186.165 352.375 4186.445 ;
        RECT 350.235 4185.545 350.515 4185.825 ;
        RECT 350.855 4185.545 351.135 4185.825 ;
        RECT 351.475 4185.545 351.755 4185.825 ;
        RECT 352.095 4185.545 352.375 4185.825 ;
        RECT 350.235 4184.925 350.515 4185.205 ;
        RECT 350.855 4184.925 351.135 4185.205 ;
        RECT 351.475 4184.925 351.755 4185.205 ;
        RECT 352.095 4184.925 352.375 4185.205 ;
        RECT 350.235 4184.305 350.515 4184.585 ;
        RECT 350.855 4184.305 351.135 4184.585 ;
        RECT 351.475 4184.305 351.755 4184.585 ;
        RECT 352.095 4184.305 352.375 4184.585 ;
        RECT 350.235 4183.685 350.515 4183.965 ;
        RECT 350.855 4183.685 351.135 4183.965 ;
        RECT 351.475 4183.685 351.755 4183.965 ;
        RECT 352.095 4183.685 352.375 4183.965 ;
        RECT 350.235 4183.065 350.515 4183.345 ;
        RECT 350.855 4183.065 351.135 4183.345 ;
        RECT 351.475 4183.065 351.755 4183.345 ;
        RECT 352.095 4183.065 352.375 4183.345 ;
        RECT 350.235 4182.445 350.515 4182.725 ;
        RECT 350.855 4182.445 351.135 4182.725 ;
        RECT 351.475 4182.445 351.755 4182.725 ;
        RECT 352.095 4182.445 352.375 4182.725 ;
        RECT 350.235 4181.825 350.515 4182.105 ;
        RECT 350.855 4181.825 351.135 4182.105 ;
        RECT 351.475 4181.825 351.755 4182.105 ;
        RECT 352.095 4181.825 352.375 4182.105 ;
        RECT 350.235 4181.205 350.515 4181.485 ;
        RECT 350.855 4181.205 351.135 4181.485 ;
        RECT 351.475 4181.205 351.755 4181.485 ;
        RECT 352.095 4181.205 352.375 4181.485 ;
        RECT 350.235 4180.585 350.515 4180.865 ;
        RECT 350.855 4180.585 351.135 4180.865 ;
        RECT 351.475 4180.585 351.755 4180.865 ;
        RECT 352.095 4180.585 352.375 4180.865 ;
        RECT 350.235 4179.965 350.515 4180.245 ;
        RECT 350.855 4179.965 351.135 4180.245 ;
        RECT 351.475 4179.965 351.755 4180.245 ;
        RECT 352.095 4179.965 352.375 4180.245 ;
        RECT 350.235 4179.345 350.515 4179.625 ;
        RECT 350.855 4179.345 351.135 4179.625 ;
        RECT 351.475 4179.345 351.755 4179.625 ;
        RECT 352.095 4179.345 352.375 4179.625 ;
        RECT 350.235 4175.625 350.515 4175.905 ;
        RECT 350.855 4175.625 351.135 4175.905 ;
        RECT 351.475 4175.625 351.755 4175.905 ;
        RECT 352.095 4175.625 352.375 4175.905 ;
        RECT 350.235 4175.005 350.515 4175.285 ;
        RECT 350.855 4175.005 351.135 4175.285 ;
        RECT 351.475 4175.005 351.755 4175.285 ;
        RECT 352.095 4175.005 352.375 4175.285 ;
        RECT 350.235 4174.385 350.515 4174.665 ;
        RECT 350.855 4174.385 351.135 4174.665 ;
        RECT 351.475 4174.385 351.755 4174.665 ;
        RECT 352.095 4174.385 352.375 4174.665 ;
        RECT 350.235 4173.765 350.515 4174.045 ;
        RECT 350.855 4173.765 351.135 4174.045 ;
        RECT 351.475 4173.765 351.755 4174.045 ;
        RECT 352.095 4173.765 352.375 4174.045 ;
        RECT 350.235 4173.145 350.515 4173.425 ;
        RECT 350.855 4173.145 351.135 4173.425 ;
        RECT 351.475 4173.145 351.755 4173.425 ;
        RECT 352.095 4173.145 352.375 4173.425 ;
        RECT 350.235 4172.525 350.515 4172.805 ;
        RECT 350.855 4172.525 351.135 4172.805 ;
        RECT 351.475 4172.525 351.755 4172.805 ;
        RECT 352.095 4172.525 352.375 4172.805 ;
        RECT 350.235 4171.905 350.515 4172.185 ;
        RECT 350.855 4171.905 351.135 4172.185 ;
        RECT 351.475 4171.905 351.755 4172.185 ;
        RECT 352.095 4171.905 352.375 4172.185 ;
        RECT 350.235 4171.285 350.515 4171.565 ;
        RECT 350.855 4171.285 351.135 4171.565 ;
        RECT 351.475 4171.285 351.755 4171.565 ;
        RECT 352.095 4171.285 352.375 4171.565 ;
        RECT 350.235 4170.665 350.515 4170.945 ;
        RECT 350.855 4170.665 351.135 4170.945 ;
        RECT 351.475 4170.665 351.755 4170.945 ;
        RECT 352.095 4170.665 352.375 4170.945 ;
        RECT 350.235 4170.045 350.515 4170.325 ;
        RECT 350.855 4170.045 351.135 4170.325 ;
        RECT 351.475 4170.045 351.755 4170.325 ;
        RECT 352.095 4170.045 352.375 4170.325 ;
        RECT 350.235 4169.425 350.515 4169.705 ;
        RECT 350.855 4169.425 351.135 4169.705 ;
        RECT 351.475 4169.425 351.755 4169.705 ;
        RECT 352.095 4169.425 352.375 4169.705 ;
        RECT 350.235 4168.805 350.515 4169.085 ;
        RECT 350.855 4168.805 351.135 4169.085 ;
        RECT 351.475 4168.805 351.755 4169.085 ;
        RECT 352.095 4168.805 352.375 4169.085 ;
        RECT 350.235 4168.185 350.515 4168.465 ;
        RECT 350.855 4168.185 351.135 4168.465 ;
        RECT 351.475 4168.185 351.755 4168.465 ;
        RECT 352.095 4168.185 352.375 4168.465 ;
        RECT 350.235 4167.565 350.515 4167.845 ;
        RECT 350.855 4167.565 351.135 4167.845 ;
        RECT 351.475 4167.565 351.755 4167.845 ;
        RECT 352.095 4167.565 352.375 4167.845 ;
        RECT 350.235 4166.945 350.515 4167.225 ;
        RECT 350.855 4166.945 351.135 4167.225 ;
        RECT 351.475 4166.945 351.755 4167.225 ;
        RECT 352.095 4166.945 352.375 4167.225 ;
        RECT 350.235 4166.325 350.515 4166.605 ;
        RECT 350.855 4166.325 351.135 4166.605 ;
        RECT 351.475 4166.325 351.755 4166.605 ;
        RECT 352.095 4166.325 352.375 4166.605 ;
        RECT 350.235 4163.775 350.515 4164.055 ;
        RECT 350.855 4163.775 351.135 4164.055 ;
        RECT 351.475 4163.775 351.755 4164.055 ;
        RECT 352.095 4163.775 352.375 4164.055 ;
        RECT 350.235 4163.155 350.515 4163.435 ;
        RECT 350.855 4163.155 351.135 4163.435 ;
        RECT 351.475 4163.155 351.755 4163.435 ;
        RECT 352.095 4163.155 352.375 4163.435 ;
        RECT 350.235 4162.535 350.515 4162.815 ;
        RECT 350.855 4162.535 351.135 4162.815 ;
        RECT 351.475 4162.535 351.755 4162.815 ;
        RECT 352.095 4162.535 352.375 4162.815 ;
        RECT 350.235 4161.915 350.515 4162.195 ;
        RECT 350.855 4161.915 351.135 4162.195 ;
        RECT 351.475 4161.915 351.755 4162.195 ;
        RECT 352.095 4161.915 352.375 4162.195 ;
        RECT 350.235 4161.295 350.515 4161.575 ;
        RECT 350.855 4161.295 351.135 4161.575 ;
        RECT 351.475 4161.295 351.755 4161.575 ;
        RECT 352.095 4161.295 352.375 4161.575 ;
        RECT 350.235 4160.675 350.515 4160.955 ;
        RECT 350.855 4160.675 351.135 4160.955 ;
        RECT 351.475 4160.675 351.755 4160.955 ;
        RECT 352.095 4160.675 352.375 4160.955 ;
        RECT 350.235 4160.055 350.515 4160.335 ;
        RECT 350.855 4160.055 351.135 4160.335 ;
        RECT 351.475 4160.055 351.755 4160.335 ;
        RECT 352.095 4160.055 352.375 4160.335 ;
        RECT 350.235 4159.435 350.515 4159.715 ;
        RECT 350.855 4159.435 351.135 4159.715 ;
        RECT 351.475 4159.435 351.755 4159.715 ;
        RECT 352.095 4159.435 352.375 4159.715 ;
        RECT 350.235 4158.815 350.515 4159.095 ;
        RECT 350.855 4158.815 351.135 4159.095 ;
        RECT 351.475 4158.815 351.755 4159.095 ;
        RECT 352.095 4158.815 352.375 4159.095 ;
        RECT 350.235 4158.195 350.515 4158.475 ;
        RECT 350.855 4158.195 351.135 4158.475 ;
        RECT 351.475 4158.195 351.755 4158.475 ;
        RECT 352.095 4158.195 352.375 4158.475 ;
        RECT 350.235 4157.575 350.515 4157.855 ;
        RECT 350.855 4157.575 351.135 4157.855 ;
        RECT 351.475 4157.575 351.755 4157.855 ;
        RECT 352.095 4157.575 352.375 4157.855 ;
        RECT 350.235 4156.955 350.515 4157.235 ;
        RECT 350.855 4156.955 351.135 4157.235 ;
        RECT 351.475 4156.955 351.755 4157.235 ;
        RECT 352.095 4156.955 352.375 4157.235 ;
        RECT 350.235 4156.335 350.515 4156.615 ;
        RECT 350.855 4156.335 351.135 4156.615 ;
        RECT 351.475 4156.335 351.755 4156.615 ;
        RECT 352.095 4156.335 352.375 4156.615 ;
        RECT 350.235 4155.715 350.515 4155.995 ;
        RECT 350.855 4155.715 351.135 4155.995 ;
        RECT 351.475 4155.715 351.755 4155.995 ;
        RECT 352.095 4155.715 352.375 4155.995 ;
        RECT 350.235 4155.095 350.515 4155.375 ;
        RECT 350.855 4155.095 351.135 4155.375 ;
        RECT 351.475 4155.095 351.755 4155.375 ;
        RECT 352.095 4155.095 352.375 4155.375 ;
        RECT 350.235 4154.475 350.515 4154.755 ;
        RECT 350.855 4154.475 351.135 4154.755 ;
        RECT 351.475 4154.475 351.755 4154.755 ;
        RECT 352.095 4154.475 352.375 4154.755 ;
        RECT 350.235 4150.245 350.515 4150.525 ;
        RECT 350.855 4150.245 351.135 4150.525 ;
        RECT 351.475 4150.245 351.755 4150.525 ;
        RECT 352.095 4150.245 352.375 4150.525 ;
        RECT 350.235 4149.625 350.515 4149.905 ;
        RECT 350.855 4149.625 351.135 4149.905 ;
        RECT 351.475 4149.625 351.755 4149.905 ;
        RECT 352.095 4149.625 352.375 4149.905 ;
        RECT 350.235 4149.005 350.515 4149.285 ;
        RECT 350.855 4149.005 351.135 4149.285 ;
        RECT 351.475 4149.005 351.755 4149.285 ;
        RECT 352.095 4149.005 352.375 4149.285 ;
        RECT 350.235 4148.385 350.515 4148.665 ;
        RECT 350.855 4148.385 351.135 4148.665 ;
        RECT 351.475 4148.385 351.755 4148.665 ;
        RECT 352.095 4148.385 352.375 4148.665 ;
        RECT 350.235 4147.765 350.515 4148.045 ;
        RECT 350.855 4147.765 351.135 4148.045 ;
        RECT 351.475 4147.765 351.755 4148.045 ;
        RECT 352.095 4147.765 352.375 4148.045 ;
        RECT 350.235 4147.145 350.515 4147.425 ;
        RECT 350.855 4147.145 351.135 4147.425 ;
        RECT 351.475 4147.145 351.755 4147.425 ;
        RECT 352.095 4147.145 352.375 4147.425 ;
        RECT 350.235 4146.525 350.515 4146.805 ;
        RECT 350.855 4146.525 351.135 4146.805 ;
        RECT 351.475 4146.525 351.755 4146.805 ;
        RECT 352.095 4146.525 352.375 4146.805 ;
        RECT 350.235 4145.905 350.515 4146.185 ;
        RECT 350.855 4145.905 351.135 4146.185 ;
        RECT 351.475 4145.905 351.755 4146.185 ;
        RECT 352.095 4145.905 352.375 4146.185 ;
        RECT 350.235 4145.285 350.515 4145.565 ;
        RECT 350.855 4145.285 351.135 4145.565 ;
        RECT 351.475 4145.285 351.755 4145.565 ;
        RECT 352.095 4145.285 352.375 4145.565 ;
        RECT 350.235 4144.665 350.515 4144.945 ;
        RECT 350.855 4144.665 351.135 4144.945 ;
        RECT 351.475 4144.665 351.755 4144.945 ;
        RECT 352.095 4144.665 352.375 4144.945 ;
        RECT 350.235 4144.045 350.515 4144.325 ;
        RECT 350.855 4144.045 351.135 4144.325 ;
        RECT 351.475 4144.045 351.755 4144.325 ;
        RECT 352.095 4144.045 352.375 4144.325 ;
        RECT 350.235 4143.425 350.515 4143.705 ;
        RECT 350.855 4143.425 351.135 4143.705 ;
        RECT 351.475 4143.425 351.755 4143.705 ;
        RECT 352.095 4143.425 352.375 4143.705 ;
        RECT 350.235 4142.805 350.515 4143.085 ;
        RECT 350.855 4142.805 351.135 4143.085 ;
        RECT 351.475 4142.805 351.755 4143.085 ;
        RECT 352.095 4142.805 352.375 4143.085 ;
        RECT 350.235 4142.185 350.515 4142.465 ;
        RECT 350.855 4142.185 351.135 4142.465 ;
        RECT 351.475 4142.185 351.755 4142.465 ;
        RECT 352.095 4142.185 352.375 4142.465 ;
        RECT 350.235 4141.565 350.515 4141.845 ;
        RECT 350.855 4141.565 351.135 4141.845 ;
        RECT 351.475 4141.565 351.755 4141.845 ;
        RECT 352.095 4141.565 352.375 4141.845 ;
        RECT 350.235 4140.945 350.515 4141.225 ;
        RECT 350.855 4140.945 351.135 4141.225 ;
        RECT 351.475 4140.945 351.755 4141.225 ;
        RECT 352.095 4140.945 352.375 4141.225 ;
        RECT 350.235 4138.395 350.515 4138.675 ;
        RECT 350.855 4138.395 351.135 4138.675 ;
        RECT 351.475 4138.395 351.755 4138.675 ;
        RECT 352.095 4138.395 352.375 4138.675 ;
        RECT 350.235 4137.775 350.515 4138.055 ;
        RECT 350.855 4137.775 351.135 4138.055 ;
        RECT 351.475 4137.775 351.755 4138.055 ;
        RECT 352.095 4137.775 352.375 4138.055 ;
        RECT 350.235 4137.155 350.515 4137.435 ;
        RECT 350.855 4137.155 351.135 4137.435 ;
        RECT 351.475 4137.155 351.755 4137.435 ;
        RECT 352.095 4137.155 352.375 4137.435 ;
        RECT 350.235 4136.535 350.515 4136.815 ;
        RECT 350.855 4136.535 351.135 4136.815 ;
        RECT 351.475 4136.535 351.755 4136.815 ;
        RECT 352.095 4136.535 352.375 4136.815 ;
        RECT 350.235 4135.915 350.515 4136.195 ;
        RECT 350.855 4135.915 351.135 4136.195 ;
        RECT 351.475 4135.915 351.755 4136.195 ;
        RECT 352.095 4135.915 352.375 4136.195 ;
        RECT 350.235 4135.295 350.515 4135.575 ;
        RECT 350.855 4135.295 351.135 4135.575 ;
        RECT 351.475 4135.295 351.755 4135.575 ;
        RECT 352.095 4135.295 352.375 4135.575 ;
        RECT 350.235 4134.675 350.515 4134.955 ;
        RECT 350.855 4134.675 351.135 4134.955 ;
        RECT 351.475 4134.675 351.755 4134.955 ;
        RECT 352.095 4134.675 352.375 4134.955 ;
        RECT 350.235 4134.055 350.515 4134.335 ;
        RECT 350.855 4134.055 351.135 4134.335 ;
        RECT 351.475 4134.055 351.755 4134.335 ;
        RECT 352.095 4134.055 352.375 4134.335 ;
        RECT 350.235 4133.435 350.515 4133.715 ;
        RECT 350.855 4133.435 351.135 4133.715 ;
        RECT 351.475 4133.435 351.755 4133.715 ;
        RECT 352.095 4133.435 352.375 4133.715 ;
        RECT 350.235 4132.815 350.515 4133.095 ;
        RECT 350.855 4132.815 351.135 4133.095 ;
        RECT 351.475 4132.815 351.755 4133.095 ;
        RECT 352.095 4132.815 352.375 4133.095 ;
        RECT 350.235 4132.195 350.515 4132.475 ;
        RECT 350.855 4132.195 351.135 4132.475 ;
        RECT 351.475 4132.195 351.755 4132.475 ;
        RECT 352.095 4132.195 352.375 4132.475 ;
        RECT 350.235 4131.575 350.515 4131.855 ;
        RECT 350.855 4131.575 351.135 4131.855 ;
        RECT 351.475 4131.575 351.755 4131.855 ;
        RECT 352.095 4131.575 352.375 4131.855 ;
        RECT 350.235 4130.955 350.515 4131.235 ;
        RECT 350.855 4130.955 351.135 4131.235 ;
        RECT 351.475 4130.955 351.755 4131.235 ;
        RECT 352.095 4130.955 352.375 4131.235 ;
        RECT 350.235 4130.335 350.515 4130.615 ;
        RECT 350.855 4130.335 351.135 4130.615 ;
        RECT 351.475 4130.335 351.755 4130.615 ;
        RECT 352.095 4130.335 352.375 4130.615 ;
        RECT 350.235 4129.715 350.515 4129.995 ;
        RECT 350.855 4129.715 351.135 4129.995 ;
        RECT 351.475 4129.715 351.755 4129.995 ;
        RECT 352.095 4129.715 352.375 4129.995 ;
        RECT 350.235 4129.095 350.515 4129.375 ;
        RECT 350.855 4129.095 351.135 4129.375 ;
        RECT 351.475 4129.095 351.755 4129.375 ;
        RECT 352.095 4129.095 352.375 4129.375 ;
        RECT 350.235 4125.245 350.515 4125.525 ;
        RECT 350.855 4125.245 351.135 4125.525 ;
        RECT 351.475 4125.245 351.755 4125.525 ;
        RECT 352.095 4125.245 352.375 4125.525 ;
        RECT 350.235 4124.625 350.515 4124.905 ;
        RECT 350.855 4124.625 351.135 4124.905 ;
        RECT 351.475 4124.625 351.755 4124.905 ;
        RECT 352.095 4124.625 352.375 4124.905 ;
        RECT 350.235 4124.005 350.515 4124.285 ;
        RECT 350.855 4124.005 351.135 4124.285 ;
        RECT 351.475 4124.005 351.755 4124.285 ;
        RECT 352.095 4124.005 352.375 4124.285 ;
        RECT 350.235 4123.385 350.515 4123.665 ;
        RECT 350.855 4123.385 351.135 4123.665 ;
        RECT 351.475 4123.385 351.755 4123.665 ;
        RECT 352.095 4123.385 352.375 4123.665 ;
        RECT 350.235 4122.765 350.515 4123.045 ;
        RECT 350.855 4122.765 351.135 4123.045 ;
        RECT 351.475 4122.765 351.755 4123.045 ;
        RECT 352.095 4122.765 352.375 4123.045 ;
        RECT 350.235 4122.145 350.515 4122.425 ;
        RECT 350.855 4122.145 351.135 4122.425 ;
        RECT 351.475 4122.145 351.755 4122.425 ;
        RECT 352.095 4122.145 352.375 4122.425 ;
        RECT 350.235 4121.525 350.515 4121.805 ;
        RECT 350.855 4121.525 351.135 4121.805 ;
        RECT 351.475 4121.525 351.755 4121.805 ;
        RECT 352.095 4121.525 352.375 4121.805 ;
        RECT 350.235 4120.905 350.515 4121.185 ;
        RECT 350.855 4120.905 351.135 4121.185 ;
        RECT 351.475 4120.905 351.755 4121.185 ;
        RECT 352.095 4120.905 352.375 4121.185 ;
        RECT 350.235 4120.285 350.515 4120.565 ;
        RECT 350.855 4120.285 351.135 4120.565 ;
        RECT 351.475 4120.285 351.755 4120.565 ;
        RECT 352.095 4120.285 352.375 4120.565 ;
        RECT 350.235 4119.665 350.515 4119.945 ;
        RECT 350.855 4119.665 351.135 4119.945 ;
        RECT 351.475 4119.665 351.755 4119.945 ;
        RECT 352.095 4119.665 352.375 4119.945 ;
        RECT 350.235 4119.045 350.515 4119.325 ;
        RECT 350.855 4119.045 351.135 4119.325 ;
        RECT 351.475 4119.045 351.755 4119.325 ;
        RECT 352.095 4119.045 352.375 4119.325 ;
        RECT 350.235 4118.425 350.515 4118.705 ;
        RECT 350.855 4118.425 351.135 4118.705 ;
        RECT 351.475 4118.425 351.755 4118.705 ;
        RECT 352.095 4118.425 352.375 4118.705 ;
        RECT 350.235 4117.805 350.515 4118.085 ;
        RECT 350.855 4117.805 351.135 4118.085 ;
        RECT 351.475 4117.805 351.755 4118.085 ;
        RECT 352.095 4117.805 352.375 4118.085 ;
        RECT 350.235 4117.185 350.515 4117.465 ;
        RECT 350.855 4117.185 351.135 4117.465 ;
        RECT 351.475 4117.185 351.755 4117.465 ;
        RECT 352.095 4117.185 352.375 4117.465 ;
        RECT 350.235 4116.565 350.515 4116.845 ;
        RECT 350.855 4116.565 351.135 4116.845 ;
        RECT 351.475 4116.565 351.755 4116.845 ;
        RECT 352.095 4116.565 352.375 4116.845 ;
        RECT 350.235 3983.025 350.515 3983.305 ;
        RECT 350.855 3983.025 351.135 3983.305 ;
        RECT 351.475 3983.025 351.755 3983.305 ;
        RECT 352.095 3983.025 352.375 3983.305 ;
        RECT 350.235 3982.405 350.515 3982.685 ;
        RECT 350.855 3982.405 351.135 3982.685 ;
        RECT 351.475 3982.405 351.755 3982.685 ;
        RECT 352.095 3982.405 352.375 3982.685 ;
        RECT 350.235 3981.785 350.515 3982.065 ;
        RECT 350.855 3981.785 351.135 3982.065 ;
        RECT 351.475 3981.785 351.755 3982.065 ;
        RECT 352.095 3981.785 352.375 3982.065 ;
        RECT 350.235 3981.165 350.515 3981.445 ;
        RECT 350.855 3981.165 351.135 3981.445 ;
        RECT 351.475 3981.165 351.755 3981.445 ;
        RECT 352.095 3981.165 352.375 3981.445 ;
        RECT 350.235 3980.545 350.515 3980.825 ;
        RECT 350.855 3980.545 351.135 3980.825 ;
        RECT 351.475 3980.545 351.755 3980.825 ;
        RECT 352.095 3980.545 352.375 3980.825 ;
        RECT 350.235 3979.925 350.515 3980.205 ;
        RECT 350.855 3979.925 351.135 3980.205 ;
        RECT 351.475 3979.925 351.755 3980.205 ;
        RECT 352.095 3979.925 352.375 3980.205 ;
        RECT 350.235 3979.305 350.515 3979.585 ;
        RECT 350.855 3979.305 351.135 3979.585 ;
        RECT 351.475 3979.305 351.755 3979.585 ;
        RECT 352.095 3979.305 352.375 3979.585 ;
        RECT 350.235 3978.685 350.515 3978.965 ;
        RECT 350.855 3978.685 351.135 3978.965 ;
        RECT 351.475 3978.685 351.755 3978.965 ;
        RECT 352.095 3978.685 352.375 3978.965 ;
        RECT 350.235 3978.065 350.515 3978.345 ;
        RECT 350.855 3978.065 351.135 3978.345 ;
        RECT 351.475 3978.065 351.755 3978.345 ;
        RECT 352.095 3978.065 352.375 3978.345 ;
        RECT 350.235 3977.445 350.515 3977.725 ;
        RECT 350.855 3977.445 351.135 3977.725 ;
        RECT 351.475 3977.445 351.755 3977.725 ;
        RECT 352.095 3977.445 352.375 3977.725 ;
        RECT 350.235 3976.825 350.515 3977.105 ;
        RECT 350.855 3976.825 351.135 3977.105 ;
        RECT 351.475 3976.825 351.755 3977.105 ;
        RECT 352.095 3976.825 352.375 3977.105 ;
        RECT 350.235 3976.205 350.515 3976.485 ;
        RECT 350.855 3976.205 351.135 3976.485 ;
        RECT 351.475 3976.205 351.755 3976.485 ;
        RECT 352.095 3976.205 352.375 3976.485 ;
        RECT 350.235 3975.585 350.515 3975.865 ;
        RECT 350.855 3975.585 351.135 3975.865 ;
        RECT 351.475 3975.585 351.755 3975.865 ;
        RECT 352.095 3975.585 352.375 3975.865 ;
        RECT 350.235 3974.965 350.515 3975.245 ;
        RECT 350.855 3974.965 351.135 3975.245 ;
        RECT 351.475 3974.965 351.755 3975.245 ;
        RECT 352.095 3974.965 352.375 3975.245 ;
        RECT 350.235 3974.345 350.515 3974.625 ;
        RECT 350.855 3974.345 351.135 3974.625 ;
        RECT 351.475 3974.345 351.755 3974.625 ;
        RECT 352.095 3974.345 352.375 3974.625 ;
        RECT 350.235 3970.625 350.515 3970.905 ;
        RECT 350.855 3970.625 351.135 3970.905 ;
        RECT 351.475 3970.625 351.755 3970.905 ;
        RECT 352.095 3970.625 352.375 3970.905 ;
        RECT 350.235 3970.005 350.515 3970.285 ;
        RECT 350.855 3970.005 351.135 3970.285 ;
        RECT 351.475 3970.005 351.755 3970.285 ;
        RECT 352.095 3970.005 352.375 3970.285 ;
        RECT 350.235 3969.385 350.515 3969.665 ;
        RECT 350.855 3969.385 351.135 3969.665 ;
        RECT 351.475 3969.385 351.755 3969.665 ;
        RECT 352.095 3969.385 352.375 3969.665 ;
        RECT 350.235 3968.765 350.515 3969.045 ;
        RECT 350.855 3968.765 351.135 3969.045 ;
        RECT 351.475 3968.765 351.755 3969.045 ;
        RECT 352.095 3968.765 352.375 3969.045 ;
        RECT 350.235 3968.145 350.515 3968.425 ;
        RECT 350.855 3968.145 351.135 3968.425 ;
        RECT 351.475 3968.145 351.755 3968.425 ;
        RECT 352.095 3968.145 352.375 3968.425 ;
        RECT 350.235 3967.525 350.515 3967.805 ;
        RECT 350.855 3967.525 351.135 3967.805 ;
        RECT 351.475 3967.525 351.755 3967.805 ;
        RECT 352.095 3967.525 352.375 3967.805 ;
        RECT 350.235 3966.905 350.515 3967.185 ;
        RECT 350.855 3966.905 351.135 3967.185 ;
        RECT 351.475 3966.905 351.755 3967.185 ;
        RECT 352.095 3966.905 352.375 3967.185 ;
        RECT 350.235 3966.285 350.515 3966.565 ;
        RECT 350.855 3966.285 351.135 3966.565 ;
        RECT 351.475 3966.285 351.755 3966.565 ;
        RECT 352.095 3966.285 352.375 3966.565 ;
        RECT 350.235 3965.665 350.515 3965.945 ;
        RECT 350.855 3965.665 351.135 3965.945 ;
        RECT 351.475 3965.665 351.755 3965.945 ;
        RECT 352.095 3965.665 352.375 3965.945 ;
        RECT 350.235 3965.045 350.515 3965.325 ;
        RECT 350.855 3965.045 351.135 3965.325 ;
        RECT 351.475 3965.045 351.755 3965.325 ;
        RECT 352.095 3965.045 352.375 3965.325 ;
        RECT 350.235 3964.425 350.515 3964.705 ;
        RECT 350.855 3964.425 351.135 3964.705 ;
        RECT 351.475 3964.425 351.755 3964.705 ;
        RECT 352.095 3964.425 352.375 3964.705 ;
        RECT 350.235 3963.805 350.515 3964.085 ;
        RECT 350.855 3963.805 351.135 3964.085 ;
        RECT 351.475 3963.805 351.755 3964.085 ;
        RECT 352.095 3963.805 352.375 3964.085 ;
        RECT 350.235 3963.185 350.515 3963.465 ;
        RECT 350.855 3963.185 351.135 3963.465 ;
        RECT 351.475 3963.185 351.755 3963.465 ;
        RECT 352.095 3963.185 352.375 3963.465 ;
        RECT 350.235 3962.565 350.515 3962.845 ;
        RECT 350.855 3962.565 351.135 3962.845 ;
        RECT 351.475 3962.565 351.755 3962.845 ;
        RECT 352.095 3962.565 352.375 3962.845 ;
        RECT 350.235 3961.945 350.515 3962.225 ;
        RECT 350.855 3961.945 351.135 3962.225 ;
        RECT 351.475 3961.945 351.755 3962.225 ;
        RECT 352.095 3961.945 352.375 3962.225 ;
        RECT 350.235 3961.325 350.515 3961.605 ;
        RECT 350.855 3961.325 351.135 3961.605 ;
        RECT 351.475 3961.325 351.755 3961.605 ;
        RECT 352.095 3961.325 352.375 3961.605 ;
        RECT 350.235 3958.775 350.515 3959.055 ;
        RECT 350.855 3958.775 351.135 3959.055 ;
        RECT 351.475 3958.775 351.755 3959.055 ;
        RECT 352.095 3958.775 352.375 3959.055 ;
        RECT 350.235 3958.155 350.515 3958.435 ;
        RECT 350.855 3958.155 351.135 3958.435 ;
        RECT 351.475 3958.155 351.755 3958.435 ;
        RECT 352.095 3958.155 352.375 3958.435 ;
        RECT 350.235 3957.535 350.515 3957.815 ;
        RECT 350.855 3957.535 351.135 3957.815 ;
        RECT 351.475 3957.535 351.755 3957.815 ;
        RECT 352.095 3957.535 352.375 3957.815 ;
        RECT 350.235 3956.915 350.515 3957.195 ;
        RECT 350.855 3956.915 351.135 3957.195 ;
        RECT 351.475 3956.915 351.755 3957.195 ;
        RECT 352.095 3956.915 352.375 3957.195 ;
        RECT 350.235 3956.295 350.515 3956.575 ;
        RECT 350.855 3956.295 351.135 3956.575 ;
        RECT 351.475 3956.295 351.755 3956.575 ;
        RECT 352.095 3956.295 352.375 3956.575 ;
        RECT 350.235 3955.675 350.515 3955.955 ;
        RECT 350.855 3955.675 351.135 3955.955 ;
        RECT 351.475 3955.675 351.755 3955.955 ;
        RECT 352.095 3955.675 352.375 3955.955 ;
        RECT 350.235 3955.055 350.515 3955.335 ;
        RECT 350.855 3955.055 351.135 3955.335 ;
        RECT 351.475 3955.055 351.755 3955.335 ;
        RECT 352.095 3955.055 352.375 3955.335 ;
        RECT 350.235 3954.435 350.515 3954.715 ;
        RECT 350.855 3954.435 351.135 3954.715 ;
        RECT 351.475 3954.435 351.755 3954.715 ;
        RECT 352.095 3954.435 352.375 3954.715 ;
        RECT 350.235 3953.815 350.515 3954.095 ;
        RECT 350.855 3953.815 351.135 3954.095 ;
        RECT 351.475 3953.815 351.755 3954.095 ;
        RECT 352.095 3953.815 352.375 3954.095 ;
        RECT 350.235 3953.195 350.515 3953.475 ;
        RECT 350.855 3953.195 351.135 3953.475 ;
        RECT 351.475 3953.195 351.755 3953.475 ;
        RECT 352.095 3953.195 352.375 3953.475 ;
        RECT 350.235 3952.575 350.515 3952.855 ;
        RECT 350.855 3952.575 351.135 3952.855 ;
        RECT 351.475 3952.575 351.755 3952.855 ;
        RECT 352.095 3952.575 352.375 3952.855 ;
        RECT 350.235 3951.955 350.515 3952.235 ;
        RECT 350.855 3951.955 351.135 3952.235 ;
        RECT 351.475 3951.955 351.755 3952.235 ;
        RECT 352.095 3951.955 352.375 3952.235 ;
        RECT 350.235 3951.335 350.515 3951.615 ;
        RECT 350.855 3951.335 351.135 3951.615 ;
        RECT 351.475 3951.335 351.755 3951.615 ;
        RECT 352.095 3951.335 352.375 3951.615 ;
        RECT 350.235 3950.715 350.515 3950.995 ;
        RECT 350.855 3950.715 351.135 3950.995 ;
        RECT 351.475 3950.715 351.755 3950.995 ;
        RECT 352.095 3950.715 352.375 3950.995 ;
        RECT 350.235 3950.095 350.515 3950.375 ;
        RECT 350.855 3950.095 351.135 3950.375 ;
        RECT 351.475 3950.095 351.755 3950.375 ;
        RECT 352.095 3950.095 352.375 3950.375 ;
        RECT 350.235 3949.475 350.515 3949.755 ;
        RECT 350.855 3949.475 351.135 3949.755 ;
        RECT 351.475 3949.475 351.755 3949.755 ;
        RECT 352.095 3949.475 352.375 3949.755 ;
        RECT 3527.625 3958.155 3527.905 3958.435 ;
        RECT 3528.245 3958.155 3528.525 3958.435 ;
        RECT 3528.865 3958.155 3529.145 3958.435 ;
        RECT 3529.485 3958.155 3529.765 3958.435 ;
        RECT 3527.625 3957.535 3527.905 3957.815 ;
        RECT 3528.245 3957.535 3528.525 3957.815 ;
        RECT 3528.865 3957.535 3529.145 3957.815 ;
        RECT 3529.485 3957.535 3529.765 3957.815 ;
        RECT 3527.625 3956.915 3527.905 3957.195 ;
        RECT 3528.245 3956.915 3528.525 3957.195 ;
        RECT 3528.865 3956.915 3529.145 3957.195 ;
        RECT 3529.485 3956.915 3529.765 3957.195 ;
        RECT 3527.625 3956.295 3527.905 3956.575 ;
        RECT 3528.245 3956.295 3528.525 3956.575 ;
        RECT 3528.865 3956.295 3529.145 3956.575 ;
        RECT 3529.485 3956.295 3529.765 3956.575 ;
        RECT 3527.625 3955.675 3527.905 3955.955 ;
        RECT 3528.245 3955.675 3528.525 3955.955 ;
        RECT 3528.865 3955.675 3529.145 3955.955 ;
        RECT 3529.485 3955.675 3529.765 3955.955 ;
        RECT 3527.625 3955.055 3527.905 3955.335 ;
        RECT 3528.245 3955.055 3528.525 3955.335 ;
        RECT 3528.865 3955.055 3529.145 3955.335 ;
        RECT 3529.485 3955.055 3529.765 3955.335 ;
        RECT 3527.625 3954.435 3527.905 3954.715 ;
        RECT 3528.245 3954.435 3528.525 3954.715 ;
        RECT 3528.865 3954.435 3529.145 3954.715 ;
        RECT 3529.485 3954.435 3529.765 3954.715 ;
        RECT 3527.625 3953.815 3527.905 3954.095 ;
        RECT 3528.245 3953.815 3528.525 3954.095 ;
        RECT 3528.865 3953.815 3529.145 3954.095 ;
        RECT 3529.485 3953.815 3529.765 3954.095 ;
        RECT 3527.625 3953.195 3527.905 3953.475 ;
        RECT 3528.245 3953.195 3528.525 3953.475 ;
        RECT 3528.865 3953.195 3529.145 3953.475 ;
        RECT 3529.485 3953.195 3529.765 3953.475 ;
        RECT 3527.625 3952.575 3527.905 3952.855 ;
        RECT 3528.245 3952.575 3528.525 3952.855 ;
        RECT 3528.865 3952.575 3529.145 3952.855 ;
        RECT 3529.485 3952.575 3529.765 3952.855 ;
        RECT 3527.625 3951.955 3527.905 3952.235 ;
        RECT 3528.245 3951.955 3528.525 3952.235 ;
        RECT 3528.865 3951.955 3529.145 3952.235 ;
        RECT 3529.485 3951.955 3529.765 3952.235 ;
        RECT 3527.625 3951.335 3527.905 3951.615 ;
        RECT 3528.245 3951.335 3528.525 3951.615 ;
        RECT 3528.865 3951.335 3529.145 3951.615 ;
        RECT 3529.485 3951.335 3529.765 3951.615 ;
        RECT 3527.625 3950.715 3527.905 3950.995 ;
        RECT 3528.245 3950.715 3528.525 3950.995 ;
        RECT 3528.865 3950.715 3529.145 3950.995 ;
        RECT 3529.485 3950.715 3529.765 3950.995 ;
        RECT 3527.625 3950.095 3527.905 3950.375 ;
        RECT 3528.245 3950.095 3528.525 3950.375 ;
        RECT 3528.865 3950.095 3529.145 3950.375 ;
        RECT 3529.485 3950.095 3529.765 3950.375 ;
        RECT 3527.625 3949.475 3527.905 3949.755 ;
        RECT 3528.245 3949.475 3528.525 3949.755 ;
        RECT 3528.865 3949.475 3529.145 3949.755 ;
        RECT 3529.485 3949.475 3529.765 3949.755 ;
        RECT 350.235 3945.245 350.515 3945.525 ;
        RECT 350.855 3945.245 351.135 3945.525 ;
        RECT 351.475 3945.245 351.755 3945.525 ;
        RECT 352.095 3945.245 352.375 3945.525 ;
        RECT 350.235 3944.625 350.515 3944.905 ;
        RECT 350.855 3944.625 351.135 3944.905 ;
        RECT 351.475 3944.625 351.755 3944.905 ;
        RECT 352.095 3944.625 352.375 3944.905 ;
        RECT 350.235 3944.005 350.515 3944.285 ;
        RECT 350.855 3944.005 351.135 3944.285 ;
        RECT 351.475 3944.005 351.755 3944.285 ;
        RECT 352.095 3944.005 352.375 3944.285 ;
        RECT 350.235 3943.385 350.515 3943.665 ;
        RECT 350.855 3943.385 351.135 3943.665 ;
        RECT 351.475 3943.385 351.755 3943.665 ;
        RECT 352.095 3943.385 352.375 3943.665 ;
        RECT 350.235 3942.765 350.515 3943.045 ;
        RECT 350.855 3942.765 351.135 3943.045 ;
        RECT 351.475 3942.765 351.755 3943.045 ;
        RECT 352.095 3942.765 352.375 3943.045 ;
        RECT 350.235 3942.145 350.515 3942.425 ;
        RECT 350.855 3942.145 351.135 3942.425 ;
        RECT 351.475 3942.145 351.755 3942.425 ;
        RECT 352.095 3942.145 352.375 3942.425 ;
        RECT 350.235 3941.525 350.515 3941.805 ;
        RECT 350.855 3941.525 351.135 3941.805 ;
        RECT 351.475 3941.525 351.755 3941.805 ;
        RECT 352.095 3941.525 352.375 3941.805 ;
        RECT 350.235 3940.905 350.515 3941.185 ;
        RECT 350.855 3940.905 351.135 3941.185 ;
        RECT 351.475 3940.905 351.755 3941.185 ;
        RECT 352.095 3940.905 352.375 3941.185 ;
        RECT 350.235 3940.285 350.515 3940.565 ;
        RECT 350.855 3940.285 351.135 3940.565 ;
        RECT 351.475 3940.285 351.755 3940.565 ;
        RECT 352.095 3940.285 352.375 3940.565 ;
        RECT 350.235 3939.665 350.515 3939.945 ;
        RECT 350.855 3939.665 351.135 3939.945 ;
        RECT 351.475 3939.665 351.755 3939.945 ;
        RECT 352.095 3939.665 352.375 3939.945 ;
        RECT 350.235 3939.045 350.515 3939.325 ;
        RECT 350.855 3939.045 351.135 3939.325 ;
        RECT 351.475 3939.045 351.755 3939.325 ;
        RECT 352.095 3939.045 352.375 3939.325 ;
        RECT 350.235 3938.425 350.515 3938.705 ;
        RECT 350.855 3938.425 351.135 3938.705 ;
        RECT 351.475 3938.425 351.755 3938.705 ;
        RECT 352.095 3938.425 352.375 3938.705 ;
        RECT 350.235 3937.805 350.515 3938.085 ;
        RECT 350.855 3937.805 351.135 3938.085 ;
        RECT 351.475 3937.805 351.755 3938.085 ;
        RECT 352.095 3937.805 352.375 3938.085 ;
        RECT 350.235 3937.185 350.515 3937.465 ;
        RECT 350.855 3937.185 351.135 3937.465 ;
        RECT 351.475 3937.185 351.755 3937.465 ;
        RECT 352.095 3937.185 352.375 3937.465 ;
        RECT 350.235 3936.565 350.515 3936.845 ;
        RECT 350.855 3936.565 351.135 3936.845 ;
        RECT 351.475 3936.565 351.755 3936.845 ;
        RECT 352.095 3936.565 352.375 3936.845 ;
        RECT 350.235 3935.945 350.515 3936.225 ;
        RECT 350.855 3935.945 351.135 3936.225 ;
        RECT 351.475 3935.945 351.755 3936.225 ;
        RECT 352.095 3935.945 352.375 3936.225 ;
        RECT 3527.625 3945.625 3527.905 3945.905 ;
        RECT 3528.245 3945.625 3528.525 3945.905 ;
        RECT 3528.865 3945.625 3529.145 3945.905 ;
        RECT 3529.485 3945.625 3529.765 3945.905 ;
        RECT 3527.625 3945.005 3527.905 3945.285 ;
        RECT 3528.245 3945.005 3528.525 3945.285 ;
        RECT 3528.865 3945.005 3529.145 3945.285 ;
        RECT 3529.485 3945.005 3529.765 3945.285 ;
        RECT 3527.625 3944.385 3527.905 3944.665 ;
        RECT 3528.245 3944.385 3528.525 3944.665 ;
        RECT 3528.865 3944.385 3529.145 3944.665 ;
        RECT 3529.485 3944.385 3529.765 3944.665 ;
        RECT 3527.625 3943.765 3527.905 3944.045 ;
        RECT 3528.245 3943.765 3528.525 3944.045 ;
        RECT 3528.865 3943.765 3529.145 3944.045 ;
        RECT 3529.485 3943.765 3529.765 3944.045 ;
        RECT 3527.625 3943.145 3527.905 3943.425 ;
        RECT 3528.245 3943.145 3528.525 3943.425 ;
        RECT 3528.865 3943.145 3529.145 3943.425 ;
        RECT 3529.485 3943.145 3529.765 3943.425 ;
        RECT 3527.625 3942.525 3527.905 3942.805 ;
        RECT 3528.245 3942.525 3528.525 3942.805 ;
        RECT 3528.865 3942.525 3529.145 3942.805 ;
        RECT 3529.485 3942.525 3529.765 3942.805 ;
        RECT 3527.625 3941.905 3527.905 3942.185 ;
        RECT 3528.245 3941.905 3528.525 3942.185 ;
        RECT 3528.865 3941.905 3529.145 3942.185 ;
        RECT 3529.485 3941.905 3529.765 3942.185 ;
        RECT 3527.625 3941.285 3527.905 3941.565 ;
        RECT 3528.245 3941.285 3528.525 3941.565 ;
        RECT 3528.865 3941.285 3529.145 3941.565 ;
        RECT 3529.485 3941.285 3529.765 3941.565 ;
        RECT 3527.625 3940.665 3527.905 3940.945 ;
        RECT 3528.245 3940.665 3528.525 3940.945 ;
        RECT 3528.865 3940.665 3529.145 3940.945 ;
        RECT 3529.485 3940.665 3529.765 3940.945 ;
        RECT 3527.625 3940.045 3527.905 3940.325 ;
        RECT 3528.245 3940.045 3528.525 3940.325 ;
        RECT 3528.865 3940.045 3529.145 3940.325 ;
        RECT 3529.485 3940.045 3529.765 3940.325 ;
        RECT 3527.625 3939.425 3527.905 3939.705 ;
        RECT 3528.245 3939.425 3528.525 3939.705 ;
        RECT 3528.865 3939.425 3529.145 3939.705 ;
        RECT 3529.485 3939.425 3529.765 3939.705 ;
        RECT 3527.625 3938.805 3527.905 3939.085 ;
        RECT 3528.245 3938.805 3528.525 3939.085 ;
        RECT 3528.865 3938.805 3529.145 3939.085 ;
        RECT 3529.485 3938.805 3529.765 3939.085 ;
        RECT 3527.625 3938.185 3527.905 3938.465 ;
        RECT 3528.245 3938.185 3528.525 3938.465 ;
        RECT 3528.865 3938.185 3529.145 3938.465 ;
        RECT 3529.485 3938.185 3529.765 3938.465 ;
        RECT 3527.625 3937.565 3527.905 3937.845 ;
        RECT 3528.245 3937.565 3528.525 3937.845 ;
        RECT 3528.865 3937.565 3529.145 3937.845 ;
        RECT 3529.485 3937.565 3529.765 3937.845 ;
        RECT 3527.625 3936.945 3527.905 3937.225 ;
        RECT 3528.245 3936.945 3528.525 3937.225 ;
        RECT 3528.865 3936.945 3529.145 3937.225 ;
        RECT 3529.485 3936.945 3529.765 3937.225 ;
        RECT 3527.625 3936.325 3527.905 3936.605 ;
        RECT 3528.245 3936.325 3528.525 3936.605 ;
        RECT 3528.865 3936.325 3529.145 3936.605 ;
        RECT 3529.485 3936.325 3529.765 3936.605 ;
        RECT 350.235 3933.395 350.515 3933.675 ;
        RECT 350.855 3933.395 351.135 3933.675 ;
        RECT 351.475 3933.395 351.755 3933.675 ;
        RECT 352.095 3933.395 352.375 3933.675 ;
        RECT 350.235 3932.775 350.515 3933.055 ;
        RECT 350.855 3932.775 351.135 3933.055 ;
        RECT 351.475 3932.775 351.755 3933.055 ;
        RECT 352.095 3932.775 352.375 3933.055 ;
        RECT 350.235 3932.155 350.515 3932.435 ;
        RECT 350.855 3932.155 351.135 3932.435 ;
        RECT 351.475 3932.155 351.755 3932.435 ;
        RECT 352.095 3932.155 352.375 3932.435 ;
        RECT 350.235 3931.535 350.515 3931.815 ;
        RECT 350.855 3931.535 351.135 3931.815 ;
        RECT 351.475 3931.535 351.755 3931.815 ;
        RECT 352.095 3931.535 352.375 3931.815 ;
        RECT 350.235 3930.915 350.515 3931.195 ;
        RECT 350.855 3930.915 351.135 3931.195 ;
        RECT 351.475 3930.915 351.755 3931.195 ;
        RECT 352.095 3930.915 352.375 3931.195 ;
        RECT 350.235 3930.295 350.515 3930.575 ;
        RECT 350.855 3930.295 351.135 3930.575 ;
        RECT 351.475 3930.295 351.755 3930.575 ;
        RECT 352.095 3930.295 352.375 3930.575 ;
        RECT 350.235 3929.675 350.515 3929.955 ;
        RECT 350.855 3929.675 351.135 3929.955 ;
        RECT 351.475 3929.675 351.755 3929.955 ;
        RECT 352.095 3929.675 352.375 3929.955 ;
        RECT 350.235 3929.055 350.515 3929.335 ;
        RECT 350.855 3929.055 351.135 3929.335 ;
        RECT 351.475 3929.055 351.755 3929.335 ;
        RECT 352.095 3929.055 352.375 3929.335 ;
        RECT 350.235 3928.435 350.515 3928.715 ;
        RECT 350.855 3928.435 351.135 3928.715 ;
        RECT 351.475 3928.435 351.755 3928.715 ;
        RECT 352.095 3928.435 352.375 3928.715 ;
        RECT 350.235 3927.815 350.515 3928.095 ;
        RECT 350.855 3927.815 351.135 3928.095 ;
        RECT 351.475 3927.815 351.755 3928.095 ;
        RECT 352.095 3927.815 352.375 3928.095 ;
        RECT 350.235 3927.195 350.515 3927.475 ;
        RECT 350.855 3927.195 351.135 3927.475 ;
        RECT 351.475 3927.195 351.755 3927.475 ;
        RECT 352.095 3927.195 352.375 3927.475 ;
        RECT 350.235 3926.575 350.515 3926.855 ;
        RECT 350.855 3926.575 351.135 3926.855 ;
        RECT 351.475 3926.575 351.755 3926.855 ;
        RECT 352.095 3926.575 352.375 3926.855 ;
        RECT 350.235 3925.955 350.515 3926.235 ;
        RECT 350.855 3925.955 351.135 3926.235 ;
        RECT 351.475 3925.955 351.755 3926.235 ;
        RECT 352.095 3925.955 352.375 3926.235 ;
        RECT 350.235 3925.335 350.515 3925.615 ;
        RECT 350.855 3925.335 351.135 3925.615 ;
        RECT 351.475 3925.335 351.755 3925.615 ;
        RECT 352.095 3925.335 352.375 3925.615 ;
        RECT 350.235 3924.715 350.515 3924.995 ;
        RECT 350.855 3924.715 351.135 3924.995 ;
        RECT 351.475 3924.715 351.755 3924.995 ;
        RECT 352.095 3924.715 352.375 3924.995 ;
        RECT 350.235 3924.095 350.515 3924.375 ;
        RECT 350.855 3924.095 351.135 3924.375 ;
        RECT 351.475 3924.095 351.755 3924.375 ;
        RECT 352.095 3924.095 352.375 3924.375 ;
        RECT 3527.625 3933.775 3527.905 3934.055 ;
        RECT 3528.245 3933.775 3528.525 3934.055 ;
        RECT 3528.865 3933.775 3529.145 3934.055 ;
        RECT 3529.485 3933.775 3529.765 3934.055 ;
        RECT 3527.625 3933.155 3527.905 3933.435 ;
        RECT 3528.245 3933.155 3528.525 3933.435 ;
        RECT 3528.865 3933.155 3529.145 3933.435 ;
        RECT 3529.485 3933.155 3529.765 3933.435 ;
        RECT 3527.625 3932.535 3527.905 3932.815 ;
        RECT 3528.245 3932.535 3528.525 3932.815 ;
        RECT 3528.865 3932.535 3529.145 3932.815 ;
        RECT 3529.485 3932.535 3529.765 3932.815 ;
        RECT 3527.625 3931.915 3527.905 3932.195 ;
        RECT 3528.245 3931.915 3528.525 3932.195 ;
        RECT 3528.865 3931.915 3529.145 3932.195 ;
        RECT 3529.485 3931.915 3529.765 3932.195 ;
        RECT 3527.625 3931.295 3527.905 3931.575 ;
        RECT 3528.245 3931.295 3528.525 3931.575 ;
        RECT 3528.865 3931.295 3529.145 3931.575 ;
        RECT 3529.485 3931.295 3529.765 3931.575 ;
        RECT 3527.625 3930.675 3527.905 3930.955 ;
        RECT 3528.245 3930.675 3528.525 3930.955 ;
        RECT 3528.865 3930.675 3529.145 3930.955 ;
        RECT 3529.485 3930.675 3529.765 3930.955 ;
        RECT 3527.625 3930.055 3527.905 3930.335 ;
        RECT 3528.245 3930.055 3528.525 3930.335 ;
        RECT 3528.865 3930.055 3529.145 3930.335 ;
        RECT 3529.485 3930.055 3529.765 3930.335 ;
        RECT 3527.625 3929.435 3527.905 3929.715 ;
        RECT 3528.245 3929.435 3528.525 3929.715 ;
        RECT 3528.865 3929.435 3529.145 3929.715 ;
        RECT 3529.485 3929.435 3529.765 3929.715 ;
        RECT 3527.625 3928.815 3527.905 3929.095 ;
        RECT 3528.245 3928.815 3528.525 3929.095 ;
        RECT 3528.865 3928.815 3529.145 3929.095 ;
        RECT 3529.485 3928.815 3529.765 3929.095 ;
        RECT 3527.625 3928.195 3527.905 3928.475 ;
        RECT 3528.245 3928.195 3528.525 3928.475 ;
        RECT 3528.865 3928.195 3529.145 3928.475 ;
        RECT 3529.485 3928.195 3529.765 3928.475 ;
        RECT 3527.625 3927.575 3527.905 3927.855 ;
        RECT 3528.245 3927.575 3528.525 3927.855 ;
        RECT 3528.865 3927.575 3529.145 3927.855 ;
        RECT 3529.485 3927.575 3529.765 3927.855 ;
        RECT 3527.625 3926.955 3527.905 3927.235 ;
        RECT 3528.245 3926.955 3528.525 3927.235 ;
        RECT 3528.865 3926.955 3529.145 3927.235 ;
        RECT 3529.485 3926.955 3529.765 3927.235 ;
        RECT 3527.625 3926.335 3527.905 3926.615 ;
        RECT 3528.245 3926.335 3528.525 3926.615 ;
        RECT 3528.865 3926.335 3529.145 3926.615 ;
        RECT 3529.485 3926.335 3529.765 3926.615 ;
        RECT 3527.625 3925.715 3527.905 3925.995 ;
        RECT 3528.245 3925.715 3528.525 3925.995 ;
        RECT 3528.865 3925.715 3529.145 3925.995 ;
        RECT 3529.485 3925.715 3529.765 3925.995 ;
        RECT 3527.625 3925.095 3527.905 3925.375 ;
        RECT 3528.245 3925.095 3528.525 3925.375 ;
        RECT 3528.865 3925.095 3529.145 3925.375 ;
        RECT 3529.485 3925.095 3529.765 3925.375 ;
        RECT 3527.625 3924.475 3527.905 3924.755 ;
        RECT 3528.245 3924.475 3528.525 3924.755 ;
        RECT 3528.865 3924.475 3529.145 3924.755 ;
        RECT 3529.485 3924.475 3529.765 3924.755 ;
        RECT 350.235 3920.245 350.515 3920.525 ;
        RECT 350.855 3920.245 351.135 3920.525 ;
        RECT 351.475 3920.245 351.755 3920.525 ;
        RECT 352.095 3920.245 352.375 3920.525 ;
        RECT 350.235 3919.625 350.515 3919.905 ;
        RECT 350.855 3919.625 351.135 3919.905 ;
        RECT 351.475 3919.625 351.755 3919.905 ;
        RECT 352.095 3919.625 352.375 3919.905 ;
        RECT 350.235 3919.005 350.515 3919.285 ;
        RECT 350.855 3919.005 351.135 3919.285 ;
        RECT 351.475 3919.005 351.755 3919.285 ;
        RECT 352.095 3919.005 352.375 3919.285 ;
        RECT 350.235 3918.385 350.515 3918.665 ;
        RECT 350.855 3918.385 351.135 3918.665 ;
        RECT 351.475 3918.385 351.755 3918.665 ;
        RECT 352.095 3918.385 352.375 3918.665 ;
        RECT 350.235 3917.765 350.515 3918.045 ;
        RECT 350.855 3917.765 351.135 3918.045 ;
        RECT 351.475 3917.765 351.755 3918.045 ;
        RECT 352.095 3917.765 352.375 3918.045 ;
        RECT 350.235 3917.145 350.515 3917.425 ;
        RECT 350.855 3917.145 351.135 3917.425 ;
        RECT 351.475 3917.145 351.755 3917.425 ;
        RECT 352.095 3917.145 352.375 3917.425 ;
        RECT 350.235 3916.525 350.515 3916.805 ;
        RECT 350.855 3916.525 351.135 3916.805 ;
        RECT 351.475 3916.525 351.755 3916.805 ;
        RECT 352.095 3916.525 352.375 3916.805 ;
        RECT 350.235 3915.905 350.515 3916.185 ;
        RECT 350.855 3915.905 351.135 3916.185 ;
        RECT 351.475 3915.905 351.755 3916.185 ;
        RECT 352.095 3915.905 352.375 3916.185 ;
        RECT 350.235 3915.285 350.515 3915.565 ;
        RECT 350.855 3915.285 351.135 3915.565 ;
        RECT 351.475 3915.285 351.755 3915.565 ;
        RECT 352.095 3915.285 352.375 3915.565 ;
        RECT 350.235 3914.665 350.515 3914.945 ;
        RECT 350.855 3914.665 351.135 3914.945 ;
        RECT 351.475 3914.665 351.755 3914.945 ;
        RECT 352.095 3914.665 352.375 3914.945 ;
        RECT 350.235 3914.045 350.515 3914.325 ;
        RECT 350.855 3914.045 351.135 3914.325 ;
        RECT 351.475 3914.045 351.755 3914.325 ;
        RECT 352.095 3914.045 352.375 3914.325 ;
        RECT 350.235 3913.425 350.515 3913.705 ;
        RECT 350.855 3913.425 351.135 3913.705 ;
        RECT 351.475 3913.425 351.755 3913.705 ;
        RECT 352.095 3913.425 352.375 3913.705 ;
        RECT 350.235 3912.805 350.515 3913.085 ;
        RECT 350.855 3912.805 351.135 3913.085 ;
        RECT 351.475 3912.805 351.755 3913.085 ;
        RECT 352.095 3912.805 352.375 3913.085 ;
        RECT 350.235 3912.185 350.515 3912.465 ;
        RECT 350.855 3912.185 351.135 3912.465 ;
        RECT 351.475 3912.185 351.755 3912.465 ;
        RECT 352.095 3912.185 352.375 3912.465 ;
        RECT 350.235 3911.565 350.515 3911.845 ;
        RECT 350.855 3911.565 351.135 3911.845 ;
        RECT 351.475 3911.565 351.755 3911.845 ;
        RECT 352.095 3911.565 352.375 3911.845 ;
        RECT 3527.625 3920.245 3527.905 3920.525 ;
        RECT 3528.245 3920.245 3528.525 3920.525 ;
        RECT 3528.865 3920.245 3529.145 3920.525 ;
        RECT 3529.485 3920.245 3529.765 3920.525 ;
        RECT 3527.625 3919.625 3527.905 3919.905 ;
        RECT 3528.245 3919.625 3528.525 3919.905 ;
        RECT 3528.865 3919.625 3529.145 3919.905 ;
        RECT 3529.485 3919.625 3529.765 3919.905 ;
        RECT 3527.625 3919.005 3527.905 3919.285 ;
        RECT 3528.245 3919.005 3528.525 3919.285 ;
        RECT 3528.865 3919.005 3529.145 3919.285 ;
        RECT 3529.485 3919.005 3529.765 3919.285 ;
        RECT 3527.625 3918.385 3527.905 3918.665 ;
        RECT 3528.245 3918.385 3528.525 3918.665 ;
        RECT 3528.865 3918.385 3529.145 3918.665 ;
        RECT 3529.485 3918.385 3529.765 3918.665 ;
        RECT 3527.625 3917.765 3527.905 3918.045 ;
        RECT 3528.245 3917.765 3528.525 3918.045 ;
        RECT 3528.865 3917.765 3529.145 3918.045 ;
        RECT 3529.485 3917.765 3529.765 3918.045 ;
        RECT 3527.625 3917.145 3527.905 3917.425 ;
        RECT 3528.245 3917.145 3528.525 3917.425 ;
        RECT 3528.865 3917.145 3529.145 3917.425 ;
        RECT 3529.485 3917.145 3529.765 3917.425 ;
        RECT 3527.625 3916.525 3527.905 3916.805 ;
        RECT 3528.245 3916.525 3528.525 3916.805 ;
        RECT 3528.865 3916.525 3529.145 3916.805 ;
        RECT 3529.485 3916.525 3529.765 3916.805 ;
        RECT 3527.625 3915.905 3527.905 3916.185 ;
        RECT 3528.245 3915.905 3528.525 3916.185 ;
        RECT 3528.865 3915.905 3529.145 3916.185 ;
        RECT 3529.485 3915.905 3529.765 3916.185 ;
        RECT 3527.625 3915.285 3527.905 3915.565 ;
        RECT 3528.245 3915.285 3528.525 3915.565 ;
        RECT 3528.865 3915.285 3529.145 3915.565 ;
        RECT 3529.485 3915.285 3529.765 3915.565 ;
        RECT 3527.625 3914.665 3527.905 3914.945 ;
        RECT 3528.245 3914.665 3528.525 3914.945 ;
        RECT 3528.865 3914.665 3529.145 3914.945 ;
        RECT 3529.485 3914.665 3529.765 3914.945 ;
        RECT 3527.625 3914.045 3527.905 3914.325 ;
        RECT 3528.245 3914.045 3528.525 3914.325 ;
        RECT 3528.865 3914.045 3529.145 3914.325 ;
        RECT 3529.485 3914.045 3529.765 3914.325 ;
        RECT 3527.625 3913.425 3527.905 3913.705 ;
        RECT 3528.245 3913.425 3528.525 3913.705 ;
        RECT 3528.865 3913.425 3529.145 3913.705 ;
        RECT 3529.485 3913.425 3529.765 3913.705 ;
        RECT 3527.625 3912.805 3527.905 3913.085 ;
        RECT 3528.245 3912.805 3528.525 3913.085 ;
        RECT 3528.865 3912.805 3529.145 3913.085 ;
        RECT 3529.485 3912.805 3529.765 3913.085 ;
        RECT 3527.625 3912.185 3527.905 3912.465 ;
        RECT 3528.245 3912.185 3528.525 3912.465 ;
        RECT 3528.865 3912.185 3529.145 3912.465 ;
        RECT 3529.485 3912.185 3529.765 3912.465 ;
        RECT 3527.625 3911.565 3527.905 3911.845 ;
        RECT 3528.245 3911.565 3528.525 3911.845 ;
        RECT 3528.865 3911.565 3529.145 3911.845 ;
        RECT 3529.485 3911.565 3529.765 3911.845 ;
        RECT 3527.625 3910.945 3527.905 3911.225 ;
        RECT 3528.245 3910.945 3528.525 3911.225 ;
        RECT 3528.865 3910.945 3529.145 3911.225 ;
        RECT 3529.485 3910.945 3529.765 3911.225 ;
        RECT 3527.625 3908.395 3527.905 3908.675 ;
        RECT 3528.245 3908.395 3528.525 3908.675 ;
        RECT 3528.865 3908.395 3529.145 3908.675 ;
        RECT 3529.485 3908.395 3529.765 3908.675 ;
        RECT 3527.625 3907.775 3527.905 3908.055 ;
        RECT 3528.245 3907.775 3528.525 3908.055 ;
        RECT 3528.865 3907.775 3529.145 3908.055 ;
        RECT 3529.485 3907.775 3529.765 3908.055 ;
        RECT 3527.625 3907.155 3527.905 3907.435 ;
        RECT 3528.245 3907.155 3528.525 3907.435 ;
        RECT 3528.865 3907.155 3529.145 3907.435 ;
        RECT 3529.485 3907.155 3529.765 3907.435 ;
        RECT 3527.625 3906.535 3527.905 3906.815 ;
        RECT 3528.245 3906.535 3528.525 3906.815 ;
        RECT 3528.865 3906.535 3529.145 3906.815 ;
        RECT 3529.485 3906.535 3529.765 3906.815 ;
        RECT 3527.625 3905.915 3527.905 3906.195 ;
        RECT 3528.245 3905.915 3528.525 3906.195 ;
        RECT 3528.865 3905.915 3529.145 3906.195 ;
        RECT 3529.485 3905.915 3529.765 3906.195 ;
        RECT 3527.625 3905.295 3527.905 3905.575 ;
        RECT 3528.245 3905.295 3528.525 3905.575 ;
        RECT 3528.865 3905.295 3529.145 3905.575 ;
        RECT 3529.485 3905.295 3529.765 3905.575 ;
        RECT 3527.625 3904.675 3527.905 3904.955 ;
        RECT 3528.245 3904.675 3528.525 3904.955 ;
        RECT 3528.865 3904.675 3529.145 3904.955 ;
        RECT 3529.485 3904.675 3529.765 3904.955 ;
        RECT 3527.625 3904.055 3527.905 3904.335 ;
        RECT 3528.245 3904.055 3528.525 3904.335 ;
        RECT 3528.865 3904.055 3529.145 3904.335 ;
        RECT 3529.485 3904.055 3529.765 3904.335 ;
        RECT 3527.625 3903.435 3527.905 3903.715 ;
        RECT 3528.245 3903.435 3528.525 3903.715 ;
        RECT 3528.865 3903.435 3529.145 3903.715 ;
        RECT 3529.485 3903.435 3529.765 3903.715 ;
        RECT 3527.625 3902.815 3527.905 3903.095 ;
        RECT 3528.245 3902.815 3528.525 3903.095 ;
        RECT 3528.865 3902.815 3529.145 3903.095 ;
        RECT 3529.485 3902.815 3529.765 3903.095 ;
        RECT 3527.625 3902.195 3527.905 3902.475 ;
        RECT 3528.245 3902.195 3528.525 3902.475 ;
        RECT 3528.865 3902.195 3529.145 3902.475 ;
        RECT 3529.485 3902.195 3529.765 3902.475 ;
        RECT 3527.625 3901.575 3527.905 3901.855 ;
        RECT 3528.245 3901.575 3528.525 3901.855 ;
        RECT 3528.865 3901.575 3529.145 3901.855 ;
        RECT 3529.485 3901.575 3529.765 3901.855 ;
        RECT 3527.625 3900.955 3527.905 3901.235 ;
        RECT 3528.245 3900.955 3528.525 3901.235 ;
        RECT 3528.865 3900.955 3529.145 3901.235 ;
        RECT 3529.485 3900.955 3529.765 3901.235 ;
        RECT 3527.625 3900.335 3527.905 3900.615 ;
        RECT 3528.245 3900.335 3528.525 3900.615 ;
        RECT 3528.865 3900.335 3529.145 3900.615 ;
        RECT 3529.485 3900.335 3529.765 3900.615 ;
        RECT 3527.625 3899.715 3527.905 3899.995 ;
        RECT 3528.245 3899.715 3528.525 3899.995 ;
        RECT 3528.865 3899.715 3529.145 3899.995 ;
        RECT 3529.485 3899.715 3529.765 3899.995 ;
        RECT 3527.625 3899.095 3527.905 3899.375 ;
        RECT 3528.245 3899.095 3528.525 3899.375 ;
        RECT 3528.865 3899.095 3529.145 3899.375 ;
        RECT 3529.485 3899.095 3529.765 3899.375 ;
        RECT 3527.625 3895.375 3527.905 3895.655 ;
        RECT 3528.245 3895.375 3528.525 3895.655 ;
        RECT 3528.865 3895.375 3529.145 3895.655 ;
        RECT 3529.485 3895.375 3529.765 3895.655 ;
        RECT 3527.625 3894.755 3527.905 3895.035 ;
        RECT 3528.245 3894.755 3528.525 3895.035 ;
        RECT 3528.865 3894.755 3529.145 3895.035 ;
        RECT 3529.485 3894.755 3529.765 3895.035 ;
        RECT 3527.625 3894.135 3527.905 3894.415 ;
        RECT 3528.245 3894.135 3528.525 3894.415 ;
        RECT 3528.865 3894.135 3529.145 3894.415 ;
        RECT 3529.485 3894.135 3529.765 3894.415 ;
        RECT 3527.625 3893.515 3527.905 3893.795 ;
        RECT 3528.245 3893.515 3528.525 3893.795 ;
        RECT 3528.865 3893.515 3529.145 3893.795 ;
        RECT 3529.485 3893.515 3529.765 3893.795 ;
        RECT 3527.625 3892.895 3527.905 3893.175 ;
        RECT 3528.245 3892.895 3528.525 3893.175 ;
        RECT 3528.865 3892.895 3529.145 3893.175 ;
        RECT 3529.485 3892.895 3529.765 3893.175 ;
        RECT 3527.625 3892.275 3527.905 3892.555 ;
        RECT 3528.245 3892.275 3528.525 3892.555 ;
        RECT 3528.865 3892.275 3529.145 3892.555 ;
        RECT 3529.485 3892.275 3529.765 3892.555 ;
        RECT 3527.625 3891.655 3527.905 3891.935 ;
        RECT 3528.245 3891.655 3528.525 3891.935 ;
        RECT 3528.865 3891.655 3529.145 3891.935 ;
        RECT 3529.485 3891.655 3529.765 3891.935 ;
        RECT 3527.625 3891.035 3527.905 3891.315 ;
        RECT 3528.245 3891.035 3528.525 3891.315 ;
        RECT 3528.865 3891.035 3529.145 3891.315 ;
        RECT 3529.485 3891.035 3529.765 3891.315 ;
        RECT 3527.625 3890.415 3527.905 3890.695 ;
        RECT 3528.245 3890.415 3528.525 3890.695 ;
        RECT 3528.865 3890.415 3529.145 3890.695 ;
        RECT 3529.485 3890.415 3529.765 3890.695 ;
        RECT 3527.625 3889.795 3527.905 3890.075 ;
        RECT 3528.245 3889.795 3528.525 3890.075 ;
        RECT 3528.865 3889.795 3529.145 3890.075 ;
        RECT 3529.485 3889.795 3529.765 3890.075 ;
        RECT 3527.625 3889.175 3527.905 3889.455 ;
        RECT 3528.245 3889.175 3528.525 3889.455 ;
        RECT 3528.865 3889.175 3529.145 3889.455 ;
        RECT 3529.485 3889.175 3529.765 3889.455 ;
        RECT 3527.625 3888.555 3527.905 3888.835 ;
        RECT 3528.245 3888.555 3528.525 3888.835 ;
        RECT 3528.865 3888.555 3529.145 3888.835 ;
        RECT 3529.485 3888.555 3529.765 3888.835 ;
        RECT 3527.625 3887.935 3527.905 3888.215 ;
        RECT 3528.245 3887.935 3528.525 3888.215 ;
        RECT 3528.865 3887.935 3529.145 3888.215 ;
        RECT 3529.485 3887.935 3529.765 3888.215 ;
        RECT 3527.625 3887.315 3527.905 3887.595 ;
        RECT 3528.245 3887.315 3528.525 3887.595 ;
        RECT 3528.865 3887.315 3529.145 3887.595 ;
        RECT 3529.485 3887.315 3529.765 3887.595 ;
        RECT 3527.625 3886.695 3527.905 3886.975 ;
        RECT 3528.245 3886.695 3528.525 3886.975 ;
        RECT 3528.865 3886.695 3529.145 3886.975 ;
        RECT 3529.485 3886.695 3529.765 3886.975 ;
        RECT 3527.625 2453.155 3527.905 2453.435 ;
        RECT 3528.245 2453.155 3528.525 2453.435 ;
        RECT 3528.865 2453.155 3529.145 2453.435 ;
        RECT 3529.485 2453.155 3529.765 2453.435 ;
        RECT 3527.625 2452.535 3527.905 2452.815 ;
        RECT 3528.245 2452.535 3528.525 2452.815 ;
        RECT 3528.865 2452.535 3529.145 2452.815 ;
        RECT 3529.485 2452.535 3529.765 2452.815 ;
        RECT 3527.625 2451.915 3527.905 2452.195 ;
        RECT 3528.245 2451.915 3528.525 2452.195 ;
        RECT 3528.865 2451.915 3529.145 2452.195 ;
        RECT 3529.485 2451.915 3529.765 2452.195 ;
        RECT 3527.625 2451.295 3527.905 2451.575 ;
        RECT 3528.245 2451.295 3528.525 2451.575 ;
        RECT 3528.865 2451.295 3529.145 2451.575 ;
        RECT 3529.485 2451.295 3529.765 2451.575 ;
        RECT 3527.625 2450.675 3527.905 2450.955 ;
        RECT 3528.245 2450.675 3528.525 2450.955 ;
        RECT 3528.865 2450.675 3529.145 2450.955 ;
        RECT 3529.485 2450.675 3529.765 2450.955 ;
        RECT 3527.625 2450.055 3527.905 2450.335 ;
        RECT 3528.245 2450.055 3528.525 2450.335 ;
        RECT 3528.865 2450.055 3529.145 2450.335 ;
        RECT 3529.485 2450.055 3529.765 2450.335 ;
        RECT 3527.625 2449.435 3527.905 2449.715 ;
        RECT 3528.245 2449.435 3528.525 2449.715 ;
        RECT 3528.865 2449.435 3529.145 2449.715 ;
        RECT 3529.485 2449.435 3529.765 2449.715 ;
        RECT 3527.625 2448.815 3527.905 2449.095 ;
        RECT 3528.245 2448.815 3528.525 2449.095 ;
        RECT 3528.865 2448.815 3529.145 2449.095 ;
        RECT 3529.485 2448.815 3529.765 2449.095 ;
        RECT 3527.625 2448.195 3527.905 2448.475 ;
        RECT 3528.245 2448.195 3528.525 2448.475 ;
        RECT 3528.865 2448.195 3529.145 2448.475 ;
        RECT 3529.485 2448.195 3529.765 2448.475 ;
        RECT 3527.625 2447.575 3527.905 2447.855 ;
        RECT 3528.245 2447.575 3528.525 2447.855 ;
        RECT 3528.865 2447.575 3529.145 2447.855 ;
        RECT 3529.485 2447.575 3529.765 2447.855 ;
        RECT 3527.625 2446.955 3527.905 2447.235 ;
        RECT 3528.245 2446.955 3528.525 2447.235 ;
        RECT 3528.865 2446.955 3529.145 2447.235 ;
        RECT 3529.485 2446.955 3529.765 2447.235 ;
        RECT 3527.625 2446.335 3527.905 2446.615 ;
        RECT 3528.245 2446.335 3528.525 2446.615 ;
        RECT 3528.865 2446.335 3529.145 2446.615 ;
        RECT 3529.485 2446.335 3529.765 2446.615 ;
        RECT 3527.625 2445.715 3527.905 2445.995 ;
        RECT 3528.245 2445.715 3528.525 2445.995 ;
        RECT 3528.865 2445.715 3529.145 2445.995 ;
        RECT 3529.485 2445.715 3529.765 2445.995 ;
        RECT 3527.625 2445.095 3527.905 2445.375 ;
        RECT 3528.245 2445.095 3528.525 2445.375 ;
        RECT 3528.865 2445.095 3529.145 2445.375 ;
        RECT 3529.485 2445.095 3529.765 2445.375 ;
        RECT 3527.625 2444.475 3527.905 2444.755 ;
        RECT 3528.245 2444.475 3528.525 2444.755 ;
        RECT 3528.865 2444.475 3529.145 2444.755 ;
        RECT 3529.485 2444.475 3529.765 2444.755 ;
        RECT 3527.625 2440.625 3527.905 2440.905 ;
        RECT 3528.245 2440.625 3528.525 2440.905 ;
        RECT 3528.865 2440.625 3529.145 2440.905 ;
        RECT 3529.485 2440.625 3529.765 2440.905 ;
        RECT 3527.625 2440.005 3527.905 2440.285 ;
        RECT 3528.245 2440.005 3528.525 2440.285 ;
        RECT 3528.865 2440.005 3529.145 2440.285 ;
        RECT 3529.485 2440.005 3529.765 2440.285 ;
        RECT 3527.625 2439.385 3527.905 2439.665 ;
        RECT 3528.245 2439.385 3528.525 2439.665 ;
        RECT 3528.865 2439.385 3529.145 2439.665 ;
        RECT 3529.485 2439.385 3529.765 2439.665 ;
        RECT 3527.625 2438.765 3527.905 2439.045 ;
        RECT 3528.245 2438.765 3528.525 2439.045 ;
        RECT 3528.865 2438.765 3529.145 2439.045 ;
        RECT 3529.485 2438.765 3529.765 2439.045 ;
        RECT 3527.625 2438.145 3527.905 2438.425 ;
        RECT 3528.245 2438.145 3528.525 2438.425 ;
        RECT 3528.865 2438.145 3529.145 2438.425 ;
        RECT 3529.485 2438.145 3529.765 2438.425 ;
        RECT 3527.625 2437.525 3527.905 2437.805 ;
        RECT 3528.245 2437.525 3528.525 2437.805 ;
        RECT 3528.865 2437.525 3529.145 2437.805 ;
        RECT 3529.485 2437.525 3529.765 2437.805 ;
        RECT 3527.625 2436.905 3527.905 2437.185 ;
        RECT 3528.245 2436.905 3528.525 2437.185 ;
        RECT 3528.865 2436.905 3529.145 2437.185 ;
        RECT 3529.485 2436.905 3529.765 2437.185 ;
        RECT 3527.625 2436.285 3527.905 2436.565 ;
        RECT 3528.245 2436.285 3528.525 2436.565 ;
        RECT 3528.865 2436.285 3529.145 2436.565 ;
        RECT 3529.485 2436.285 3529.765 2436.565 ;
        RECT 3527.625 2435.665 3527.905 2435.945 ;
        RECT 3528.245 2435.665 3528.525 2435.945 ;
        RECT 3528.865 2435.665 3529.145 2435.945 ;
        RECT 3529.485 2435.665 3529.765 2435.945 ;
        RECT 3527.625 2435.045 3527.905 2435.325 ;
        RECT 3528.245 2435.045 3528.525 2435.325 ;
        RECT 3528.865 2435.045 3529.145 2435.325 ;
        RECT 3529.485 2435.045 3529.765 2435.325 ;
        RECT 3527.625 2434.425 3527.905 2434.705 ;
        RECT 3528.245 2434.425 3528.525 2434.705 ;
        RECT 3528.865 2434.425 3529.145 2434.705 ;
        RECT 3529.485 2434.425 3529.765 2434.705 ;
        RECT 3527.625 2433.805 3527.905 2434.085 ;
        RECT 3528.245 2433.805 3528.525 2434.085 ;
        RECT 3528.865 2433.805 3529.145 2434.085 ;
        RECT 3529.485 2433.805 3529.765 2434.085 ;
        RECT 3527.625 2433.185 3527.905 2433.465 ;
        RECT 3528.245 2433.185 3528.525 2433.465 ;
        RECT 3528.865 2433.185 3529.145 2433.465 ;
        RECT 3529.485 2433.185 3529.765 2433.465 ;
        RECT 3527.625 2432.565 3527.905 2432.845 ;
        RECT 3528.245 2432.565 3528.525 2432.845 ;
        RECT 3528.865 2432.565 3529.145 2432.845 ;
        RECT 3529.485 2432.565 3529.765 2432.845 ;
        RECT 3527.625 2431.945 3527.905 2432.225 ;
        RECT 3528.245 2431.945 3528.525 2432.225 ;
        RECT 3528.865 2431.945 3529.145 2432.225 ;
        RECT 3529.485 2431.945 3529.765 2432.225 ;
        RECT 3527.625 2431.325 3527.905 2431.605 ;
        RECT 3528.245 2431.325 3528.525 2431.605 ;
        RECT 3528.865 2431.325 3529.145 2431.605 ;
        RECT 3529.485 2431.325 3529.765 2431.605 ;
        RECT 3527.625 2428.775 3527.905 2429.055 ;
        RECT 3528.245 2428.775 3528.525 2429.055 ;
        RECT 3528.865 2428.775 3529.145 2429.055 ;
        RECT 3529.485 2428.775 3529.765 2429.055 ;
        RECT 3527.625 2428.155 3527.905 2428.435 ;
        RECT 3528.245 2428.155 3528.525 2428.435 ;
        RECT 3528.865 2428.155 3529.145 2428.435 ;
        RECT 3529.485 2428.155 3529.765 2428.435 ;
        RECT 3527.625 2427.535 3527.905 2427.815 ;
        RECT 3528.245 2427.535 3528.525 2427.815 ;
        RECT 3528.865 2427.535 3529.145 2427.815 ;
        RECT 3529.485 2427.535 3529.765 2427.815 ;
        RECT 3527.625 2426.915 3527.905 2427.195 ;
        RECT 3528.245 2426.915 3528.525 2427.195 ;
        RECT 3528.865 2426.915 3529.145 2427.195 ;
        RECT 3529.485 2426.915 3529.765 2427.195 ;
        RECT 3527.625 2426.295 3527.905 2426.575 ;
        RECT 3528.245 2426.295 3528.525 2426.575 ;
        RECT 3528.865 2426.295 3529.145 2426.575 ;
        RECT 3529.485 2426.295 3529.765 2426.575 ;
        RECT 3527.625 2425.675 3527.905 2425.955 ;
        RECT 3528.245 2425.675 3528.525 2425.955 ;
        RECT 3528.865 2425.675 3529.145 2425.955 ;
        RECT 3529.485 2425.675 3529.765 2425.955 ;
        RECT 3527.625 2425.055 3527.905 2425.335 ;
        RECT 3528.245 2425.055 3528.525 2425.335 ;
        RECT 3528.865 2425.055 3529.145 2425.335 ;
        RECT 3529.485 2425.055 3529.765 2425.335 ;
        RECT 3527.625 2424.435 3527.905 2424.715 ;
        RECT 3528.245 2424.435 3528.525 2424.715 ;
        RECT 3528.865 2424.435 3529.145 2424.715 ;
        RECT 3529.485 2424.435 3529.765 2424.715 ;
        RECT 3527.625 2423.815 3527.905 2424.095 ;
        RECT 3528.245 2423.815 3528.525 2424.095 ;
        RECT 3528.865 2423.815 3529.145 2424.095 ;
        RECT 3529.485 2423.815 3529.765 2424.095 ;
        RECT 3527.625 2423.195 3527.905 2423.475 ;
        RECT 3528.245 2423.195 3528.525 2423.475 ;
        RECT 3528.865 2423.195 3529.145 2423.475 ;
        RECT 3529.485 2423.195 3529.765 2423.475 ;
        RECT 3527.625 2422.575 3527.905 2422.855 ;
        RECT 3528.245 2422.575 3528.525 2422.855 ;
        RECT 3528.865 2422.575 3529.145 2422.855 ;
        RECT 3529.485 2422.575 3529.765 2422.855 ;
        RECT 3527.625 2421.955 3527.905 2422.235 ;
        RECT 3528.245 2421.955 3528.525 2422.235 ;
        RECT 3528.865 2421.955 3529.145 2422.235 ;
        RECT 3529.485 2421.955 3529.765 2422.235 ;
        RECT 3527.625 2421.335 3527.905 2421.615 ;
        RECT 3528.245 2421.335 3528.525 2421.615 ;
        RECT 3528.865 2421.335 3529.145 2421.615 ;
        RECT 3529.485 2421.335 3529.765 2421.615 ;
        RECT 3527.625 2420.715 3527.905 2420.995 ;
        RECT 3528.245 2420.715 3528.525 2420.995 ;
        RECT 3528.865 2420.715 3529.145 2420.995 ;
        RECT 3529.485 2420.715 3529.765 2420.995 ;
        RECT 3527.625 2420.095 3527.905 2420.375 ;
        RECT 3528.245 2420.095 3528.525 2420.375 ;
        RECT 3528.865 2420.095 3529.145 2420.375 ;
        RECT 3529.485 2420.095 3529.765 2420.375 ;
        RECT 3527.625 2419.475 3527.905 2419.755 ;
        RECT 3528.245 2419.475 3528.525 2419.755 ;
        RECT 3528.865 2419.475 3529.145 2419.755 ;
        RECT 3529.485 2419.475 3529.765 2419.755 ;
        RECT 3527.625 2415.245 3527.905 2415.525 ;
        RECT 3528.245 2415.245 3528.525 2415.525 ;
        RECT 3528.865 2415.245 3529.145 2415.525 ;
        RECT 3529.485 2415.245 3529.765 2415.525 ;
        RECT 3527.625 2414.625 3527.905 2414.905 ;
        RECT 3528.245 2414.625 3528.525 2414.905 ;
        RECT 3528.865 2414.625 3529.145 2414.905 ;
        RECT 3529.485 2414.625 3529.765 2414.905 ;
        RECT 3527.625 2414.005 3527.905 2414.285 ;
        RECT 3528.245 2414.005 3528.525 2414.285 ;
        RECT 3528.865 2414.005 3529.145 2414.285 ;
        RECT 3529.485 2414.005 3529.765 2414.285 ;
        RECT 3527.625 2413.385 3527.905 2413.665 ;
        RECT 3528.245 2413.385 3528.525 2413.665 ;
        RECT 3528.865 2413.385 3529.145 2413.665 ;
        RECT 3529.485 2413.385 3529.765 2413.665 ;
        RECT 3527.625 2412.765 3527.905 2413.045 ;
        RECT 3528.245 2412.765 3528.525 2413.045 ;
        RECT 3528.865 2412.765 3529.145 2413.045 ;
        RECT 3529.485 2412.765 3529.765 2413.045 ;
        RECT 3527.625 2412.145 3527.905 2412.425 ;
        RECT 3528.245 2412.145 3528.525 2412.425 ;
        RECT 3528.865 2412.145 3529.145 2412.425 ;
        RECT 3529.485 2412.145 3529.765 2412.425 ;
        RECT 3527.625 2411.525 3527.905 2411.805 ;
        RECT 3528.245 2411.525 3528.525 2411.805 ;
        RECT 3528.865 2411.525 3529.145 2411.805 ;
        RECT 3529.485 2411.525 3529.765 2411.805 ;
        RECT 3527.625 2410.905 3527.905 2411.185 ;
        RECT 3528.245 2410.905 3528.525 2411.185 ;
        RECT 3528.865 2410.905 3529.145 2411.185 ;
        RECT 3529.485 2410.905 3529.765 2411.185 ;
        RECT 3527.625 2410.285 3527.905 2410.565 ;
        RECT 3528.245 2410.285 3528.525 2410.565 ;
        RECT 3528.865 2410.285 3529.145 2410.565 ;
        RECT 3529.485 2410.285 3529.765 2410.565 ;
        RECT 3527.625 2409.665 3527.905 2409.945 ;
        RECT 3528.245 2409.665 3528.525 2409.945 ;
        RECT 3528.865 2409.665 3529.145 2409.945 ;
        RECT 3529.485 2409.665 3529.765 2409.945 ;
        RECT 3527.625 2409.045 3527.905 2409.325 ;
        RECT 3528.245 2409.045 3528.525 2409.325 ;
        RECT 3528.865 2409.045 3529.145 2409.325 ;
        RECT 3529.485 2409.045 3529.765 2409.325 ;
        RECT 3527.625 2408.425 3527.905 2408.705 ;
        RECT 3528.245 2408.425 3528.525 2408.705 ;
        RECT 3528.865 2408.425 3529.145 2408.705 ;
        RECT 3529.485 2408.425 3529.765 2408.705 ;
        RECT 3527.625 2407.805 3527.905 2408.085 ;
        RECT 3528.245 2407.805 3528.525 2408.085 ;
        RECT 3528.865 2407.805 3529.145 2408.085 ;
        RECT 3529.485 2407.805 3529.765 2408.085 ;
        RECT 3527.625 2407.185 3527.905 2407.465 ;
        RECT 3528.245 2407.185 3528.525 2407.465 ;
        RECT 3528.865 2407.185 3529.145 2407.465 ;
        RECT 3529.485 2407.185 3529.765 2407.465 ;
        RECT 3527.625 2406.565 3527.905 2406.845 ;
        RECT 3528.245 2406.565 3528.525 2406.845 ;
        RECT 3528.865 2406.565 3529.145 2406.845 ;
        RECT 3529.485 2406.565 3529.765 2406.845 ;
        RECT 3527.625 2405.945 3527.905 2406.225 ;
        RECT 3528.245 2405.945 3528.525 2406.225 ;
        RECT 3528.865 2405.945 3529.145 2406.225 ;
        RECT 3529.485 2405.945 3529.765 2406.225 ;
        RECT 3527.625 2403.395 3527.905 2403.675 ;
        RECT 3528.245 2403.395 3528.525 2403.675 ;
        RECT 3528.865 2403.395 3529.145 2403.675 ;
        RECT 3529.485 2403.395 3529.765 2403.675 ;
        RECT 3527.625 2402.775 3527.905 2403.055 ;
        RECT 3528.245 2402.775 3528.525 2403.055 ;
        RECT 3528.865 2402.775 3529.145 2403.055 ;
        RECT 3529.485 2402.775 3529.765 2403.055 ;
        RECT 3527.625 2402.155 3527.905 2402.435 ;
        RECT 3528.245 2402.155 3528.525 2402.435 ;
        RECT 3528.865 2402.155 3529.145 2402.435 ;
        RECT 3529.485 2402.155 3529.765 2402.435 ;
        RECT 3527.625 2401.535 3527.905 2401.815 ;
        RECT 3528.245 2401.535 3528.525 2401.815 ;
        RECT 3528.865 2401.535 3529.145 2401.815 ;
        RECT 3529.485 2401.535 3529.765 2401.815 ;
        RECT 3527.625 2400.915 3527.905 2401.195 ;
        RECT 3528.245 2400.915 3528.525 2401.195 ;
        RECT 3528.865 2400.915 3529.145 2401.195 ;
        RECT 3529.485 2400.915 3529.765 2401.195 ;
        RECT 3527.625 2400.295 3527.905 2400.575 ;
        RECT 3528.245 2400.295 3528.525 2400.575 ;
        RECT 3528.865 2400.295 3529.145 2400.575 ;
        RECT 3529.485 2400.295 3529.765 2400.575 ;
        RECT 3527.625 2399.675 3527.905 2399.955 ;
        RECT 3528.245 2399.675 3528.525 2399.955 ;
        RECT 3528.865 2399.675 3529.145 2399.955 ;
        RECT 3529.485 2399.675 3529.765 2399.955 ;
        RECT 3527.625 2399.055 3527.905 2399.335 ;
        RECT 3528.245 2399.055 3528.525 2399.335 ;
        RECT 3528.865 2399.055 3529.145 2399.335 ;
        RECT 3529.485 2399.055 3529.765 2399.335 ;
        RECT 3527.625 2398.435 3527.905 2398.715 ;
        RECT 3528.245 2398.435 3528.525 2398.715 ;
        RECT 3528.865 2398.435 3529.145 2398.715 ;
        RECT 3529.485 2398.435 3529.765 2398.715 ;
        RECT 3527.625 2397.815 3527.905 2398.095 ;
        RECT 3528.245 2397.815 3528.525 2398.095 ;
        RECT 3528.865 2397.815 3529.145 2398.095 ;
        RECT 3529.485 2397.815 3529.765 2398.095 ;
        RECT 3527.625 2397.195 3527.905 2397.475 ;
        RECT 3528.245 2397.195 3528.525 2397.475 ;
        RECT 3528.865 2397.195 3529.145 2397.475 ;
        RECT 3529.485 2397.195 3529.765 2397.475 ;
        RECT 3527.625 2396.575 3527.905 2396.855 ;
        RECT 3528.245 2396.575 3528.525 2396.855 ;
        RECT 3528.865 2396.575 3529.145 2396.855 ;
        RECT 3529.485 2396.575 3529.765 2396.855 ;
        RECT 3527.625 2395.955 3527.905 2396.235 ;
        RECT 3528.245 2395.955 3528.525 2396.235 ;
        RECT 3528.865 2395.955 3529.145 2396.235 ;
        RECT 3529.485 2395.955 3529.765 2396.235 ;
        RECT 3527.625 2395.335 3527.905 2395.615 ;
        RECT 3528.245 2395.335 3528.525 2395.615 ;
        RECT 3528.865 2395.335 3529.145 2395.615 ;
        RECT 3529.485 2395.335 3529.765 2395.615 ;
        RECT 3527.625 2394.715 3527.905 2394.995 ;
        RECT 3528.245 2394.715 3528.525 2394.995 ;
        RECT 3528.865 2394.715 3529.145 2394.995 ;
        RECT 3529.485 2394.715 3529.765 2394.995 ;
        RECT 3527.625 2394.095 3527.905 2394.375 ;
        RECT 3528.245 2394.095 3528.525 2394.375 ;
        RECT 3528.865 2394.095 3529.145 2394.375 ;
        RECT 3529.485 2394.095 3529.765 2394.375 ;
        RECT 3527.625 2390.375 3527.905 2390.655 ;
        RECT 3528.245 2390.375 3528.525 2390.655 ;
        RECT 3528.865 2390.375 3529.145 2390.655 ;
        RECT 3529.485 2390.375 3529.765 2390.655 ;
        RECT 3527.625 2389.755 3527.905 2390.035 ;
        RECT 3528.245 2389.755 3528.525 2390.035 ;
        RECT 3528.865 2389.755 3529.145 2390.035 ;
        RECT 3529.485 2389.755 3529.765 2390.035 ;
        RECT 3527.625 2389.135 3527.905 2389.415 ;
        RECT 3528.245 2389.135 3528.525 2389.415 ;
        RECT 3528.865 2389.135 3529.145 2389.415 ;
        RECT 3529.485 2389.135 3529.765 2389.415 ;
        RECT 3527.625 2388.515 3527.905 2388.795 ;
        RECT 3528.245 2388.515 3528.525 2388.795 ;
        RECT 3528.865 2388.515 3529.145 2388.795 ;
        RECT 3529.485 2388.515 3529.765 2388.795 ;
        RECT 3527.625 2387.895 3527.905 2388.175 ;
        RECT 3528.245 2387.895 3528.525 2388.175 ;
        RECT 3528.865 2387.895 3529.145 2388.175 ;
        RECT 3529.485 2387.895 3529.765 2388.175 ;
        RECT 3527.625 2387.275 3527.905 2387.555 ;
        RECT 3528.245 2387.275 3528.525 2387.555 ;
        RECT 3528.865 2387.275 3529.145 2387.555 ;
        RECT 3529.485 2387.275 3529.765 2387.555 ;
        RECT 3527.625 2386.655 3527.905 2386.935 ;
        RECT 3528.245 2386.655 3528.525 2386.935 ;
        RECT 3528.865 2386.655 3529.145 2386.935 ;
        RECT 3529.485 2386.655 3529.765 2386.935 ;
        RECT 3527.625 2386.035 3527.905 2386.315 ;
        RECT 3528.245 2386.035 3528.525 2386.315 ;
        RECT 3528.865 2386.035 3529.145 2386.315 ;
        RECT 3529.485 2386.035 3529.765 2386.315 ;
        RECT 3527.625 2385.415 3527.905 2385.695 ;
        RECT 3528.245 2385.415 3528.525 2385.695 ;
        RECT 3528.865 2385.415 3529.145 2385.695 ;
        RECT 3529.485 2385.415 3529.765 2385.695 ;
        RECT 3527.625 2384.795 3527.905 2385.075 ;
        RECT 3528.245 2384.795 3528.525 2385.075 ;
        RECT 3528.865 2384.795 3529.145 2385.075 ;
        RECT 3529.485 2384.795 3529.765 2385.075 ;
        RECT 3527.625 2384.175 3527.905 2384.455 ;
        RECT 3528.245 2384.175 3528.525 2384.455 ;
        RECT 3528.865 2384.175 3529.145 2384.455 ;
        RECT 3529.485 2384.175 3529.765 2384.455 ;
        RECT 3527.625 2383.555 3527.905 2383.835 ;
        RECT 3528.245 2383.555 3528.525 2383.835 ;
        RECT 3528.865 2383.555 3529.145 2383.835 ;
        RECT 3529.485 2383.555 3529.765 2383.835 ;
        RECT 3527.625 2382.935 3527.905 2383.215 ;
        RECT 3528.245 2382.935 3528.525 2383.215 ;
        RECT 3528.865 2382.935 3529.145 2383.215 ;
        RECT 3529.485 2382.935 3529.765 2383.215 ;
        RECT 3527.625 2382.315 3527.905 2382.595 ;
        RECT 3528.245 2382.315 3528.525 2382.595 ;
        RECT 3528.865 2382.315 3529.145 2382.595 ;
        RECT 3529.485 2382.315 3529.765 2382.595 ;
        RECT 3527.625 2381.695 3527.905 2381.975 ;
        RECT 3528.245 2381.695 3528.525 2381.975 ;
        RECT 3528.865 2381.695 3529.145 2381.975 ;
        RECT 3529.485 2381.695 3529.765 2381.975 ;
        RECT 350.235 2343.025 350.515 2343.305 ;
        RECT 350.855 2343.025 351.135 2343.305 ;
        RECT 351.475 2343.025 351.755 2343.305 ;
        RECT 352.095 2343.025 352.375 2343.305 ;
        RECT 350.235 2342.405 350.515 2342.685 ;
        RECT 350.855 2342.405 351.135 2342.685 ;
        RECT 351.475 2342.405 351.755 2342.685 ;
        RECT 352.095 2342.405 352.375 2342.685 ;
        RECT 350.235 2341.785 350.515 2342.065 ;
        RECT 350.855 2341.785 351.135 2342.065 ;
        RECT 351.475 2341.785 351.755 2342.065 ;
        RECT 352.095 2341.785 352.375 2342.065 ;
        RECT 350.235 2341.165 350.515 2341.445 ;
        RECT 350.855 2341.165 351.135 2341.445 ;
        RECT 351.475 2341.165 351.755 2341.445 ;
        RECT 352.095 2341.165 352.375 2341.445 ;
        RECT 350.235 2340.545 350.515 2340.825 ;
        RECT 350.855 2340.545 351.135 2340.825 ;
        RECT 351.475 2340.545 351.755 2340.825 ;
        RECT 352.095 2340.545 352.375 2340.825 ;
        RECT 350.235 2339.925 350.515 2340.205 ;
        RECT 350.855 2339.925 351.135 2340.205 ;
        RECT 351.475 2339.925 351.755 2340.205 ;
        RECT 352.095 2339.925 352.375 2340.205 ;
        RECT 350.235 2339.305 350.515 2339.585 ;
        RECT 350.855 2339.305 351.135 2339.585 ;
        RECT 351.475 2339.305 351.755 2339.585 ;
        RECT 352.095 2339.305 352.375 2339.585 ;
        RECT 350.235 2338.685 350.515 2338.965 ;
        RECT 350.855 2338.685 351.135 2338.965 ;
        RECT 351.475 2338.685 351.755 2338.965 ;
        RECT 352.095 2338.685 352.375 2338.965 ;
        RECT 350.235 2338.065 350.515 2338.345 ;
        RECT 350.855 2338.065 351.135 2338.345 ;
        RECT 351.475 2338.065 351.755 2338.345 ;
        RECT 352.095 2338.065 352.375 2338.345 ;
        RECT 350.235 2337.445 350.515 2337.725 ;
        RECT 350.855 2337.445 351.135 2337.725 ;
        RECT 351.475 2337.445 351.755 2337.725 ;
        RECT 352.095 2337.445 352.375 2337.725 ;
        RECT 350.235 2336.825 350.515 2337.105 ;
        RECT 350.855 2336.825 351.135 2337.105 ;
        RECT 351.475 2336.825 351.755 2337.105 ;
        RECT 352.095 2336.825 352.375 2337.105 ;
        RECT 350.235 2336.205 350.515 2336.485 ;
        RECT 350.855 2336.205 351.135 2336.485 ;
        RECT 351.475 2336.205 351.755 2336.485 ;
        RECT 352.095 2336.205 352.375 2336.485 ;
        RECT 350.235 2335.585 350.515 2335.865 ;
        RECT 350.855 2335.585 351.135 2335.865 ;
        RECT 351.475 2335.585 351.755 2335.865 ;
        RECT 352.095 2335.585 352.375 2335.865 ;
        RECT 350.235 2334.965 350.515 2335.245 ;
        RECT 350.855 2334.965 351.135 2335.245 ;
        RECT 351.475 2334.965 351.755 2335.245 ;
        RECT 352.095 2334.965 352.375 2335.245 ;
        RECT 350.235 2334.345 350.515 2334.625 ;
        RECT 350.855 2334.345 351.135 2334.625 ;
        RECT 351.475 2334.345 351.755 2334.625 ;
        RECT 352.095 2334.345 352.375 2334.625 ;
        RECT 350.235 2330.625 350.515 2330.905 ;
        RECT 350.855 2330.625 351.135 2330.905 ;
        RECT 351.475 2330.625 351.755 2330.905 ;
        RECT 352.095 2330.625 352.375 2330.905 ;
        RECT 350.235 2330.005 350.515 2330.285 ;
        RECT 350.855 2330.005 351.135 2330.285 ;
        RECT 351.475 2330.005 351.755 2330.285 ;
        RECT 352.095 2330.005 352.375 2330.285 ;
        RECT 350.235 2329.385 350.515 2329.665 ;
        RECT 350.855 2329.385 351.135 2329.665 ;
        RECT 351.475 2329.385 351.755 2329.665 ;
        RECT 352.095 2329.385 352.375 2329.665 ;
        RECT 350.235 2328.765 350.515 2329.045 ;
        RECT 350.855 2328.765 351.135 2329.045 ;
        RECT 351.475 2328.765 351.755 2329.045 ;
        RECT 352.095 2328.765 352.375 2329.045 ;
        RECT 350.235 2328.145 350.515 2328.425 ;
        RECT 350.855 2328.145 351.135 2328.425 ;
        RECT 351.475 2328.145 351.755 2328.425 ;
        RECT 352.095 2328.145 352.375 2328.425 ;
        RECT 350.235 2327.525 350.515 2327.805 ;
        RECT 350.855 2327.525 351.135 2327.805 ;
        RECT 351.475 2327.525 351.755 2327.805 ;
        RECT 352.095 2327.525 352.375 2327.805 ;
        RECT 350.235 2326.905 350.515 2327.185 ;
        RECT 350.855 2326.905 351.135 2327.185 ;
        RECT 351.475 2326.905 351.755 2327.185 ;
        RECT 352.095 2326.905 352.375 2327.185 ;
        RECT 350.235 2326.285 350.515 2326.565 ;
        RECT 350.855 2326.285 351.135 2326.565 ;
        RECT 351.475 2326.285 351.755 2326.565 ;
        RECT 352.095 2326.285 352.375 2326.565 ;
        RECT 350.235 2325.665 350.515 2325.945 ;
        RECT 350.855 2325.665 351.135 2325.945 ;
        RECT 351.475 2325.665 351.755 2325.945 ;
        RECT 352.095 2325.665 352.375 2325.945 ;
        RECT 350.235 2325.045 350.515 2325.325 ;
        RECT 350.855 2325.045 351.135 2325.325 ;
        RECT 351.475 2325.045 351.755 2325.325 ;
        RECT 352.095 2325.045 352.375 2325.325 ;
        RECT 350.235 2324.425 350.515 2324.705 ;
        RECT 350.855 2324.425 351.135 2324.705 ;
        RECT 351.475 2324.425 351.755 2324.705 ;
        RECT 352.095 2324.425 352.375 2324.705 ;
        RECT 350.235 2323.805 350.515 2324.085 ;
        RECT 350.855 2323.805 351.135 2324.085 ;
        RECT 351.475 2323.805 351.755 2324.085 ;
        RECT 352.095 2323.805 352.375 2324.085 ;
        RECT 350.235 2323.185 350.515 2323.465 ;
        RECT 350.855 2323.185 351.135 2323.465 ;
        RECT 351.475 2323.185 351.755 2323.465 ;
        RECT 352.095 2323.185 352.375 2323.465 ;
        RECT 350.235 2322.565 350.515 2322.845 ;
        RECT 350.855 2322.565 351.135 2322.845 ;
        RECT 351.475 2322.565 351.755 2322.845 ;
        RECT 352.095 2322.565 352.375 2322.845 ;
        RECT 350.235 2321.945 350.515 2322.225 ;
        RECT 350.855 2321.945 351.135 2322.225 ;
        RECT 351.475 2321.945 351.755 2322.225 ;
        RECT 352.095 2321.945 352.375 2322.225 ;
        RECT 350.235 2321.325 350.515 2321.605 ;
        RECT 350.855 2321.325 351.135 2321.605 ;
        RECT 351.475 2321.325 351.755 2321.605 ;
        RECT 352.095 2321.325 352.375 2321.605 ;
        RECT 350.235 2318.775 350.515 2319.055 ;
        RECT 350.855 2318.775 351.135 2319.055 ;
        RECT 351.475 2318.775 351.755 2319.055 ;
        RECT 352.095 2318.775 352.375 2319.055 ;
        RECT 350.235 2318.155 350.515 2318.435 ;
        RECT 350.855 2318.155 351.135 2318.435 ;
        RECT 351.475 2318.155 351.755 2318.435 ;
        RECT 352.095 2318.155 352.375 2318.435 ;
        RECT 350.235 2317.535 350.515 2317.815 ;
        RECT 350.855 2317.535 351.135 2317.815 ;
        RECT 351.475 2317.535 351.755 2317.815 ;
        RECT 352.095 2317.535 352.375 2317.815 ;
        RECT 350.235 2316.915 350.515 2317.195 ;
        RECT 350.855 2316.915 351.135 2317.195 ;
        RECT 351.475 2316.915 351.755 2317.195 ;
        RECT 352.095 2316.915 352.375 2317.195 ;
        RECT 350.235 2316.295 350.515 2316.575 ;
        RECT 350.855 2316.295 351.135 2316.575 ;
        RECT 351.475 2316.295 351.755 2316.575 ;
        RECT 352.095 2316.295 352.375 2316.575 ;
        RECT 350.235 2315.675 350.515 2315.955 ;
        RECT 350.855 2315.675 351.135 2315.955 ;
        RECT 351.475 2315.675 351.755 2315.955 ;
        RECT 352.095 2315.675 352.375 2315.955 ;
        RECT 350.235 2315.055 350.515 2315.335 ;
        RECT 350.855 2315.055 351.135 2315.335 ;
        RECT 351.475 2315.055 351.755 2315.335 ;
        RECT 352.095 2315.055 352.375 2315.335 ;
        RECT 350.235 2314.435 350.515 2314.715 ;
        RECT 350.855 2314.435 351.135 2314.715 ;
        RECT 351.475 2314.435 351.755 2314.715 ;
        RECT 352.095 2314.435 352.375 2314.715 ;
        RECT 350.235 2313.815 350.515 2314.095 ;
        RECT 350.855 2313.815 351.135 2314.095 ;
        RECT 351.475 2313.815 351.755 2314.095 ;
        RECT 352.095 2313.815 352.375 2314.095 ;
        RECT 350.235 2313.195 350.515 2313.475 ;
        RECT 350.855 2313.195 351.135 2313.475 ;
        RECT 351.475 2313.195 351.755 2313.475 ;
        RECT 352.095 2313.195 352.375 2313.475 ;
        RECT 350.235 2312.575 350.515 2312.855 ;
        RECT 350.855 2312.575 351.135 2312.855 ;
        RECT 351.475 2312.575 351.755 2312.855 ;
        RECT 352.095 2312.575 352.375 2312.855 ;
        RECT 350.235 2311.955 350.515 2312.235 ;
        RECT 350.855 2311.955 351.135 2312.235 ;
        RECT 351.475 2311.955 351.755 2312.235 ;
        RECT 352.095 2311.955 352.375 2312.235 ;
        RECT 350.235 2311.335 350.515 2311.615 ;
        RECT 350.855 2311.335 351.135 2311.615 ;
        RECT 351.475 2311.335 351.755 2311.615 ;
        RECT 352.095 2311.335 352.375 2311.615 ;
        RECT 350.235 2310.715 350.515 2310.995 ;
        RECT 350.855 2310.715 351.135 2310.995 ;
        RECT 351.475 2310.715 351.755 2310.995 ;
        RECT 352.095 2310.715 352.375 2310.995 ;
        RECT 350.235 2310.095 350.515 2310.375 ;
        RECT 350.855 2310.095 351.135 2310.375 ;
        RECT 351.475 2310.095 351.755 2310.375 ;
        RECT 352.095 2310.095 352.375 2310.375 ;
        RECT 350.235 2309.475 350.515 2309.755 ;
        RECT 350.855 2309.475 351.135 2309.755 ;
        RECT 351.475 2309.475 351.755 2309.755 ;
        RECT 352.095 2309.475 352.375 2309.755 ;
        RECT 350.235 2305.245 350.515 2305.525 ;
        RECT 350.855 2305.245 351.135 2305.525 ;
        RECT 351.475 2305.245 351.755 2305.525 ;
        RECT 352.095 2305.245 352.375 2305.525 ;
        RECT 350.235 2304.625 350.515 2304.905 ;
        RECT 350.855 2304.625 351.135 2304.905 ;
        RECT 351.475 2304.625 351.755 2304.905 ;
        RECT 352.095 2304.625 352.375 2304.905 ;
        RECT 350.235 2304.005 350.515 2304.285 ;
        RECT 350.855 2304.005 351.135 2304.285 ;
        RECT 351.475 2304.005 351.755 2304.285 ;
        RECT 352.095 2304.005 352.375 2304.285 ;
        RECT 350.235 2303.385 350.515 2303.665 ;
        RECT 350.855 2303.385 351.135 2303.665 ;
        RECT 351.475 2303.385 351.755 2303.665 ;
        RECT 352.095 2303.385 352.375 2303.665 ;
        RECT 350.235 2302.765 350.515 2303.045 ;
        RECT 350.855 2302.765 351.135 2303.045 ;
        RECT 351.475 2302.765 351.755 2303.045 ;
        RECT 352.095 2302.765 352.375 2303.045 ;
        RECT 350.235 2302.145 350.515 2302.425 ;
        RECT 350.855 2302.145 351.135 2302.425 ;
        RECT 351.475 2302.145 351.755 2302.425 ;
        RECT 352.095 2302.145 352.375 2302.425 ;
        RECT 350.235 2301.525 350.515 2301.805 ;
        RECT 350.855 2301.525 351.135 2301.805 ;
        RECT 351.475 2301.525 351.755 2301.805 ;
        RECT 352.095 2301.525 352.375 2301.805 ;
        RECT 350.235 2300.905 350.515 2301.185 ;
        RECT 350.855 2300.905 351.135 2301.185 ;
        RECT 351.475 2300.905 351.755 2301.185 ;
        RECT 352.095 2300.905 352.375 2301.185 ;
        RECT 350.235 2300.285 350.515 2300.565 ;
        RECT 350.855 2300.285 351.135 2300.565 ;
        RECT 351.475 2300.285 351.755 2300.565 ;
        RECT 352.095 2300.285 352.375 2300.565 ;
        RECT 350.235 2299.665 350.515 2299.945 ;
        RECT 350.855 2299.665 351.135 2299.945 ;
        RECT 351.475 2299.665 351.755 2299.945 ;
        RECT 352.095 2299.665 352.375 2299.945 ;
        RECT 350.235 2299.045 350.515 2299.325 ;
        RECT 350.855 2299.045 351.135 2299.325 ;
        RECT 351.475 2299.045 351.755 2299.325 ;
        RECT 352.095 2299.045 352.375 2299.325 ;
        RECT 350.235 2298.425 350.515 2298.705 ;
        RECT 350.855 2298.425 351.135 2298.705 ;
        RECT 351.475 2298.425 351.755 2298.705 ;
        RECT 352.095 2298.425 352.375 2298.705 ;
        RECT 350.235 2297.805 350.515 2298.085 ;
        RECT 350.855 2297.805 351.135 2298.085 ;
        RECT 351.475 2297.805 351.755 2298.085 ;
        RECT 352.095 2297.805 352.375 2298.085 ;
        RECT 350.235 2297.185 350.515 2297.465 ;
        RECT 350.855 2297.185 351.135 2297.465 ;
        RECT 351.475 2297.185 351.755 2297.465 ;
        RECT 352.095 2297.185 352.375 2297.465 ;
        RECT 350.235 2296.565 350.515 2296.845 ;
        RECT 350.855 2296.565 351.135 2296.845 ;
        RECT 351.475 2296.565 351.755 2296.845 ;
        RECT 352.095 2296.565 352.375 2296.845 ;
        RECT 350.235 2295.945 350.515 2296.225 ;
        RECT 350.855 2295.945 351.135 2296.225 ;
        RECT 351.475 2295.945 351.755 2296.225 ;
        RECT 352.095 2295.945 352.375 2296.225 ;
        RECT 350.235 2293.395 350.515 2293.675 ;
        RECT 350.855 2293.395 351.135 2293.675 ;
        RECT 351.475 2293.395 351.755 2293.675 ;
        RECT 352.095 2293.395 352.375 2293.675 ;
        RECT 350.235 2292.775 350.515 2293.055 ;
        RECT 350.855 2292.775 351.135 2293.055 ;
        RECT 351.475 2292.775 351.755 2293.055 ;
        RECT 352.095 2292.775 352.375 2293.055 ;
        RECT 350.235 2292.155 350.515 2292.435 ;
        RECT 350.855 2292.155 351.135 2292.435 ;
        RECT 351.475 2292.155 351.755 2292.435 ;
        RECT 352.095 2292.155 352.375 2292.435 ;
        RECT 350.235 2291.535 350.515 2291.815 ;
        RECT 350.855 2291.535 351.135 2291.815 ;
        RECT 351.475 2291.535 351.755 2291.815 ;
        RECT 352.095 2291.535 352.375 2291.815 ;
        RECT 350.235 2290.915 350.515 2291.195 ;
        RECT 350.855 2290.915 351.135 2291.195 ;
        RECT 351.475 2290.915 351.755 2291.195 ;
        RECT 352.095 2290.915 352.375 2291.195 ;
        RECT 350.235 2290.295 350.515 2290.575 ;
        RECT 350.855 2290.295 351.135 2290.575 ;
        RECT 351.475 2290.295 351.755 2290.575 ;
        RECT 352.095 2290.295 352.375 2290.575 ;
        RECT 350.235 2289.675 350.515 2289.955 ;
        RECT 350.855 2289.675 351.135 2289.955 ;
        RECT 351.475 2289.675 351.755 2289.955 ;
        RECT 352.095 2289.675 352.375 2289.955 ;
        RECT 350.235 2289.055 350.515 2289.335 ;
        RECT 350.855 2289.055 351.135 2289.335 ;
        RECT 351.475 2289.055 351.755 2289.335 ;
        RECT 352.095 2289.055 352.375 2289.335 ;
        RECT 350.235 2288.435 350.515 2288.715 ;
        RECT 350.855 2288.435 351.135 2288.715 ;
        RECT 351.475 2288.435 351.755 2288.715 ;
        RECT 352.095 2288.435 352.375 2288.715 ;
        RECT 350.235 2287.815 350.515 2288.095 ;
        RECT 350.855 2287.815 351.135 2288.095 ;
        RECT 351.475 2287.815 351.755 2288.095 ;
        RECT 352.095 2287.815 352.375 2288.095 ;
        RECT 350.235 2287.195 350.515 2287.475 ;
        RECT 350.855 2287.195 351.135 2287.475 ;
        RECT 351.475 2287.195 351.755 2287.475 ;
        RECT 352.095 2287.195 352.375 2287.475 ;
        RECT 350.235 2286.575 350.515 2286.855 ;
        RECT 350.855 2286.575 351.135 2286.855 ;
        RECT 351.475 2286.575 351.755 2286.855 ;
        RECT 352.095 2286.575 352.375 2286.855 ;
        RECT 350.235 2285.955 350.515 2286.235 ;
        RECT 350.855 2285.955 351.135 2286.235 ;
        RECT 351.475 2285.955 351.755 2286.235 ;
        RECT 352.095 2285.955 352.375 2286.235 ;
        RECT 350.235 2285.335 350.515 2285.615 ;
        RECT 350.855 2285.335 351.135 2285.615 ;
        RECT 351.475 2285.335 351.755 2285.615 ;
        RECT 352.095 2285.335 352.375 2285.615 ;
        RECT 350.235 2284.715 350.515 2284.995 ;
        RECT 350.855 2284.715 351.135 2284.995 ;
        RECT 351.475 2284.715 351.755 2284.995 ;
        RECT 352.095 2284.715 352.375 2284.995 ;
        RECT 350.235 2284.095 350.515 2284.375 ;
        RECT 350.855 2284.095 351.135 2284.375 ;
        RECT 351.475 2284.095 351.755 2284.375 ;
        RECT 352.095 2284.095 352.375 2284.375 ;
        RECT 350.235 2280.245 350.515 2280.525 ;
        RECT 350.855 2280.245 351.135 2280.525 ;
        RECT 351.475 2280.245 351.755 2280.525 ;
        RECT 352.095 2280.245 352.375 2280.525 ;
        RECT 350.235 2279.625 350.515 2279.905 ;
        RECT 350.855 2279.625 351.135 2279.905 ;
        RECT 351.475 2279.625 351.755 2279.905 ;
        RECT 352.095 2279.625 352.375 2279.905 ;
        RECT 350.235 2279.005 350.515 2279.285 ;
        RECT 350.855 2279.005 351.135 2279.285 ;
        RECT 351.475 2279.005 351.755 2279.285 ;
        RECT 352.095 2279.005 352.375 2279.285 ;
        RECT 350.235 2278.385 350.515 2278.665 ;
        RECT 350.855 2278.385 351.135 2278.665 ;
        RECT 351.475 2278.385 351.755 2278.665 ;
        RECT 352.095 2278.385 352.375 2278.665 ;
        RECT 350.235 2277.765 350.515 2278.045 ;
        RECT 350.855 2277.765 351.135 2278.045 ;
        RECT 351.475 2277.765 351.755 2278.045 ;
        RECT 352.095 2277.765 352.375 2278.045 ;
        RECT 350.235 2277.145 350.515 2277.425 ;
        RECT 350.855 2277.145 351.135 2277.425 ;
        RECT 351.475 2277.145 351.755 2277.425 ;
        RECT 352.095 2277.145 352.375 2277.425 ;
        RECT 350.235 2276.525 350.515 2276.805 ;
        RECT 350.855 2276.525 351.135 2276.805 ;
        RECT 351.475 2276.525 351.755 2276.805 ;
        RECT 352.095 2276.525 352.375 2276.805 ;
        RECT 350.235 2275.905 350.515 2276.185 ;
        RECT 350.855 2275.905 351.135 2276.185 ;
        RECT 351.475 2275.905 351.755 2276.185 ;
        RECT 352.095 2275.905 352.375 2276.185 ;
        RECT 350.235 2275.285 350.515 2275.565 ;
        RECT 350.855 2275.285 351.135 2275.565 ;
        RECT 351.475 2275.285 351.755 2275.565 ;
        RECT 352.095 2275.285 352.375 2275.565 ;
        RECT 350.235 2274.665 350.515 2274.945 ;
        RECT 350.855 2274.665 351.135 2274.945 ;
        RECT 351.475 2274.665 351.755 2274.945 ;
        RECT 352.095 2274.665 352.375 2274.945 ;
        RECT 350.235 2274.045 350.515 2274.325 ;
        RECT 350.855 2274.045 351.135 2274.325 ;
        RECT 351.475 2274.045 351.755 2274.325 ;
        RECT 352.095 2274.045 352.375 2274.325 ;
        RECT 350.235 2273.425 350.515 2273.705 ;
        RECT 350.855 2273.425 351.135 2273.705 ;
        RECT 351.475 2273.425 351.755 2273.705 ;
        RECT 352.095 2273.425 352.375 2273.705 ;
        RECT 350.235 2272.805 350.515 2273.085 ;
        RECT 350.855 2272.805 351.135 2273.085 ;
        RECT 351.475 2272.805 351.755 2273.085 ;
        RECT 352.095 2272.805 352.375 2273.085 ;
        RECT 350.235 2272.185 350.515 2272.465 ;
        RECT 350.855 2272.185 351.135 2272.465 ;
        RECT 351.475 2272.185 351.755 2272.465 ;
        RECT 352.095 2272.185 352.375 2272.465 ;
        RECT 350.235 2271.565 350.515 2271.845 ;
        RECT 350.855 2271.565 351.135 2271.845 ;
        RECT 351.475 2271.565 351.755 2271.845 ;
        RECT 352.095 2271.565 352.375 2271.845 ;
        RECT 3527.625 2238.155 3527.905 2238.435 ;
        RECT 3528.245 2238.155 3528.525 2238.435 ;
        RECT 3528.865 2238.155 3529.145 2238.435 ;
        RECT 3529.485 2238.155 3529.765 2238.435 ;
        RECT 3527.625 2237.535 3527.905 2237.815 ;
        RECT 3528.245 2237.535 3528.525 2237.815 ;
        RECT 3528.865 2237.535 3529.145 2237.815 ;
        RECT 3529.485 2237.535 3529.765 2237.815 ;
        RECT 3527.625 2236.915 3527.905 2237.195 ;
        RECT 3528.245 2236.915 3528.525 2237.195 ;
        RECT 3528.865 2236.915 3529.145 2237.195 ;
        RECT 3529.485 2236.915 3529.765 2237.195 ;
        RECT 3527.625 2236.295 3527.905 2236.575 ;
        RECT 3528.245 2236.295 3528.525 2236.575 ;
        RECT 3528.865 2236.295 3529.145 2236.575 ;
        RECT 3529.485 2236.295 3529.765 2236.575 ;
        RECT 3527.625 2235.675 3527.905 2235.955 ;
        RECT 3528.245 2235.675 3528.525 2235.955 ;
        RECT 3528.865 2235.675 3529.145 2235.955 ;
        RECT 3529.485 2235.675 3529.765 2235.955 ;
        RECT 3527.625 2235.055 3527.905 2235.335 ;
        RECT 3528.245 2235.055 3528.525 2235.335 ;
        RECT 3528.865 2235.055 3529.145 2235.335 ;
        RECT 3529.485 2235.055 3529.765 2235.335 ;
        RECT 3527.625 2234.435 3527.905 2234.715 ;
        RECT 3528.245 2234.435 3528.525 2234.715 ;
        RECT 3528.865 2234.435 3529.145 2234.715 ;
        RECT 3529.485 2234.435 3529.765 2234.715 ;
        RECT 3527.625 2233.815 3527.905 2234.095 ;
        RECT 3528.245 2233.815 3528.525 2234.095 ;
        RECT 3528.865 2233.815 3529.145 2234.095 ;
        RECT 3529.485 2233.815 3529.765 2234.095 ;
        RECT 3527.625 2233.195 3527.905 2233.475 ;
        RECT 3528.245 2233.195 3528.525 2233.475 ;
        RECT 3528.865 2233.195 3529.145 2233.475 ;
        RECT 3529.485 2233.195 3529.765 2233.475 ;
        RECT 3527.625 2232.575 3527.905 2232.855 ;
        RECT 3528.245 2232.575 3528.525 2232.855 ;
        RECT 3528.865 2232.575 3529.145 2232.855 ;
        RECT 3529.485 2232.575 3529.765 2232.855 ;
        RECT 3527.625 2231.955 3527.905 2232.235 ;
        RECT 3528.245 2231.955 3528.525 2232.235 ;
        RECT 3528.865 2231.955 3529.145 2232.235 ;
        RECT 3529.485 2231.955 3529.765 2232.235 ;
        RECT 3527.625 2231.335 3527.905 2231.615 ;
        RECT 3528.245 2231.335 3528.525 2231.615 ;
        RECT 3528.865 2231.335 3529.145 2231.615 ;
        RECT 3529.485 2231.335 3529.765 2231.615 ;
        RECT 3527.625 2230.715 3527.905 2230.995 ;
        RECT 3528.245 2230.715 3528.525 2230.995 ;
        RECT 3528.865 2230.715 3529.145 2230.995 ;
        RECT 3529.485 2230.715 3529.765 2230.995 ;
        RECT 3527.625 2230.095 3527.905 2230.375 ;
        RECT 3528.245 2230.095 3528.525 2230.375 ;
        RECT 3528.865 2230.095 3529.145 2230.375 ;
        RECT 3529.485 2230.095 3529.765 2230.375 ;
        RECT 3527.625 2229.475 3527.905 2229.755 ;
        RECT 3528.245 2229.475 3528.525 2229.755 ;
        RECT 3528.865 2229.475 3529.145 2229.755 ;
        RECT 3529.485 2229.475 3529.765 2229.755 ;
        RECT 3527.625 2225.625 3527.905 2225.905 ;
        RECT 3528.245 2225.625 3528.525 2225.905 ;
        RECT 3528.865 2225.625 3529.145 2225.905 ;
        RECT 3529.485 2225.625 3529.765 2225.905 ;
        RECT 3527.625 2225.005 3527.905 2225.285 ;
        RECT 3528.245 2225.005 3528.525 2225.285 ;
        RECT 3528.865 2225.005 3529.145 2225.285 ;
        RECT 3529.485 2225.005 3529.765 2225.285 ;
        RECT 3527.625 2224.385 3527.905 2224.665 ;
        RECT 3528.245 2224.385 3528.525 2224.665 ;
        RECT 3528.865 2224.385 3529.145 2224.665 ;
        RECT 3529.485 2224.385 3529.765 2224.665 ;
        RECT 3527.625 2223.765 3527.905 2224.045 ;
        RECT 3528.245 2223.765 3528.525 2224.045 ;
        RECT 3528.865 2223.765 3529.145 2224.045 ;
        RECT 3529.485 2223.765 3529.765 2224.045 ;
        RECT 3527.625 2223.145 3527.905 2223.425 ;
        RECT 3528.245 2223.145 3528.525 2223.425 ;
        RECT 3528.865 2223.145 3529.145 2223.425 ;
        RECT 3529.485 2223.145 3529.765 2223.425 ;
        RECT 3527.625 2222.525 3527.905 2222.805 ;
        RECT 3528.245 2222.525 3528.525 2222.805 ;
        RECT 3528.865 2222.525 3529.145 2222.805 ;
        RECT 3529.485 2222.525 3529.765 2222.805 ;
        RECT 3527.625 2221.905 3527.905 2222.185 ;
        RECT 3528.245 2221.905 3528.525 2222.185 ;
        RECT 3528.865 2221.905 3529.145 2222.185 ;
        RECT 3529.485 2221.905 3529.765 2222.185 ;
        RECT 3527.625 2221.285 3527.905 2221.565 ;
        RECT 3528.245 2221.285 3528.525 2221.565 ;
        RECT 3528.865 2221.285 3529.145 2221.565 ;
        RECT 3529.485 2221.285 3529.765 2221.565 ;
        RECT 3527.625 2220.665 3527.905 2220.945 ;
        RECT 3528.245 2220.665 3528.525 2220.945 ;
        RECT 3528.865 2220.665 3529.145 2220.945 ;
        RECT 3529.485 2220.665 3529.765 2220.945 ;
        RECT 3527.625 2220.045 3527.905 2220.325 ;
        RECT 3528.245 2220.045 3528.525 2220.325 ;
        RECT 3528.865 2220.045 3529.145 2220.325 ;
        RECT 3529.485 2220.045 3529.765 2220.325 ;
        RECT 3527.625 2219.425 3527.905 2219.705 ;
        RECT 3528.245 2219.425 3528.525 2219.705 ;
        RECT 3528.865 2219.425 3529.145 2219.705 ;
        RECT 3529.485 2219.425 3529.765 2219.705 ;
        RECT 3527.625 2218.805 3527.905 2219.085 ;
        RECT 3528.245 2218.805 3528.525 2219.085 ;
        RECT 3528.865 2218.805 3529.145 2219.085 ;
        RECT 3529.485 2218.805 3529.765 2219.085 ;
        RECT 3527.625 2218.185 3527.905 2218.465 ;
        RECT 3528.245 2218.185 3528.525 2218.465 ;
        RECT 3528.865 2218.185 3529.145 2218.465 ;
        RECT 3529.485 2218.185 3529.765 2218.465 ;
        RECT 3527.625 2217.565 3527.905 2217.845 ;
        RECT 3528.245 2217.565 3528.525 2217.845 ;
        RECT 3528.865 2217.565 3529.145 2217.845 ;
        RECT 3529.485 2217.565 3529.765 2217.845 ;
        RECT 3527.625 2216.945 3527.905 2217.225 ;
        RECT 3528.245 2216.945 3528.525 2217.225 ;
        RECT 3528.865 2216.945 3529.145 2217.225 ;
        RECT 3529.485 2216.945 3529.765 2217.225 ;
        RECT 3527.625 2216.325 3527.905 2216.605 ;
        RECT 3528.245 2216.325 3528.525 2216.605 ;
        RECT 3528.865 2216.325 3529.145 2216.605 ;
        RECT 3529.485 2216.325 3529.765 2216.605 ;
        RECT 3527.625 2213.775 3527.905 2214.055 ;
        RECT 3528.245 2213.775 3528.525 2214.055 ;
        RECT 3528.865 2213.775 3529.145 2214.055 ;
        RECT 3529.485 2213.775 3529.765 2214.055 ;
        RECT 3527.625 2213.155 3527.905 2213.435 ;
        RECT 3528.245 2213.155 3528.525 2213.435 ;
        RECT 3528.865 2213.155 3529.145 2213.435 ;
        RECT 3529.485 2213.155 3529.765 2213.435 ;
        RECT 3527.625 2212.535 3527.905 2212.815 ;
        RECT 3528.245 2212.535 3528.525 2212.815 ;
        RECT 3528.865 2212.535 3529.145 2212.815 ;
        RECT 3529.485 2212.535 3529.765 2212.815 ;
        RECT 3527.625 2211.915 3527.905 2212.195 ;
        RECT 3528.245 2211.915 3528.525 2212.195 ;
        RECT 3528.865 2211.915 3529.145 2212.195 ;
        RECT 3529.485 2211.915 3529.765 2212.195 ;
        RECT 3527.625 2211.295 3527.905 2211.575 ;
        RECT 3528.245 2211.295 3528.525 2211.575 ;
        RECT 3528.865 2211.295 3529.145 2211.575 ;
        RECT 3529.485 2211.295 3529.765 2211.575 ;
        RECT 3527.625 2210.675 3527.905 2210.955 ;
        RECT 3528.245 2210.675 3528.525 2210.955 ;
        RECT 3528.865 2210.675 3529.145 2210.955 ;
        RECT 3529.485 2210.675 3529.765 2210.955 ;
        RECT 3527.625 2210.055 3527.905 2210.335 ;
        RECT 3528.245 2210.055 3528.525 2210.335 ;
        RECT 3528.865 2210.055 3529.145 2210.335 ;
        RECT 3529.485 2210.055 3529.765 2210.335 ;
        RECT 3527.625 2209.435 3527.905 2209.715 ;
        RECT 3528.245 2209.435 3528.525 2209.715 ;
        RECT 3528.865 2209.435 3529.145 2209.715 ;
        RECT 3529.485 2209.435 3529.765 2209.715 ;
        RECT 3527.625 2208.815 3527.905 2209.095 ;
        RECT 3528.245 2208.815 3528.525 2209.095 ;
        RECT 3528.865 2208.815 3529.145 2209.095 ;
        RECT 3529.485 2208.815 3529.765 2209.095 ;
        RECT 3527.625 2208.195 3527.905 2208.475 ;
        RECT 3528.245 2208.195 3528.525 2208.475 ;
        RECT 3528.865 2208.195 3529.145 2208.475 ;
        RECT 3529.485 2208.195 3529.765 2208.475 ;
        RECT 3527.625 2207.575 3527.905 2207.855 ;
        RECT 3528.245 2207.575 3528.525 2207.855 ;
        RECT 3528.865 2207.575 3529.145 2207.855 ;
        RECT 3529.485 2207.575 3529.765 2207.855 ;
        RECT 3527.625 2206.955 3527.905 2207.235 ;
        RECT 3528.245 2206.955 3528.525 2207.235 ;
        RECT 3528.865 2206.955 3529.145 2207.235 ;
        RECT 3529.485 2206.955 3529.765 2207.235 ;
        RECT 3527.625 2206.335 3527.905 2206.615 ;
        RECT 3528.245 2206.335 3528.525 2206.615 ;
        RECT 3528.865 2206.335 3529.145 2206.615 ;
        RECT 3529.485 2206.335 3529.765 2206.615 ;
        RECT 3527.625 2205.715 3527.905 2205.995 ;
        RECT 3528.245 2205.715 3528.525 2205.995 ;
        RECT 3528.865 2205.715 3529.145 2205.995 ;
        RECT 3529.485 2205.715 3529.765 2205.995 ;
        RECT 3527.625 2205.095 3527.905 2205.375 ;
        RECT 3528.245 2205.095 3528.525 2205.375 ;
        RECT 3528.865 2205.095 3529.145 2205.375 ;
        RECT 3529.485 2205.095 3529.765 2205.375 ;
        RECT 3527.625 2204.475 3527.905 2204.755 ;
        RECT 3528.245 2204.475 3528.525 2204.755 ;
        RECT 3528.865 2204.475 3529.145 2204.755 ;
        RECT 3529.485 2204.475 3529.765 2204.755 ;
        RECT 3527.625 2200.245 3527.905 2200.525 ;
        RECT 3528.245 2200.245 3528.525 2200.525 ;
        RECT 3528.865 2200.245 3529.145 2200.525 ;
        RECT 3529.485 2200.245 3529.765 2200.525 ;
        RECT 3527.625 2199.625 3527.905 2199.905 ;
        RECT 3528.245 2199.625 3528.525 2199.905 ;
        RECT 3528.865 2199.625 3529.145 2199.905 ;
        RECT 3529.485 2199.625 3529.765 2199.905 ;
        RECT 3527.625 2199.005 3527.905 2199.285 ;
        RECT 3528.245 2199.005 3528.525 2199.285 ;
        RECT 3528.865 2199.005 3529.145 2199.285 ;
        RECT 3529.485 2199.005 3529.765 2199.285 ;
        RECT 3527.625 2198.385 3527.905 2198.665 ;
        RECT 3528.245 2198.385 3528.525 2198.665 ;
        RECT 3528.865 2198.385 3529.145 2198.665 ;
        RECT 3529.485 2198.385 3529.765 2198.665 ;
        RECT 3527.625 2197.765 3527.905 2198.045 ;
        RECT 3528.245 2197.765 3528.525 2198.045 ;
        RECT 3528.865 2197.765 3529.145 2198.045 ;
        RECT 3529.485 2197.765 3529.765 2198.045 ;
        RECT 3527.625 2197.145 3527.905 2197.425 ;
        RECT 3528.245 2197.145 3528.525 2197.425 ;
        RECT 3528.865 2197.145 3529.145 2197.425 ;
        RECT 3529.485 2197.145 3529.765 2197.425 ;
        RECT 3527.625 2196.525 3527.905 2196.805 ;
        RECT 3528.245 2196.525 3528.525 2196.805 ;
        RECT 3528.865 2196.525 3529.145 2196.805 ;
        RECT 3529.485 2196.525 3529.765 2196.805 ;
        RECT 3527.625 2195.905 3527.905 2196.185 ;
        RECT 3528.245 2195.905 3528.525 2196.185 ;
        RECT 3528.865 2195.905 3529.145 2196.185 ;
        RECT 3529.485 2195.905 3529.765 2196.185 ;
        RECT 3527.625 2195.285 3527.905 2195.565 ;
        RECT 3528.245 2195.285 3528.525 2195.565 ;
        RECT 3528.865 2195.285 3529.145 2195.565 ;
        RECT 3529.485 2195.285 3529.765 2195.565 ;
        RECT 3527.625 2194.665 3527.905 2194.945 ;
        RECT 3528.245 2194.665 3528.525 2194.945 ;
        RECT 3528.865 2194.665 3529.145 2194.945 ;
        RECT 3529.485 2194.665 3529.765 2194.945 ;
        RECT 3527.625 2194.045 3527.905 2194.325 ;
        RECT 3528.245 2194.045 3528.525 2194.325 ;
        RECT 3528.865 2194.045 3529.145 2194.325 ;
        RECT 3529.485 2194.045 3529.765 2194.325 ;
        RECT 3527.625 2193.425 3527.905 2193.705 ;
        RECT 3528.245 2193.425 3528.525 2193.705 ;
        RECT 3528.865 2193.425 3529.145 2193.705 ;
        RECT 3529.485 2193.425 3529.765 2193.705 ;
        RECT 3527.625 2192.805 3527.905 2193.085 ;
        RECT 3528.245 2192.805 3528.525 2193.085 ;
        RECT 3528.865 2192.805 3529.145 2193.085 ;
        RECT 3529.485 2192.805 3529.765 2193.085 ;
        RECT 3527.625 2192.185 3527.905 2192.465 ;
        RECT 3528.245 2192.185 3528.525 2192.465 ;
        RECT 3528.865 2192.185 3529.145 2192.465 ;
        RECT 3529.485 2192.185 3529.765 2192.465 ;
        RECT 3527.625 2191.565 3527.905 2191.845 ;
        RECT 3528.245 2191.565 3528.525 2191.845 ;
        RECT 3528.865 2191.565 3529.145 2191.845 ;
        RECT 3529.485 2191.565 3529.765 2191.845 ;
        RECT 3527.625 2190.945 3527.905 2191.225 ;
        RECT 3528.245 2190.945 3528.525 2191.225 ;
        RECT 3528.865 2190.945 3529.145 2191.225 ;
        RECT 3529.485 2190.945 3529.765 2191.225 ;
        RECT 3527.625 2188.395 3527.905 2188.675 ;
        RECT 3528.245 2188.395 3528.525 2188.675 ;
        RECT 3528.865 2188.395 3529.145 2188.675 ;
        RECT 3529.485 2188.395 3529.765 2188.675 ;
        RECT 3527.625 2187.775 3527.905 2188.055 ;
        RECT 3528.245 2187.775 3528.525 2188.055 ;
        RECT 3528.865 2187.775 3529.145 2188.055 ;
        RECT 3529.485 2187.775 3529.765 2188.055 ;
        RECT 3527.625 2187.155 3527.905 2187.435 ;
        RECT 3528.245 2187.155 3528.525 2187.435 ;
        RECT 3528.865 2187.155 3529.145 2187.435 ;
        RECT 3529.485 2187.155 3529.765 2187.435 ;
        RECT 3527.625 2186.535 3527.905 2186.815 ;
        RECT 3528.245 2186.535 3528.525 2186.815 ;
        RECT 3528.865 2186.535 3529.145 2186.815 ;
        RECT 3529.485 2186.535 3529.765 2186.815 ;
        RECT 3527.625 2185.915 3527.905 2186.195 ;
        RECT 3528.245 2185.915 3528.525 2186.195 ;
        RECT 3528.865 2185.915 3529.145 2186.195 ;
        RECT 3529.485 2185.915 3529.765 2186.195 ;
        RECT 3527.625 2185.295 3527.905 2185.575 ;
        RECT 3528.245 2185.295 3528.525 2185.575 ;
        RECT 3528.865 2185.295 3529.145 2185.575 ;
        RECT 3529.485 2185.295 3529.765 2185.575 ;
        RECT 3527.625 2184.675 3527.905 2184.955 ;
        RECT 3528.245 2184.675 3528.525 2184.955 ;
        RECT 3528.865 2184.675 3529.145 2184.955 ;
        RECT 3529.485 2184.675 3529.765 2184.955 ;
        RECT 3527.625 2184.055 3527.905 2184.335 ;
        RECT 3528.245 2184.055 3528.525 2184.335 ;
        RECT 3528.865 2184.055 3529.145 2184.335 ;
        RECT 3529.485 2184.055 3529.765 2184.335 ;
        RECT 3527.625 2183.435 3527.905 2183.715 ;
        RECT 3528.245 2183.435 3528.525 2183.715 ;
        RECT 3528.865 2183.435 3529.145 2183.715 ;
        RECT 3529.485 2183.435 3529.765 2183.715 ;
        RECT 3527.625 2182.815 3527.905 2183.095 ;
        RECT 3528.245 2182.815 3528.525 2183.095 ;
        RECT 3528.865 2182.815 3529.145 2183.095 ;
        RECT 3529.485 2182.815 3529.765 2183.095 ;
        RECT 3527.625 2182.195 3527.905 2182.475 ;
        RECT 3528.245 2182.195 3528.525 2182.475 ;
        RECT 3528.865 2182.195 3529.145 2182.475 ;
        RECT 3529.485 2182.195 3529.765 2182.475 ;
        RECT 3527.625 2181.575 3527.905 2181.855 ;
        RECT 3528.245 2181.575 3528.525 2181.855 ;
        RECT 3528.865 2181.575 3529.145 2181.855 ;
        RECT 3529.485 2181.575 3529.765 2181.855 ;
        RECT 3527.625 2180.955 3527.905 2181.235 ;
        RECT 3528.245 2180.955 3528.525 2181.235 ;
        RECT 3528.865 2180.955 3529.145 2181.235 ;
        RECT 3529.485 2180.955 3529.765 2181.235 ;
        RECT 3527.625 2175.375 3527.905 2175.655 ;
        RECT 3528.245 2175.375 3528.525 2175.655 ;
        RECT 3528.865 2175.375 3529.145 2175.655 ;
        RECT 3529.485 2175.375 3529.765 2175.655 ;
        RECT 3527.625 2174.755 3527.905 2175.035 ;
        RECT 3528.245 2174.755 3528.525 2175.035 ;
        RECT 3528.865 2174.755 3529.145 2175.035 ;
        RECT 3529.485 2174.755 3529.765 2175.035 ;
        RECT 3527.625 2174.135 3527.905 2174.415 ;
        RECT 3528.245 2174.135 3528.525 2174.415 ;
        RECT 3528.865 2174.135 3529.145 2174.415 ;
        RECT 3529.485 2174.135 3529.765 2174.415 ;
        RECT 3527.625 2173.515 3527.905 2173.795 ;
        RECT 3528.245 2173.515 3528.525 2173.795 ;
        RECT 3528.865 2173.515 3529.145 2173.795 ;
        RECT 3529.485 2173.515 3529.765 2173.795 ;
        RECT 3527.625 2172.895 3527.905 2173.175 ;
        RECT 3528.245 2172.895 3528.525 2173.175 ;
        RECT 3528.865 2172.895 3529.145 2173.175 ;
        RECT 3529.485 2172.895 3529.765 2173.175 ;
        RECT 3527.625 2172.275 3527.905 2172.555 ;
        RECT 3528.245 2172.275 3528.525 2172.555 ;
        RECT 3528.865 2172.275 3529.145 2172.555 ;
        RECT 3529.485 2172.275 3529.765 2172.555 ;
        RECT 3527.625 2171.655 3527.905 2171.935 ;
        RECT 3528.245 2171.655 3528.525 2171.935 ;
        RECT 3528.865 2171.655 3529.145 2171.935 ;
        RECT 3529.485 2171.655 3529.765 2171.935 ;
        RECT 3527.625 2171.035 3527.905 2171.315 ;
        RECT 3528.245 2171.035 3528.525 2171.315 ;
        RECT 3528.865 2171.035 3529.145 2171.315 ;
        RECT 3529.485 2171.035 3529.765 2171.315 ;
        RECT 3527.625 2170.415 3527.905 2170.695 ;
        RECT 3528.245 2170.415 3528.525 2170.695 ;
        RECT 3528.865 2170.415 3529.145 2170.695 ;
        RECT 3529.485 2170.415 3529.765 2170.695 ;
        RECT 3527.625 2169.795 3527.905 2170.075 ;
        RECT 3528.245 2169.795 3528.525 2170.075 ;
        RECT 3528.865 2169.795 3529.145 2170.075 ;
        RECT 3529.485 2169.795 3529.765 2170.075 ;
        RECT 3527.625 2169.175 3527.905 2169.455 ;
        RECT 3528.245 2169.175 3528.525 2169.455 ;
        RECT 3528.865 2169.175 3529.145 2169.455 ;
        RECT 3529.485 2169.175 3529.765 2169.455 ;
        RECT 3527.625 2168.555 3527.905 2168.835 ;
        RECT 3528.245 2168.555 3528.525 2168.835 ;
        RECT 3528.865 2168.555 3529.145 2168.835 ;
        RECT 3529.485 2168.555 3529.765 2168.835 ;
        RECT 3527.625 2167.935 3527.905 2168.215 ;
        RECT 3528.245 2167.935 3528.525 2168.215 ;
        RECT 3528.865 2167.935 3529.145 2168.215 ;
        RECT 3529.485 2167.935 3529.765 2168.215 ;
        RECT 3527.625 2167.315 3527.905 2167.595 ;
        RECT 3528.245 2167.315 3528.525 2167.595 ;
        RECT 3528.865 2167.315 3529.145 2167.595 ;
        RECT 3529.485 2167.315 3529.765 2167.595 ;
        RECT 3527.625 2166.695 3527.905 2166.975 ;
        RECT 3528.245 2166.695 3528.525 2166.975 ;
        RECT 3528.865 2166.695 3529.145 2166.975 ;
        RECT 3529.485 2166.695 3529.765 2166.975 ;
        RECT 350.235 2138.025 350.515 2138.305 ;
        RECT 350.855 2138.025 351.135 2138.305 ;
        RECT 351.475 2138.025 351.755 2138.305 ;
        RECT 352.095 2138.025 352.375 2138.305 ;
        RECT 350.235 2137.405 350.515 2137.685 ;
        RECT 350.855 2137.405 351.135 2137.685 ;
        RECT 351.475 2137.405 351.755 2137.685 ;
        RECT 352.095 2137.405 352.375 2137.685 ;
        RECT 350.235 2136.785 350.515 2137.065 ;
        RECT 350.855 2136.785 351.135 2137.065 ;
        RECT 351.475 2136.785 351.755 2137.065 ;
        RECT 352.095 2136.785 352.375 2137.065 ;
        RECT 350.235 2136.165 350.515 2136.445 ;
        RECT 350.855 2136.165 351.135 2136.445 ;
        RECT 351.475 2136.165 351.755 2136.445 ;
        RECT 352.095 2136.165 352.375 2136.445 ;
        RECT 350.235 2135.545 350.515 2135.825 ;
        RECT 350.855 2135.545 351.135 2135.825 ;
        RECT 351.475 2135.545 351.755 2135.825 ;
        RECT 352.095 2135.545 352.375 2135.825 ;
        RECT 350.235 2134.925 350.515 2135.205 ;
        RECT 350.855 2134.925 351.135 2135.205 ;
        RECT 351.475 2134.925 351.755 2135.205 ;
        RECT 352.095 2134.925 352.375 2135.205 ;
        RECT 350.235 2134.305 350.515 2134.585 ;
        RECT 350.855 2134.305 351.135 2134.585 ;
        RECT 351.475 2134.305 351.755 2134.585 ;
        RECT 352.095 2134.305 352.375 2134.585 ;
        RECT 350.235 2133.685 350.515 2133.965 ;
        RECT 350.855 2133.685 351.135 2133.965 ;
        RECT 351.475 2133.685 351.755 2133.965 ;
        RECT 352.095 2133.685 352.375 2133.965 ;
        RECT 350.235 2133.065 350.515 2133.345 ;
        RECT 350.855 2133.065 351.135 2133.345 ;
        RECT 351.475 2133.065 351.755 2133.345 ;
        RECT 352.095 2133.065 352.375 2133.345 ;
        RECT 350.235 2132.445 350.515 2132.725 ;
        RECT 350.855 2132.445 351.135 2132.725 ;
        RECT 351.475 2132.445 351.755 2132.725 ;
        RECT 352.095 2132.445 352.375 2132.725 ;
        RECT 350.235 2131.825 350.515 2132.105 ;
        RECT 350.855 2131.825 351.135 2132.105 ;
        RECT 351.475 2131.825 351.755 2132.105 ;
        RECT 352.095 2131.825 352.375 2132.105 ;
        RECT 350.235 2131.205 350.515 2131.485 ;
        RECT 350.855 2131.205 351.135 2131.485 ;
        RECT 351.475 2131.205 351.755 2131.485 ;
        RECT 352.095 2131.205 352.375 2131.485 ;
        RECT 350.235 2130.585 350.515 2130.865 ;
        RECT 350.855 2130.585 351.135 2130.865 ;
        RECT 351.475 2130.585 351.755 2130.865 ;
        RECT 352.095 2130.585 352.375 2130.865 ;
        RECT 350.235 2129.965 350.515 2130.245 ;
        RECT 350.855 2129.965 351.135 2130.245 ;
        RECT 351.475 2129.965 351.755 2130.245 ;
        RECT 352.095 2129.965 352.375 2130.245 ;
        RECT 350.235 2129.345 350.515 2129.625 ;
        RECT 350.855 2129.345 351.135 2129.625 ;
        RECT 351.475 2129.345 351.755 2129.625 ;
        RECT 352.095 2129.345 352.375 2129.625 ;
        RECT 350.235 2125.625 350.515 2125.905 ;
        RECT 350.855 2125.625 351.135 2125.905 ;
        RECT 351.475 2125.625 351.755 2125.905 ;
        RECT 352.095 2125.625 352.375 2125.905 ;
        RECT 350.235 2125.005 350.515 2125.285 ;
        RECT 350.855 2125.005 351.135 2125.285 ;
        RECT 351.475 2125.005 351.755 2125.285 ;
        RECT 352.095 2125.005 352.375 2125.285 ;
        RECT 350.235 2124.385 350.515 2124.665 ;
        RECT 350.855 2124.385 351.135 2124.665 ;
        RECT 351.475 2124.385 351.755 2124.665 ;
        RECT 352.095 2124.385 352.375 2124.665 ;
        RECT 350.235 2123.765 350.515 2124.045 ;
        RECT 350.855 2123.765 351.135 2124.045 ;
        RECT 351.475 2123.765 351.755 2124.045 ;
        RECT 352.095 2123.765 352.375 2124.045 ;
        RECT 350.235 2123.145 350.515 2123.425 ;
        RECT 350.855 2123.145 351.135 2123.425 ;
        RECT 351.475 2123.145 351.755 2123.425 ;
        RECT 352.095 2123.145 352.375 2123.425 ;
        RECT 350.235 2122.525 350.515 2122.805 ;
        RECT 350.855 2122.525 351.135 2122.805 ;
        RECT 351.475 2122.525 351.755 2122.805 ;
        RECT 352.095 2122.525 352.375 2122.805 ;
        RECT 350.235 2121.905 350.515 2122.185 ;
        RECT 350.855 2121.905 351.135 2122.185 ;
        RECT 351.475 2121.905 351.755 2122.185 ;
        RECT 352.095 2121.905 352.375 2122.185 ;
        RECT 350.235 2121.285 350.515 2121.565 ;
        RECT 350.855 2121.285 351.135 2121.565 ;
        RECT 351.475 2121.285 351.755 2121.565 ;
        RECT 352.095 2121.285 352.375 2121.565 ;
        RECT 350.235 2120.665 350.515 2120.945 ;
        RECT 350.855 2120.665 351.135 2120.945 ;
        RECT 351.475 2120.665 351.755 2120.945 ;
        RECT 352.095 2120.665 352.375 2120.945 ;
        RECT 350.235 2120.045 350.515 2120.325 ;
        RECT 350.855 2120.045 351.135 2120.325 ;
        RECT 351.475 2120.045 351.755 2120.325 ;
        RECT 352.095 2120.045 352.375 2120.325 ;
        RECT 350.235 2119.425 350.515 2119.705 ;
        RECT 350.855 2119.425 351.135 2119.705 ;
        RECT 351.475 2119.425 351.755 2119.705 ;
        RECT 352.095 2119.425 352.375 2119.705 ;
        RECT 350.235 2118.805 350.515 2119.085 ;
        RECT 350.855 2118.805 351.135 2119.085 ;
        RECT 351.475 2118.805 351.755 2119.085 ;
        RECT 352.095 2118.805 352.375 2119.085 ;
        RECT 350.235 2118.185 350.515 2118.465 ;
        RECT 350.855 2118.185 351.135 2118.465 ;
        RECT 351.475 2118.185 351.755 2118.465 ;
        RECT 352.095 2118.185 352.375 2118.465 ;
        RECT 350.235 2117.565 350.515 2117.845 ;
        RECT 350.855 2117.565 351.135 2117.845 ;
        RECT 351.475 2117.565 351.755 2117.845 ;
        RECT 352.095 2117.565 352.375 2117.845 ;
        RECT 350.235 2116.945 350.515 2117.225 ;
        RECT 350.855 2116.945 351.135 2117.225 ;
        RECT 351.475 2116.945 351.755 2117.225 ;
        RECT 352.095 2116.945 352.375 2117.225 ;
        RECT 350.235 2116.325 350.515 2116.605 ;
        RECT 350.855 2116.325 351.135 2116.605 ;
        RECT 351.475 2116.325 351.755 2116.605 ;
        RECT 352.095 2116.325 352.375 2116.605 ;
        RECT 350.235 2113.775 350.515 2114.055 ;
        RECT 350.855 2113.775 351.135 2114.055 ;
        RECT 351.475 2113.775 351.755 2114.055 ;
        RECT 352.095 2113.775 352.375 2114.055 ;
        RECT 350.235 2113.155 350.515 2113.435 ;
        RECT 350.855 2113.155 351.135 2113.435 ;
        RECT 351.475 2113.155 351.755 2113.435 ;
        RECT 352.095 2113.155 352.375 2113.435 ;
        RECT 350.235 2112.535 350.515 2112.815 ;
        RECT 350.855 2112.535 351.135 2112.815 ;
        RECT 351.475 2112.535 351.755 2112.815 ;
        RECT 352.095 2112.535 352.375 2112.815 ;
        RECT 350.235 2111.915 350.515 2112.195 ;
        RECT 350.855 2111.915 351.135 2112.195 ;
        RECT 351.475 2111.915 351.755 2112.195 ;
        RECT 352.095 2111.915 352.375 2112.195 ;
        RECT 350.235 2111.295 350.515 2111.575 ;
        RECT 350.855 2111.295 351.135 2111.575 ;
        RECT 351.475 2111.295 351.755 2111.575 ;
        RECT 352.095 2111.295 352.375 2111.575 ;
        RECT 350.235 2110.675 350.515 2110.955 ;
        RECT 350.855 2110.675 351.135 2110.955 ;
        RECT 351.475 2110.675 351.755 2110.955 ;
        RECT 352.095 2110.675 352.375 2110.955 ;
        RECT 350.235 2110.055 350.515 2110.335 ;
        RECT 350.855 2110.055 351.135 2110.335 ;
        RECT 351.475 2110.055 351.755 2110.335 ;
        RECT 352.095 2110.055 352.375 2110.335 ;
        RECT 350.235 2109.435 350.515 2109.715 ;
        RECT 350.855 2109.435 351.135 2109.715 ;
        RECT 351.475 2109.435 351.755 2109.715 ;
        RECT 352.095 2109.435 352.375 2109.715 ;
        RECT 350.235 2108.815 350.515 2109.095 ;
        RECT 350.855 2108.815 351.135 2109.095 ;
        RECT 351.475 2108.815 351.755 2109.095 ;
        RECT 352.095 2108.815 352.375 2109.095 ;
        RECT 350.235 2108.195 350.515 2108.475 ;
        RECT 350.855 2108.195 351.135 2108.475 ;
        RECT 351.475 2108.195 351.755 2108.475 ;
        RECT 352.095 2108.195 352.375 2108.475 ;
        RECT 350.235 2107.575 350.515 2107.855 ;
        RECT 350.855 2107.575 351.135 2107.855 ;
        RECT 351.475 2107.575 351.755 2107.855 ;
        RECT 352.095 2107.575 352.375 2107.855 ;
        RECT 350.235 2106.955 350.515 2107.235 ;
        RECT 350.855 2106.955 351.135 2107.235 ;
        RECT 351.475 2106.955 351.755 2107.235 ;
        RECT 352.095 2106.955 352.375 2107.235 ;
        RECT 350.235 2106.335 350.515 2106.615 ;
        RECT 350.855 2106.335 351.135 2106.615 ;
        RECT 351.475 2106.335 351.755 2106.615 ;
        RECT 352.095 2106.335 352.375 2106.615 ;
        RECT 350.235 2105.715 350.515 2105.995 ;
        RECT 350.855 2105.715 351.135 2105.995 ;
        RECT 351.475 2105.715 351.755 2105.995 ;
        RECT 352.095 2105.715 352.375 2105.995 ;
        RECT 350.235 2105.095 350.515 2105.375 ;
        RECT 350.855 2105.095 351.135 2105.375 ;
        RECT 351.475 2105.095 351.755 2105.375 ;
        RECT 352.095 2105.095 352.375 2105.375 ;
        RECT 350.235 2104.475 350.515 2104.755 ;
        RECT 350.855 2104.475 351.135 2104.755 ;
        RECT 351.475 2104.475 351.755 2104.755 ;
        RECT 352.095 2104.475 352.375 2104.755 ;
        RECT 350.235 2100.245 350.515 2100.525 ;
        RECT 350.855 2100.245 351.135 2100.525 ;
        RECT 351.475 2100.245 351.755 2100.525 ;
        RECT 352.095 2100.245 352.375 2100.525 ;
        RECT 350.235 2099.625 350.515 2099.905 ;
        RECT 350.855 2099.625 351.135 2099.905 ;
        RECT 351.475 2099.625 351.755 2099.905 ;
        RECT 352.095 2099.625 352.375 2099.905 ;
        RECT 350.235 2099.005 350.515 2099.285 ;
        RECT 350.855 2099.005 351.135 2099.285 ;
        RECT 351.475 2099.005 351.755 2099.285 ;
        RECT 352.095 2099.005 352.375 2099.285 ;
        RECT 350.235 2098.385 350.515 2098.665 ;
        RECT 350.855 2098.385 351.135 2098.665 ;
        RECT 351.475 2098.385 351.755 2098.665 ;
        RECT 352.095 2098.385 352.375 2098.665 ;
        RECT 350.235 2097.765 350.515 2098.045 ;
        RECT 350.855 2097.765 351.135 2098.045 ;
        RECT 351.475 2097.765 351.755 2098.045 ;
        RECT 352.095 2097.765 352.375 2098.045 ;
        RECT 350.235 2097.145 350.515 2097.425 ;
        RECT 350.855 2097.145 351.135 2097.425 ;
        RECT 351.475 2097.145 351.755 2097.425 ;
        RECT 352.095 2097.145 352.375 2097.425 ;
        RECT 350.235 2096.525 350.515 2096.805 ;
        RECT 350.855 2096.525 351.135 2096.805 ;
        RECT 351.475 2096.525 351.755 2096.805 ;
        RECT 352.095 2096.525 352.375 2096.805 ;
        RECT 350.235 2095.905 350.515 2096.185 ;
        RECT 350.855 2095.905 351.135 2096.185 ;
        RECT 351.475 2095.905 351.755 2096.185 ;
        RECT 352.095 2095.905 352.375 2096.185 ;
        RECT 350.235 2095.285 350.515 2095.565 ;
        RECT 350.855 2095.285 351.135 2095.565 ;
        RECT 351.475 2095.285 351.755 2095.565 ;
        RECT 352.095 2095.285 352.375 2095.565 ;
        RECT 350.235 2094.665 350.515 2094.945 ;
        RECT 350.855 2094.665 351.135 2094.945 ;
        RECT 351.475 2094.665 351.755 2094.945 ;
        RECT 352.095 2094.665 352.375 2094.945 ;
        RECT 350.235 2094.045 350.515 2094.325 ;
        RECT 350.855 2094.045 351.135 2094.325 ;
        RECT 351.475 2094.045 351.755 2094.325 ;
        RECT 352.095 2094.045 352.375 2094.325 ;
        RECT 350.235 2093.425 350.515 2093.705 ;
        RECT 350.855 2093.425 351.135 2093.705 ;
        RECT 351.475 2093.425 351.755 2093.705 ;
        RECT 352.095 2093.425 352.375 2093.705 ;
        RECT 350.235 2092.805 350.515 2093.085 ;
        RECT 350.855 2092.805 351.135 2093.085 ;
        RECT 351.475 2092.805 351.755 2093.085 ;
        RECT 352.095 2092.805 352.375 2093.085 ;
        RECT 350.235 2092.185 350.515 2092.465 ;
        RECT 350.855 2092.185 351.135 2092.465 ;
        RECT 351.475 2092.185 351.755 2092.465 ;
        RECT 352.095 2092.185 352.375 2092.465 ;
        RECT 350.235 2091.565 350.515 2091.845 ;
        RECT 350.855 2091.565 351.135 2091.845 ;
        RECT 351.475 2091.565 351.755 2091.845 ;
        RECT 352.095 2091.565 352.375 2091.845 ;
        RECT 350.235 2090.945 350.515 2091.225 ;
        RECT 350.855 2090.945 351.135 2091.225 ;
        RECT 351.475 2090.945 351.755 2091.225 ;
        RECT 352.095 2090.945 352.375 2091.225 ;
        RECT 350.235 2088.395 350.515 2088.675 ;
        RECT 350.855 2088.395 351.135 2088.675 ;
        RECT 351.475 2088.395 351.755 2088.675 ;
        RECT 352.095 2088.395 352.375 2088.675 ;
        RECT 350.235 2087.775 350.515 2088.055 ;
        RECT 350.855 2087.775 351.135 2088.055 ;
        RECT 351.475 2087.775 351.755 2088.055 ;
        RECT 352.095 2087.775 352.375 2088.055 ;
        RECT 350.235 2087.155 350.515 2087.435 ;
        RECT 350.855 2087.155 351.135 2087.435 ;
        RECT 351.475 2087.155 351.755 2087.435 ;
        RECT 352.095 2087.155 352.375 2087.435 ;
        RECT 350.235 2086.535 350.515 2086.815 ;
        RECT 350.855 2086.535 351.135 2086.815 ;
        RECT 351.475 2086.535 351.755 2086.815 ;
        RECT 352.095 2086.535 352.375 2086.815 ;
        RECT 350.235 2085.915 350.515 2086.195 ;
        RECT 350.855 2085.915 351.135 2086.195 ;
        RECT 351.475 2085.915 351.755 2086.195 ;
        RECT 352.095 2085.915 352.375 2086.195 ;
        RECT 350.235 2085.295 350.515 2085.575 ;
        RECT 350.855 2085.295 351.135 2085.575 ;
        RECT 351.475 2085.295 351.755 2085.575 ;
        RECT 352.095 2085.295 352.375 2085.575 ;
        RECT 350.235 2084.675 350.515 2084.955 ;
        RECT 350.855 2084.675 351.135 2084.955 ;
        RECT 351.475 2084.675 351.755 2084.955 ;
        RECT 352.095 2084.675 352.375 2084.955 ;
        RECT 350.235 2084.055 350.515 2084.335 ;
        RECT 350.855 2084.055 351.135 2084.335 ;
        RECT 351.475 2084.055 351.755 2084.335 ;
        RECT 352.095 2084.055 352.375 2084.335 ;
        RECT 350.235 2083.435 350.515 2083.715 ;
        RECT 350.855 2083.435 351.135 2083.715 ;
        RECT 351.475 2083.435 351.755 2083.715 ;
        RECT 352.095 2083.435 352.375 2083.715 ;
        RECT 350.235 2082.815 350.515 2083.095 ;
        RECT 350.855 2082.815 351.135 2083.095 ;
        RECT 351.475 2082.815 351.755 2083.095 ;
        RECT 352.095 2082.815 352.375 2083.095 ;
        RECT 350.235 2082.195 350.515 2082.475 ;
        RECT 350.855 2082.195 351.135 2082.475 ;
        RECT 351.475 2082.195 351.755 2082.475 ;
        RECT 352.095 2082.195 352.375 2082.475 ;
        RECT 350.235 2081.575 350.515 2081.855 ;
        RECT 350.855 2081.575 351.135 2081.855 ;
        RECT 351.475 2081.575 351.755 2081.855 ;
        RECT 352.095 2081.575 352.375 2081.855 ;
        RECT 350.235 2080.955 350.515 2081.235 ;
        RECT 350.855 2080.955 351.135 2081.235 ;
        RECT 351.475 2080.955 351.755 2081.235 ;
        RECT 352.095 2080.955 352.375 2081.235 ;
        RECT 350.235 2080.335 350.515 2080.615 ;
        RECT 350.855 2080.335 351.135 2080.615 ;
        RECT 351.475 2080.335 351.755 2080.615 ;
        RECT 352.095 2080.335 352.375 2080.615 ;
        RECT 350.235 2079.715 350.515 2079.995 ;
        RECT 350.855 2079.715 351.135 2079.995 ;
        RECT 351.475 2079.715 351.755 2079.995 ;
        RECT 352.095 2079.715 352.375 2079.995 ;
        RECT 350.235 2079.095 350.515 2079.375 ;
        RECT 350.855 2079.095 351.135 2079.375 ;
        RECT 351.475 2079.095 351.755 2079.375 ;
        RECT 352.095 2079.095 352.375 2079.375 ;
        RECT 350.235 2075.245 350.515 2075.525 ;
        RECT 350.855 2075.245 351.135 2075.525 ;
        RECT 351.475 2075.245 351.755 2075.525 ;
        RECT 352.095 2075.245 352.375 2075.525 ;
        RECT 350.235 2074.625 350.515 2074.905 ;
        RECT 350.855 2074.625 351.135 2074.905 ;
        RECT 351.475 2074.625 351.755 2074.905 ;
        RECT 352.095 2074.625 352.375 2074.905 ;
        RECT 350.235 2074.005 350.515 2074.285 ;
        RECT 350.855 2074.005 351.135 2074.285 ;
        RECT 351.475 2074.005 351.755 2074.285 ;
        RECT 352.095 2074.005 352.375 2074.285 ;
        RECT 350.235 2073.385 350.515 2073.665 ;
        RECT 350.855 2073.385 351.135 2073.665 ;
        RECT 351.475 2073.385 351.755 2073.665 ;
        RECT 352.095 2073.385 352.375 2073.665 ;
        RECT 350.235 2072.765 350.515 2073.045 ;
        RECT 350.855 2072.765 351.135 2073.045 ;
        RECT 351.475 2072.765 351.755 2073.045 ;
        RECT 352.095 2072.765 352.375 2073.045 ;
        RECT 350.235 2072.145 350.515 2072.425 ;
        RECT 350.855 2072.145 351.135 2072.425 ;
        RECT 351.475 2072.145 351.755 2072.425 ;
        RECT 352.095 2072.145 352.375 2072.425 ;
        RECT 350.235 2071.525 350.515 2071.805 ;
        RECT 350.855 2071.525 351.135 2071.805 ;
        RECT 351.475 2071.525 351.755 2071.805 ;
        RECT 352.095 2071.525 352.375 2071.805 ;
        RECT 350.235 2070.905 350.515 2071.185 ;
        RECT 350.855 2070.905 351.135 2071.185 ;
        RECT 351.475 2070.905 351.755 2071.185 ;
        RECT 352.095 2070.905 352.375 2071.185 ;
        RECT 350.235 2070.285 350.515 2070.565 ;
        RECT 350.855 2070.285 351.135 2070.565 ;
        RECT 351.475 2070.285 351.755 2070.565 ;
        RECT 352.095 2070.285 352.375 2070.565 ;
        RECT 350.235 2069.665 350.515 2069.945 ;
        RECT 350.855 2069.665 351.135 2069.945 ;
        RECT 351.475 2069.665 351.755 2069.945 ;
        RECT 352.095 2069.665 352.375 2069.945 ;
        RECT 350.235 2069.045 350.515 2069.325 ;
        RECT 350.855 2069.045 351.135 2069.325 ;
        RECT 351.475 2069.045 351.755 2069.325 ;
        RECT 352.095 2069.045 352.375 2069.325 ;
        RECT 350.235 2068.425 350.515 2068.705 ;
        RECT 350.855 2068.425 351.135 2068.705 ;
        RECT 351.475 2068.425 351.755 2068.705 ;
        RECT 352.095 2068.425 352.375 2068.705 ;
        RECT 350.235 2067.805 350.515 2068.085 ;
        RECT 350.855 2067.805 351.135 2068.085 ;
        RECT 351.475 2067.805 351.755 2068.085 ;
        RECT 352.095 2067.805 352.375 2068.085 ;
        RECT 350.235 2067.185 350.515 2067.465 ;
        RECT 350.855 2067.185 351.135 2067.465 ;
        RECT 351.475 2067.185 351.755 2067.465 ;
        RECT 352.095 2067.185 352.375 2067.465 ;
        RECT 350.235 2066.565 350.515 2066.845 ;
        RECT 350.855 2066.565 351.135 2066.845 ;
        RECT 351.475 2066.565 351.755 2066.845 ;
        RECT 352.095 2066.565 352.375 2066.845 ;
        RECT 3527.625 2023.155 3527.905 2023.435 ;
        RECT 3528.245 2023.155 3528.525 2023.435 ;
        RECT 3528.865 2023.155 3529.145 2023.435 ;
        RECT 3529.485 2023.155 3529.765 2023.435 ;
        RECT 3527.625 2022.535 3527.905 2022.815 ;
        RECT 3528.245 2022.535 3528.525 2022.815 ;
        RECT 3528.865 2022.535 3529.145 2022.815 ;
        RECT 3529.485 2022.535 3529.765 2022.815 ;
        RECT 3527.625 2021.915 3527.905 2022.195 ;
        RECT 3528.245 2021.915 3528.525 2022.195 ;
        RECT 3528.865 2021.915 3529.145 2022.195 ;
        RECT 3529.485 2021.915 3529.765 2022.195 ;
        RECT 3527.625 2021.295 3527.905 2021.575 ;
        RECT 3528.245 2021.295 3528.525 2021.575 ;
        RECT 3528.865 2021.295 3529.145 2021.575 ;
        RECT 3529.485 2021.295 3529.765 2021.575 ;
        RECT 3527.625 2020.675 3527.905 2020.955 ;
        RECT 3528.245 2020.675 3528.525 2020.955 ;
        RECT 3528.865 2020.675 3529.145 2020.955 ;
        RECT 3529.485 2020.675 3529.765 2020.955 ;
        RECT 3527.625 2020.055 3527.905 2020.335 ;
        RECT 3528.245 2020.055 3528.525 2020.335 ;
        RECT 3528.865 2020.055 3529.145 2020.335 ;
        RECT 3529.485 2020.055 3529.765 2020.335 ;
        RECT 3527.625 2019.435 3527.905 2019.715 ;
        RECT 3528.245 2019.435 3528.525 2019.715 ;
        RECT 3528.865 2019.435 3529.145 2019.715 ;
        RECT 3529.485 2019.435 3529.765 2019.715 ;
        RECT 3527.625 2018.815 3527.905 2019.095 ;
        RECT 3528.245 2018.815 3528.525 2019.095 ;
        RECT 3528.865 2018.815 3529.145 2019.095 ;
        RECT 3529.485 2018.815 3529.765 2019.095 ;
        RECT 3527.625 2018.195 3527.905 2018.475 ;
        RECT 3528.245 2018.195 3528.525 2018.475 ;
        RECT 3528.865 2018.195 3529.145 2018.475 ;
        RECT 3529.485 2018.195 3529.765 2018.475 ;
        RECT 3527.625 2017.575 3527.905 2017.855 ;
        RECT 3528.245 2017.575 3528.525 2017.855 ;
        RECT 3528.865 2017.575 3529.145 2017.855 ;
        RECT 3529.485 2017.575 3529.765 2017.855 ;
        RECT 3527.625 2016.955 3527.905 2017.235 ;
        RECT 3528.245 2016.955 3528.525 2017.235 ;
        RECT 3528.865 2016.955 3529.145 2017.235 ;
        RECT 3529.485 2016.955 3529.765 2017.235 ;
        RECT 3527.625 2016.335 3527.905 2016.615 ;
        RECT 3528.245 2016.335 3528.525 2016.615 ;
        RECT 3528.865 2016.335 3529.145 2016.615 ;
        RECT 3529.485 2016.335 3529.765 2016.615 ;
        RECT 3527.625 2015.715 3527.905 2015.995 ;
        RECT 3528.245 2015.715 3528.525 2015.995 ;
        RECT 3528.865 2015.715 3529.145 2015.995 ;
        RECT 3529.485 2015.715 3529.765 2015.995 ;
        RECT 3527.625 2015.095 3527.905 2015.375 ;
        RECT 3528.245 2015.095 3528.525 2015.375 ;
        RECT 3528.865 2015.095 3529.145 2015.375 ;
        RECT 3529.485 2015.095 3529.765 2015.375 ;
        RECT 3527.625 2014.475 3527.905 2014.755 ;
        RECT 3528.245 2014.475 3528.525 2014.755 ;
        RECT 3528.865 2014.475 3529.145 2014.755 ;
        RECT 3529.485 2014.475 3529.765 2014.755 ;
        RECT 3527.625 2010.625 3527.905 2010.905 ;
        RECT 3528.245 2010.625 3528.525 2010.905 ;
        RECT 3528.865 2010.625 3529.145 2010.905 ;
        RECT 3529.485 2010.625 3529.765 2010.905 ;
        RECT 3527.625 2010.005 3527.905 2010.285 ;
        RECT 3528.245 2010.005 3528.525 2010.285 ;
        RECT 3528.865 2010.005 3529.145 2010.285 ;
        RECT 3529.485 2010.005 3529.765 2010.285 ;
        RECT 3527.625 2009.385 3527.905 2009.665 ;
        RECT 3528.245 2009.385 3528.525 2009.665 ;
        RECT 3528.865 2009.385 3529.145 2009.665 ;
        RECT 3529.485 2009.385 3529.765 2009.665 ;
        RECT 3527.625 2008.765 3527.905 2009.045 ;
        RECT 3528.245 2008.765 3528.525 2009.045 ;
        RECT 3528.865 2008.765 3529.145 2009.045 ;
        RECT 3529.485 2008.765 3529.765 2009.045 ;
        RECT 3527.625 2008.145 3527.905 2008.425 ;
        RECT 3528.245 2008.145 3528.525 2008.425 ;
        RECT 3528.865 2008.145 3529.145 2008.425 ;
        RECT 3529.485 2008.145 3529.765 2008.425 ;
        RECT 3527.625 2007.525 3527.905 2007.805 ;
        RECT 3528.245 2007.525 3528.525 2007.805 ;
        RECT 3528.865 2007.525 3529.145 2007.805 ;
        RECT 3529.485 2007.525 3529.765 2007.805 ;
        RECT 3527.625 2006.905 3527.905 2007.185 ;
        RECT 3528.245 2006.905 3528.525 2007.185 ;
        RECT 3528.865 2006.905 3529.145 2007.185 ;
        RECT 3529.485 2006.905 3529.765 2007.185 ;
        RECT 3527.625 2006.285 3527.905 2006.565 ;
        RECT 3528.245 2006.285 3528.525 2006.565 ;
        RECT 3528.865 2006.285 3529.145 2006.565 ;
        RECT 3529.485 2006.285 3529.765 2006.565 ;
        RECT 3527.625 2005.665 3527.905 2005.945 ;
        RECT 3528.245 2005.665 3528.525 2005.945 ;
        RECT 3528.865 2005.665 3529.145 2005.945 ;
        RECT 3529.485 2005.665 3529.765 2005.945 ;
        RECT 3527.625 2005.045 3527.905 2005.325 ;
        RECT 3528.245 2005.045 3528.525 2005.325 ;
        RECT 3528.865 2005.045 3529.145 2005.325 ;
        RECT 3529.485 2005.045 3529.765 2005.325 ;
        RECT 3527.625 2004.425 3527.905 2004.705 ;
        RECT 3528.245 2004.425 3528.525 2004.705 ;
        RECT 3528.865 2004.425 3529.145 2004.705 ;
        RECT 3529.485 2004.425 3529.765 2004.705 ;
        RECT 3527.625 2003.805 3527.905 2004.085 ;
        RECT 3528.245 2003.805 3528.525 2004.085 ;
        RECT 3528.865 2003.805 3529.145 2004.085 ;
        RECT 3529.485 2003.805 3529.765 2004.085 ;
        RECT 3527.625 2003.185 3527.905 2003.465 ;
        RECT 3528.245 2003.185 3528.525 2003.465 ;
        RECT 3528.865 2003.185 3529.145 2003.465 ;
        RECT 3529.485 2003.185 3529.765 2003.465 ;
        RECT 3527.625 2002.565 3527.905 2002.845 ;
        RECT 3528.245 2002.565 3528.525 2002.845 ;
        RECT 3528.865 2002.565 3529.145 2002.845 ;
        RECT 3529.485 2002.565 3529.765 2002.845 ;
        RECT 3527.625 2001.945 3527.905 2002.225 ;
        RECT 3528.245 2001.945 3528.525 2002.225 ;
        RECT 3528.865 2001.945 3529.145 2002.225 ;
        RECT 3529.485 2001.945 3529.765 2002.225 ;
        RECT 3527.625 2001.325 3527.905 2001.605 ;
        RECT 3528.245 2001.325 3528.525 2001.605 ;
        RECT 3528.865 2001.325 3529.145 2001.605 ;
        RECT 3529.485 2001.325 3529.765 2001.605 ;
        RECT 3527.625 1998.775 3527.905 1999.055 ;
        RECT 3528.245 1998.775 3528.525 1999.055 ;
        RECT 3528.865 1998.775 3529.145 1999.055 ;
        RECT 3529.485 1998.775 3529.765 1999.055 ;
        RECT 3527.625 1998.155 3527.905 1998.435 ;
        RECT 3528.245 1998.155 3528.525 1998.435 ;
        RECT 3528.865 1998.155 3529.145 1998.435 ;
        RECT 3529.485 1998.155 3529.765 1998.435 ;
        RECT 3527.625 1997.535 3527.905 1997.815 ;
        RECT 3528.245 1997.535 3528.525 1997.815 ;
        RECT 3528.865 1997.535 3529.145 1997.815 ;
        RECT 3529.485 1997.535 3529.765 1997.815 ;
        RECT 3527.625 1996.915 3527.905 1997.195 ;
        RECT 3528.245 1996.915 3528.525 1997.195 ;
        RECT 3528.865 1996.915 3529.145 1997.195 ;
        RECT 3529.485 1996.915 3529.765 1997.195 ;
        RECT 3527.625 1996.295 3527.905 1996.575 ;
        RECT 3528.245 1996.295 3528.525 1996.575 ;
        RECT 3528.865 1996.295 3529.145 1996.575 ;
        RECT 3529.485 1996.295 3529.765 1996.575 ;
        RECT 3527.625 1995.675 3527.905 1995.955 ;
        RECT 3528.245 1995.675 3528.525 1995.955 ;
        RECT 3528.865 1995.675 3529.145 1995.955 ;
        RECT 3529.485 1995.675 3529.765 1995.955 ;
        RECT 3527.625 1995.055 3527.905 1995.335 ;
        RECT 3528.245 1995.055 3528.525 1995.335 ;
        RECT 3528.865 1995.055 3529.145 1995.335 ;
        RECT 3529.485 1995.055 3529.765 1995.335 ;
        RECT 3527.625 1994.435 3527.905 1994.715 ;
        RECT 3528.245 1994.435 3528.525 1994.715 ;
        RECT 3528.865 1994.435 3529.145 1994.715 ;
        RECT 3529.485 1994.435 3529.765 1994.715 ;
        RECT 3527.625 1993.815 3527.905 1994.095 ;
        RECT 3528.245 1993.815 3528.525 1994.095 ;
        RECT 3528.865 1993.815 3529.145 1994.095 ;
        RECT 3529.485 1993.815 3529.765 1994.095 ;
        RECT 3527.625 1993.195 3527.905 1993.475 ;
        RECT 3528.245 1993.195 3528.525 1993.475 ;
        RECT 3528.865 1993.195 3529.145 1993.475 ;
        RECT 3529.485 1993.195 3529.765 1993.475 ;
        RECT 3527.625 1992.575 3527.905 1992.855 ;
        RECT 3528.245 1992.575 3528.525 1992.855 ;
        RECT 3528.865 1992.575 3529.145 1992.855 ;
        RECT 3529.485 1992.575 3529.765 1992.855 ;
        RECT 3527.625 1991.955 3527.905 1992.235 ;
        RECT 3528.245 1991.955 3528.525 1992.235 ;
        RECT 3528.865 1991.955 3529.145 1992.235 ;
        RECT 3529.485 1991.955 3529.765 1992.235 ;
        RECT 3527.625 1991.335 3527.905 1991.615 ;
        RECT 3528.245 1991.335 3528.525 1991.615 ;
        RECT 3528.865 1991.335 3529.145 1991.615 ;
        RECT 3529.485 1991.335 3529.765 1991.615 ;
        RECT 3527.625 1990.715 3527.905 1990.995 ;
        RECT 3528.245 1990.715 3528.525 1990.995 ;
        RECT 3528.865 1990.715 3529.145 1990.995 ;
        RECT 3529.485 1990.715 3529.765 1990.995 ;
        RECT 3527.625 1990.095 3527.905 1990.375 ;
        RECT 3528.245 1990.095 3528.525 1990.375 ;
        RECT 3528.865 1990.095 3529.145 1990.375 ;
        RECT 3529.485 1990.095 3529.765 1990.375 ;
        RECT 3527.625 1989.475 3527.905 1989.755 ;
        RECT 3528.245 1989.475 3528.525 1989.755 ;
        RECT 3528.865 1989.475 3529.145 1989.755 ;
        RECT 3529.485 1989.475 3529.765 1989.755 ;
        RECT 3527.625 1985.245 3527.905 1985.525 ;
        RECT 3528.245 1985.245 3528.525 1985.525 ;
        RECT 3528.865 1985.245 3529.145 1985.525 ;
        RECT 3529.485 1985.245 3529.765 1985.525 ;
        RECT 3527.625 1984.625 3527.905 1984.905 ;
        RECT 3528.245 1984.625 3528.525 1984.905 ;
        RECT 3528.865 1984.625 3529.145 1984.905 ;
        RECT 3529.485 1984.625 3529.765 1984.905 ;
        RECT 3527.625 1984.005 3527.905 1984.285 ;
        RECT 3528.245 1984.005 3528.525 1984.285 ;
        RECT 3528.865 1984.005 3529.145 1984.285 ;
        RECT 3529.485 1984.005 3529.765 1984.285 ;
        RECT 3527.625 1983.385 3527.905 1983.665 ;
        RECT 3528.245 1983.385 3528.525 1983.665 ;
        RECT 3528.865 1983.385 3529.145 1983.665 ;
        RECT 3529.485 1983.385 3529.765 1983.665 ;
        RECT 3527.625 1982.765 3527.905 1983.045 ;
        RECT 3528.245 1982.765 3528.525 1983.045 ;
        RECT 3528.865 1982.765 3529.145 1983.045 ;
        RECT 3529.485 1982.765 3529.765 1983.045 ;
        RECT 3527.625 1982.145 3527.905 1982.425 ;
        RECT 3528.245 1982.145 3528.525 1982.425 ;
        RECT 3528.865 1982.145 3529.145 1982.425 ;
        RECT 3529.485 1982.145 3529.765 1982.425 ;
        RECT 3527.625 1981.525 3527.905 1981.805 ;
        RECT 3528.245 1981.525 3528.525 1981.805 ;
        RECT 3528.865 1981.525 3529.145 1981.805 ;
        RECT 3529.485 1981.525 3529.765 1981.805 ;
        RECT 3527.625 1980.905 3527.905 1981.185 ;
        RECT 3528.245 1980.905 3528.525 1981.185 ;
        RECT 3528.865 1980.905 3529.145 1981.185 ;
        RECT 3529.485 1980.905 3529.765 1981.185 ;
        RECT 3527.625 1980.285 3527.905 1980.565 ;
        RECT 3528.245 1980.285 3528.525 1980.565 ;
        RECT 3528.865 1980.285 3529.145 1980.565 ;
        RECT 3529.485 1980.285 3529.765 1980.565 ;
        RECT 3527.625 1979.665 3527.905 1979.945 ;
        RECT 3528.245 1979.665 3528.525 1979.945 ;
        RECT 3528.865 1979.665 3529.145 1979.945 ;
        RECT 3529.485 1979.665 3529.765 1979.945 ;
        RECT 3527.625 1979.045 3527.905 1979.325 ;
        RECT 3528.245 1979.045 3528.525 1979.325 ;
        RECT 3528.865 1979.045 3529.145 1979.325 ;
        RECT 3529.485 1979.045 3529.765 1979.325 ;
        RECT 3527.625 1978.425 3527.905 1978.705 ;
        RECT 3528.245 1978.425 3528.525 1978.705 ;
        RECT 3528.865 1978.425 3529.145 1978.705 ;
        RECT 3529.485 1978.425 3529.765 1978.705 ;
        RECT 3527.625 1977.805 3527.905 1978.085 ;
        RECT 3528.245 1977.805 3528.525 1978.085 ;
        RECT 3528.865 1977.805 3529.145 1978.085 ;
        RECT 3529.485 1977.805 3529.765 1978.085 ;
        RECT 3527.625 1977.185 3527.905 1977.465 ;
        RECT 3528.245 1977.185 3528.525 1977.465 ;
        RECT 3528.865 1977.185 3529.145 1977.465 ;
        RECT 3529.485 1977.185 3529.765 1977.465 ;
        RECT 3527.625 1976.565 3527.905 1976.845 ;
        RECT 3528.245 1976.565 3528.525 1976.845 ;
        RECT 3528.865 1976.565 3529.145 1976.845 ;
        RECT 3529.485 1976.565 3529.765 1976.845 ;
        RECT 3527.625 1975.945 3527.905 1976.225 ;
        RECT 3528.245 1975.945 3528.525 1976.225 ;
        RECT 3528.865 1975.945 3529.145 1976.225 ;
        RECT 3529.485 1975.945 3529.765 1976.225 ;
        RECT 3527.625 1973.395 3527.905 1973.675 ;
        RECT 3528.245 1973.395 3528.525 1973.675 ;
        RECT 3528.865 1973.395 3529.145 1973.675 ;
        RECT 3529.485 1973.395 3529.765 1973.675 ;
        RECT 3527.625 1972.775 3527.905 1973.055 ;
        RECT 3528.245 1972.775 3528.525 1973.055 ;
        RECT 3528.865 1972.775 3529.145 1973.055 ;
        RECT 3529.485 1972.775 3529.765 1973.055 ;
        RECT 3527.625 1972.155 3527.905 1972.435 ;
        RECT 3528.245 1972.155 3528.525 1972.435 ;
        RECT 3528.865 1972.155 3529.145 1972.435 ;
        RECT 3529.485 1972.155 3529.765 1972.435 ;
        RECT 3527.625 1971.535 3527.905 1971.815 ;
        RECT 3528.245 1971.535 3528.525 1971.815 ;
        RECT 3528.865 1971.535 3529.145 1971.815 ;
        RECT 3529.485 1971.535 3529.765 1971.815 ;
        RECT 3527.625 1970.915 3527.905 1971.195 ;
        RECT 3528.245 1970.915 3528.525 1971.195 ;
        RECT 3528.865 1970.915 3529.145 1971.195 ;
        RECT 3529.485 1970.915 3529.765 1971.195 ;
        RECT 3527.625 1970.295 3527.905 1970.575 ;
        RECT 3528.245 1970.295 3528.525 1970.575 ;
        RECT 3528.865 1970.295 3529.145 1970.575 ;
        RECT 3529.485 1970.295 3529.765 1970.575 ;
        RECT 3527.625 1969.675 3527.905 1969.955 ;
        RECT 3528.245 1969.675 3528.525 1969.955 ;
        RECT 3528.865 1969.675 3529.145 1969.955 ;
        RECT 3529.485 1969.675 3529.765 1969.955 ;
        RECT 3527.625 1969.055 3527.905 1969.335 ;
        RECT 3528.245 1969.055 3528.525 1969.335 ;
        RECT 3528.865 1969.055 3529.145 1969.335 ;
        RECT 3529.485 1969.055 3529.765 1969.335 ;
        RECT 3527.625 1968.435 3527.905 1968.715 ;
        RECT 3528.245 1968.435 3528.525 1968.715 ;
        RECT 3528.865 1968.435 3529.145 1968.715 ;
        RECT 3529.485 1968.435 3529.765 1968.715 ;
        RECT 3527.625 1967.815 3527.905 1968.095 ;
        RECT 3528.245 1967.815 3528.525 1968.095 ;
        RECT 3528.865 1967.815 3529.145 1968.095 ;
        RECT 3529.485 1967.815 3529.765 1968.095 ;
        RECT 3527.625 1967.195 3527.905 1967.475 ;
        RECT 3528.245 1967.195 3528.525 1967.475 ;
        RECT 3528.865 1967.195 3529.145 1967.475 ;
        RECT 3529.485 1967.195 3529.765 1967.475 ;
        RECT 3527.625 1966.575 3527.905 1966.855 ;
        RECT 3528.245 1966.575 3528.525 1966.855 ;
        RECT 3528.865 1966.575 3529.145 1966.855 ;
        RECT 3529.485 1966.575 3529.765 1966.855 ;
        RECT 3527.625 1965.955 3527.905 1966.235 ;
        RECT 3528.245 1965.955 3528.525 1966.235 ;
        RECT 3528.865 1965.955 3529.145 1966.235 ;
        RECT 3529.485 1965.955 3529.765 1966.235 ;
        RECT 3527.625 1965.335 3527.905 1965.615 ;
        RECT 3528.245 1965.335 3528.525 1965.615 ;
        RECT 3528.865 1965.335 3529.145 1965.615 ;
        RECT 3529.485 1965.335 3529.765 1965.615 ;
        RECT 3527.625 1964.715 3527.905 1964.995 ;
        RECT 3528.245 1964.715 3528.525 1964.995 ;
        RECT 3528.865 1964.715 3529.145 1964.995 ;
        RECT 3529.485 1964.715 3529.765 1964.995 ;
        RECT 3527.625 1964.095 3527.905 1964.375 ;
        RECT 3528.245 1964.095 3528.525 1964.375 ;
        RECT 3528.865 1964.095 3529.145 1964.375 ;
        RECT 3529.485 1964.095 3529.765 1964.375 ;
        RECT 3527.625 1960.375 3527.905 1960.655 ;
        RECT 3528.245 1960.375 3528.525 1960.655 ;
        RECT 3528.865 1960.375 3529.145 1960.655 ;
        RECT 3529.485 1960.375 3529.765 1960.655 ;
        RECT 3527.625 1959.755 3527.905 1960.035 ;
        RECT 3528.245 1959.755 3528.525 1960.035 ;
        RECT 3528.865 1959.755 3529.145 1960.035 ;
        RECT 3529.485 1959.755 3529.765 1960.035 ;
        RECT 3527.625 1959.135 3527.905 1959.415 ;
        RECT 3528.245 1959.135 3528.525 1959.415 ;
        RECT 3528.865 1959.135 3529.145 1959.415 ;
        RECT 3529.485 1959.135 3529.765 1959.415 ;
        RECT 3527.625 1958.515 3527.905 1958.795 ;
        RECT 3528.245 1958.515 3528.525 1958.795 ;
        RECT 3528.865 1958.515 3529.145 1958.795 ;
        RECT 3529.485 1958.515 3529.765 1958.795 ;
        RECT 3527.625 1957.895 3527.905 1958.175 ;
        RECT 3528.245 1957.895 3528.525 1958.175 ;
        RECT 3528.865 1957.895 3529.145 1958.175 ;
        RECT 3529.485 1957.895 3529.765 1958.175 ;
        RECT 3527.625 1957.275 3527.905 1957.555 ;
        RECT 3528.245 1957.275 3528.525 1957.555 ;
        RECT 3528.865 1957.275 3529.145 1957.555 ;
        RECT 3529.485 1957.275 3529.765 1957.555 ;
        RECT 3527.625 1956.655 3527.905 1956.935 ;
        RECT 3528.245 1956.655 3528.525 1956.935 ;
        RECT 3528.865 1956.655 3529.145 1956.935 ;
        RECT 3529.485 1956.655 3529.765 1956.935 ;
        RECT 3527.625 1956.035 3527.905 1956.315 ;
        RECT 3528.245 1956.035 3528.525 1956.315 ;
        RECT 3528.865 1956.035 3529.145 1956.315 ;
        RECT 3529.485 1956.035 3529.765 1956.315 ;
        RECT 3527.625 1955.415 3527.905 1955.695 ;
        RECT 3528.245 1955.415 3528.525 1955.695 ;
        RECT 3528.865 1955.415 3529.145 1955.695 ;
        RECT 3529.485 1955.415 3529.765 1955.695 ;
        RECT 3527.625 1954.795 3527.905 1955.075 ;
        RECT 3528.245 1954.795 3528.525 1955.075 ;
        RECT 3528.865 1954.795 3529.145 1955.075 ;
        RECT 3529.485 1954.795 3529.765 1955.075 ;
        RECT 3527.625 1954.175 3527.905 1954.455 ;
        RECT 3528.245 1954.175 3528.525 1954.455 ;
        RECT 3528.865 1954.175 3529.145 1954.455 ;
        RECT 3529.485 1954.175 3529.765 1954.455 ;
        RECT 3527.625 1953.555 3527.905 1953.835 ;
        RECT 3528.245 1953.555 3528.525 1953.835 ;
        RECT 3528.865 1953.555 3529.145 1953.835 ;
        RECT 3529.485 1953.555 3529.765 1953.835 ;
        RECT 3527.625 1952.935 3527.905 1953.215 ;
        RECT 3528.245 1952.935 3528.525 1953.215 ;
        RECT 3528.865 1952.935 3529.145 1953.215 ;
        RECT 3529.485 1952.935 3529.765 1953.215 ;
        RECT 3527.625 1952.315 3527.905 1952.595 ;
        RECT 3528.245 1952.315 3528.525 1952.595 ;
        RECT 3528.865 1952.315 3529.145 1952.595 ;
        RECT 3529.485 1952.315 3529.765 1952.595 ;
        RECT 3527.625 1951.695 3527.905 1951.975 ;
        RECT 3528.245 1951.695 3528.525 1951.975 ;
        RECT 3528.865 1951.695 3529.145 1951.975 ;
        RECT 3529.485 1951.695 3529.765 1951.975 ;
        RECT 350.235 703.025 350.515 703.305 ;
        RECT 350.855 703.025 351.135 703.305 ;
        RECT 351.475 703.025 351.755 703.305 ;
        RECT 352.095 703.025 352.375 703.305 ;
        RECT 350.235 702.405 350.515 702.685 ;
        RECT 350.855 702.405 351.135 702.685 ;
        RECT 351.475 702.405 351.755 702.685 ;
        RECT 352.095 702.405 352.375 702.685 ;
        RECT 350.235 701.785 350.515 702.065 ;
        RECT 350.855 701.785 351.135 702.065 ;
        RECT 351.475 701.785 351.755 702.065 ;
        RECT 352.095 701.785 352.375 702.065 ;
        RECT 350.235 701.165 350.515 701.445 ;
        RECT 350.855 701.165 351.135 701.445 ;
        RECT 351.475 701.165 351.755 701.445 ;
        RECT 352.095 701.165 352.375 701.445 ;
        RECT 350.235 700.545 350.515 700.825 ;
        RECT 350.855 700.545 351.135 700.825 ;
        RECT 351.475 700.545 351.755 700.825 ;
        RECT 352.095 700.545 352.375 700.825 ;
        RECT 350.235 699.925 350.515 700.205 ;
        RECT 350.855 699.925 351.135 700.205 ;
        RECT 351.475 699.925 351.755 700.205 ;
        RECT 352.095 699.925 352.375 700.205 ;
        RECT 350.235 699.305 350.515 699.585 ;
        RECT 350.855 699.305 351.135 699.585 ;
        RECT 351.475 699.305 351.755 699.585 ;
        RECT 352.095 699.305 352.375 699.585 ;
        RECT 350.235 698.685 350.515 698.965 ;
        RECT 350.855 698.685 351.135 698.965 ;
        RECT 351.475 698.685 351.755 698.965 ;
        RECT 352.095 698.685 352.375 698.965 ;
        RECT 350.235 698.065 350.515 698.345 ;
        RECT 350.855 698.065 351.135 698.345 ;
        RECT 351.475 698.065 351.755 698.345 ;
        RECT 352.095 698.065 352.375 698.345 ;
        RECT 350.235 697.445 350.515 697.725 ;
        RECT 350.855 697.445 351.135 697.725 ;
        RECT 351.475 697.445 351.755 697.725 ;
        RECT 352.095 697.445 352.375 697.725 ;
        RECT 350.235 696.825 350.515 697.105 ;
        RECT 350.855 696.825 351.135 697.105 ;
        RECT 351.475 696.825 351.755 697.105 ;
        RECT 352.095 696.825 352.375 697.105 ;
        RECT 350.235 696.205 350.515 696.485 ;
        RECT 350.855 696.205 351.135 696.485 ;
        RECT 351.475 696.205 351.755 696.485 ;
        RECT 352.095 696.205 352.375 696.485 ;
        RECT 350.235 695.585 350.515 695.865 ;
        RECT 350.855 695.585 351.135 695.865 ;
        RECT 351.475 695.585 351.755 695.865 ;
        RECT 352.095 695.585 352.375 695.865 ;
        RECT 350.235 694.965 350.515 695.245 ;
        RECT 350.855 694.965 351.135 695.245 ;
        RECT 351.475 694.965 351.755 695.245 ;
        RECT 352.095 694.965 352.375 695.245 ;
        RECT 350.235 694.345 350.515 694.625 ;
        RECT 350.855 694.345 351.135 694.625 ;
        RECT 351.475 694.345 351.755 694.625 ;
        RECT 352.095 694.345 352.375 694.625 ;
        RECT 350.235 690.625 350.515 690.905 ;
        RECT 350.855 690.625 351.135 690.905 ;
        RECT 351.475 690.625 351.755 690.905 ;
        RECT 352.095 690.625 352.375 690.905 ;
        RECT 350.235 690.005 350.515 690.285 ;
        RECT 350.855 690.005 351.135 690.285 ;
        RECT 351.475 690.005 351.755 690.285 ;
        RECT 352.095 690.005 352.375 690.285 ;
        RECT 350.235 689.385 350.515 689.665 ;
        RECT 350.855 689.385 351.135 689.665 ;
        RECT 351.475 689.385 351.755 689.665 ;
        RECT 352.095 689.385 352.375 689.665 ;
        RECT 350.235 688.765 350.515 689.045 ;
        RECT 350.855 688.765 351.135 689.045 ;
        RECT 351.475 688.765 351.755 689.045 ;
        RECT 352.095 688.765 352.375 689.045 ;
        RECT 350.235 688.145 350.515 688.425 ;
        RECT 350.855 688.145 351.135 688.425 ;
        RECT 351.475 688.145 351.755 688.425 ;
        RECT 352.095 688.145 352.375 688.425 ;
        RECT 350.235 687.525 350.515 687.805 ;
        RECT 350.855 687.525 351.135 687.805 ;
        RECT 351.475 687.525 351.755 687.805 ;
        RECT 352.095 687.525 352.375 687.805 ;
        RECT 350.235 686.905 350.515 687.185 ;
        RECT 350.855 686.905 351.135 687.185 ;
        RECT 351.475 686.905 351.755 687.185 ;
        RECT 352.095 686.905 352.375 687.185 ;
        RECT 350.235 686.285 350.515 686.565 ;
        RECT 350.855 686.285 351.135 686.565 ;
        RECT 351.475 686.285 351.755 686.565 ;
        RECT 352.095 686.285 352.375 686.565 ;
        RECT 350.235 685.665 350.515 685.945 ;
        RECT 350.855 685.665 351.135 685.945 ;
        RECT 351.475 685.665 351.755 685.945 ;
        RECT 352.095 685.665 352.375 685.945 ;
        RECT 350.235 685.045 350.515 685.325 ;
        RECT 350.855 685.045 351.135 685.325 ;
        RECT 351.475 685.045 351.755 685.325 ;
        RECT 352.095 685.045 352.375 685.325 ;
        RECT 350.235 684.425 350.515 684.705 ;
        RECT 350.855 684.425 351.135 684.705 ;
        RECT 351.475 684.425 351.755 684.705 ;
        RECT 352.095 684.425 352.375 684.705 ;
        RECT 350.235 683.805 350.515 684.085 ;
        RECT 350.855 683.805 351.135 684.085 ;
        RECT 351.475 683.805 351.755 684.085 ;
        RECT 352.095 683.805 352.375 684.085 ;
        RECT 350.235 683.185 350.515 683.465 ;
        RECT 350.855 683.185 351.135 683.465 ;
        RECT 351.475 683.185 351.755 683.465 ;
        RECT 352.095 683.185 352.375 683.465 ;
        RECT 350.235 682.565 350.515 682.845 ;
        RECT 350.855 682.565 351.135 682.845 ;
        RECT 351.475 682.565 351.755 682.845 ;
        RECT 352.095 682.565 352.375 682.845 ;
        RECT 350.235 681.945 350.515 682.225 ;
        RECT 350.855 681.945 351.135 682.225 ;
        RECT 351.475 681.945 351.755 682.225 ;
        RECT 352.095 681.945 352.375 682.225 ;
        RECT 350.235 681.325 350.515 681.605 ;
        RECT 350.855 681.325 351.135 681.605 ;
        RECT 351.475 681.325 351.755 681.605 ;
        RECT 352.095 681.325 352.375 681.605 ;
        RECT 350.235 678.775 350.515 679.055 ;
        RECT 350.855 678.775 351.135 679.055 ;
        RECT 351.475 678.775 351.755 679.055 ;
        RECT 352.095 678.775 352.375 679.055 ;
        RECT 350.235 678.155 350.515 678.435 ;
        RECT 350.855 678.155 351.135 678.435 ;
        RECT 351.475 678.155 351.755 678.435 ;
        RECT 352.095 678.155 352.375 678.435 ;
        RECT 350.235 677.535 350.515 677.815 ;
        RECT 350.855 677.535 351.135 677.815 ;
        RECT 351.475 677.535 351.755 677.815 ;
        RECT 352.095 677.535 352.375 677.815 ;
        RECT 350.235 676.915 350.515 677.195 ;
        RECT 350.855 676.915 351.135 677.195 ;
        RECT 351.475 676.915 351.755 677.195 ;
        RECT 352.095 676.915 352.375 677.195 ;
        RECT 350.235 676.295 350.515 676.575 ;
        RECT 350.855 676.295 351.135 676.575 ;
        RECT 351.475 676.295 351.755 676.575 ;
        RECT 352.095 676.295 352.375 676.575 ;
        RECT 350.235 675.675 350.515 675.955 ;
        RECT 350.855 675.675 351.135 675.955 ;
        RECT 351.475 675.675 351.755 675.955 ;
        RECT 352.095 675.675 352.375 675.955 ;
        RECT 350.235 675.055 350.515 675.335 ;
        RECT 350.855 675.055 351.135 675.335 ;
        RECT 351.475 675.055 351.755 675.335 ;
        RECT 352.095 675.055 352.375 675.335 ;
        RECT 350.235 674.435 350.515 674.715 ;
        RECT 350.855 674.435 351.135 674.715 ;
        RECT 351.475 674.435 351.755 674.715 ;
        RECT 352.095 674.435 352.375 674.715 ;
        RECT 350.235 673.815 350.515 674.095 ;
        RECT 350.855 673.815 351.135 674.095 ;
        RECT 351.475 673.815 351.755 674.095 ;
        RECT 352.095 673.815 352.375 674.095 ;
        RECT 350.235 673.195 350.515 673.475 ;
        RECT 350.855 673.195 351.135 673.475 ;
        RECT 351.475 673.195 351.755 673.475 ;
        RECT 352.095 673.195 352.375 673.475 ;
        RECT 350.235 672.575 350.515 672.855 ;
        RECT 350.855 672.575 351.135 672.855 ;
        RECT 351.475 672.575 351.755 672.855 ;
        RECT 352.095 672.575 352.375 672.855 ;
        RECT 350.235 671.955 350.515 672.235 ;
        RECT 350.855 671.955 351.135 672.235 ;
        RECT 351.475 671.955 351.755 672.235 ;
        RECT 352.095 671.955 352.375 672.235 ;
        RECT 350.235 671.335 350.515 671.615 ;
        RECT 350.855 671.335 351.135 671.615 ;
        RECT 351.475 671.335 351.755 671.615 ;
        RECT 352.095 671.335 352.375 671.615 ;
        RECT 350.235 670.715 350.515 670.995 ;
        RECT 350.855 670.715 351.135 670.995 ;
        RECT 351.475 670.715 351.755 670.995 ;
        RECT 352.095 670.715 352.375 670.995 ;
        RECT 350.235 670.095 350.515 670.375 ;
        RECT 350.855 670.095 351.135 670.375 ;
        RECT 351.475 670.095 351.755 670.375 ;
        RECT 352.095 670.095 352.375 670.375 ;
        RECT 350.235 669.475 350.515 669.755 ;
        RECT 350.855 669.475 351.135 669.755 ;
        RECT 351.475 669.475 351.755 669.755 ;
        RECT 352.095 669.475 352.375 669.755 ;
        RECT 350.235 665.245 350.515 665.525 ;
        RECT 350.855 665.245 351.135 665.525 ;
        RECT 351.475 665.245 351.755 665.525 ;
        RECT 352.095 665.245 352.375 665.525 ;
        RECT 350.235 664.625 350.515 664.905 ;
        RECT 350.855 664.625 351.135 664.905 ;
        RECT 351.475 664.625 351.755 664.905 ;
        RECT 352.095 664.625 352.375 664.905 ;
        RECT 350.235 664.005 350.515 664.285 ;
        RECT 350.855 664.005 351.135 664.285 ;
        RECT 351.475 664.005 351.755 664.285 ;
        RECT 352.095 664.005 352.375 664.285 ;
        RECT 350.235 663.385 350.515 663.665 ;
        RECT 350.855 663.385 351.135 663.665 ;
        RECT 351.475 663.385 351.755 663.665 ;
        RECT 352.095 663.385 352.375 663.665 ;
        RECT 350.235 662.765 350.515 663.045 ;
        RECT 350.855 662.765 351.135 663.045 ;
        RECT 351.475 662.765 351.755 663.045 ;
        RECT 352.095 662.765 352.375 663.045 ;
        RECT 350.235 662.145 350.515 662.425 ;
        RECT 350.855 662.145 351.135 662.425 ;
        RECT 351.475 662.145 351.755 662.425 ;
        RECT 352.095 662.145 352.375 662.425 ;
        RECT 350.235 661.525 350.515 661.805 ;
        RECT 350.855 661.525 351.135 661.805 ;
        RECT 351.475 661.525 351.755 661.805 ;
        RECT 352.095 661.525 352.375 661.805 ;
        RECT 350.235 660.905 350.515 661.185 ;
        RECT 350.855 660.905 351.135 661.185 ;
        RECT 351.475 660.905 351.755 661.185 ;
        RECT 352.095 660.905 352.375 661.185 ;
        RECT 350.235 660.285 350.515 660.565 ;
        RECT 350.855 660.285 351.135 660.565 ;
        RECT 351.475 660.285 351.755 660.565 ;
        RECT 352.095 660.285 352.375 660.565 ;
        RECT 350.235 659.665 350.515 659.945 ;
        RECT 350.855 659.665 351.135 659.945 ;
        RECT 351.475 659.665 351.755 659.945 ;
        RECT 352.095 659.665 352.375 659.945 ;
        RECT 350.235 659.045 350.515 659.325 ;
        RECT 350.855 659.045 351.135 659.325 ;
        RECT 351.475 659.045 351.755 659.325 ;
        RECT 352.095 659.045 352.375 659.325 ;
        RECT 350.235 658.425 350.515 658.705 ;
        RECT 350.855 658.425 351.135 658.705 ;
        RECT 351.475 658.425 351.755 658.705 ;
        RECT 352.095 658.425 352.375 658.705 ;
        RECT 350.235 657.805 350.515 658.085 ;
        RECT 350.855 657.805 351.135 658.085 ;
        RECT 351.475 657.805 351.755 658.085 ;
        RECT 352.095 657.805 352.375 658.085 ;
        RECT 350.235 657.185 350.515 657.465 ;
        RECT 350.855 657.185 351.135 657.465 ;
        RECT 351.475 657.185 351.755 657.465 ;
        RECT 352.095 657.185 352.375 657.465 ;
        RECT 350.235 656.565 350.515 656.845 ;
        RECT 350.855 656.565 351.135 656.845 ;
        RECT 351.475 656.565 351.755 656.845 ;
        RECT 352.095 656.565 352.375 656.845 ;
        RECT 350.235 655.945 350.515 656.225 ;
        RECT 350.855 655.945 351.135 656.225 ;
        RECT 351.475 655.945 351.755 656.225 ;
        RECT 352.095 655.945 352.375 656.225 ;
        RECT 350.235 653.395 350.515 653.675 ;
        RECT 350.855 653.395 351.135 653.675 ;
        RECT 351.475 653.395 351.755 653.675 ;
        RECT 352.095 653.395 352.375 653.675 ;
        RECT 350.235 652.775 350.515 653.055 ;
        RECT 350.855 652.775 351.135 653.055 ;
        RECT 351.475 652.775 351.755 653.055 ;
        RECT 352.095 652.775 352.375 653.055 ;
        RECT 350.235 652.155 350.515 652.435 ;
        RECT 350.855 652.155 351.135 652.435 ;
        RECT 351.475 652.155 351.755 652.435 ;
        RECT 352.095 652.155 352.375 652.435 ;
        RECT 350.235 651.535 350.515 651.815 ;
        RECT 350.855 651.535 351.135 651.815 ;
        RECT 351.475 651.535 351.755 651.815 ;
        RECT 352.095 651.535 352.375 651.815 ;
        RECT 350.235 650.915 350.515 651.195 ;
        RECT 350.855 650.915 351.135 651.195 ;
        RECT 351.475 650.915 351.755 651.195 ;
        RECT 352.095 650.915 352.375 651.195 ;
        RECT 350.235 650.295 350.515 650.575 ;
        RECT 350.855 650.295 351.135 650.575 ;
        RECT 351.475 650.295 351.755 650.575 ;
        RECT 352.095 650.295 352.375 650.575 ;
        RECT 350.235 649.675 350.515 649.955 ;
        RECT 350.855 649.675 351.135 649.955 ;
        RECT 351.475 649.675 351.755 649.955 ;
        RECT 352.095 649.675 352.375 649.955 ;
        RECT 350.235 649.055 350.515 649.335 ;
        RECT 350.855 649.055 351.135 649.335 ;
        RECT 351.475 649.055 351.755 649.335 ;
        RECT 352.095 649.055 352.375 649.335 ;
        RECT 350.235 648.435 350.515 648.715 ;
        RECT 350.855 648.435 351.135 648.715 ;
        RECT 351.475 648.435 351.755 648.715 ;
        RECT 352.095 648.435 352.375 648.715 ;
        RECT 350.235 647.815 350.515 648.095 ;
        RECT 350.855 647.815 351.135 648.095 ;
        RECT 351.475 647.815 351.755 648.095 ;
        RECT 352.095 647.815 352.375 648.095 ;
        RECT 350.235 647.195 350.515 647.475 ;
        RECT 350.855 647.195 351.135 647.475 ;
        RECT 351.475 647.195 351.755 647.475 ;
        RECT 352.095 647.195 352.375 647.475 ;
        RECT 350.235 646.575 350.515 646.855 ;
        RECT 350.855 646.575 351.135 646.855 ;
        RECT 351.475 646.575 351.755 646.855 ;
        RECT 352.095 646.575 352.375 646.855 ;
        RECT 350.235 645.955 350.515 646.235 ;
        RECT 350.855 645.955 351.135 646.235 ;
        RECT 351.475 645.955 351.755 646.235 ;
        RECT 352.095 645.955 352.375 646.235 ;
        RECT 350.235 645.335 350.515 645.615 ;
        RECT 350.855 645.335 351.135 645.615 ;
        RECT 351.475 645.335 351.755 645.615 ;
        RECT 352.095 645.335 352.375 645.615 ;
        RECT 350.235 644.715 350.515 644.995 ;
        RECT 350.855 644.715 351.135 644.995 ;
        RECT 351.475 644.715 351.755 644.995 ;
        RECT 352.095 644.715 352.375 644.995 ;
        RECT 350.235 644.095 350.515 644.375 ;
        RECT 350.855 644.095 351.135 644.375 ;
        RECT 351.475 644.095 351.755 644.375 ;
        RECT 352.095 644.095 352.375 644.375 ;
        RECT 350.235 640.245 350.515 640.525 ;
        RECT 350.855 640.245 351.135 640.525 ;
        RECT 351.475 640.245 351.755 640.525 ;
        RECT 352.095 640.245 352.375 640.525 ;
        RECT 350.235 639.625 350.515 639.905 ;
        RECT 350.855 639.625 351.135 639.905 ;
        RECT 351.475 639.625 351.755 639.905 ;
        RECT 352.095 639.625 352.375 639.905 ;
        RECT 350.235 639.005 350.515 639.285 ;
        RECT 350.855 639.005 351.135 639.285 ;
        RECT 351.475 639.005 351.755 639.285 ;
        RECT 352.095 639.005 352.375 639.285 ;
        RECT 350.235 638.385 350.515 638.665 ;
        RECT 350.855 638.385 351.135 638.665 ;
        RECT 351.475 638.385 351.755 638.665 ;
        RECT 352.095 638.385 352.375 638.665 ;
        RECT 350.235 637.765 350.515 638.045 ;
        RECT 350.855 637.765 351.135 638.045 ;
        RECT 351.475 637.765 351.755 638.045 ;
        RECT 352.095 637.765 352.375 638.045 ;
        RECT 350.235 637.145 350.515 637.425 ;
        RECT 350.855 637.145 351.135 637.425 ;
        RECT 351.475 637.145 351.755 637.425 ;
        RECT 352.095 637.145 352.375 637.425 ;
        RECT 350.235 636.525 350.515 636.805 ;
        RECT 350.855 636.525 351.135 636.805 ;
        RECT 351.475 636.525 351.755 636.805 ;
        RECT 352.095 636.525 352.375 636.805 ;
        RECT 350.235 635.905 350.515 636.185 ;
        RECT 350.855 635.905 351.135 636.185 ;
        RECT 351.475 635.905 351.755 636.185 ;
        RECT 352.095 635.905 352.375 636.185 ;
        RECT 350.235 635.285 350.515 635.565 ;
        RECT 350.855 635.285 351.135 635.565 ;
        RECT 351.475 635.285 351.755 635.565 ;
        RECT 352.095 635.285 352.375 635.565 ;
        RECT 350.235 634.665 350.515 634.945 ;
        RECT 350.855 634.665 351.135 634.945 ;
        RECT 351.475 634.665 351.755 634.945 ;
        RECT 352.095 634.665 352.375 634.945 ;
        RECT 350.235 634.045 350.515 634.325 ;
        RECT 350.855 634.045 351.135 634.325 ;
        RECT 351.475 634.045 351.755 634.325 ;
        RECT 352.095 634.045 352.375 634.325 ;
        RECT 350.235 633.425 350.515 633.705 ;
        RECT 350.855 633.425 351.135 633.705 ;
        RECT 351.475 633.425 351.755 633.705 ;
        RECT 352.095 633.425 352.375 633.705 ;
        RECT 350.235 632.805 350.515 633.085 ;
        RECT 350.855 632.805 351.135 633.085 ;
        RECT 351.475 632.805 351.755 633.085 ;
        RECT 352.095 632.805 352.375 633.085 ;
        RECT 350.235 632.185 350.515 632.465 ;
        RECT 350.855 632.185 351.135 632.465 ;
        RECT 351.475 632.185 351.755 632.465 ;
        RECT 352.095 632.185 352.375 632.465 ;
        RECT 350.235 631.565 350.515 631.845 ;
        RECT 350.855 631.565 351.135 631.845 ;
        RECT 351.475 631.565 351.755 631.845 ;
        RECT 352.095 631.565 352.375 631.845 ;
        RECT 350.235 498.025 350.515 498.305 ;
        RECT 350.855 498.025 351.135 498.305 ;
        RECT 351.475 498.025 351.755 498.305 ;
        RECT 352.095 498.025 352.375 498.305 ;
        RECT 350.235 497.405 350.515 497.685 ;
        RECT 350.855 497.405 351.135 497.685 ;
        RECT 351.475 497.405 351.755 497.685 ;
        RECT 352.095 497.405 352.375 497.685 ;
        RECT 350.235 496.785 350.515 497.065 ;
        RECT 350.855 496.785 351.135 497.065 ;
        RECT 351.475 496.785 351.755 497.065 ;
        RECT 352.095 496.785 352.375 497.065 ;
        RECT 350.235 496.165 350.515 496.445 ;
        RECT 350.855 496.165 351.135 496.445 ;
        RECT 351.475 496.165 351.755 496.445 ;
        RECT 352.095 496.165 352.375 496.445 ;
        RECT 350.235 495.545 350.515 495.825 ;
        RECT 350.855 495.545 351.135 495.825 ;
        RECT 351.475 495.545 351.755 495.825 ;
        RECT 352.095 495.545 352.375 495.825 ;
        RECT 350.235 494.925 350.515 495.205 ;
        RECT 350.855 494.925 351.135 495.205 ;
        RECT 351.475 494.925 351.755 495.205 ;
        RECT 352.095 494.925 352.375 495.205 ;
        RECT 350.235 494.305 350.515 494.585 ;
        RECT 350.855 494.305 351.135 494.585 ;
        RECT 351.475 494.305 351.755 494.585 ;
        RECT 352.095 494.305 352.375 494.585 ;
        RECT 350.235 493.685 350.515 493.965 ;
        RECT 350.855 493.685 351.135 493.965 ;
        RECT 351.475 493.685 351.755 493.965 ;
        RECT 352.095 493.685 352.375 493.965 ;
        RECT 350.235 493.065 350.515 493.345 ;
        RECT 350.855 493.065 351.135 493.345 ;
        RECT 351.475 493.065 351.755 493.345 ;
        RECT 352.095 493.065 352.375 493.345 ;
        RECT 350.235 492.445 350.515 492.725 ;
        RECT 350.855 492.445 351.135 492.725 ;
        RECT 351.475 492.445 351.755 492.725 ;
        RECT 352.095 492.445 352.375 492.725 ;
        RECT 350.235 491.825 350.515 492.105 ;
        RECT 350.855 491.825 351.135 492.105 ;
        RECT 351.475 491.825 351.755 492.105 ;
        RECT 352.095 491.825 352.375 492.105 ;
        RECT 350.235 491.205 350.515 491.485 ;
        RECT 350.855 491.205 351.135 491.485 ;
        RECT 351.475 491.205 351.755 491.485 ;
        RECT 352.095 491.205 352.375 491.485 ;
        RECT 350.235 490.585 350.515 490.865 ;
        RECT 350.855 490.585 351.135 490.865 ;
        RECT 351.475 490.585 351.755 490.865 ;
        RECT 352.095 490.585 352.375 490.865 ;
        RECT 350.235 489.965 350.515 490.245 ;
        RECT 350.855 489.965 351.135 490.245 ;
        RECT 351.475 489.965 351.755 490.245 ;
        RECT 352.095 489.965 352.375 490.245 ;
        RECT 350.235 489.345 350.515 489.625 ;
        RECT 350.855 489.345 351.135 489.625 ;
        RECT 351.475 489.345 351.755 489.625 ;
        RECT 352.095 489.345 352.375 489.625 ;
        RECT 350.235 485.625 350.515 485.905 ;
        RECT 350.855 485.625 351.135 485.905 ;
        RECT 351.475 485.625 351.755 485.905 ;
        RECT 352.095 485.625 352.375 485.905 ;
        RECT 350.235 485.005 350.515 485.285 ;
        RECT 350.855 485.005 351.135 485.285 ;
        RECT 351.475 485.005 351.755 485.285 ;
        RECT 352.095 485.005 352.375 485.285 ;
        RECT 350.235 484.385 350.515 484.665 ;
        RECT 350.855 484.385 351.135 484.665 ;
        RECT 351.475 484.385 351.755 484.665 ;
        RECT 352.095 484.385 352.375 484.665 ;
        RECT 350.235 483.765 350.515 484.045 ;
        RECT 350.855 483.765 351.135 484.045 ;
        RECT 351.475 483.765 351.755 484.045 ;
        RECT 352.095 483.765 352.375 484.045 ;
        RECT 350.235 483.145 350.515 483.425 ;
        RECT 350.855 483.145 351.135 483.425 ;
        RECT 351.475 483.145 351.755 483.425 ;
        RECT 352.095 483.145 352.375 483.425 ;
        RECT 350.235 482.525 350.515 482.805 ;
        RECT 350.855 482.525 351.135 482.805 ;
        RECT 351.475 482.525 351.755 482.805 ;
        RECT 352.095 482.525 352.375 482.805 ;
        RECT 350.235 481.905 350.515 482.185 ;
        RECT 350.855 481.905 351.135 482.185 ;
        RECT 351.475 481.905 351.755 482.185 ;
        RECT 352.095 481.905 352.375 482.185 ;
        RECT 350.235 481.285 350.515 481.565 ;
        RECT 350.855 481.285 351.135 481.565 ;
        RECT 351.475 481.285 351.755 481.565 ;
        RECT 352.095 481.285 352.375 481.565 ;
        RECT 350.235 480.665 350.515 480.945 ;
        RECT 350.855 480.665 351.135 480.945 ;
        RECT 351.475 480.665 351.755 480.945 ;
        RECT 352.095 480.665 352.375 480.945 ;
        RECT 350.235 480.045 350.515 480.325 ;
        RECT 350.855 480.045 351.135 480.325 ;
        RECT 351.475 480.045 351.755 480.325 ;
        RECT 352.095 480.045 352.375 480.325 ;
        RECT 350.235 479.425 350.515 479.705 ;
        RECT 350.855 479.425 351.135 479.705 ;
        RECT 351.475 479.425 351.755 479.705 ;
        RECT 352.095 479.425 352.375 479.705 ;
        RECT 350.235 478.805 350.515 479.085 ;
        RECT 350.855 478.805 351.135 479.085 ;
        RECT 351.475 478.805 351.755 479.085 ;
        RECT 352.095 478.805 352.375 479.085 ;
        RECT 350.235 478.185 350.515 478.465 ;
        RECT 350.855 478.185 351.135 478.465 ;
        RECT 351.475 478.185 351.755 478.465 ;
        RECT 352.095 478.185 352.375 478.465 ;
        RECT 350.235 477.565 350.515 477.845 ;
        RECT 350.855 477.565 351.135 477.845 ;
        RECT 351.475 477.565 351.755 477.845 ;
        RECT 352.095 477.565 352.375 477.845 ;
        RECT 350.235 476.945 350.515 477.225 ;
        RECT 350.855 476.945 351.135 477.225 ;
        RECT 351.475 476.945 351.755 477.225 ;
        RECT 352.095 476.945 352.375 477.225 ;
        RECT 350.235 476.325 350.515 476.605 ;
        RECT 350.855 476.325 351.135 476.605 ;
        RECT 351.475 476.325 351.755 476.605 ;
        RECT 352.095 476.325 352.375 476.605 ;
        RECT 350.235 473.775 350.515 474.055 ;
        RECT 350.855 473.775 351.135 474.055 ;
        RECT 351.475 473.775 351.755 474.055 ;
        RECT 352.095 473.775 352.375 474.055 ;
        RECT 350.235 473.155 350.515 473.435 ;
        RECT 350.855 473.155 351.135 473.435 ;
        RECT 351.475 473.155 351.755 473.435 ;
        RECT 352.095 473.155 352.375 473.435 ;
        RECT 350.235 472.535 350.515 472.815 ;
        RECT 350.855 472.535 351.135 472.815 ;
        RECT 351.475 472.535 351.755 472.815 ;
        RECT 352.095 472.535 352.375 472.815 ;
        RECT 350.235 471.915 350.515 472.195 ;
        RECT 350.855 471.915 351.135 472.195 ;
        RECT 351.475 471.915 351.755 472.195 ;
        RECT 352.095 471.915 352.375 472.195 ;
        RECT 350.235 471.295 350.515 471.575 ;
        RECT 350.855 471.295 351.135 471.575 ;
        RECT 351.475 471.295 351.755 471.575 ;
        RECT 352.095 471.295 352.375 471.575 ;
        RECT 350.235 470.675 350.515 470.955 ;
        RECT 350.855 470.675 351.135 470.955 ;
        RECT 351.475 470.675 351.755 470.955 ;
        RECT 352.095 470.675 352.375 470.955 ;
        RECT 350.235 470.055 350.515 470.335 ;
        RECT 350.855 470.055 351.135 470.335 ;
        RECT 351.475 470.055 351.755 470.335 ;
        RECT 352.095 470.055 352.375 470.335 ;
        RECT 350.235 469.435 350.515 469.715 ;
        RECT 350.855 469.435 351.135 469.715 ;
        RECT 351.475 469.435 351.755 469.715 ;
        RECT 352.095 469.435 352.375 469.715 ;
        RECT 350.235 468.815 350.515 469.095 ;
        RECT 350.855 468.815 351.135 469.095 ;
        RECT 351.475 468.815 351.755 469.095 ;
        RECT 352.095 468.815 352.375 469.095 ;
        RECT 350.235 468.195 350.515 468.475 ;
        RECT 350.855 468.195 351.135 468.475 ;
        RECT 351.475 468.195 351.755 468.475 ;
        RECT 352.095 468.195 352.375 468.475 ;
        RECT 350.235 467.575 350.515 467.855 ;
        RECT 350.855 467.575 351.135 467.855 ;
        RECT 351.475 467.575 351.755 467.855 ;
        RECT 352.095 467.575 352.375 467.855 ;
        RECT 350.235 466.955 350.515 467.235 ;
        RECT 350.855 466.955 351.135 467.235 ;
        RECT 351.475 466.955 351.755 467.235 ;
        RECT 352.095 466.955 352.375 467.235 ;
        RECT 350.235 466.335 350.515 466.615 ;
        RECT 350.855 466.335 351.135 466.615 ;
        RECT 351.475 466.335 351.755 466.615 ;
        RECT 352.095 466.335 352.375 466.615 ;
        RECT 350.235 465.715 350.515 465.995 ;
        RECT 350.855 465.715 351.135 465.995 ;
        RECT 351.475 465.715 351.755 465.995 ;
        RECT 352.095 465.715 352.375 465.995 ;
        RECT 350.235 465.095 350.515 465.375 ;
        RECT 350.855 465.095 351.135 465.375 ;
        RECT 351.475 465.095 351.755 465.375 ;
        RECT 352.095 465.095 352.375 465.375 ;
        RECT 350.235 464.475 350.515 464.755 ;
        RECT 350.855 464.475 351.135 464.755 ;
        RECT 351.475 464.475 351.755 464.755 ;
        RECT 352.095 464.475 352.375 464.755 ;
        RECT 350.235 460.245 350.515 460.525 ;
        RECT 350.855 460.245 351.135 460.525 ;
        RECT 351.475 460.245 351.755 460.525 ;
        RECT 352.095 460.245 352.375 460.525 ;
        RECT 350.235 459.625 350.515 459.905 ;
        RECT 350.855 459.625 351.135 459.905 ;
        RECT 351.475 459.625 351.755 459.905 ;
        RECT 352.095 459.625 352.375 459.905 ;
        RECT 350.235 459.005 350.515 459.285 ;
        RECT 350.855 459.005 351.135 459.285 ;
        RECT 351.475 459.005 351.755 459.285 ;
        RECT 352.095 459.005 352.375 459.285 ;
        RECT 350.235 458.385 350.515 458.665 ;
        RECT 350.855 458.385 351.135 458.665 ;
        RECT 351.475 458.385 351.755 458.665 ;
        RECT 352.095 458.385 352.375 458.665 ;
        RECT 350.235 457.765 350.515 458.045 ;
        RECT 350.855 457.765 351.135 458.045 ;
        RECT 351.475 457.765 351.755 458.045 ;
        RECT 352.095 457.765 352.375 458.045 ;
        RECT 350.235 457.145 350.515 457.425 ;
        RECT 350.855 457.145 351.135 457.425 ;
        RECT 351.475 457.145 351.755 457.425 ;
        RECT 352.095 457.145 352.375 457.425 ;
        RECT 350.235 456.525 350.515 456.805 ;
        RECT 350.855 456.525 351.135 456.805 ;
        RECT 351.475 456.525 351.755 456.805 ;
        RECT 352.095 456.525 352.375 456.805 ;
        RECT 350.235 455.905 350.515 456.185 ;
        RECT 350.855 455.905 351.135 456.185 ;
        RECT 351.475 455.905 351.755 456.185 ;
        RECT 352.095 455.905 352.375 456.185 ;
        RECT 350.235 455.285 350.515 455.565 ;
        RECT 350.855 455.285 351.135 455.565 ;
        RECT 351.475 455.285 351.755 455.565 ;
        RECT 352.095 455.285 352.375 455.565 ;
        RECT 350.235 454.665 350.515 454.945 ;
        RECT 350.855 454.665 351.135 454.945 ;
        RECT 351.475 454.665 351.755 454.945 ;
        RECT 352.095 454.665 352.375 454.945 ;
        RECT 350.235 454.045 350.515 454.325 ;
        RECT 350.855 454.045 351.135 454.325 ;
        RECT 351.475 454.045 351.755 454.325 ;
        RECT 352.095 454.045 352.375 454.325 ;
        RECT 350.235 453.425 350.515 453.705 ;
        RECT 350.855 453.425 351.135 453.705 ;
        RECT 351.475 453.425 351.755 453.705 ;
        RECT 352.095 453.425 352.375 453.705 ;
        RECT 350.235 452.805 350.515 453.085 ;
        RECT 350.855 452.805 351.135 453.085 ;
        RECT 351.475 452.805 351.755 453.085 ;
        RECT 352.095 452.805 352.375 453.085 ;
        RECT 350.235 452.185 350.515 452.465 ;
        RECT 350.855 452.185 351.135 452.465 ;
        RECT 351.475 452.185 351.755 452.465 ;
        RECT 352.095 452.185 352.375 452.465 ;
        RECT 350.235 451.565 350.515 451.845 ;
        RECT 350.855 451.565 351.135 451.845 ;
        RECT 351.475 451.565 351.755 451.845 ;
        RECT 352.095 451.565 352.375 451.845 ;
        RECT 350.235 450.945 350.515 451.225 ;
        RECT 350.855 450.945 351.135 451.225 ;
        RECT 351.475 450.945 351.755 451.225 ;
        RECT 352.095 450.945 352.375 451.225 ;
        RECT 350.235 448.395 350.515 448.675 ;
        RECT 350.855 448.395 351.135 448.675 ;
        RECT 351.475 448.395 351.755 448.675 ;
        RECT 352.095 448.395 352.375 448.675 ;
        RECT 350.235 447.775 350.515 448.055 ;
        RECT 350.855 447.775 351.135 448.055 ;
        RECT 351.475 447.775 351.755 448.055 ;
        RECT 352.095 447.775 352.375 448.055 ;
        RECT 350.235 447.155 350.515 447.435 ;
        RECT 350.855 447.155 351.135 447.435 ;
        RECT 351.475 447.155 351.755 447.435 ;
        RECT 352.095 447.155 352.375 447.435 ;
        RECT 350.235 446.535 350.515 446.815 ;
        RECT 350.855 446.535 351.135 446.815 ;
        RECT 351.475 446.535 351.755 446.815 ;
        RECT 352.095 446.535 352.375 446.815 ;
        RECT 350.235 445.915 350.515 446.195 ;
        RECT 350.855 445.915 351.135 446.195 ;
        RECT 351.475 445.915 351.755 446.195 ;
        RECT 352.095 445.915 352.375 446.195 ;
        RECT 350.235 445.295 350.515 445.575 ;
        RECT 350.855 445.295 351.135 445.575 ;
        RECT 351.475 445.295 351.755 445.575 ;
        RECT 352.095 445.295 352.375 445.575 ;
        RECT 350.235 444.675 350.515 444.955 ;
        RECT 350.855 444.675 351.135 444.955 ;
        RECT 351.475 444.675 351.755 444.955 ;
        RECT 352.095 444.675 352.375 444.955 ;
        RECT 350.235 444.055 350.515 444.335 ;
        RECT 350.855 444.055 351.135 444.335 ;
        RECT 351.475 444.055 351.755 444.335 ;
        RECT 352.095 444.055 352.375 444.335 ;
        RECT 350.235 443.435 350.515 443.715 ;
        RECT 350.855 443.435 351.135 443.715 ;
        RECT 351.475 443.435 351.755 443.715 ;
        RECT 352.095 443.435 352.375 443.715 ;
        RECT 350.235 442.815 350.515 443.095 ;
        RECT 350.855 442.815 351.135 443.095 ;
        RECT 351.475 442.815 351.755 443.095 ;
        RECT 352.095 442.815 352.375 443.095 ;
        RECT 350.235 442.195 350.515 442.475 ;
        RECT 350.855 442.195 351.135 442.475 ;
        RECT 351.475 442.195 351.755 442.475 ;
        RECT 352.095 442.195 352.375 442.475 ;
        RECT 350.235 441.575 350.515 441.855 ;
        RECT 350.855 441.575 351.135 441.855 ;
        RECT 351.475 441.575 351.755 441.855 ;
        RECT 352.095 441.575 352.375 441.855 ;
        RECT 350.235 440.955 350.515 441.235 ;
        RECT 350.855 440.955 351.135 441.235 ;
        RECT 351.475 440.955 351.755 441.235 ;
        RECT 352.095 440.955 352.375 441.235 ;
        RECT 350.235 440.335 350.515 440.615 ;
        RECT 350.855 440.335 351.135 440.615 ;
        RECT 351.475 440.335 351.755 440.615 ;
        RECT 352.095 440.335 352.375 440.615 ;
        RECT 350.235 439.715 350.515 439.995 ;
        RECT 350.855 439.715 351.135 439.995 ;
        RECT 351.475 439.715 351.755 439.995 ;
        RECT 352.095 439.715 352.375 439.995 ;
        RECT 350.235 439.095 350.515 439.375 ;
        RECT 350.855 439.095 351.135 439.375 ;
        RECT 351.475 439.095 351.755 439.375 ;
        RECT 352.095 439.095 352.375 439.375 ;
        RECT 350.235 435.245 350.515 435.525 ;
        RECT 350.855 435.245 351.135 435.525 ;
        RECT 351.475 435.245 351.755 435.525 ;
        RECT 352.095 435.245 352.375 435.525 ;
        RECT 350.235 434.625 350.515 434.905 ;
        RECT 350.855 434.625 351.135 434.905 ;
        RECT 351.475 434.625 351.755 434.905 ;
        RECT 352.095 434.625 352.375 434.905 ;
        RECT 350.235 434.005 350.515 434.285 ;
        RECT 350.855 434.005 351.135 434.285 ;
        RECT 351.475 434.005 351.755 434.285 ;
        RECT 352.095 434.005 352.375 434.285 ;
        RECT 350.235 433.385 350.515 433.665 ;
        RECT 350.855 433.385 351.135 433.665 ;
        RECT 351.475 433.385 351.755 433.665 ;
        RECT 352.095 433.385 352.375 433.665 ;
        RECT 350.235 432.765 350.515 433.045 ;
        RECT 350.855 432.765 351.135 433.045 ;
        RECT 351.475 432.765 351.755 433.045 ;
        RECT 352.095 432.765 352.375 433.045 ;
        RECT 350.235 432.145 350.515 432.425 ;
        RECT 350.855 432.145 351.135 432.425 ;
        RECT 351.475 432.145 351.755 432.425 ;
        RECT 352.095 432.145 352.375 432.425 ;
        RECT 350.235 431.525 350.515 431.805 ;
        RECT 350.855 431.525 351.135 431.805 ;
        RECT 351.475 431.525 351.755 431.805 ;
        RECT 352.095 431.525 352.375 431.805 ;
        RECT 350.235 430.905 350.515 431.185 ;
        RECT 350.855 430.905 351.135 431.185 ;
        RECT 351.475 430.905 351.755 431.185 ;
        RECT 352.095 430.905 352.375 431.185 ;
        RECT 350.235 430.285 350.515 430.565 ;
        RECT 350.855 430.285 351.135 430.565 ;
        RECT 351.475 430.285 351.755 430.565 ;
        RECT 352.095 430.285 352.375 430.565 ;
        RECT 350.235 429.665 350.515 429.945 ;
        RECT 350.855 429.665 351.135 429.945 ;
        RECT 351.475 429.665 351.755 429.945 ;
        RECT 352.095 429.665 352.375 429.945 ;
        RECT 350.235 429.045 350.515 429.325 ;
        RECT 350.855 429.045 351.135 429.325 ;
        RECT 351.475 429.045 351.755 429.325 ;
        RECT 352.095 429.045 352.375 429.325 ;
        RECT 350.235 428.425 350.515 428.705 ;
        RECT 350.855 428.425 351.135 428.705 ;
        RECT 351.475 428.425 351.755 428.705 ;
        RECT 352.095 428.425 352.375 428.705 ;
        RECT 350.235 427.805 350.515 428.085 ;
        RECT 350.855 427.805 351.135 428.085 ;
        RECT 351.475 427.805 351.755 428.085 ;
        RECT 352.095 427.805 352.375 428.085 ;
        RECT 350.235 427.185 350.515 427.465 ;
        RECT 350.855 427.185 351.135 427.465 ;
        RECT 351.475 427.185 351.755 427.465 ;
        RECT 352.095 427.185 352.375 427.465 ;
        RECT 350.235 426.565 350.515 426.845 ;
        RECT 350.855 426.565 351.135 426.845 ;
        RECT 351.475 426.565 351.755 426.845 ;
        RECT 352.095 426.565 352.375 426.845 ;
        RECT 3276.630 379.445 3276.910 379.725 ;
        RECT 3277.250 379.445 3277.530 379.725 ;
        RECT 3277.870 379.445 3278.150 379.725 ;
        RECT 3278.490 379.445 3278.770 379.725 ;
        RECT 3279.110 379.445 3279.390 379.725 ;
        RECT 3279.730 379.445 3280.010 379.725 ;
        RECT 3280.350 379.445 3280.630 379.725 ;
        RECT 3280.970 379.445 3281.250 379.725 ;
        RECT 3281.590 379.445 3281.870 379.725 ;
        RECT 3276.630 378.825 3276.910 379.105 ;
        RECT 3277.250 378.825 3277.530 379.105 ;
        RECT 3277.870 378.825 3278.150 379.105 ;
        RECT 3278.490 378.825 3278.770 379.105 ;
        RECT 3279.110 378.825 3279.390 379.105 ;
        RECT 3279.730 378.825 3280.010 379.105 ;
        RECT 3280.350 378.825 3280.630 379.105 ;
        RECT 3280.970 378.825 3281.250 379.105 ;
        RECT 3281.590 378.825 3281.870 379.105 ;
        RECT 3276.630 378.205 3276.910 378.485 ;
        RECT 3277.250 378.205 3277.530 378.485 ;
        RECT 3277.870 378.205 3278.150 378.485 ;
        RECT 3278.490 378.205 3278.770 378.485 ;
        RECT 3279.110 378.205 3279.390 378.485 ;
        RECT 3279.730 378.205 3280.010 378.485 ;
        RECT 3280.350 378.205 3280.630 378.485 ;
        RECT 3280.970 378.205 3281.250 378.485 ;
        RECT 3281.590 378.205 3281.870 378.485 ;
        RECT 3276.630 377.585 3276.910 377.865 ;
        RECT 3277.250 377.585 3277.530 377.865 ;
        RECT 3277.870 377.585 3278.150 377.865 ;
        RECT 3278.490 377.585 3278.770 377.865 ;
        RECT 3279.110 377.585 3279.390 377.865 ;
        RECT 3279.730 377.585 3280.010 377.865 ;
        RECT 3280.350 377.585 3280.630 377.865 ;
        RECT 3280.970 377.585 3281.250 377.865 ;
        RECT 3281.590 377.585 3281.870 377.865 ;
        RECT 3276.630 376.965 3276.910 377.245 ;
        RECT 3277.250 376.965 3277.530 377.245 ;
        RECT 3277.870 376.965 3278.150 377.245 ;
        RECT 3278.490 376.965 3278.770 377.245 ;
        RECT 3279.110 376.965 3279.390 377.245 ;
        RECT 3279.730 376.965 3280.010 377.245 ;
        RECT 3280.350 376.965 3280.630 377.245 ;
        RECT 3280.970 376.965 3281.250 377.245 ;
        RECT 3281.590 376.965 3281.870 377.245 ;
        RECT 3276.630 376.345 3276.910 376.625 ;
        RECT 3277.250 376.345 3277.530 376.625 ;
        RECT 3277.870 376.345 3278.150 376.625 ;
        RECT 3278.490 376.345 3278.770 376.625 ;
        RECT 3279.110 376.345 3279.390 376.625 ;
        RECT 3279.730 376.345 3280.010 376.625 ;
        RECT 3280.350 376.345 3280.630 376.625 ;
        RECT 3280.970 376.345 3281.250 376.625 ;
        RECT 3281.590 376.345 3281.870 376.625 ;
        RECT 3276.630 375.725 3276.910 376.005 ;
        RECT 3277.250 375.725 3277.530 376.005 ;
        RECT 3277.870 375.725 3278.150 376.005 ;
        RECT 3278.490 375.725 3278.770 376.005 ;
        RECT 3279.110 375.725 3279.390 376.005 ;
        RECT 3279.730 375.725 3280.010 376.005 ;
        RECT 3280.350 375.725 3280.630 376.005 ;
        RECT 3280.970 375.725 3281.250 376.005 ;
        RECT 3281.590 375.725 3281.870 376.005 ;
        RECT 3276.630 375.105 3276.910 375.385 ;
        RECT 3277.250 375.105 3277.530 375.385 ;
        RECT 3277.870 375.105 3278.150 375.385 ;
        RECT 3278.490 375.105 3278.770 375.385 ;
        RECT 3279.110 375.105 3279.390 375.385 ;
        RECT 3279.730 375.105 3280.010 375.385 ;
        RECT 3280.350 375.105 3280.630 375.385 ;
        RECT 3280.970 375.105 3281.250 375.385 ;
        RECT 3281.590 375.105 3281.870 375.385 ;
        RECT 3276.630 374.485 3276.910 374.765 ;
        RECT 3277.250 374.485 3277.530 374.765 ;
        RECT 3277.870 374.485 3278.150 374.765 ;
        RECT 3278.490 374.485 3278.770 374.765 ;
        RECT 3279.110 374.485 3279.390 374.765 ;
        RECT 3279.730 374.485 3280.010 374.765 ;
        RECT 3280.350 374.485 3280.630 374.765 ;
        RECT 3280.970 374.485 3281.250 374.765 ;
        RECT 3281.590 374.485 3281.870 374.765 ;
        RECT 3276.630 373.865 3276.910 374.145 ;
        RECT 3277.250 373.865 3277.530 374.145 ;
        RECT 3277.870 373.865 3278.150 374.145 ;
        RECT 3278.490 373.865 3278.770 374.145 ;
        RECT 3279.110 373.865 3279.390 374.145 ;
        RECT 3279.730 373.865 3280.010 374.145 ;
        RECT 3280.350 373.865 3280.630 374.145 ;
        RECT 3280.970 373.865 3281.250 374.145 ;
        RECT 3281.590 373.865 3281.870 374.145 ;
        RECT 3276.630 373.245 3276.910 373.525 ;
        RECT 3277.250 373.245 3277.530 373.525 ;
        RECT 3277.870 373.245 3278.150 373.525 ;
        RECT 3278.490 373.245 3278.770 373.525 ;
        RECT 3279.110 373.245 3279.390 373.525 ;
        RECT 3279.730 373.245 3280.010 373.525 ;
        RECT 3280.350 373.245 3280.630 373.525 ;
        RECT 3280.970 373.245 3281.250 373.525 ;
        RECT 3281.590 373.245 3281.870 373.525 ;
        RECT 3276.630 372.625 3276.910 372.905 ;
        RECT 3277.250 372.625 3277.530 372.905 ;
        RECT 3277.870 372.625 3278.150 372.905 ;
        RECT 3278.490 372.625 3278.770 372.905 ;
        RECT 3279.110 372.625 3279.390 372.905 ;
        RECT 3279.730 372.625 3280.010 372.905 ;
        RECT 3280.350 372.625 3280.630 372.905 ;
        RECT 3280.970 372.625 3281.250 372.905 ;
        RECT 3281.590 372.625 3281.870 372.905 ;
        RECT 526.630 369.445 526.910 369.725 ;
        RECT 527.250 369.445 527.530 369.725 ;
        RECT 527.870 369.445 528.150 369.725 ;
        RECT 528.490 369.445 528.770 369.725 ;
        RECT 529.110 369.445 529.390 369.725 ;
        RECT 529.730 369.445 530.010 369.725 ;
        RECT 530.350 369.445 530.630 369.725 ;
        RECT 530.970 369.445 531.250 369.725 ;
        RECT 531.590 369.445 531.870 369.725 ;
        RECT 532.210 369.445 532.490 369.725 ;
        RECT 532.830 369.445 533.110 369.725 ;
        RECT 533.450 369.445 533.730 369.725 ;
        RECT 534.070 369.445 534.350 369.725 ;
        RECT 534.690 369.445 534.970 369.725 ;
        RECT 535.310 369.445 535.590 369.725 ;
        RECT 526.630 368.825 526.910 369.105 ;
        RECT 527.250 368.825 527.530 369.105 ;
        RECT 527.870 368.825 528.150 369.105 ;
        RECT 528.490 368.825 528.770 369.105 ;
        RECT 529.110 368.825 529.390 369.105 ;
        RECT 529.730 368.825 530.010 369.105 ;
        RECT 530.350 368.825 530.630 369.105 ;
        RECT 530.970 368.825 531.250 369.105 ;
        RECT 531.590 368.825 531.870 369.105 ;
        RECT 532.210 368.825 532.490 369.105 ;
        RECT 532.830 368.825 533.110 369.105 ;
        RECT 533.450 368.825 533.730 369.105 ;
        RECT 534.070 368.825 534.350 369.105 ;
        RECT 534.690 368.825 534.970 369.105 ;
        RECT 535.310 368.825 535.590 369.105 ;
        RECT 526.630 368.205 526.910 368.485 ;
        RECT 527.250 368.205 527.530 368.485 ;
        RECT 527.870 368.205 528.150 368.485 ;
        RECT 528.490 368.205 528.770 368.485 ;
        RECT 529.110 368.205 529.390 368.485 ;
        RECT 529.730 368.205 530.010 368.485 ;
        RECT 530.350 368.205 530.630 368.485 ;
        RECT 530.970 368.205 531.250 368.485 ;
        RECT 531.590 368.205 531.870 368.485 ;
        RECT 532.210 368.205 532.490 368.485 ;
        RECT 532.830 368.205 533.110 368.485 ;
        RECT 533.450 368.205 533.730 368.485 ;
        RECT 534.070 368.205 534.350 368.485 ;
        RECT 534.690 368.205 534.970 368.485 ;
        RECT 535.310 368.205 535.590 368.485 ;
        RECT 526.630 367.585 526.910 367.865 ;
        RECT 527.250 367.585 527.530 367.865 ;
        RECT 527.870 367.585 528.150 367.865 ;
        RECT 528.490 367.585 528.770 367.865 ;
        RECT 529.110 367.585 529.390 367.865 ;
        RECT 529.730 367.585 530.010 367.865 ;
        RECT 530.350 367.585 530.630 367.865 ;
        RECT 530.970 367.585 531.250 367.865 ;
        RECT 531.590 367.585 531.870 367.865 ;
        RECT 532.210 367.585 532.490 367.865 ;
        RECT 532.830 367.585 533.110 367.865 ;
        RECT 533.450 367.585 533.730 367.865 ;
        RECT 534.070 367.585 534.350 367.865 ;
        RECT 534.690 367.585 534.970 367.865 ;
        RECT 535.310 367.585 535.590 367.865 ;
        RECT 526.630 366.965 526.910 367.245 ;
        RECT 527.250 366.965 527.530 367.245 ;
        RECT 527.870 366.965 528.150 367.245 ;
        RECT 528.490 366.965 528.770 367.245 ;
        RECT 529.110 366.965 529.390 367.245 ;
        RECT 529.730 366.965 530.010 367.245 ;
        RECT 530.350 366.965 530.630 367.245 ;
        RECT 530.970 366.965 531.250 367.245 ;
        RECT 531.590 366.965 531.870 367.245 ;
        RECT 532.210 366.965 532.490 367.245 ;
        RECT 532.830 366.965 533.110 367.245 ;
        RECT 533.450 366.965 533.730 367.245 ;
        RECT 534.070 366.965 534.350 367.245 ;
        RECT 534.690 366.965 534.970 367.245 ;
        RECT 535.310 366.965 535.590 367.245 ;
        RECT 526.630 366.345 526.910 366.625 ;
        RECT 527.250 366.345 527.530 366.625 ;
        RECT 527.870 366.345 528.150 366.625 ;
        RECT 528.490 366.345 528.770 366.625 ;
        RECT 529.110 366.345 529.390 366.625 ;
        RECT 529.730 366.345 530.010 366.625 ;
        RECT 530.350 366.345 530.630 366.625 ;
        RECT 530.970 366.345 531.250 366.625 ;
        RECT 531.590 366.345 531.870 366.625 ;
        RECT 532.210 366.345 532.490 366.625 ;
        RECT 532.830 366.345 533.110 366.625 ;
        RECT 533.450 366.345 533.730 366.625 ;
        RECT 534.070 366.345 534.350 366.625 ;
        RECT 534.690 366.345 534.970 366.625 ;
        RECT 535.310 366.345 535.590 366.625 ;
        RECT 526.630 365.725 526.910 366.005 ;
        RECT 527.250 365.725 527.530 366.005 ;
        RECT 527.870 365.725 528.150 366.005 ;
        RECT 528.490 365.725 528.770 366.005 ;
        RECT 529.110 365.725 529.390 366.005 ;
        RECT 529.730 365.725 530.010 366.005 ;
        RECT 530.350 365.725 530.630 366.005 ;
        RECT 530.970 365.725 531.250 366.005 ;
        RECT 531.590 365.725 531.870 366.005 ;
        RECT 532.210 365.725 532.490 366.005 ;
        RECT 532.830 365.725 533.110 366.005 ;
        RECT 533.450 365.725 533.730 366.005 ;
        RECT 534.070 365.725 534.350 366.005 ;
        RECT 534.690 365.725 534.970 366.005 ;
        RECT 535.310 365.725 535.590 366.005 ;
        RECT 526.630 365.105 526.910 365.385 ;
        RECT 527.250 365.105 527.530 365.385 ;
        RECT 527.870 365.105 528.150 365.385 ;
        RECT 528.490 365.105 528.770 365.385 ;
        RECT 529.110 365.105 529.390 365.385 ;
        RECT 529.730 365.105 530.010 365.385 ;
        RECT 530.350 365.105 530.630 365.385 ;
        RECT 530.970 365.105 531.250 365.385 ;
        RECT 531.590 365.105 531.870 365.385 ;
        RECT 532.210 365.105 532.490 365.385 ;
        RECT 532.830 365.105 533.110 365.385 ;
        RECT 533.450 365.105 533.730 365.385 ;
        RECT 534.070 365.105 534.350 365.385 ;
        RECT 534.690 365.105 534.970 365.385 ;
        RECT 535.310 365.105 535.590 365.385 ;
        RECT 526.630 364.485 526.910 364.765 ;
        RECT 527.250 364.485 527.530 364.765 ;
        RECT 527.870 364.485 528.150 364.765 ;
        RECT 528.490 364.485 528.770 364.765 ;
        RECT 529.110 364.485 529.390 364.765 ;
        RECT 529.730 364.485 530.010 364.765 ;
        RECT 530.350 364.485 530.630 364.765 ;
        RECT 530.970 364.485 531.250 364.765 ;
        RECT 531.590 364.485 531.870 364.765 ;
        RECT 532.210 364.485 532.490 364.765 ;
        RECT 532.830 364.485 533.110 364.765 ;
        RECT 533.450 364.485 533.730 364.765 ;
        RECT 534.070 364.485 534.350 364.765 ;
        RECT 534.690 364.485 534.970 364.765 ;
        RECT 535.310 364.485 535.590 364.765 ;
        RECT 526.630 363.865 526.910 364.145 ;
        RECT 527.250 363.865 527.530 364.145 ;
        RECT 527.870 363.865 528.150 364.145 ;
        RECT 528.490 363.865 528.770 364.145 ;
        RECT 529.110 363.865 529.390 364.145 ;
        RECT 529.730 363.865 530.010 364.145 ;
        RECT 530.350 363.865 530.630 364.145 ;
        RECT 530.970 363.865 531.250 364.145 ;
        RECT 531.590 363.865 531.870 364.145 ;
        RECT 532.210 363.865 532.490 364.145 ;
        RECT 532.830 363.865 533.110 364.145 ;
        RECT 533.450 363.865 533.730 364.145 ;
        RECT 534.070 363.865 534.350 364.145 ;
        RECT 534.690 363.865 534.970 364.145 ;
        RECT 535.310 363.865 535.590 364.145 ;
        RECT 526.630 363.245 526.910 363.525 ;
        RECT 527.250 363.245 527.530 363.525 ;
        RECT 527.870 363.245 528.150 363.525 ;
        RECT 528.490 363.245 528.770 363.525 ;
        RECT 529.110 363.245 529.390 363.525 ;
        RECT 529.730 363.245 530.010 363.525 ;
        RECT 530.350 363.245 530.630 363.525 ;
        RECT 530.970 363.245 531.250 363.525 ;
        RECT 531.590 363.245 531.870 363.525 ;
        RECT 532.210 363.245 532.490 363.525 ;
        RECT 532.830 363.245 533.110 363.525 ;
        RECT 533.450 363.245 533.730 363.525 ;
        RECT 534.070 363.245 534.350 363.525 ;
        RECT 534.690 363.245 534.970 363.525 ;
        RECT 535.310 363.245 535.590 363.525 ;
        RECT 526.630 362.625 526.910 362.905 ;
        RECT 527.250 362.625 527.530 362.905 ;
        RECT 527.870 362.625 528.150 362.905 ;
        RECT 528.490 362.625 528.770 362.905 ;
        RECT 529.110 362.625 529.390 362.905 ;
        RECT 529.730 362.625 530.010 362.905 ;
        RECT 530.350 362.625 530.630 362.905 ;
        RECT 530.970 362.625 531.250 362.905 ;
        RECT 531.590 362.625 531.870 362.905 ;
        RECT 532.210 362.625 532.490 362.905 ;
        RECT 532.830 362.625 533.110 362.905 ;
        RECT 533.450 362.625 533.730 362.905 ;
        RECT 534.070 362.625 534.350 362.905 ;
        RECT 534.690 362.625 534.970 362.905 ;
        RECT 535.310 362.625 535.590 362.905 ;
        RECT 526.630 362.005 526.910 362.285 ;
        RECT 527.250 362.005 527.530 362.285 ;
        RECT 527.870 362.005 528.150 362.285 ;
        RECT 528.490 362.005 528.770 362.285 ;
        RECT 529.110 362.005 529.390 362.285 ;
        RECT 529.730 362.005 530.010 362.285 ;
        RECT 530.350 362.005 530.630 362.285 ;
        RECT 530.970 362.005 531.250 362.285 ;
        RECT 531.590 362.005 531.870 362.285 ;
        RECT 532.210 362.005 532.490 362.285 ;
        RECT 532.830 362.005 533.110 362.285 ;
        RECT 533.450 362.005 533.730 362.285 ;
        RECT 534.070 362.005 534.350 362.285 ;
        RECT 534.690 362.005 534.970 362.285 ;
        RECT 535.310 362.005 535.590 362.285 ;
        RECT 526.630 361.385 526.910 361.665 ;
        RECT 527.250 361.385 527.530 361.665 ;
        RECT 527.870 361.385 528.150 361.665 ;
        RECT 528.490 361.385 528.770 361.665 ;
        RECT 529.110 361.385 529.390 361.665 ;
        RECT 529.730 361.385 530.010 361.665 ;
        RECT 530.350 361.385 530.630 361.665 ;
        RECT 530.970 361.385 531.250 361.665 ;
        RECT 531.590 361.385 531.870 361.665 ;
        RECT 532.210 361.385 532.490 361.665 ;
        RECT 532.830 361.385 533.110 361.665 ;
        RECT 533.450 361.385 533.730 361.665 ;
        RECT 534.070 361.385 534.350 361.665 ;
        RECT 534.690 361.385 534.970 361.665 ;
        RECT 535.310 361.385 535.590 361.665 ;
        RECT 526.630 360.765 526.910 361.045 ;
        RECT 527.250 360.765 527.530 361.045 ;
        RECT 527.870 360.765 528.150 361.045 ;
        RECT 528.490 360.765 528.770 361.045 ;
        RECT 529.110 360.765 529.390 361.045 ;
        RECT 529.730 360.765 530.010 361.045 ;
        RECT 530.350 360.765 530.630 361.045 ;
        RECT 530.970 360.765 531.250 361.045 ;
        RECT 531.590 360.765 531.870 361.045 ;
        RECT 532.210 360.765 532.490 361.045 ;
        RECT 532.830 360.765 533.110 361.045 ;
        RECT 533.450 360.765 533.730 361.045 ;
        RECT 534.070 360.765 534.350 361.045 ;
        RECT 534.690 360.765 534.970 361.045 ;
        RECT 535.310 360.765 535.590 361.045 ;
        RECT 545.230 369.445 545.510 369.725 ;
        RECT 545.850 369.445 546.130 369.725 ;
        RECT 546.470 369.445 546.750 369.725 ;
        RECT 547.090 369.445 547.370 369.725 ;
        RECT 547.710 369.445 547.990 369.725 ;
        RECT 548.330 369.445 548.610 369.725 ;
        RECT 545.230 368.825 545.510 369.105 ;
        RECT 545.850 368.825 546.130 369.105 ;
        RECT 546.470 368.825 546.750 369.105 ;
        RECT 547.090 368.825 547.370 369.105 ;
        RECT 547.710 368.825 547.990 369.105 ;
        RECT 548.330 368.825 548.610 369.105 ;
        RECT 545.230 368.205 545.510 368.485 ;
        RECT 545.850 368.205 546.130 368.485 ;
        RECT 546.470 368.205 546.750 368.485 ;
        RECT 547.090 368.205 547.370 368.485 ;
        RECT 547.710 368.205 547.990 368.485 ;
        RECT 548.330 368.205 548.610 368.485 ;
        RECT 545.230 367.585 545.510 367.865 ;
        RECT 545.850 367.585 546.130 367.865 ;
        RECT 546.470 367.585 546.750 367.865 ;
        RECT 547.090 367.585 547.370 367.865 ;
        RECT 547.710 367.585 547.990 367.865 ;
        RECT 548.330 367.585 548.610 367.865 ;
        RECT 545.230 366.965 545.510 367.245 ;
        RECT 545.850 366.965 546.130 367.245 ;
        RECT 546.470 366.965 546.750 367.245 ;
        RECT 547.090 366.965 547.370 367.245 ;
        RECT 547.710 366.965 547.990 367.245 ;
        RECT 548.330 366.965 548.610 367.245 ;
        RECT 545.230 366.345 545.510 366.625 ;
        RECT 545.850 366.345 546.130 366.625 ;
        RECT 546.470 366.345 546.750 366.625 ;
        RECT 547.090 366.345 547.370 366.625 ;
        RECT 547.710 366.345 547.990 366.625 ;
        RECT 548.330 366.345 548.610 366.625 ;
        RECT 545.230 365.725 545.510 366.005 ;
        RECT 545.850 365.725 546.130 366.005 ;
        RECT 546.470 365.725 546.750 366.005 ;
        RECT 547.090 365.725 547.370 366.005 ;
        RECT 547.710 365.725 547.990 366.005 ;
        RECT 548.330 365.725 548.610 366.005 ;
        RECT 545.230 365.105 545.510 365.385 ;
        RECT 545.850 365.105 546.130 365.385 ;
        RECT 546.470 365.105 546.750 365.385 ;
        RECT 547.090 365.105 547.370 365.385 ;
        RECT 547.710 365.105 547.990 365.385 ;
        RECT 548.330 365.105 548.610 365.385 ;
        RECT 545.230 364.485 545.510 364.765 ;
        RECT 545.850 364.485 546.130 364.765 ;
        RECT 546.470 364.485 546.750 364.765 ;
        RECT 547.090 364.485 547.370 364.765 ;
        RECT 547.710 364.485 547.990 364.765 ;
        RECT 548.330 364.485 548.610 364.765 ;
        RECT 545.230 363.865 545.510 364.145 ;
        RECT 545.850 363.865 546.130 364.145 ;
        RECT 546.470 363.865 546.750 364.145 ;
        RECT 547.090 363.865 547.370 364.145 ;
        RECT 547.710 363.865 547.990 364.145 ;
        RECT 548.330 363.865 548.610 364.145 ;
        RECT 545.230 363.245 545.510 363.525 ;
        RECT 545.850 363.245 546.130 363.525 ;
        RECT 546.470 363.245 546.750 363.525 ;
        RECT 547.090 363.245 547.370 363.525 ;
        RECT 547.710 363.245 547.990 363.525 ;
        RECT 548.330 363.245 548.610 363.525 ;
        RECT 545.230 362.625 545.510 362.905 ;
        RECT 545.850 362.625 546.130 362.905 ;
        RECT 546.470 362.625 546.750 362.905 ;
        RECT 547.090 362.625 547.370 362.905 ;
        RECT 547.710 362.625 547.990 362.905 ;
        RECT 548.330 362.625 548.610 362.905 ;
        RECT 545.230 362.005 545.510 362.285 ;
        RECT 545.850 362.005 546.130 362.285 ;
        RECT 546.470 362.005 546.750 362.285 ;
        RECT 547.090 362.005 547.370 362.285 ;
        RECT 547.710 362.005 547.990 362.285 ;
        RECT 548.330 362.005 548.610 362.285 ;
        RECT 545.230 361.385 545.510 361.665 ;
        RECT 545.850 361.385 546.130 361.665 ;
        RECT 546.470 361.385 546.750 361.665 ;
        RECT 547.090 361.385 547.370 361.665 ;
        RECT 547.710 361.385 547.990 361.665 ;
        RECT 548.330 361.385 548.610 361.665 ;
        RECT 545.230 360.765 545.510 361.045 ;
        RECT 545.850 360.765 546.130 361.045 ;
        RECT 546.470 360.765 546.750 361.045 ;
        RECT 547.090 360.765 547.370 361.045 ;
        RECT 547.710 360.765 547.990 361.045 ;
        RECT 548.330 360.765 548.610 361.045 ;
        RECT 550.880 369.445 551.160 369.725 ;
        RECT 551.500 369.445 551.780 369.725 ;
        RECT 552.120 369.445 552.400 369.725 ;
        RECT 552.740 369.445 553.020 369.725 ;
        RECT 553.360 369.445 553.640 369.725 ;
        RECT 553.980 369.445 554.260 369.725 ;
        RECT 554.600 369.445 554.880 369.725 ;
        RECT 555.220 369.445 555.500 369.725 ;
        RECT 555.840 369.445 556.120 369.725 ;
        RECT 556.460 369.445 556.740 369.725 ;
        RECT 557.080 369.445 557.360 369.725 ;
        RECT 557.700 369.445 557.980 369.725 ;
        RECT 558.320 369.445 558.600 369.725 ;
        RECT 558.940 369.445 559.220 369.725 ;
        RECT 559.560 369.445 559.840 369.725 ;
        RECT 560.180 369.445 560.460 369.725 ;
        RECT 550.880 368.825 551.160 369.105 ;
        RECT 551.500 368.825 551.780 369.105 ;
        RECT 552.120 368.825 552.400 369.105 ;
        RECT 552.740 368.825 553.020 369.105 ;
        RECT 553.360 368.825 553.640 369.105 ;
        RECT 553.980 368.825 554.260 369.105 ;
        RECT 554.600 368.825 554.880 369.105 ;
        RECT 555.220 368.825 555.500 369.105 ;
        RECT 555.840 368.825 556.120 369.105 ;
        RECT 556.460 368.825 556.740 369.105 ;
        RECT 557.080 368.825 557.360 369.105 ;
        RECT 557.700 368.825 557.980 369.105 ;
        RECT 558.320 368.825 558.600 369.105 ;
        RECT 558.940 368.825 559.220 369.105 ;
        RECT 559.560 368.825 559.840 369.105 ;
        RECT 560.180 368.825 560.460 369.105 ;
        RECT 550.880 368.205 551.160 368.485 ;
        RECT 551.500 368.205 551.780 368.485 ;
        RECT 552.120 368.205 552.400 368.485 ;
        RECT 552.740 368.205 553.020 368.485 ;
        RECT 553.360 368.205 553.640 368.485 ;
        RECT 553.980 368.205 554.260 368.485 ;
        RECT 554.600 368.205 554.880 368.485 ;
        RECT 555.220 368.205 555.500 368.485 ;
        RECT 555.840 368.205 556.120 368.485 ;
        RECT 556.460 368.205 556.740 368.485 ;
        RECT 557.080 368.205 557.360 368.485 ;
        RECT 557.700 368.205 557.980 368.485 ;
        RECT 558.320 368.205 558.600 368.485 ;
        RECT 558.940 368.205 559.220 368.485 ;
        RECT 559.560 368.205 559.840 368.485 ;
        RECT 560.180 368.205 560.460 368.485 ;
        RECT 550.880 367.585 551.160 367.865 ;
        RECT 551.500 367.585 551.780 367.865 ;
        RECT 552.120 367.585 552.400 367.865 ;
        RECT 552.740 367.585 553.020 367.865 ;
        RECT 553.360 367.585 553.640 367.865 ;
        RECT 553.980 367.585 554.260 367.865 ;
        RECT 554.600 367.585 554.880 367.865 ;
        RECT 555.220 367.585 555.500 367.865 ;
        RECT 555.840 367.585 556.120 367.865 ;
        RECT 556.460 367.585 556.740 367.865 ;
        RECT 557.080 367.585 557.360 367.865 ;
        RECT 557.700 367.585 557.980 367.865 ;
        RECT 558.320 367.585 558.600 367.865 ;
        RECT 558.940 367.585 559.220 367.865 ;
        RECT 559.560 367.585 559.840 367.865 ;
        RECT 560.180 367.585 560.460 367.865 ;
        RECT 550.880 366.965 551.160 367.245 ;
        RECT 551.500 366.965 551.780 367.245 ;
        RECT 552.120 366.965 552.400 367.245 ;
        RECT 552.740 366.965 553.020 367.245 ;
        RECT 553.360 366.965 553.640 367.245 ;
        RECT 553.980 366.965 554.260 367.245 ;
        RECT 554.600 366.965 554.880 367.245 ;
        RECT 555.220 366.965 555.500 367.245 ;
        RECT 555.840 366.965 556.120 367.245 ;
        RECT 556.460 366.965 556.740 367.245 ;
        RECT 557.080 366.965 557.360 367.245 ;
        RECT 557.700 366.965 557.980 367.245 ;
        RECT 558.320 366.965 558.600 367.245 ;
        RECT 558.940 366.965 559.220 367.245 ;
        RECT 559.560 366.965 559.840 367.245 ;
        RECT 560.180 366.965 560.460 367.245 ;
        RECT 550.880 366.345 551.160 366.625 ;
        RECT 551.500 366.345 551.780 366.625 ;
        RECT 552.120 366.345 552.400 366.625 ;
        RECT 552.740 366.345 553.020 366.625 ;
        RECT 553.360 366.345 553.640 366.625 ;
        RECT 553.980 366.345 554.260 366.625 ;
        RECT 554.600 366.345 554.880 366.625 ;
        RECT 555.220 366.345 555.500 366.625 ;
        RECT 555.840 366.345 556.120 366.625 ;
        RECT 556.460 366.345 556.740 366.625 ;
        RECT 557.080 366.345 557.360 366.625 ;
        RECT 557.700 366.345 557.980 366.625 ;
        RECT 558.320 366.345 558.600 366.625 ;
        RECT 558.940 366.345 559.220 366.625 ;
        RECT 559.560 366.345 559.840 366.625 ;
        RECT 560.180 366.345 560.460 366.625 ;
        RECT 550.880 365.725 551.160 366.005 ;
        RECT 551.500 365.725 551.780 366.005 ;
        RECT 552.120 365.725 552.400 366.005 ;
        RECT 552.740 365.725 553.020 366.005 ;
        RECT 553.360 365.725 553.640 366.005 ;
        RECT 553.980 365.725 554.260 366.005 ;
        RECT 554.600 365.725 554.880 366.005 ;
        RECT 555.220 365.725 555.500 366.005 ;
        RECT 555.840 365.725 556.120 366.005 ;
        RECT 556.460 365.725 556.740 366.005 ;
        RECT 557.080 365.725 557.360 366.005 ;
        RECT 557.700 365.725 557.980 366.005 ;
        RECT 558.320 365.725 558.600 366.005 ;
        RECT 558.940 365.725 559.220 366.005 ;
        RECT 559.560 365.725 559.840 366.005 ;
        RECT 560.180 365.725 560.460 366.005 ;
        RECT 550.880 365.105 551.160 365.385 ;
        RECT 551.500 365.105 551.780 365.385 ;
        RECT 552.120 365.105 552.400 365.385 ;
        RECT 552.740 365.105 553.020 365.385 ;
        RECT 553.360 365.105 553.640 365.385 ;
        RECT 553.980 365.105 554.260 365.385 ;
        RECT 554.600 365.105 554.880 365.385 ;
        RECT 555.220 365.105 555.500 365.385 ;
        RECT 555.840 365.105 556.120 365.385 ;
        RECT 556.460 365.105 556.740 365.385 ;
        RECT 557.080 365.105 557.360 365.385 ;
        RECT 557.700 365.105 557.980 365.385 ;
        RECT 558.320 365.105 558.600 365.385 ;
        RECT 558.940 365.105 559.220 365.385 ;
        RECT 559.560 365.105 559.840 365.385 ;
        RECT 560.180 365.105 560.460 365.385 ;
        RECT 550.880 364.485 551.160 364.765 ;
        RECT 551.500 364.485 551.780 364.765 ;
        RECT 552.120 364.485 552.400 364.765 ;
        RECT 552.740 364.485 553.020 364.765 ;
        RECT 553.360 364.485 553.640 364.765 ;
        RECT 553.980 364.485 554.260 364.765 ;
        RECT 554.600 364.485 554.880 364.765 ;
        RECT 555.220 364.485 555.500 364.765 ;
        RECT 555.840 364.485 556.120 364.765 ;
        RECT 556.460 364.485 556.740 364.765 ;
        RECT 557.080 364.485 557.360 364.765 ;
        RECT 557.700 364.485 557.980 364.765 ;
        RECT 558.320 364.485 558.600 364.765 ;
        RECT 558.940 364.485 559.220 364.765 ;
        RECT 559.560 364.485 559.840 364.765 ;
        RECT 560.180 364.485 560.460 364.765 ;
        RECT 550.880 363.865 551.160 364.145 ;
        RECT 551.500 363.865 551.780 364.145 ;
        RECT 552.120 363.865 552.400 364.145 ;
        RECT 552.740 363.865 553.020 364.145 ;
        RECT 553.360 363.865 553.640 364.145 ;
        RECT 553.980 363.865 554.260 364.145 ;
        RECT 554.600 363.865 554.880 364.145 ;
        RECT 555.220 363.865 555.500 364.145 ;
        RECT 555.840 363.865 556.120 364.145 ;
        RECT 556.460 363.865 556.740 364.145 ;
        RECT 557.080 363.865 557.360 364.145 ;
        RECT 557.700 363.865 557.980 364.145 ;
        RECT 558.320 363.865 558.600 364.145 ;
        RECT 558.940 363.865 559.220 364.145 ;
        RECT 559.560 363.865 559.840 364.145 ;
        RECT 560.180 363.865 560.460 364.145 ;
        RECT 550.880 363.245 551.160 363.525 ;
        RECT 551.500 363.245 551.780 363.525 ;
        RECT 552.120 363.245 552.400 363.525 ;
        RECT 552.740 363.245 553.020 363.525 ;
        RECT 553.360 363.245 553.640 363.525 ;
        RECT 553.980 363.245 554.260 363.525 ;
        RECT 554.600 363.245 554.880 363.525 ;
        RECT 555.220 363.245 555.500 363.525 ;
        RECT 555.840 363.245 556.120 363.525 ;
        RECT 556.460 363.245 556.740 363.525 ;
        RECT 557.080 363.245 557.360 363.525 ;
        RECT 557.700 363.245 557.980 363.525 ;
        RECT 558.320 363.245 558.600 363.525 ;
        RECT 558.940 363.245 559.220 363.525 ;
        RECT 559.560 363.245 559.840 363.525 ;
        RECT 560.180 363.245 560.460 363.525 ;
        RECT 550.880 362.625 551.160 362.905 ;
        RECT 551.500 362.625 551.780 362.905 ;
        RECT 552.120 362.625 552.400 362.905 ;
        RECT 552.740 362.625 553.020 362.905 ;
        RECT 553.360 362.625 553.640 362.905 ;
        RECT 553.980 362.625 554.260 362.905 ;
        RECT 554.600 362.625 554.880 362.905 ;
        RECT 555.220 362.625 555.500 362.905 ;
        RECT 555.840 362.625 556.120 362.905 ;
        RECT 556.460 362.625 556.740 362.905 ;
        RECT 557.080 362.625 557.360 362.905 ;
        RECT 557.700 362.625 557.980 362.905 ;
        RECT 558.320 362.625 558.600 362.905 ;
        RECT 558.940 362.625 559.220 362.905 ;
        RECT 559.560 362.625 559.840 362.905 ;
        RECT 560.180 362.625 560.460 362.905 ;
        RECT 550.880 362.005 551.160 362.285 ;
        RECT 551.500 362.005 551.780 362.285 ;
        RECT 552.120 362.005 552.400 362.285 ;
        RECT 552.740 362.005 553.020 362.285 ;
        RECT 553.360 362.005 553.640 362.285 ;
        RECT 553.980 362.005 554.260 362.285 ;
        RECT 554.600 362.005 554.880 362.285 ;
        RECT 555.220 362.005 555.500 362.285 ;
        RECT 555.840 362.005 556.120 362.285 ;
        RECT 556.460 362.005 556.740 362.285 ;
        RECT 557.080 362.005 557.360 362.285 ;
        RECT 557.700 362.005 557.980 362.285 ;
        RECT 558.320 362.005 558.600 362.285 ;
        RECT 558.940 362.005 559.220 362.285 ;
        RECT 559.560 362.005 559.840 362.285 ;
        RECT 560.180 362.005 560.460 362.285 ;
        RECT 550.880 361.385 551.160 361.665 ;
        RECT 551.500 361.385 551.780 361.665 ;
        RECT 552.120 361.385 552.400 361.665 ;
        RECT 552.740 361.385 553.020 361.665 ;
        RECT 553.360 361.385 553.640 361.665 ;
        RECT 553.980 361.385 554.260 361.665 ;
        RECT 554.600 361.385 554.880 361.665 ;
        RECT 555.220 361.385 555.500 361.665 ;
        RECT 555.840 361.385 556.120 361.665 ;
        RECT 556.460 361.385 556.740 361.665 ;
        RECT 557.080 361.385 557.360 361.665 ;
        RECT 557.700 361.385 557.980 361.665 ;
        RECT 558.320 361.385 558.600 361.665 ;
        RECT 558.940 361.385 559.220 361.665 ;
        RECT 559.560 361.385 559.840 361.665 ;
        RECT 560.180 361.385 560.460 361.665 ;
        RECT 550.880 360.765 551.160 361.045 ;
        RECT 551.500 360.765 551.780 361.045 ;
        RECT 552.120 360.765 552.400 361.045 ;
        RECT 552.740 360.765 553.020 361.045 ;
        RECT 553.360 360.765 553.640 361.045 ;
        RECT 553.980 360.765 554.260 361.045 ;
        RECT 554.600 360.765 554.880 361.045 ;
        RECT 555.220 360.765 555.500 361.045 ;
        RECT 555.840 360.765 556.120 361.045 ;
        RECT 556.460 360.765 556.740 361.045 ;
        RECT 557.080 360.765 557.360 361.045 ;
        RECT 557.700 360.765 557.980 361.045 ;
        RECT 558.320 360.765 558.600 361.045 ;
        RECT 558.940 360.765 559.220 361.045 ;
        RECT 559.560 360.765 559.840 361.045 ;
        RECT 560.180 360.765 560.460 361.045 ;
        RECT 564.410 369.445 564.690 369.725 ;
        RECT 565.030 369.445 565.310 369.725 ;
        RECT 565.650 369.445 565.930 369.725 ;
        RECT 566.270 369.445 566.550 369.725 ;
        RECT 566.890 369.445 567.170 369.725 ;
        RECT 567.510 369.445 567.790 369.725 ;
        RECT 568.130 369.445 568.410 369.725 ;
        RECT 568.750 369.445 569.030 369.725 ;
        RECT 569.370 369.445 569.650 369.725 ;
        RECT 569.990 369.445 570.270 369.725 ;
        RECT 570.610 369.445 570.890 369.725 ;
        RECT 571.230 369.445 571.510 369.725 ;
        RECT 571.850 369.445 572.130 369.725 ;
        RECT 572.470 369.445 572.750 369.725 ;
        RECT 573.090 369.445 573.370 369.725 ;
        RECT 573.710 369.445 573.990 369.725 ;
        RECT 564.410 368.825 564.690 369.105 ;
        RECT 565.030 368.825 565.310 369.105 ;
        RECT 565.650 368.825 565.930 369.105 ;
        RECT 566.270 368.825 566.550 369.105 ;
        RECT 566.890 368.825 567.170 369.105 ;
        RECT 567.510 368.825 567.790 369.105 ;
        RECT 568.130 368.825 568.410 369.105 ;
        RECT 568.750 368.825 569.030 369.105 ;
        RECT 569.370 368.825 569.650 369.105 ;
        RECT 569.990 368.825 570.270 369.105 ;
        RECT 570.610 368.825 570.890 369.105 ;
        RECT 571.230 368.825 571.510 369.105 ;
        RECT 571.850 368.825 572.130 369.105 ;
        RECT 572.470 368.825 572.750 369.105 ;
        RECT 573.090 368.825 573.370 369.105 ;
        RECT 573.710 368.825 573.990 369.105 ;
        RECT 564.410 368.205 564.690 368.485 ;
        RECT 565.030 368.205 565.310 368.485 ;
        RECT 565.650 368.205 565.930 368.485 ;
        RECT 566.270 368.205 566.550 368.485 ;
        RECT 566.890 368.205 567.170 368.485 ;
        RECT 567.510 368.205 567.790 368.485 ;
        RECT 568.130 368.205 568.410 368.485 ;
        RECT 568.750 368.205 569.030 368.485 ;
        RECT 569.370 368.205 569.650 368.485 ;
        RECT 569.990 368.205 570.270 368.485 ;
        RECT 570.610 368.205 570.890 368.485 ;
        RECT 571.230 368.205 571.510 368.485 ;
        RECT 571.850 368.205 572.130 368.485 ;
        RECT 572.470 368.205 572.750 368.485 ;
        RECT 573.090 368.205 573.370 368.485 ;
        RECT 573.710 368.205 573.990 368.485 ;
        RECT 564.410 367.585 564.690 367.865 ;
        RECT 565.030 367.585 565.310 367.865 ;
        RECT 565.650 367.585 565.930 367.865 ;
        RECT 566.270 367.585 566.550 367.865 ;
        RECT 566.890 367.585 567.170 367.865 ;
        RECT 567.510 367.585 567.790 367.865 ;
        RECT 568.130 367.585 568.410 367.865 ;
        RECT 568.750 367.585 569.030 367.865 ;
        RECT 569.370 367.585 569.650 367.865 ;
        RECT 569.990 367.585 570.270 367.865 ;
        RECT 570.610 367.585 570.890 367.865 ;
        RECT 571.230 367.585 571.510 367.865 ;
        RECT 571.850 367.585 572.130 367.865 ;
        RECT 572.470 367.585 572.750 367.865 ;
        RECT 573.090 367.585 573.370 367.865 ;
        RECT 573.710 367.585 573.990 367.865 ;
        RECT 564.410 366.965 564.690 367.245 ;
        RECT 565.030 366.965 565.310 367.245 ;
        RECT 565.650 366.965 565.930 367.245 ;
        RECT 566.270 366.965 566.550 367.245 ;
        RECT 566.890 366.965 567.170 367.245 ;
        RECT 567.510 366.965 567.790 367.245 ;
        RECT 568.130 366.965 568.410 367.245 ;
        RECT 568.750 366.965 569.030 367.245 ;
        RECT 569.370 366.965 569.650 367.245 ;
        RECT 569.990 366.965 570.270 367.245 ;
        RECT 570.610 366.965 570.890 367.245 ;
        RECT 571.230 366.965 571.510 367.245 ;
        RECT 571.850 366.965 572.130 367.245 ;
        RECT 572.470 366.965 572.750 367.245 ;
        RECT 573.090 366.965 573.370 367.245 ;
        RECT 573.710 366.965 573.990 367.245 ;
        RECT 564.410 366.345 564.690 366.625 ;
        RECT 565.030 366.345 565.310 366.625 ;
        RECT 565.650 366.345 565.930 366.625 ;
        RECT 566.270 366.345 566.550 366.625 ;
        RECT 566.890 366.345 567.170 366.625 ;
        RECT 567.510 366.345 567.790 366.625 ;
        RECT 568.130 366.345 568.410 366.625 ;
        RECT 568.750 366.345 569.030 366.625 ;
        RECT 569.370 366.345 569.650 366.625 ;
        RECT 569.990 366.345 570.270 366.625 ;
        RECT 570.610 366.345 570.890 366.625 ;
        RECT 571.230 366.345 571.510 366.625 ;
        RECT 571.850 366.345 572.130 366.625 ;
        RECT 572.470 366.345 572.750 366.625 ;
        RECT 573.090 366.345 573.370 366.625 ;
        RECT 573.710 366.345 573.990 366.625 ;
        RECT 564.410 365.725 564.690 366.005 ;
        RECT 565.030 365.725 565.310 366.005 ;
        RECT 565.650 365.725 565.930 366.005 ;
        RECT 566.270 365.725 566.550 366.005 ;
        RECT 566.890 365.725 567.170 366.005 ;
        RECT 567.510 365.725 567.790 366.005 ;
        RECT 568.130 365.725 568.410 366.005 ;
        RECT 568.750 365.725 569.030 366.005 ;
        RECT 569.370 365.725 569.650 366.005 ;
        RECT 569.990 365.725 570.270 366.005 ;
        RECT 570.610 365.725 570.890 366.005 ;
        RECT 571.230 365.725 571.510 366.005 ;
        RECT 571.850 365.725 572.130 366.005 ;
        RECT 572.470 365.725 572.750 366.005 ;
        RECT 573.090 365.725 573.370 366.005 ;
        RECT 573.710 365.725 573.990 366.005 ;
        RECT 564.410 365.105 564.690 365.385 ;
        RECT 565.030 365.105 565.310 365.385 ;
        RECT 565.650 365.105 565.930 365.385 ;
        RECT 566.270 365.105 566.550 365.385 ;
        RECT 566.890 365.105 567.170 365.385 ;
        RECT 567.510 365.105 567.790 365.385 ;
        RECT 568.130 365.105 568.410 365.385 ;
        RECT 568.750 365.105 569.030 365.385 ;
        RECT 569.370 365.105 569.650 365.385 ;
        RECT 569.990 365.105 570.270 365.385 ;
        RECT 570.610 365.105 570.890 365.385 ;
        RECT 571.230 365.105 571.510 365.385 ;
        RECT 571.850 365.105 572.130 365.385 ;
        RECT 572.470 365.105 572.750 365.385 ;
        RECT 573.090 365.105 573.370 365.385 ;
        RECT 573.710 365.105 573.990 365.385 ;
        RECT 564.410 364.485 564.690 364.765 ;
        RECT 565.030 364.485 565.310 364.765 ;
        RECT 565.650 364.485 565.930 364.765 ;
        RECT 566.270 364.485 566.550 364.765 ;
        RECT 566.890 364.485 567.170 364.765 ;
        RECT 567.510 364.485 567.790 364.765 ;
        RECT 568.130 364.485 568.410 364.765 ;
        RECT 568.750 364.485 569.030 364.765 ;
        RECT 569.370 364.485 569.650 364.765 ;
        RECT 569.990 364.485 570.270 364.765 ;
        RECT 570.610 364.485 570.890 364.765 ;
        RECT 571.230 364.485 571.510 364.765 ;
        RECT 571.850 364.485 572.130 364.765 ;
        RECT 572.470 364.485 572.750 364.765 ;
        RECT 573.090 364.485 573.370 364.765 ;
        RECT 573.710 364.485 573.990 364.765 ;
        RECT 564.410 363.865 564.690 364.145 ;
        RECT 565.030 363.865 565.310 364.145 ;
        RECT 565.650 363.865 565.930 364.145 ;
        RECT 566.270 363.865 566.550 364.145 ;
        RECT 566.890 363.865 567.170 364.145 ;
        RECT 567.510 363.865 567.790 364.145 ;
        RECT 568.130 363.865 568.410 364.145 ;
        RECT 568.750 363.865 569.030 364.145 ;
        RECT 569.370 363.865 569.650 364.145 ;
        RECT 569.990 363.865 570.270 364.145 ;
        RECT 570.610 363.865 570.890 364.145 ;
        RECT 571.230 363.865 571.510 364.145 ;
        RECT 571.850 363.865 572.130 364.145 ;
        RECT 572.470 363.865 572.750 364.145 ;
        RECT 573.090 363.865 573.370 364.145 ;
        RECT 573.710 363.865 573.990 364.145 ;
        RECT 564.410 363.245 564.690 363.525 ;
        RECT 565.030 363.245 565.310 363.525 ;
        RECT 565.650 363.245 565.930 363.525 ;
        RECT 566.270 363.245 566.550 363.525 ;
        RECT 566.890 363.245 567.170 363.525 ;
        RECT 567.510 363.245 567.790 363.525 ;
        RECT 568.130 363.245 568.410 363.525 ;
        RECT 568.750 363.245 569.030 363.525 ;
        RECT 569.370 363.245 569.650 363.525 ;
        RECT 569.990 363.245 570.270 363.525 ;
        RECT 570.610 363.245 570.890 363.525 ;
        RECT 571.230 363.245 571.510 363.525 ;
        RECT 571.850 363.245 572.130 363.525 ;
        RECT 572.470 363.245 572.750 363.525 ;
        RECT 573.090 363.245 573.370 363.525 ;
        RECT 573.710 363.245 573.990 363.525 ;
        RECT 564.410 362.625 564.690 362.905 ;
        RECT 565.030 362.625 565.310 362.905 ;
        RECT 565.650 362.625 565.930 362.905 ;
        RECT 566.270 362.625 566.550 362.905 ;
        RECT 566.890 362.625 567.170 362.905 ;
        RECT 567.510 362.625 567.790 362.905 ;
        RECT 568.130 362.625 568.410 362.905 ;
        RECT 568.750 362.625 569.030 362.905 ;
        RECT 569.370 362.625 569.650 362.905 ;
        RECT 569.990 362.625 570.270 362.905 ;
        RECT 570.610 362.625 570.890 362.905 ;
        RECT 571.230 362.625 571.510 362.905 ;
        RECT 571.850 362.625 572.130 362.905 ;
        RECT 572.470 362.625 572.750 362.905 ;
        RECT 573.090 362.625 573.370 362.905 ;
        RECT 573.710 362.625 573.990 362.905 ;
        RECT 564.410 362.005 564.690 362.285 ;
        RECT 565.030 362.005 565.310 362.285 ;
        RECT 565.650 362.005 565.930 362.285 ;
        RECT 566.270 362.005 566.550 362.285 ;
        RECT 566.890 362.005 567.170 362.285 ;
        RECT 567.510 362.005 567.790 362.285 ;
        RECT 568.130 362.005 568.410 362.285 ;
        RECT 568.750 362.005 569.030 362.285 ;
        RECT 569.370 362.005 569.650 362.285 ;
        RECT 569.990 362.005 570.270 362.285 ;
        RECT 570.610 362.005 570.890 362.285 ;
        RECT 571.230 362.005 571.510 362.285 ;
        RECT 571.850 362.005 572.130 362.285 ;
        RECT 572.470 362.005 572.750 362.285 ;
        RECT 573.090 362.005 573.370 362.285 ;
        RECT 573.710 362.005 573.990 362.285 ;
        RECT 564.410 361.385 564.690 361.665 ;
        RECT 565.030 361.385 565.310 361.665 ;
        RECT 565.650 361.385 565.930 361.665 ;
        RECT 566.270 361.385 566.550 361.665 ;
        RECT 566.890 361.385 567.170 361.665 ;
        RECT 567.510 361.385 567.790 361.665 ;
        RECT 568.130 361.385 568.410 361.665 ;
        RECT 568.750 361.385 569.030 361.665 ;
        RECT 569.370 361.385 569.650 361.665 ;
        RECT 569.990 361.385 570.270 361.665 ;
        RECT 570.610 361.385 570.890 361.665 ;
        RECT 571.230 361.385 571.510 361.665 ;
        RECT 571.850 361.385 572.130 361.665 ;
        RECT 572.470 361.385 572.750 361.665 ;
        RECT 573.090 361.385 573.370 361.665 ;
        RECT 573.710 361.385 573.990 361.665 ;
        RECT 564.410 360.765 564.690 361.045 ;
        RECT 565.030 360.765 565.310 361.045 ;
        RECT 565.650 360.765 565.930 361.045 ;
        RECT 566.270 360.765 566.550 361.045 ;
        RECT 566.890 360.765 567.170 361.045 ;
        RECT 567.510 360.765 567.790 361.045 ;
        RECT 568.130 360.765 568.410 361.045 ;
        RECT 568.750 360.765 569.030 361.045 ;
        RECT 569.370 360.765 569.650 361.045 ;
        RECT 569.990 360.765 570.270 361.045 ;
        RECT 570.610 360.765 570.890 361.045 ;
        RECT 571.230 360.765 571.510 361.045 ;
        RECT 571.850 360.765 572.130 361.045 ;
        RECT 572.470 360.765 572.750 361.045 ;
        RECT 573.090 360.765 573.370 361.045 ;
        RECT 573.710 360.765 573.990 361.045 ;
        RECT 576.260 369.445 576.540 369.725 ;
        RECT 576.880 369.445 577.160 369.725 ;
        RECT 577.500 369.445 577.780 369.725 ;
        RECT 578.120 369.445 578.400 369.725 ;
        RECT 578.740 369.445 579.020 369.725 ;
        RECT 579.360 369.445 579.640 369.725 ;
        RECT 579.980 369.445 580.260 369.725 ;
        RECT 580.600 369.445 580.880 369.725 ;
        RECT 581.220 369.445 581.500 369.725 ;
        RECT 581.840 369.445 582.120 369.725 ;
        RECT 582.460 369.445 582.740 369.725 ;
        RECT 583.080 369.445 583.360 369.725 ;
        RECT 583.700 369.445 583.980 369.725 ;
        RECT 584.320 369.445 584.600 369.725 ;
        RECT 584.940 369.445 585.220 369.725 ;
        RECT 585.560 369.445 585.840 369.725 ;
        RECT 576.260 368.825 576.540 369.105 ;
        RECT 576.880 368.825 577.160 369.105 ;
        RECT 577.500 368.825 577.780 369.105 ;
        RECT 578.120 368.825 578.400 369.105 ;
        RECT 578.740 368.825 579.020 369.105 ;
        RECT 579.360 368.825 579.640 369.105 ;
        RECT 579.980 368.825 580.260 369.105 ;
        RECT 580.600 368.825 580.880 369.105 ;
        RECT 581.220 368.825 581.500 369.105 ;
        RECT 581.840 368.825 582.120 369.105 ;
        RECT 582.460 368.825 582.740 369.105 ;
        RECT 583.080 368.825 583.360 369.105 ;
        RECT 583.700 368.825 583.980 369.105 ;
        RECT 584.320 368.825 584.600 369.105 ;
        RECT 584.940 368.825 585.220 369.105 ;
        RECT 585.560 368.825 585.840 369.105 ;
        RECT 576.260 368.205 576.540 368.485 ;
        RECT 576.880 368.205 577.160 368.485 ;
        RECT 577.500 368.205 577.780 368.485 ;
        RECT 578.120 368.205 578.400 368.485 ;
        RECT 578.740 368.205 579.020 368.485 ;
        RECT 579.360 368.205 579.640 368.485 ;
        RECT 579.980 368.205 580.260 368.485 ;
        RECT 580.600 368.205 580.880 368.485 ;
        RECT 581.220 368.205 581.500 368.485 ;
        RECT 581.840 368.205 582.120 368.485 ;
        RECT 582.460 368.205 582.740 368.485 ;
        RECT 583.080 368.205 583.360 368.485 ;
        RECT 583.700 368.205 583.980 368.485 ;
        RECT 584.320 368.205 584.600 368.485 ;
        RECT 584.940 368.205 585.220 368.485 ;
        RECT 585.560 368.205 585.840 368.485 ;
        RECT 576.260 367.585 576.540 367.865 ;
        RECT 576.880 367.585 577.160 367.865 ;
        RECT 577.500 367.585 577.780 367.865 ;
        RECT 578.120 367.585 578.400 367.865 ;
        RECT 578.740 367.585 579.020 367.865 ;
        RECT 579.360 367.585 579.640 367.865 ;
        RECT 579.980 367.585 580.260 367.865 ;
        RECT 580.600 367.585 580.880 367.865 ;
        RECT 581.220 367.585 581.500 367.865 ;
        RECT 581.840 367.585 582.120 367.865 ;
        RECT 582.460 367.585 582.740 367.865 ;
        RECT 583.080 367.585 583.360 367.865 ;
        RECT 583.700 367.585 583.980 367.865 ;
        RECT 584.320 367.585 584.600 367.865 ;
        RECT 584.940 367.585 585.220 367.865 ;
        RECT 585.560 367.585 585.840 367.865 ;
        RECT 576.260 366.965 576.540 367.245 ;
        RECT 576.880 366.965 577.160 367.245 ;
        RECT 577.500 366.965 577.780 367.245 ;
        RECT 578.120 366.965 578.400 367.245 ;
        RECT 578.740 366.965 579.020 367.245 ;
        RECT 579.360 366.965 579.640 367.245 ;
        RECT 579.980 366.965 580.260 367.245 ;
        RECT 580.600 366.965 580.880 367.245 ;
        RECT 581.220 366.965 581.500 367.245 ;
        RECT 581.840 366.965 582.120 367.245 ;
        RECT 582.460 366.965 582.740 367.245 ;
        RECT 583.080 366.965 583.360 367.245 ;
        RECT 583.700 366.965 583.980 367.245 ;
        RECT 584.320 366.965 584.600 367.245 ;
        RECT 584.940 366.965 585.220 367.245 ;
        RECT 585.560 366.965 585.840 367.245 ;
        RECT 576.260 366.345 576.540 366.625 ;
        RECT 576.880 366.345 577.160 366.625 ;
        RECT 577.500 366.345 577.780 366.625 ;
        RECT 578.120 366.345 578.400 366.625 ;
        RECT 578.740 366.345 579.020 366.625 ;
        RECT 579.360 366.345 579.640 366.625 ;
        RECT 579.980 366.345 580.260 366.625 ;
        RECT 580.600 366.345 580.880 366.625 ;
        RECT 581.220 366.345 581.500 366.625 ;
        RECT 581.840 366.345 582.120 366.625 ;
        RECT 582.460 366.345 582.740 366.625 ;
        RECT 583.080 366.345 583.360 366.625 ;
        RECT 583.700 366.345 583.980 366.625 ;
        RECT 584.320 366.345 584.600 366.625 ;
        RECT 584.940 366.345 585.220 366.625 ;
        RECT 585.560 366.345 585.840 366.625 ;
        RECT 576.260 365.725 576.540 366.005 ;
        RECT 576.880 365.725 577.160 366.005 ;
        RECT 577.500 365.725 577.780 366.005 ;
        RECT 578.120 365.725 578.400 366.005 ;
        RECT 578.740 365.725 579.020 366.005 ;
        RECT 579.360 365.725 579.640 366.005 ;
        RECT 579.980 365.725 580.260 366.005 ;
        RECT 580.600 365.725 580.880 366.005 ;
        RECT 581.220 365.725 581.500 366.005 ;
        RECT 581.840 365.725 582.120 366.005 ;
        RECT 582.460 365.725 582.740 366.005 ;
        RECT 583.080 365.725 583.360 366.005 ;
        RECT 583.700 365.725 583.980 366.005 ;
        RECT 584.320 365.725 584.600 366.005 ;
        RECT 584.940 365.725 585.220 366.005 ;
        RECT 585.560 365.725 585.840 366.005 ;
        RECT 576.260 365.105 576.540 365.385 ;
        RECT 576.880 365.105 577.160 365.385 ;
        RECT 577.500 365.105 577.780 365.385 ;
        RECT 578.120 365.105 578.400 365.385 ;
        RECT 578.740 365.105 579.020 365.385 ;
        RECT 579.360 365.105 579.640 365.385 ;
        RECT 579.980 365.105 580.260 365.385 ;
        RECT 580.600 365.105 580.880 365.385 ;
        RECT 581.220 365.105 581.500 365.385 ;
        RECT 581.840 365.105 582.120 365.385 ;
        RECT 582.460 365.105 582.740 365.385 ;
        RECT 583.080 365.105 583.360 365.385 ;
        RECT 583.700 365.105 583.980 365.385 ;
        RECT 584.320 365.105 584.600 365.385 ;
        RECT 584.940 365.105 585.220 365.385 ;
        RECT 585.560 365.105 585.840 365.385 ;
        RECT 576.260 364.485 576.540 364.765 ;
        RECT 576.880 364.485 577.160 364.765 ;
        RECT 577.500 364.485 577.780 364.765 ;
        RECT 578.120 364.485 578.400 364.765 ;
        RECT 578.740 364.485 579.020 364.765 ;
        RECT 579.360 364.485 579.640 364.765 ;
        RECT 579.980 364.485 580.260 364.765 ;
        RECT 580.600 364.485 580.880 364.765 ;
        RECT 581.220 364.485 581.500 364.765 ;
        RECT 581.840 364.485 582.120 364.765 ;
        RECT 582.460 364.485 582.740 364.765 ;
        RECT 583.080 364.485 583.360 364.765 ;
        RECT 583.700 364.485 583.980 364.765 ;
        RECT 584.320 364.485 584.600 364.765 ;
        RECT 584.940 364.485 585.220 364.765 ;
        RECT 585.560 364.485 585.840 364.765 ;
        RECT 576.260 363.865 576.540 364.145 ;
        RECT 576.880 363.865 577.160 364.145 ;
        RECT 577.500 363.865 577.780 364.145 ;
        RECT 578.120 363.865 578.400 364.145 ;
        RECT 578.740 363.865 579.020 364.145 ;
        RECT 579.360 363.865 579.640 364.145 ;
        RECT 579.980 363.865 580.260 364.145 ;
        RECT 580.600 363.865 580.880 364.145 ;
        RECT 581.220 363.865 581.500 364.145 ;
        RECT 581.840 363.865 582.120 364.145 ;
        RECT 582.460 363.865 582.740 364.145 ;
        RECT 583.080 363.865 583.360 364.145 ;
        RECT 583.700 363.865 583.980 364.145 ;
        RECT 584.320 363.865 584.600 364.145 ;
        RECT 584.940 363.865 585.220 364.145 ;
        RECT 585.560 363.865 585.840 364.145 ;
        RECT 576.260 363.245 576.540 363.525 ;
        RECT 576.880 363.245 577.160 363.525 ;
        RECT 577.500 363.245 577.780 363.525 ;
        RECT 578.120 363.245 578.400 363.525 ;
        RECT 578.740 363.245 579.020 363.525 ;
        RECT 579.360 363.245 579.640 363.525 ;
        RECT 579.980 363.245 580.260 363.525 ;
        RECT 580.600 363.245 580.880 363.525 ;
        RECT 581.220 363.245 581.500 363.525 ;
        RECT 581.840 363.245 582.120 363.525 ;
        RECT 582.460 363.245 582.740 363.525 ;
        RECT 583.080 363.245 583.360 363.525 ;
        RECT 583.700 363.245 583.980 363.525 ;
        RECT 584.320 363.245 584.600 363.525 ;
        RECT 584.940 363.245 585.220 363.525 ;
        RECT 585.560 363.245 585.840 363.525 ;
        RECT 576.260 362.625 576.540 362.905 ;
        RECT 576.880 362.625 577.160 362.905 ;
        RECT 577.500 362.625 577.780 362.905 ;
        RECT 578.120 362.625 578.400 362.905 ;
        RECT 578.740 362.625 579.020 362.905 ;
        RECT 579.360 362.625 579.640 362.905 ;
        RECT 579.980 362.625 580.260 362.905 ;
        RECT 580.600 362.625 580.880 362.905 ;
        RECT 581.220 362.625 581.500 362.905 ;
        RECT 581.840 362.625 582.120 362.905 ;
        RECT 582.460 362.625 582.740 362.905 ;
        RECT 583.080 362.625 583.360 362.905 ;
        RECT 583.700 362.625 583.980 362.905 ;
        RECT 584.320 362.625 584.600 362.905 ;
        RECT 584.940 362.625 585.220 362.905 ;
        RECT 585.560 362.625 585.840 362.905 ;
        RECT 576.260 362.005 576.540 362.285 ;
        RECT 576.880 362.005 577.160 362.285 ;
        RECT 577.500 362.005 577.780 362.285 ;
        RECT 578.120 362.005 578.400 362.285 ;
        RECT 578.740 362.005 579.020 362.285 ;
        RECT 579.360 362.005 579.640 362.285 ;
        RECT 579.980 362.005 580.260 362.285 ;
        RECT 580.600 362.005 580.880 362.285 ;
        RECT 581.220 362.005 581.500 362.285 ;
        RECT 581.840 362.005 582.120 362.285 ;
        RECT 582.460 362.005 582.740 362.285 ;
        RECT 583.080 362.005 583.360 362.285 ;
        RECT 583.700 362.005 583.980 362.285 ;
        RECT 584.320 362.005 584.600 362.285 ;
        RECT 584.940 362.005 585.220 362.285 ;
        RECT 585.560 362.005 585.840 362.285 ;
        RECT 576.260 361.385 576.540 361.665 ;
        RECT 576.880 361.385 577.160 361.665 ;
        RECT 577.500 361.385 577.780 361.665 ;
        RECT 578.120 361.385 578.400 361.665 ;
        RECT 578.740 361.385 579.020 361.665 ;
        RECT 579.360 361.385 579.640 361.665 ;
        RECT 579.980 361.385 580.260 361.665 ;
        RECT 580.600 361.385 580.880 361.665 ;
        RECT 581.220 361.385 581.500 361.665 ;
        RECT 581.840 361.385 582.120 361.665 ;
        RECT 582.460 361.385 582.740 361.665 ;
        RECT 583.080 361.385 583.360 361.665 ;
        RECT 583.700 361.385 583.980 361.665 ;
        RECT 584.320 361.385 584.600 361.665 ;
        RECT 584.940 361.385 585.220 361.665 ;
        RECT 585.560 361.385 585.840 361.665 ;
        RECT 576.260 360.765 576.540 361.045 ;
        RECT 576.880 360.765 577.160 361.045 ;
        RECT 577.500 360.765 577.780 361.045 ;
        RECT 578.120 360.765 578.400 361.045 ;
        RECT 578.740 360.765 579.020 361.045 ;
        RECT 579.360 360.765 579.640 361.045 ;
        RECT 579.980 360.765 580.260 361.045 ;
        RECT 580.600 360.765 580.880 361.045 ;
        RECT 581.220 360.765 581.500 361.045 ;
        RECT 581.840 360.765 582.120 361.045 ;
        RECT 582.460 360.765 582.740 361.045 ;
        RECT 583.080 360.765 583.360 361.045 ;
        RECT 583.700 360.765 583.980 361.045 ;
        RECT 584.320 360.765 584.600 361.045 ;
        RECT 584.940 360.765 585.220 361.045 ;
        RECT 585.560 360.765 585.840 361.045 ;
        RECT 589.410 369.445 589.690 369.725 ;
        RECT 590.030 369.445 590.310 369.725 ;
        RECT 590.650 369.445 590.930 369.725 ;
        RECT 591.270 369.445 591.550 369.725 ;
        RECT 591.890 369.445 592.170 369.725 ;
        RECT 592.510 369.445 592.790 369.725 ;
        RECT 593.130 369.445 593.410 369.725 ;
        RECT 593.750 369.445 594.030 369.725 ;
        RECT 594.370 369.445 594.650 369.725 ;
        RECT 594.990 369.445 595.270 369.725 ;
        RECT 595.610 369.445 595.890 369.725 ;
        RECT 596.230 369.445 596.510 369.725 ;
        RECT 596.850 369.445 597.130 369.725 ;
        RECT 597.470 369.445 597.750 369.725 ;
        RECT 598.090 369.445 598.370 369.725 ;
        RECT 589.410 368.825 589.690 369.105 ;
        RECT 590.030 368.825 590.310 369.105 ;
        RECT 590.650 368.825 590.930 369.105 ;
        RECT 591.270 368.825 591.550 369.105 ;
        RECT 591.890 368.825 592.170 369.105 ;
        RECT 592.510 368.825 592.790 369.105 ;
        RECT 593.130 368.825 593.410 369.105 ;
        RECT 593.750 368.825 594.030 369.105 ;
        RECT 594.370 368.825 594.650 369.105 ;
        RECT 594.990 368.825 595.270 369.105 ;
        RECT 595.610 368.825 595.890 369.105 ;
        RECT 596.230 368.825 596.510 369.105 ;
        RECT 596.850 368.825 597.130 369.105 ;
        RECT 597.470 368.825 597.750 369.105 ;
        RECT 598.090 368.825 598.370 369.105 ;
        RECT 589.410 368.205 589.690 368.485 ;
        RECT 590.030 368.205 590.310 368.485 ;
        RECT 590.650 368.205 590.930 368.485 ;
        RECT 591.270 368.205 591.550 368.485 ;
        RECT 591.890 368.205 592.170 368.485 ;
        RECT 592.510 368.205 592.790 368.485 ;
        RECT 593.130 368.205 593.410 368.485 ;
        RECT 593.750 368.205 594.030 368.485 ;
        RECT 594.370 368.205 594.650 368.485 ;
        RECT 594.990 368.205 595.270 368.485 ;
        RECT 595.610 368.205 595.890 368.485 ;
        RECT 596.230 368.205 596.510 368.485 ;
        RECT 596.850 368.205 597.130 368.485 ;
        RECT 597.470 368.205 597.750 368.485 ;
        RECT 598.090 368.205 598.370 368.485 ;
        RECT 589.410 367.585 589.690 367.865 ;
        RECT 590.030 367.585 590.310 367.865 ;
        RECT 590.650 367.585 590.930 367.865 ;
        RECT 591.270 367.585 591.550 367.865 ;
        RECT 591.890 367.585 592.170 367.865 ;
        RECT 592.510 367.585 592.790 367.865 ;
        RECT 593.130 367.585 593.410 367.865 ;
        RECT 593.750 367.585 594.030 367.865 ;
        RECT 594.370 367.585 594.650 367.865 ;
        RECT 594.990 367.585 595.270 367.865 ;
        RECT 595.610 367.585 595.890 367.865 ;
        RECT 596.230 367.585 596.510 367.865 ;
        RECT 596.850 367.585 597.130 367.865 ;
        RECT 597.470 367.585 597.750 367.865 ;
        RECT 598.090 367.585 598.370 367.865 ;
        RECT 589.410 366.965 589.690 367.245 ;
        RECT 590.030 366.965 590.310 367.245 ;
        RECT 590.650 366.965 590.930 367.245 ;
        RECT 591.270 366.965 591.550 367.245 ;
        RECT 591.890 366.965 592.170 367.245 ;
        RECT 592.510 366.965 592.790 367.245 ;
        RECT 593.130 366.965 593.410 367.245 ;
        RECT 593.750 366.965 594.030 367.245 ;
        RECT 594.370 366.965 594.650 367.245 ;
        RECT 594.990 366.965 595.270 367.245 ;
        RECT 595.610 366.965 595.890 367.245 ;
        RECT 596.230 366.965 596.510 367.245 ;
        RECT 596.850 366.965 597.130 367.245 ;
        RECT 597.470 366.965 597.750 367.245 ;
        RECT 598.090 366.965 598.370 367.245 ;
        RECT 589.410 366.345 589.690 366.625 ;
        RECT 590.030 366.345 590.310 366.625 ;
        RECT 590.650 366.345 590.930 366.625 ;
        RECT 591.270 366.345 591.550 366.625 ;
        RECT 591.890 366.345 592.170 366.625 ;
        RECT 592.510 366.345 592.790 366.625 ;
        RECT 593.130 366.345 593.410 366.625 ;
        RECT 593.750 366.345 594.030 366.625 ;
        RECT 594.370 366.345 594.650 366.625 ;
        RECT 594.990 366.345 595.270 366.625 ;
        RECT 595.610 366.345 595.890 366.625 ;
        RECT 596.230 366.345 596.510 366.625 ;
        RECT 596.850 366.345 597.130 366.625 ;
        RECT 597.470 366.345 597.750 366.625 ;
        RECT 598.090 366.345 598.370 366.625 ;
        RECT 589.410 365.725 589.690 366.005 ;
        RECT 590.030 365.725 590.310 366.005 ;
        RECT 590.650 365.725 590.930 366.005 ;
        RECT 591.270 365.725 591.550 366.005 ;
        RECT 591.890 365.725 592.170 366.005 ;
        RECT 592.510 365.725 592.790 366.005 ;
        RECT 593.130 365.725 593.410 366.005 ;
        RECT 593.750 365.725 594.030 366.005 ;
        RECT 594.370 365.725 594.650 366.005 ;
        RECT 594.990 365.725 595.270 366.005 ;
        RECT 595.610 365.725 595.890 366.005 ;
        RECT 596.230 365.725 596.510 366.005 ;
        RECT 596.850 365.725 597.130 366.005 ;
        RECT 597.470 365.725 597.750 366.005 ;
        RECT 598.090 365.725 598.370 366.005 ;
        RECT 589.410 365.105 589.690 365.385 ;
        RECT 590.030 365.105 590.310 365.385 ;
        RECT 590.650 365.105 590.930 365.385 ;
        RECT 591.270 365.105 591.550 365.385 ;
        RECT 591.890 365.105 592.170 365.385 ;
        RECT 592.510 365.105 592.790 365.385 ;
        RECT 593.130 365.105 593.410 365.385 ;
        RECT 593.750 365.105 594.030 365.385 ;
        RECT 594.370 365.105 594.650 365.385 ;
        RECT 594.990 365.105 595.270 365.385 ;
        RECT 595.610 365.105 595.890 365.385 ;
        RECT 596.230 365.105 596.510 365.385 ;
        RECT 596.850 365.105 597.130 365.385 ;
        RECT 597.470 365.105 597.750 365.385 ;
        RECT 598.090 365.105 598.370 365.385 ;
        RECT 589.410 364.485 589.690 364.765 ;
        RECT 590.030 364.485 590.310 364.765 ;
        RECT 590.650 364.485 590.930 364.765 ;
        RECT 591.270 364.485 591.550 364.765 ;
        RECT 591.890 364.485 592.170 364.765 ;
        RECT 592.510 364.485 592.790 364.765 ;
        RECT 593.130 364.485 593.410 364.765 ;
        RECT 593.750 364.485 594.030 364.765 ;
        RECT 594.370 364.485 594.650 364.765 ;
        RECT 594.990 364.485 595.270 364.765 ;
        RECT 595.610 364.485 595.890 364.765 ;
        RECT 596.230 364.485 596.510 364.765 ;
        RECT 596.850 364.485 597.130 364.765 ;
        RECT 597.470 364.485 597.750 364.765 ;
        RECT 598.090 364.485 598.370 364.765 ;
        RECT 589.410 363.865 589.690 364.145 ;
        RECT 590.030 363.865 590.310 364.145 ;
        RECT 590.650 363.865 590.930 364.145 ;
        RECT 591.270 363.865 591.550 364.145 ;
        RECT 591.890 363.865 592.170 364.145 ;
        RECT 592.510 363.865 592.790 364.145 ;
        RECT 593.130 363.865 593.410 364.145 ;
        RECT 593.750 363.865 594.030 364.145 ;
        RECT 594.370 363.865 594.650 364.145 ;
        RECT 594.990 363.865 595.270 364.145 ;
        RECT 595.610 363.865 595.890 364.145 ;
        RECT 596.230 363.865 596.510 364.145 ;
        RECT 596.850 363.865 597.130 364.145 ;
        RECT 597.470 363.865 597.750 364.145 ;
        RECT 598.090 363.865 598.370 364.145 ;
        RECT 589.410 363.245 589.690 363.525 ;
        RECT 590.030 363.245 590.310 363.525 ;
        RECT 590.650 363.245 590.930 363.525 ;
        RECT 591.270 363.245 591.550 363.525 ;
        RECT 591.890 363.245 592.170 363.525 ;
        RECT 592.510 363.245 592.790 363.525 ;
        RECT 593.130 363.245 593.410 363.525 ;
        RECT 593.750 363.245 594.030 363.525 ;
        RECT 594.370 363.245 594.650 363.525 ;
        RECT 594.990 363.245 595.270 363.525 ;
        RECT 595.610 363.245 595.890 363.525 ;
        RECT 596.230 363.245 596.510 363.525 ;
        RECT 596.850 363.245 597.130 363.525 ;
        RECT 597.470 363.245 597.750 363.525 ;
        RECT 598.090 363.245 598.370 363.525 ;
        RECT 589.410 362.625 589.690 362.905 ;
        RECT 590.030 362.625 590.310 362.905 ;
        RECT 590.650 362.625 590.930 362.905 ;
        RECT 591.270 362.625 591.550 362.905 ;
        RECT 591.890 362.625 592.170 362.905 ;
        RECT 592.510 362.625 592.790 362.905 ;
        RECT 593.130 362.625 593.410 362.905 ;
        RECT 593.750 362.625 594.030 362.905 ;
        RECT 594.370 362.625 594.650 362.905 ;
        RECT 594.990 362.625 595.270 362.905 ;
        RECT 595.610 362.625 595.890 362.905 ;
        RECT 596.230 362.625 596.510 362.905 ;
        RECT 596.850 362.625 597.130 362.905 ;
        RECT 597.470 362.625 597.750 362.905 ;
        RECT 598.090 362.625 598.370 362.905 ;
        RECT 589.410 362.005 589.690 362.285 ;
        RECT 590.030 362.005 590.310 362.285 ;
        RECT 590.650 362.005 590.930 362.285 ;
        RECT 591.270 362.005 591.550 362.285 ;
        RECT 591.890 362.005 592.170 362.285 ;
        RECT 592.510 362.005 592.790 362.285 ;
        RECT 593.130 362.005 593.410 362.285 ;
        RECT 593.750 362.005 594.030 362.285 ;
        RECT 594.370 362.005 594.650 362.285 ;
        RECT 594.990 362.005 595.270 362.285 ;
        RECT 595.610 362.005 595.890 362.285 ;
        RECT 596.230 362.005 596.510 362.285 ;
        RECT 596.850 362.005 597.130 362.285 ;
        RECT 597.470 362.005 597.750 362.285 ;
        RECT 598.090 362.005 598.370 362.285 ;
        RECT 589.410 361.385 589.690 361.665 ;
        RECT 590.030 361.385 590.310 361.665 ;
        RECT 590.650 361.385 590.930 361.665 ;
        RECT 591.270 361.385 591.550 361.665 ;
        RECT 591.890 361.385 592.170 361.665 ;
        RECT 592.510 361.385 592.790 361.665 ;
        RECT 593.130 361.385 593.410 361.665 ;
        RECT 593.750 361.385 594.030 361.665 ;
        RECT 594.370 361.385 594.650 361.665 ;
        RECT 594.990 361.385 595.270 361.665 ;
        RECT 595.610 361.385 595.890 361.665 ;
        RECT 596.230 361.385 596.510 361.665 ;
        RECT 596.850 361.385 597.130 361.665 ;
        RECT 597.470 361.385 597.750 361.665 ;
        RECT 598.090 361.385 598.370 361.665 ;
        RECT 589.410 360.765 589.690 361.045 ;
        RECT 590.030 360.765 590.310 361.045 ;
        RECT 590.650 360.765 590.930 361.045 ;
        RECT 591.270 360.765 591.550 361.045 ;
        RECT 591.890 360.765 592.170 361.045 ;
        RECT 592.510 360.765 592.790 361.045 ;
        RECT 593.130 360.765 593.410 361.045 ;
        RECT 593.750 360.765 594.030 361.045 ;
        RECT 594.370 360.765 594.650 361.045 ;
        RECT 594.990 360.765 595.270 361.045 ;
        RECT 595.610 360.765 595.890 361.045 ;
        RECT 596.230 360.765 596.510 361.045 ;
        RECT 596.850 360.765 597.130 361.045 ;
        RECT 597.470 360.765 597.750 361.045 ;
        RECT 598.090 360.765 598.370 361.045 ;
        RECT 1351.630 369.445 1351.910 369.725 ;
        RECT 1352.250 369.445 1352.530 369.725 ;
        RECT 1352.870 369.445 1353.150 369.725 ;
        RECT 1353.490 369.445 1353.770 369.725 ;
        RECT 1354.110 369.445 1354.390 369.725 ;
        RECT 1354.730 369.445 1355.010 369.725 ;
        RECT 1355.350 369.445 1355.630 369.725 ;
        RECT 1355.970 369.445 1356.250 369.725 ;
        RECT 1356.590 369.445 1356.870 369.725 ;
        RECT 1357.210 369.445 1357.490 369.725 ;
        RECT 1357.830 369.445 1358.110 369.725 ;
        RECT 1358.450 369.445 1358.730 369.725 ;
        RECT 1359.070 369.445 1359.350 369.725 ;
        RECT 1359.690 369.445 1359.970 369.725 ;
        RECT 1360.310 369.445 1360.590 369.725 ;
        RECT 1351.630 368.825 1351.910 369.105 ;
        RECT 1352.250 368.825 1352.530 369.105 ;
        RECT 1352.870 368.825 1353.150 369.105 ;
        RECT 1353.490 368.825 1353.770 369.105 ;
        RECT 1354.110 368.825 1354.390 369.105 ;
        RECT 1354.730 368.825 1355.010 369.105 ;
        RECT 1355.350 368.825 1355.630 369.105 ;
        RECT 1355.970 368.825 1356.250 369.105 ;
        RECT 1356.590 368.825 1356.870 369.105 ;
        RECT 1357.210 368.825 1357.490 369.105 ;
        RECT 1357.830 368.825 1358.110 369.105 ;
        RECT 1358.450 368.825 1358.730 369.105 ;
        RECT 1359.070 368.825 1359.350 369.105 ;
        RECT 1359.690 368.825 1359.970 369.105 ;
        RECT 1360.310 368.825 1360.590 369.105 ;
        RECT 1351.630 368.205 1351.910 368.485 ;
        RECT 1352.250 368.205 1352.530 368.485 ;
        RECT 1352.870 368.205 1353.150 368.485 ;
        RECT 1353.490 368.205 1353.770 368.485 ;
        RECT 1354.110 368.205 1354.390 368.485 ;
        RECT 1354.730 368.205 1355.010 368.485 ;
        RECT 1355.350 368.205 1355.630 368.485 ;
        RECT 1355.970 368.205 1356.250 368.485 ;
        RECT 1356.590 368.205 1356.870 368.485 ;
        RECT 1357.210 368.205 1357.490 368.485 ;
        RECT 1357.830 368.205 1358.110 368.485 ;
        RECT 1358.450 368.205 1358.730 368.485 ;
        RECT 1359.070 368.205 1359.350 368.485 ;
        RECT 1359.690 368.205 1359.970 368.485 ;
        RECT 1360.310 368.205 1360.590 368.485 ;
        RECT 1351.630 367.585 1351.910 367.865 ;
        RECT 1352.250 367.585 1352.530 367.865 ;
        RECT 1352.870 367.585 1353.150 367.865 ;
        RECT 1353.490 367.585 1353.770 367.865 ;
        RECT 1354.110 367.585 1354.390 367.865 ;
        RECT 1354.730 367.585 1355.010 367.865 ;
        RECT 1355.350 367.585 1355.630 367.865 ;
        RECT 1355.970 367.585 1356.250 367.865 ;
        RECT 1356.590 367.585 1356.870 367.865 ;
        RECT 1357.210 367.585 1357.490 367.865 ;
        RECT 1357.830 367.585 1358.110 367.865 ;
        RECT 1358.450 367.585 1358.730 367.865 ;
        RECT 1359.070 367.585 1359.350 367.865 ;
        RECT 1359.690 367.585 1359.970 367.865 ;
        RECT 1360.310 367.585 1360.590 367.865 ;
        RECT 1351.630 366.965 1351.910 367.245 ;
        RECT 1352.250 366.965 1352.530 367.245 ;
        RECT 1352.870 366.965 1353.150 367.245 ;
        RECT 1353.490 366.965 1353.770 367.245 ;
        RECT 1354.110 366.965 1354.390 367.245 ;
        RECT 1354.730 366.965 1355.010 367.245 ;
        RECT 1355.350 366.965 1355.630 367.245 ;
        RECT 1355.970 366.965 1356.250 367.245 ;
        RECT 1356.590 366.965 1356.870 367.245 ;
        RECT 1357.210 366.965 1357.490 367.245 ;
        RECT 1357.830 366.965 1358.110 367.245 ;
        RECT 1358.450 366.965 1358.730 367.245 ;
        RECT 1359.070 366.965 1359.350 367.245 ;
        RECT 1359.690 366.965 1359.970 367.245 ;
        RECT 1360.310 366.965 1360.590 367.245 ;
        RECT 1351.630 366.345 1351.910 366.625 ;
        RECT 1352.250 366.345 1352.530 366.625 ;
        RECT 1352.870 366.345 1353.150 366.625 ;
        RECT 1353.490 366.345 1353.770 366.625 ;
        RECT 1354.110 366.345 1354.390 366.625 ;
        RECT 1354.730 366.345 1355.010 366.625 ;
        RECT 1355.350 366.345 1355.630 366.625 ;
        RECT 1355.970 366.345 1356.250 366.625 ;
        RECT 1356.590 366.345 1356.870 366.625 ;
        RECT 1357.210 366.345 1357.490 366.625 ;
        RECT 1357.830 366.345 1358.110 366.625 ;
        RECT 1358.450 366.345 1358.730 366.625 ;
        RECT 1359.070 366.345 1359.350 366.625 ;
        RECT 1359.690 366.345 1359.970 366.625 ;
        RECT 1360.310 366.345 1360.590 366.625 ;
        RECT 1351.630 365.725 1351.910 366.005 ;
        RECT 1352.250 365.725 1352.530 366.005 ;
        RECT 1352.870 365.725 1353.150 366.005 ;
        RECT 1353.490 365.725 1353.770 366.005 ;
        RECT 1354.110 365.725 1354.390 366.005 ;
        RECT 1354.730 365.725 1355.010 366.005 ;
        RECT 1355.350 365.725 1355.630 366.005 ;
        RECT 1355.970 365.725 1356.250 366.005 ;
        RECT 1356.590 365.725 1356.870 366.005 ;
        RECT 1357.210 365.725 1357.490 366.005 ;
        RECT 1357.830 365.725 1358.110 366.005 ;
        RECT 1358.450 365.725 1358.730 366.005 ;
        RECT 1359.070 365.725 1359.350 366.005 ;
        RECT 1359.690 365.725 1359.970 366.005 ;
        RECT 1360.310 365.725 1360.590 366.005 ;
        RECT 1351.630 365.105 1351.910 365.385 ;
        RECT 1352.250 365.105 1352.530 365.385 ;
        RECT 1352.870 365.105 1353.150 365.385 ;
        RECT 1353.490 365.105 1353.770 365.385 ;
        RECT 1354.110 365.105 1354.390 365.385 ;
        RECT 1354.730 365.105 1355.010 365.385 ;
        RECT 1355.350 365.105 1355.630 365.385 ;
        RECT 1355.970 365.105 1356.250 365.385 ;
        RECT 1356.590 365.105 1356.870 365.385 ;
        RECT 1357.210 365.105 1357.490 365.385 ;
        RECT 1357.830 365.105 1358.110 365.385 ;
        RECT 1358.450 365.105 1358.730 365.385 ;
        RECT 1359.070 365.105 1359.350 365.385 ;
        RECT 1359.690 365.105 1359.970 365.385 ;
        RECT 1360.310 365.105 1360.590 365.385 ;
        RECT 1351.630 364.485 1351.910 364.765 ;
        RECT 1352.250 364.485 1352.530 364.765 ;
        RECT 1352.870 364.485 1353.150 364.765 ;
        RECT 1353.490 364.485 1353.770 364.765 ;
        RECT 1354.110 364.485 1354.390 364.765 ;
        RECT 1354.730 364.485 1355.010 364.765 ;
        RECT 1355.350 364.485 1355.630 364.765 ;
        RECT 1355.970 364.485 1356.250 364.765 ;
        RECT 1356.590 364.485 1356.870 364.765 ;
        RECT 1357.210 364.485 1357.490 364.765 ;
        RECT 1357.830 364.485 1358.110 364.765 ;
        RECT 1358.450 364.485 1358.730 364.765 ;
        RECT 1359.070 364.485 1359.350 364.765 ;
        RECT 1359.690 364.485 1359.970 364.765 ;
        RECT 1360.310 364.485 1360.590 364.765 ;
        RECT 1351.630 363.865 1351.910 364.145 ;
        RECT 1352.250 363.865 1352.530 364.145 ;
        RECT 1352.870 363.865 1353.150 364.145 ;
        RECT 1353.490 363.865 1353.770 364.145 ;
        RECT 1354.110 363.865 1354.390 364.145 ;
        RECT 1354.730 363.865 1355.010 364.145 ;
        RECT 1355.350 363.865 1355.630 364.145 ;
        RECT 1355.970 363.865 1356.250 364.145 ;
        RECT 1356.590 363.865 1356.870 364.145 ;
        RECT 1357.210 363.865 1357.490 364.145 ;
        RECT 1357.830 363.865 1358.110 364.145 ;
        RECT 1358.450 363.865 1358.730 364.145 ;
        RECT 1359.070 363.865 1359.350 364.145 ;
        RECT 1359.690 363.865 1359.970 364.145 ;
        RECT 1360.310 363.865 1360.590 364.145 ;
        RECT 1351.630 363.245 1351.910 363.525 ;
        RECT 1352.250 363.245 1352.530 363.525 ;
        RECT 1352.870 363.245 1353.150 363.525 ;
        RECT 1353.490 363.245 1353.770 363.525 ;
        RECT 1354.110 363.245 1354.390 363.525 ;
        RECT 1354.730 363.245 1355.010 363.525 ;
        RECT 1355.350 363.245 1355.630 363.525 ;
        RECT 1355.970 363.245 1356.250 363.525 ;
        RECT 1356.590 363.245 1356.870 363.525 ;
        RECT 1357.210 363.245 1357.490 363.525 ;
        RECT 1357.830 363.245 1358.110 363.525 ;
        RECT 1358.450 363.245 1358.730 363.525 ;
        RECT 1359.070 363.245 1359.350 363.525 ;
        RECT 1359.690 363.245 1359.970 363.525 ;
        RECT 1360.310 363.245 1360.590 363.525 ;
        RECT 1351.630 362.625 1351.910 362.905 ;
        RECT 1352.250 362.625 1352.530 362.905 ;
        RECT 1352.870 362.625 1353.150 362.905 ;
        RECT 1353.490 362.625 1353.770 362.905 ;
        RECT 1354.110 362.625 1354.390 362.905 ;
        RECT 1354.730 362.625 1355.010 362.905 ;
        RECT 1355.350 362.625 1355.630 362.905 ;
        RECT 1355.970 362.625 1356.250 362.905 ;
        RECT 1356.590 362.625 1356.870 362.905 ;
        RECT 1357.210 362.625 1357.490 362.905 ;
        RECT 1357.830 362.625 1358.110 362.905 ;
        RECT 1358.450 362.625 1358.730 362.905 ;
        RECT 1359.070 362.625 1359.350 362.905 ;
        RECT 1359.690 362.625 1359.970 362.905 ;
        RECT 1360.310 362.625 1360.590 362.905 ;
        RECT 1351.630 362.005 1351.910 362.285 ;
        RECT 1352.250 362.005 1352.530 362.285 ;
        RECT 1352.870 362.005 1353.150 362.285 ;
        RECT 1353.490 362.005 1353.770 362.285 ;
        RECT 1354.110 362.005 1354.390 362.285 ;
        RECT 1354.730 362.005 1355.010 362.285 ;
        RECT 1355.350 362.005 1355.630 362.285 ;
        RECT 1355.970 362.005 1356.250 362.285 ;
        RECT 1356.590 362.005 1356.870 362.285 ;
        RECT 1357.210 362.005 1357.490 362.285 ;
        RECT 1357.830 362.005 1358.110 362.285 ;
        RECT 1358.450 362.005 1358.730 362.285 ;
        RECT 1359.070 362.005 1359.350 362.285 ;
        RECT 1359.690 362.005 1359.970 362.285 ;
        RECT 1360.310 362.005 1360.590 362.285 ;
        RECT 1351.630 361.385 1351.910 361.665 ;
        RECT 1352.250 361.385 1352.530 361.665 ;
        RECT 1352.870 361.385 1353.150 361.665 ;
        RECT 1353.490 361.385 1353.770 361.665 ;
        RECT 1354.110 361.385 1354.390 361.665 ;
        RECT 1354.730 361.385 1355.010 361.665 ;
        RECT 1355.350 361.385 1355.630 361.665 ;
        RECT 1355.970 361.385 1356.250 361.665 ;
        RECT 1356.590 361.385 1356.870 361.665 ;
        RECT 1357.210 361.385 1357.490 361.665 ;
        RECT 1357.830 361.385 1358.110 361.665 ;
        RECT 1358.450 361.385 1358.730 361.665 ;
        RECT 1359.070 361.385 1359.350 361.665 ;
        RECT 1359.690 361.385 1359.970 361.665 ;
        RECT 1360.310 361.385 1360.590 361.665 ;
        RECT 1351.630 360.765 1351.910 361.045 ;
        RECT 1352.250 360.765 1352.530 361.045 ;
        RECT 1352.870 360.765 1353.150 361.045 ;
        RECT 1353.490 360.765 1353.770 361.045 ;
        RECT 1354.110 360.765 1354.390 361.045 ;
        RECT 1354.730 360.765 1355.010 361.045 ;
        RECT 1355.350 360.765 1355.630 361.045 ;
        RECT 1355.970 360.765 1356.250 361.045 ;
        RECT 1356.590 360.765 1356.870 361.045 ;
        RECT 1357.210 360.765 1357.490 361.045 ;
        RECT 1357.830 360.765 1358.110 361.045 ;
        RECT 1358.450 360.765 1358.730 361.045 ;
        RECT 1359.070 360.765 1359.350 361.045 ;
        RECT 1359.690 360.765 1359.970 361.045 ;
        RECT 1360.310 360.765 1360.590 361.045 ;
        RECT 1364.030 369.445 1364.310 369.725 ;
        RECT 1364.650 369.445 1364.930 369.725 ;
        RECT 1365.270 369.445 1365.550 369.725 ;
        RECT 1365.890 369.445 1366.170 369.725 ;
        RECT 1366.510 369.445 1366.790 369.725 ;
        RECT 1367.130 369.445 1367.410 369.725 ;
        RECT 1367.750 369.445 1368.030 369.725 ;
        RECT 1368.370 369.445 1368.650 369.725 ;
        RECT 1368.990 369.445 1369.270 369.725 ;
        RECT 1369.610 369.445 1369.890 369.725 ;
        RECT 1370.230 369.445 1370.510 369.725 ;
        RECT 1370.850 369.445 1371.130 369.725 ;
        RECT 1371.470 369.445 1371.750 369.725 ;
        RECT 1372.090 369.445 1372.370 369.725 ;
        RECT 1372.710 369.445 1372.990 369.725 ;
        RECT 1373.330 369.445 1373.610 369.725 ;
        RECT 1364.030 368.825 1364.310 369.105 ;
        RECT 1364.650 368.825 1364.930 369.105 ;
        RECT 1365.270 368.825 1365.550 369.105 ;
        RECT 1365.890 368.825 1366.170 369.105 ;
        RECT 1366.510 368.825 1366.790 369.105 ;
        RECT 1367.130 368.825 1367.410 369.105 ;
        RECT 1367.750 368.825 1368.030 369.105 ;
        RECT 1368.370 368.825 1368.650 369.105 ;
        RECT 1368.990 368.825 1369.270 369.105 ;
        RECT 1369.610 368.825 1369.890 369.105 ;
        RECT 1370.230 368.825 1370.510 369.105 ;
        RECT 1370.850 368.825 1371.130 369.105 ;
        RECT 1371.470 368.825 1371.750 369.105 ;
        RECT 1372.090 368.825 1372.370 369.105 ;
        RECT 1372.710 368.825 1372.990 369.105 ;
        RECT 1373.330 368.825 1373.610 369.105 ;
        RECT 1364.030 368.205 1364.310 368.485 ;
        RECT 1364.650 368.205 1364.930 368.485 ;
        RECT 1365.270 368.205 1365.550 368.485 ;
        RECT 1365.890 368.205 1366.170 368.485 ;
        RECT 1366.510 368.205 1366.790 368.485 ;
        RECT 1367.130 368.205 1367.410 368.485 ;
        RECT 1367.750 368.205 1368.030 368.485 ;
        RECT 1368.370 368.205 1368.650 368.485 ;
        RECT 1368.990 368.205 1369.270 368.485 ;
        RECT 1369.610 368.205 1369.890 368.485 ;
        RECT 1370.230 368.205 1370.510 368.485 ;
        RECT 1370.850 368.205 1371.130 368.485 ;
        RECT 1371.470 368.205 1371.750 368.485 ;
        RECT 1372.090 368.205 1372.370 368.485 ;
        RECT 1372.710 368.205 1372.990 368.485 ;
        RECT 1373.330 368.205 1373.610 368.485 ;
        RECT 1364.030 367.585 1364.310 367.865 ;
        RECT 1364.650 367.585 1364.930 367.865 ;
        RECT 1365.270 367.585 1365.550 367.865 ;
        RECT 1365.890 367.585 1366.170 367.865 ;
        RECT 1366.510 367.585 1366.790 367.865 ;
        RECT 1367.130 367.585 1367.410 367.865 ;
        RECT 1367.750 367.585 1368.030 367.865 ;
        RECT 1368.370 367.585 1368.650 367.865 ;
        RECT 1368.990 367.585 1369.270 367.865 ;
        RECT 1369.610 367.585 1369.890 367.865 ;
        RECT 1370.230 367.585 1370.510 367.865 ;
        RECT 1370.850 367.585 1371.130 367.865 ;
        RECT 1371.470 367.585 1371.750 367.865 ;
        RECT 1372.090 367.585 1372.370 367.865 ;
        RECT 1372.710 367.585 1372.990 367.865 ;
        RECT 1373.330 367.585 1373.610 367.865 ;
        RECT 1364.030 366.965 1364.310 367.245 ;
        RECT 1364.650 366.965 1364.930 367.245 ;
        RECT 1365.270 366.965 1365.550 367.245 ;
        RECT 1365.890 366.965 1366.170 367.245 ;
        RECT 1366.510 366.965 1366.790 367.245 ;
        RECT 1367.130 366.965 1367.410 367.245 ;
        RECT 1367.750 366.965 1368.030 367.245 ;
        RECT 1368.370 366.965 1368.650 367.245 ;
        RECT 1368.990 366.965 1369.270 367.245 ;
        RECT 1369.610 366.965 1369.890 367.245 ;
        RECT 1370.230 366.965 1370.510 367.245 ;
        RECT 1370.850 366.965 1371.130 367.245 ;
        RECT 1371.470 366.965 1371.750 367.245 ;
        RECT 1372.090 366.965 1372.370 367.245 ;
        RECT 1372.710 366.965 1372.990 367.245 ;
        RECT 1373.330 366.965 1373.610 367.245 ;
        RECT 1364.030 366.345 1364.310 366.625 ;
        RECT 1364.650 366.345 1364.930 366.625 ;
        RECT 1365.270 366.345 1365.550 366.625 ;
        RECT 1365.890 366.345 1366.170 366.625 ;
        RECT 1366.510 366.345 1366.790 366.625 ;
        RECT 1367.130 366.345 1367.410 366.625 ;
        RECT 1367.750 366.345 1368.030 366.625 ;
        RECT 1368.370 366.345 1368.650 366.625 ;
        RECT 1368.990 366.345 1369.270 366.625 ;
        RECT 1369.610 366.345 1369.890 366.625 ;
        RECT 1370.230 366.345 1370.510 366.625 ;
        RECT 1370.850 366.345 1371.130 366.625 ;
        RECT 1371.470 366.345 1371.750 366.625 ;
        RECT 1372.090 366.345 1372.370 366.625 ;
        RECT 1372.710 366.345 1372.990 366.625 ;
        RECT 1373.330 366.345 1373.610 366.625 ;
        RECT 1364.030 365.725 1364.310 366.005 ;
        RECT 1364.650 365.725 1364.930 366.005 ;
        RECT 1365.270 365.725 1365.550 366.005 ;
        RECT 1365.890 365.725 1366.170 366.005 ;
        RECT 1366.510 365.725 1366.790 366.005 ;
        RECT 1367.130 365.725 1367.410 366.005 ;
        RECT 1367.750 365.725 1368.030 366.005 ;
        RECT 1368.370 365.725 1368.650 366.005 ;
        RECT 1368.990 365.725 1369.270 366.005 ;
        RECT 1369.610 365.725 1369.890 366.005 ;
        RECT 1370.230 365.725 1370.510 366.005 ;
        RECT 1370.850 365.725 1371.130 366.005 ;
        RECT 1371.470 365.725 1371.750 366.005 ;
        RECT 1372.090 365.725 1372.370 366.005 ;
        RECT 1372.710 365.725 1372.990 366.005 ;
        RECT 1373.330 365.725 1373.610 366.005 ;
        RECT 1364.030 365.105 1364.310 365.385 ;
        RECT 1364.650 365.105 1364.930 365.385 ;
        RECT 1365.270 365.105 1365.550 365.385 ;
        RECT 1365.890 365.105 1366.170 365.385 ;
        RECT 1366.510 365.105 1366.790 365.385 ;
        RECT 1367.130 365.105 1367.410 365.385 ;
        RECT 1367.750 365.105 1368.030 365.385 ;
        RECT 1368.370 365.105 1368.650 365.385 ;
        RECT 1368.990 365.105 1369.270 365.385 ;
        RECT 1369.610 365.105 1369.890 365.385 ;
        RECT 1370.230 365.105 1370.510 365.385 ;
        RECT 1370.850 365.105 1371.130 365.385 ;
        RECT 1371.470 365.105 1371.750 365.385 ;
        RECT 1372.090 365.105 1372.370 365.385 ;
        RECT 1372.710 365.105 1372.990 365.385 ;
        RECT 1373.330 365.105 1373.610 365.385 ;
        RECT 1364.030 364.485 1364.310 364.765 ;
        RECT 1364.650 364.485 1364.930 364.765 ;
        RECT 1365.270 364.485 1365.550 364.765 ;
        RECT 1365.890 364.485 1366.170 364.765 ;
        RECT 1366.510 364.485 1366.790 364.765 ;
        RECT 1367.130 364.485 1367.410 364.765 ;
        RECT 1367.750 364.485 1368.030 364.765 ;
        RECT 1368.370 364.485 1368.650 364.765 ;
        RECT 1368.990 364.485 1369.270 364.765 ;
        RECT 1369.610 364.485 1369.890 364.765 ;
        RECT 1370.230 364.485 1370.510 364.765 ;
        RECT 1370.850 364.485 1371.130 364.765 ;
        RECT 1371.470 364.485 1371.750 364.765 ;
        RECT 1372.090 364.485 1372.370 364.765 ;
        RECT 1372.710 364.485 1372.990 364.765 ;
        RECT 1373.330 364.485 1373.610 364.765 ;
        RECT 1364.030 363.865 1364.310 364.145 ;
        RECT 1364.650 363.865 1364.930 364.145 ;
        RECT 1365.270 363.865 1365.550 364.145 ;
        RECT 1365.890 363.865 1366.170 364.145 ;
        RECT 1366.510 363.865 1366.790 364.145 ;
        RECT 1367.130 363.865 1367.410 364.145 ;
        RECT 1367.750 363.865 1368.030 364.145 ;
        RECT 1368.370 363.865 1368.650 364.145 ;
        RECT 1368.990 363.865 1369.270 364.145 ;
        RECT 1369.610 363.865 1369.890 364.145 ;
        RECT 1370.230 363.865 1370.510 364.145 ;
        RECT 1370.850 363.865 1371.130 364.145 ;
        RECT 1371.470 363.865 1371.750 364.145 ;
        RECT 1372.090 363.865 1372.370 364.145 ;
        RECT 1372.710 363.865 1372.990 364.145 ;
        RECT 1373.330 363.865 1373.610 364.145 ;
        RECT 1364.030 363.245 1364.310 363.525 ;
        RECT 1364.650 363.245 1364.930 363.525 ;
        RECT 1365.270 363.245 1365.550 363.525 ;
        RECT 1365.890 363.245 1366.170 363.525 ;
        RECT 1366.510 363.245 1366.790 363.525 ;
        RECT 1367.130 363.245 1367.410 363.525 ;
        RECT 1367.750 363.245 1368.030 363.525 ;
        RECT 1368.370 363.245 1368.650 363.525 ;
        RECT 1368.990 363.245 1369.270 363.525 ;
        RECT 1369.610 363.245 1369.890 363.525 ;
        RECT 1370.230 363.245 1370.510 363.525 ;
        RECT 1370.850 363.245 1371.130 363.525 ;
        RECT 1371.470 363.245 1371.750 363.525 ;
        RECT 1372.090 363.245 1372.370 363.525 ;
        RECT 1372.710 363.245 1372.990 363.525 ;
        RECT 1373.330 363.245 1373.610 363.525 ;
        RECT 1364.030 362.625 1364.310 362.905 ;
        RECT 1364.650 362.625 1364.930 362.905 ;
        RECT 1365.270 362.625 1365.550 362.905 ;
        RECT 1365.890 362.625 1366.170 362.905 ;
        RECT 1366.510 362.625 1366.790 362.905 ;
        RECT 1367.130 362.625 1367.410 362.905 ;
        RECT 1367.750 362.625 1368.030 362.905 ;
        RECT 1368.370 362.625 1368.650 362.905 ;
        RECT 1368.990 362.625 1369.270 362.905 ;
        RECT 1369.610 362.625 1369.890 362.905 ;
        RECT 1370.230 362.625 1370.510 362.905 ;
        RECT 1370.850 362.625 1371.130 362.905 ;
        RECT 1371.470 362.625 1371.750 362.905 ;
        RECT 1372.090 362.625 1372.370 362.905 ;
        RECT 1372.710 362.625 1372.990 362.905 ;
        RECT 1373.330 362.625 1373.610 362.905 ;
        RECT 1364.030 362.005 1364.310 362.285 ;
        RECT 1364.650 362.005 1364.930 362.285 ;
        RECT 1365.270 362.005 1365.550 362.285 ;
        RECT 1365.890 362.005 1366.170 362.285 ;
        RECT 1366.510 362.005 1366.790 362.285 ;
        RECT 1367.130 362.005 1367.410 362.285 ;
        RECT 1367.750 362.005 1368.030 362.285 ;
        RECT 1368.370 362.005 1368.650 362.285 ;
        RECT 1368.990 362.005 1369.270 362.285 ;
        RECT 1369.610 362.005 1369.890 362.285 ;
        RECT 1370.230 362.005 1370.510 362.285 ;
        RECT 1370.850 362.005 1371.130 362.285 ;
        RECT 1371.470 362.005 1371.750 362.285 ;
        RECT 1372.090 362.005 1372.370 362.285 ;
        RECT 1372.710 362.005 1372.990 362.285 ;
        RECT 1373.330 362.005 1373.610 362.285 ;
        RECT 1364.030 361.385 1364.310 361.665 ;
        RECT 1364.650 361.385 1364.930 361.665 ;
        RECT 1365.270 361.385 1365.550 361.665 ;
        RECT 1365.890 361.385 1366.170 361.665 ;
        RECT 1366.510 361.385 1366.790 361.665 ;
        RECT 1367.130 361.385 1367.410 361.665 ;
        RECT 1367.750 361.385 1368.030 361.665 ;
        RECT 1368.370 361.385 1368.650 361.665 ;
        RECT 1368.990 361.385 1369.270 361.665 ;
        RECT 1369.610 361.385 1369.890 361.665 ;
        RECT 1370.230 361.385 1370.510 361.665 ;
        RECT 1370.850 361.385 1371.130 361.665 ;
        RECT 1371.470 361.385 1371.750 361.665 ;
        RECT 1372.090 361.385 1372.370 361.665 ;
        RECT 1372.710 361.385 1372.990 361.665 ;
        RECT 1373.330 361.385 1373.610 361.665 ;
        RECT 1364.030 360.765 1364.310 361.045 ;
        RECT 1364.650 360.765 1364.930 361.045 ;
        RECT 1365.270 360.765 1365.550 361.045 ;
        RECT 1365.890 360.765 1366.170 361.045 ;
        RECT 1366.510 360.765 1366.790 361.045 ;
        RECT 1367.130 360.765 1367.410 361.045 ;
        RECT 1367.750 360.765 1368.030 361.045 ;
        RECT 1368.370 360.765 1368.650 361.045 ;
        RECT 1368.990 360.765 1369.270 361.045 ;
        RECT 1369.610 360.765 1369.890 361.045 ;
        RECT 1370.230 360.765 1370.510 361.045 ;
        RECT 1370.850 360.765 1371.130 361.045 ;
        RECT 1371.470 360.765 1371.750 361.045 ;
        RECT 1372.090 360.765 1372.370 361.045 ;
        RECT 1372.710 360.765 1372.990 361.045 ;
        RECT 1373.330 360.765 1373.610 361.045 ;
        RECT 1375.880 369.445 1376.160 369.725 ;
        RECT 1376.500 369.445 1376.780 369.725 ;
        RECT 1377.120 369.445 1377.400 369.725 ;
        RECT 1377.740 369.445 1378.020 369.725 ;
        RECT 1378.360 369.445 1378.640 369.725 ;
        RECT 1378.980 369.445 1379.260 369.725 ;
        RECT 1379.600 369.445 1379.880 369.725 ;
        RECT 1380.220 369.445 1380.500 369.725 ;
        RECT 1380.840 369.445 1381.120 369.725 ;
        RECT 1381.460 369.445 1381.740 369.725 ;
        RECT 1382.080 369.445 1382.360 369.725 ;
        RECT 1382.700 369.445 1382.980 369.725 ;
        RECT 1383.320 369.445 1383.600 369.725 ;
        RECT 1383.940 369.445 1384.220 369.725 ;
        RECT 1384.560 369.445 1384.840 369.725 ;
        RECT 1385.180 369.445 1385.460 369.725 ;
        RECT 1375.880 368.825 1376.160 369.105 ;
        RECT 1376.500 368.825 1376.780 369.105 ;
        RECT 1377.120 368.825 1377.400 369.105 ;
        RECT 1377.740 368.825 1378.020 369.105 ;
        RECT 1378.360 368.825 1378.640 369.105 ;
        RECT 1378.980 368.825 1379.260 369.105 ;
        RECT 1379.600 368.825 1379.880 369.105 ;
        RECT 1380.220 368.825 1380.500 369.105 ;
        RECT 1380.840 368.825 1381.120 369.105 ;
        RECT 1381.460 368.825 1381.740 369.105 ;
        RECT 1382.080 368.825 1382.360 369.105 ;
        RECT 1382.700 368.825 1382.980 369.105 ;
        RECT 1383.320 368.825 1383.600 369.105 ;
        RECT 1383.940 368.825 1384.220 369.105 ;
        RECT 1384.560 368.825 1384.840 369.105 ;
        RECT 1385.180 368.825 1385.460 369.105 ;
        RECT 1375.880 368.205 1376.160 368.485 ;
        RECT 1376.500 368.205 1376.780 368.485 ;
        RECT 1377.120 368.205 1377.400 368.485 ;
        RECT 1377.740 368.205 1378.020 368.485 ;
        RECT 1378.360 368.205 1378.640 368.485 ;
        RECT 1378.980 368.205 1379.260 368.485 ;
        RECT 1379.600 368.205 1379.880 368.485 ;
        RECT 1380.220 368.205 1380.500 368.485 ;
        RECT 1380.840 368.205 1381.120 368.485 ;
        RECT 1381.460 368.205 1381.740 368.485 ;
        RECT 1382.080 368.205 1382.360 368.485 ;
        RECT 1382.700 368.205 1382.980 368.485 ;
        RECT 1383.320 368.205 1383.600 368.485 ;
        RECT 1383.940 368.205 1384.220 368.485 ;
        RECT 1384.560 368.205 1384.840 368.485 ;
        RECT 1385.180 368.205 1385.460 368.485 ;
        RECT 1375.880 367.585 1376.160 367.865 ;
        RECT 1376.500 367.585 1376.780 367.865 ;
        RECT 1377.120 367.585 1377.400 367.865 ;
        RECT 1377.740 367.585 1378.020 367.865 ;
        RECT 1378.360 367.585 1378.640 367.865 ;
        RECT 1378.980 367.585 1379.260 367.865 ;
        RECT 1379.600 367.585 1379.880 367.865 ;
        RECT 1380.220 367.585 1380.500 367.865 ;
        RECT 1380.840 367.585 1381.120 367.865 ;
        RECT 1381.460 367.585 1381.740 367.865 ;
        RECT 1382.080 367.585 1382.360 367.865 ;
        RECT 1382.700 367.585 1382.980 367.865 ;
        RECT 1383.320 367.585 1383.600 367.865 ;
        RECT 1383.940 367.585 1384.220 367.865 ;
        RECT 1384.560 367.585 1384.840 367.865 ;
        RECT 1385.180 367.585 1385.460 367.865 ;
        RECT 1375.880 366.965 1376.160 367.245 ;
        RECT 1376.500 366.965 1376.780 367.245 ;
        RECT 1377.120 366.965 1377.400 367.245 ;
        RECT 1377.740 366.965 1378.020 367.245 ;
        RECT 1378.360 366.965 1378.640 367.245 ;
        RECT 1378.980 366.965 1379.260 367.245 ;
        RECT 1379.600 366.965 1379.880 367.245 ;
        RECT 1380.220 366.965 1380.500 367.245 ;
        RECT 1380.840 366.965 1381.120 367.245 ;
        RECT 1381.460 366.965 1381.740 367.245 ;
        RECT 1382.080 366.965 1382.360 367.245 ;
        RECT 1382.700 366.965 1382.980 367.245 ;
        RECT 1383.320 366.965 1383.600 367.245 ;
        RECT 1383.940 366.965 1384.220 367.245 ;
        RECT 1384.560 366.965 1384.840 367.245 ;
        RECT 1385.180 366.965 1385.460 367.245 ;
        RECT 1375.880 366.345 1376.160 366.625 ;
        RECT 1376.500 366.345 1376.780 366.625 ;
        RECT 1377.120 366.345 1377.400 366.625 ;
        RECT 1377.740 366.345 1378.020 366.625 ;
        RECT 1378.360 366.345 1378.640 366.625 ;
        RECT 1378.980 366.345 1379.260 366.625 ;
        RECT 1379.600 366.345 1379.880 366.625 ;
        RECT 1380.220 366.345 1380.500 366.625 ;
        RECT 1380.840 366.345 1381.120 366.625 ;
        RECT 1381.460 366.345 1381.740 366.625 ;
        RECT 1382.080 366.345 1382.360 366.625 ;
        RECT 1382.700 366.345 1382.980 366.625 ;
        RECT 1383.320 366.345 1383.600 366.625 ;
        RECT 1383.940 366.345 1384.220 366.625 ;
        RECT 1384.560 366.345 1384.840 366.625 ;
        RECT 1385.180 366.345 1385.460 366.625 ;
        RECT 1375.880 365.725 1376.160 366.005 ;
        RECT 1376.500 365.725 1376.780 366.005 ;
        RECT 1377.120 365.725 1377.400 366.005 ;
        RECT 1377.740 365.725 1378.020 366.005 ;
        RECT 1378.360 365.725 1378.640 366.005 ;
        RECT 1378.980 365.725 1379.260 366.005 ;
        RECT 1379.600 365.725 1379.880 366.005 ;
        RECT 1380.220 365.725 1380.500 366.005 ;
        RECT 1380.840 365.725 1381.120 366.005 ;
        RECT 1381.460 365.725 1381.740 366.005 ;
        RECT 1382.080 365.725 1382.360 366.005 ;
        RECT 1382.700 365.725 1382.980 366.005 ;
        RECT 1383.320 365.725 1383.600 366.005 ;
        RECT 1383.940 365.725 1384.220 366.005 ;
        RECT 1384.560 365.725 1384.840 366.005 ;
        RECT 1385.180 365.725 1385.460 366.005 ;
        RECT 1375.880 365.105 1376.160 365.385 ;
        RECT 1376.500 365.105 1376.780 365.385 ;
        RECT 1377.120 365.105 1377.400 365.385 ;
        RECT 1377.740 365.105 1378.020 365.385 ;
        RECT 1378.360 365.105 1378.640 365.385 ;
        RECT 1378.980 365.105 1379.260 365.385 ;
        RECT 1379.600 365.105 1379.880 365.385 ;
        RECT 1380.220 365.105 1380.500 365.385 ;
        RECT 1380.840 365.105 1381.120 365.385 ;
        RECT 1381.460 365.105 1381.740 365.385 ;
        RECT 1382.080 365.105 1382.360 365.385 ;
        RECT 1382.700 365.105 1382.980 365.385 ;
        RECT 1383.320 365.105 1383.600 365.385 ;
        RECT 1383.940 365.105 1384.220 365.385 ;
        RECT 1384.560 365.105 1384.840 365.385 ;
        RECT 1385.180 365.105 1385.460 365.385 ;
        RECT 1375.880 364.485 1376.160 364.765 ;
        RECT 1376.500 364.485 1376.780 364.765 ;
        RECT 1377.120 364.485 1377.400 364.765 ;
        RECT 1377.740 364.485 1378.020 364.765 ;
        RECT 1378.360 364.485 1378.640 364.765 ;
        RECT 1378.980 364.485 1379.260 364.765 ;
        RECT 1379.600 364.485 1379.880 364.765 ;
        RECT 1380.220 364.485 1380.500 364.765 ;
        RECT 1380.840 364.485 1381.120 364.765 ;
        RECT 1381.460 364.485 1381.740 364.765 ;
        RECT 1382.080 364.485 1382.360 364.765 ;
        RECT 1382.700 364.485 1382.980 364.765 ;
        RECT 1383.320 364.485 1383.600 364.765 ;
        RECT 1383.940 364.485 1384.220 364.765 ;
        RECT 1384.560 364.485 1384.840 364.765 ;
        RECT 1385.180 364.485 1385.460 364.765 ;
        RECT 1375.880 363.865 1376.160 364.145 ;
        RECT 1376.500 363.865 1376.780 364.145 ;
        RECT 1377.120 363.865 1377.400 364.145 ;
        RECT 1377.740 363.865 1378.020 364.145 ;
        RECT 1378.360 363.865 1378.640 364.145 ;
        RECT 1378.980 363.865 1379.260 364.145 ;
        RECT 1379.600 363.865 1379.880 364.145 ;
        RECT 1380.220 363.865 1380.500 364.145 ;
        RECT 1380.840 363.865 1381.120 364.145 ;
        RECT 1381.460 363.865 1381.740 364.145 ;
        RECT 1382.080 363.865 1382.360 364.145 ;
        RECT 1382.700 363.865 1382.980 364.145 ;
        RECT 1383.320 363.865 1383.600 364.145 ;
        RECT 1383.940 363.865 1384.220 364.145 ;
        RECT 1384.560 363.865 1384.840 364.145 ;
        RECT 1385.180 363.865 1385.460 364.145 ;
        RECT 1375.880 363.245 1376.160 363.525 ;
        RECT 1376.500 363.245 1376.780 363.525 ;
        RECT 1377.120 363.245 1377.400 363.525 ;
        RECT 1377.740 363.245 1378.020 363.525 ;
        RECT 1378.360 363.245 1378.640 363.525 ;
        RECT 1378.980 363.245 1379.260 363.525 ;
        RECT 1379.600 363.245 1379.880 363.525 ;
        RECT 1380.220 363.245 1380.500 363.525 ;
        RECT 1380.840 363.245 1381.120 363.525 ;
        RECT 1381.460 363.245 1381.740 363.525 ;
        RECT 1382.080 363.245 1382.360 363.525 ;
        RECT 1382.700 363.245 1382.980 363.525 ;
        RECT 1383.320 363.245 1383.600 363.525 ;
        RECT 1383.940 363.245 1384.220 363.525 ;
        RECT 1384.560 363.245 1384.840 363.525 ;
        RECT 1385.180 363.245 1385.460 363.525 ;
        RECT 1375.880 362.625 1376.160 362.905 ;
        RECT 1376.500 362.625 1376.780 362.905 ;
        RECT 1377.120 362.625 1377.400 362.905 ;
        RECT 1377.740 362.625 1378.020 362.905 ;
        RECT 1378.360 362.625 1378.640 362.905 ;
        RECT 1378.980 362.625 1379.260 362.905 ;
        RECT 1379.600 362.625 1379.880 362.905 ;
        RECT 1380.220 362.625 1380.500 362.905 ;
        RECT 1380.840 362.625 1381.120 362.905 ;
        RECT 1381.460 362.625 1381.740 362.905 ;
        RECT 1382.080 362.625 1382.360 362.905 ;
        RECT 1382.700 362.625 1382.980 362.905 ;
        RECT 1383.320 362.625 1383.600 362.905 ;
        RECT 1383.940 362.625 1384.220 362.905 ;
        RECT 1384.560 362.625 1384.840 362.905 ;
        RECT 1385.180 362.625 1385.460 362.905 ;
        RECT 1375.880 362.005 1376.160 362.285 ;
        RECT 1376.500 362.005 1376.780 362.285 ;
        RECT 1377.120 362.005 1377.400 362.285 ;
        RECT 1377.740 362.005 1378.020 362.285 ;
        RECT 1378.360 362.005 1378.640 362.285 ;
        RECT 1378.980 362.005 1379.260 362.285 ;
        RECT 1379.600 362.005 1379.880 362.285 ;
        RECT 1380.220 362.005 1380.500 362.285 ;
        RECT 1380.840 362.005 1381.120 362.285 ;
        RECT 1381.460 362.005 1381.740 362.285 ;
        RECT 1382.080 362.005 1382.360 362.285 ;
        RECT 1382.700 362.005 1382.980 362.285 ;
        RECT 1383.320 362.005 1383.600 362.285 ;
        RECT 1383.940 362.005 1384.220 362.285 ;
        RECT 1384.560 362.005 1384.840 362.285 ;
        RECT 1385.180 362.005 1385.460 362.285 ;
        RECT 1375.880 361.385 1376.160 361.665 ;
        RECT 1376.500 361.385 1376.780 361.665 ;
        RECT 1377.120 361.385 1377.400 361.665 ;
        RECT 1377.740 361.385 1378.020 361.665 ;
        RECT 1378.360 361.385 1378.640 361.665 ;
        RECT 1378.980 361.385 1379.260 361.665 ;
        RECT 1379.600 361.385 1379.880 361.665 ;
        RECT 1380.220 361.385 1380.500 361.665 ;
        RECT 1380.840 361.385 1381.120 361.665 ;
        RECT 1381.460 361.385 1381.740 361.665 ;
        RECT 1382.080 361.385 1382.360 361.665 ;
        RECT 1382.700 361.385 1382.980 361.665 ;
        RECT 1383.320 361.385 1383.600 361.665 ;
        RECT 1383.940 361.385 1384.220 361.665 ;
        RECT 1384.560 361.385 1384.840 361.665 ;
        RECT 1385.180 361.385 1385.460 361.665 ;
        RECT 1375.880 360.765 1376.160 361.045 ;
        RECT 1376.500 360.765 1376.780 361.045 ;
        RECT 1377.120 360.765 1377.400 361.045 ;
        RECT 1377.740 360.765 1378.020 361.045 ;
        RECT 1378.360 360.765 1378.640 361.045 ;
        RECT 1378.980 360.765 1379.260 361.045 ;
        RECT 1379.600 360.765 1379.880 361.045 ;
        RECT 1380.220 360.765 1380.500 361.045 ;
        RECT 1380.840 360.765 1381.120 361.045 ;
        RECT 1381.460 360.765 1381.740 361.045 ;
        RECT 1382.080 360.765 1382.360 361.045 ;
        RECT 1382.700 360.765 1382.980 361.045 ;
        RECT 1383.320 360.765 1383.600 361.045 ;
        RECT 1383.940 360.765 1384.220 361.045 ;
        RECT 1384.560 360.765 1384.840 361.045 ;
        RECT 1385.180 360.765 1385.460 361.045 ;
        RECT 1389.410 369.445 1389.690 369.725 ;
        RECT 1390.030 369.445 1390.310 369.725 ;
        RECT 1390.650 369.445 1390.930 369.725 ;
        RECT 1391.270 369.445 1391.550 369.725 ;
        RECT 1391.890 369.445 1392.170 369.725 ;
        RECT 1392.510 369.445 1392.790 369.725 ;
        RECT 1393.130 369.445 1393.410 369.725 ;
        RECT 1393.750 369.445 1394.030 369.725 ;
        RECT 1394.370 369.445 1394.650 369.725 ;
        RECT 1394.990 369.445 1395.270 369.725 ;
        RECT 1395.610 369.445 1395.890 369.725 ;
        RECT 1396.230 369.445 1396.510 369.725 ;
        RECT 1396.850 369.445 1397.130 369.725 ;
        RECT 1397.470 369.445 1397.750 369.725 ;
        RECT 1398.090 369.445 1398.370 369.725 ;
        RECT 1398.710 369.445 1398.990 369.725 ;
        RECT 1389.410 368.825 1389.690 369.105 ;
        RECT 1390.030 368.825 1390.310 369.105 ;
        RECT 1390.650 368.825 1390.930 369.105 ;
        RECT 1391.270 368.825 1391.550 369.105 ;
        RECT 1391.890 368.825 1392.170 369.105 ;
        RECT 1392.510 368.825 1392.790 369.105 ;
        RECT 1393.130 368.825 1393.410 369.105 ;
        RECT 1393.750 368.825 1394.030 369.105 ;
        RECT 1394.370 368.825 1394.650 369.105 ;
        RECT 1394.990 368.825 1395.270 369.105 ;
        RECT 1395.610 368.825 1395.890 369.105 ;
        RECT 1396.230 368.825 1396.510 369.105 ;
        RECT 1396.850 368.825 1397.130 369.105 ;
        RECT 1397.470 368.825 1397.750 369.105 ;
        RECT 1398.090 368.825 1398.370 369.105 ;
        RECT 1398.710 368.825 1398.990 369.105 ;
        RECT 1389.410 368.205 1389.690 368.485 ;
        RECT 1390.030 368.205 1390.310 368.485 ;
        RECT 1390.650 368.205 1390.930 368.485 ;
        RECT 1391.270 368.205 1391.550 368.485 ;
        RECT 1391.890 368.205 1392.170 368.485 ;
        RECT 1392.510 368.205 1392.790 368.485 ;
        RECT 1393.130 368.205 1393.410 368.485 ;
        RECT 1393.750 368.205 1394.030 368.485 ;
        RECT 1394.370 368.205 1394.650 368.485 ;
        RECT 1394.990 368.205 1395.270 368.485 ;
        RECT 1395.610 368.205 1395.890 368.485 ;
        RECT 1396.230 368.205 1396.510 368.485 ;
        RECT 1396.850 368.205 1397.130 368.485 ;
        RECT 1397.470 368.205 1397.750 368.485 ;
        RECT 1398.090 368.205 1398.370 368.485 ;
        RECT 1398.710 368.205 1398.990 368.485 ;
        RECT 1389.410 367.585 1389.690 367.865 ;
        RECT 1390.030 367.585 1390.310 367.865 ;
        RECT 1390.650 367.585 1390.930 367.865 ;
        RECT 1391.270 367.585 1391.550 367.865 ;
        RECT 1391.890 367.585 1392.170 367.865 ;
        RECT 1392.510 367.585 1392.790 367.865 ;
        RECT 1393.130 367.585 1393.410 367.865 ;
        RECT 1393.750 367.585 1394.030 367.865 ;
        RECT 1394.370 367.585 1394.650 367.865 ;
        RECT 1394.990 367.585 1395.270 367.865 ;
        RECT 1395.610 367.585 1395.890 367.865 ;
        RECT 1396.230 367.585 1396.510 367.865 ;
        RECT 1396.850 367.585 1397.130 367.865 ;
        RECT 1397.470 367.585 1397.750 367.865 ;
        RECT 1398.090 367.585 1398.370 367.865 ;
        RECT 1398.710 367.585 1398.990 367.865 ;
        RECT 1389.410 366.965 1389.690 367.245 ;
        RECT 1390.030 366.965 1390.310 367.245 ;
        RECT 1390.650 366.965 1390.930 367.245 ;
        RECT 1391.270 366.965 1391.550 367.245 ;
        RECT 1391.890 366.965 1392.170 367.245 ;
        RECT 1392.510 366.965 1392.790 367.245 ;
        RECT 1393.130 366.965 1393.410 367.245 ;
        RECT 1393.750 366.965 1394.030 367.245 ;
        RECT 1394.370 366.965 1394.650 367.245 ;
        RECT 1394.990 366.965 1395.270 367.245 ;
        RECT 1395.610 366.965 1395.890 367.245 ;
        RECT 1396.230 366.965 1396.510 367.245 ;
        RECT 1396.850 366.965 1397.130 367.245 ;
        RECT 1397.470 366.965 1397.750 367.245 ;
        RECT 1398.090 366.965 1398.370 367.245 ;
        RECT 1398.710 366.965 1398.990 367.245 ;
        RECT 1389.410 366.345 1389.690 366.625 ;
        RECT 1390.030 366.345 1390.310 366.625 ;
        RECT 1390.650 366.345 1390.930 366.625 ;
        RECT 1391.270 366.345 1391.550 366.625 ;
        RECT 1391.890 366.345 1392.170 366.625 ;
        RECT 1392.510 366.345 1392.790 366.625 ;
        RECT 1393.130 366.345 1393.410 366.625 ;
        RECT 1393.750 366.345 1394.030 366.625 ;
        RECT 1394.370 366.345 1394.650 366.625 ;
        RECT 1394.990 366.345 1395.270 366.625 ;
        RECT 1395.610 366.345 1395.890 366.625 ;
        RECT 1396.230 366.345 1396.510 366.625 ;
        RECT 1396.850 366.345 1397.130 366.625 ;
        RECT 1397.470 366.345 1397.750 366.625 ;
        RECT 1398.090 366.345 1398.370 366.625 ;
        RECT 1398.710 366.345 1398.990 366.625 ;
        RECT 1389.410 365.725 1389.690 366.005 ;
        RECT 1390.030 365.725 1390.310 366.005 ;
        RECT 1390.650 365.725 1390.930 366.005 ;
        RECT 1391.270 365.725 1391.550 366.005 ;
        RECT 1391.890 365.725 1392.170 366.005 ;
        RECT 1392.510 365.725 1392.790 366.005 ;
        RECT 1393.130 365.725 1393.410 366.005 ;
        RECT 1393.750 365.725 1394.030 366.005 ;
        RECT 1394.370 365.725 1394.650 366.005 ;
        RECT 1394.990 365.725 1395.270 366.005 ;
        RECT 1395.610 365.725 1395.890 366.005 ;
        RECT 1396.230 365.725 1396.510 366.005 ;
        RECT 1396.850 365.725 1397.130 366.005 ;
        RECT 1397.470 365.725 1397.750 366.005 ;
        RECT 1398.090 365.725 1398.370 366.005 ;
        RECT 1398.710 365.725 1398.990 366.005 ;
        RECT 1389.410 365.105 1389.690 365.385 ;
        RECT 1390.030 365.105 1390.310 365.385 ;
        RECT 1390.650 365.105 1390.930 365.385 ;
        RECT 1391.270 365.105 1391.550 365.385 ;
        RECT 1391.890 365.105 1392.170 365.385 ;
        RECT 1392.510 365.105 1392.790 365.385 ;
        RECT 1393.130 365.105 1393.410 365.385 ;
        RECT 1393.750 365.105 1394.030 365.385 ;
        RECT 1394.370 365.105 1394.650 365.385 ;
        RECT 1394.990 365.105 1395.270 365.385 ;
        RECT 1395.610 365.105 1395.890 365.385 ;
        RECT 1396.230 365.105 1396.510 365.385 ;
        RECT 1396.850 365.105 1397.130 365.385 ;
        RECT 1397.470 365.105 1397.750 365.385 ;
        RECT 1398.090 365.105 1398.370 365.385 ;
        RECT 1398.710 365.105 1398.990 365.385 ;
        RECT 1389.410 364.485 1389.690 364.765 ;
        RECT 1390.030 364.485 1390.310 364.765 ;
        RECT 1390.650 364.485 1390.930 364.765 ;
        RECT 1391.270 364.485 1391.550 364.765 ;
        RECT 1391.890 364.485 1392.170 364.765 ;
        RECT 1392.510 364.485 1392.790 364.765 ;
        RECT 1393.130 364.485 1393.410 364.765 ;
        RECT 1393.750 364.485 1394.030 364.765 ;
        RECT 1394.370 364.485 1394.650 364.765 ;
        RECT 1394.990 364.485 1395.270 364.765 ;
        RECT 1395.610 364.485 1395.890 364.765 ;
        RECT 1396.230 364.485 1396.510 364.765 ;
        RECT 1396.850 364.485 1397.130 364.765 ;
        RECT 1397.470 364.485 1397.750 364.765 ;
        RECT 1398.090 364.485 1398.370 364.765 ;
        RECT 1398.710 364.485 1398.990 364.765 ;
        RECT 1389.410 363.865 1389.690 364.145 ;
        RECT 1390.030 363.865 1390.310 364.145 ;
        RECT 1390.650 363.865 1390.930 364.145 ;
        RECT 1391.270 363.865 1391.550 364.145 ;
        RECT 1391.890 363.865 1392.170 364.145 ;
        RECT 1392.510 363.865 1392.790 364.145 ;
        RECT 1393.130 363.865 1393.410 364.145 ;
        RECT 1393.750 363.865 1394.030 364.145 ;
        RECT 1394.370 363.865 1394.650 364.145 ;
        RECT 1394.990 363.865 1395.270 364.145 ;
        RECT 1395.610 363.865 1395.890 364.145 ;
        RECT 1396.230 363.865 1396.510 364.145 ;
        RECT 1396.850 363.865 1397.130 364.145 ;
        RECT 1397.470 363.865 1397.750 364.145 ;
        RECT 1398.090 363.865 1398.370 364.145 ;
        RECT 1398.710 363.865 1398.990 364.145 ;
        RECT 1389.410 363.245 1389.690 363.525 ;
        RECT 1390.030 363.245 1390.310 363.525 ;
        RECT 1390.650 363.245 1390.930 363.525 ;
        RECT 1391.270 363.245 1391.550 363.525 ;
        RECT 1391.890 363.245 1392.170 363.525 ;
        RECT 1392.510 363.245 1392.790 363.525 ;
        RECT 1393.130 363.245 1393.410 363.525 ;
        RECT 1393.750 363.245 1394.030 363.525 ;
        RECT 1394.370 363.245 1394.650 363.525 ;
        RECT 1394.990 363.245 1395.270 363.525 ;
        RECT 1395.610 363.245 1395.890 363.525 ;
        RECT 1396.230 363.245 1396.510 363.525 ;
        RECT 1396.850 363.245 1397.130 363.525 ;
        RECT 1397.470 363.245 1397.750 363.525 ;
        RECT 1398.090 363.245 1398.370 363.525 ;
        RECT 1398.710 363.245 1398.990 363.525 ;
        RECT 1389.410 362.625 1389.690 362.905 ;
        RECT 1390.030 362.625 1390.310 362.905 ;
        RECT 1390.650 362.625 1390.930 362.905 ;
        RECT 1391.270 362.625 1391.550 362.905 ;
        RECT 1391.890 362.625 1392.170 362.905 ;
        RECT 1392.510 362.625 1392.790 362.905 ;
        RECT 1393.130 362.625 1393.410 362.905 ;
        RECT 1393.750 362.625 1394.030 362.905 ;
        RECT 1394.370 362.625 1394.650 362.905 ;
        RECT 1394.990 362.625 1395.270 362.905 ;
        RECT 1395.610 362.625 1395.890 362.905 ;
        RECT 1396.230 362.625 1396.510 362.905 ;
        RECT 1396.850 362.625 1397.130 362.905 ;
        RECT 1397.470 362.625 1397.750 362.905 ;
        RECT 1398.090 362.625 1398.370 362.905 ;
        RECT 1398.710 362.625 1398.990 362.905 ;
        RECT 1389.410 362.005 1389.690 362.285 ;
        RECT 1390.030 362.005 1390.310 362.285 ;
        RECT 1390.650 362.005 1390.930 362.285 ;
        RECT 1391.270 362.005 1391.550 362.285 ;
        RECT 1391.890 362.005 1392.170 362.285 ;
        RECT 1392.510 362.005 1392.790 362.285 ;
        RECT 1393.130 362.005 1393.410 362.285 ;
        RECT 1393.750 362.005 1394.030 362.285 ;
        RECT 1394.370 362.005 1394.650 362.285 ;
        RECT 1394.990 362.005 1395.270 362.285 ;
        RECT 1395.610 362.005 1395.890 362.285 ;
        RECT 1396.230 362.005 1396.510 362.285 ;
        RECT 1396.850 362.005 1397.130 362.285 ;
        RECT 1397.470 362.005 1397.750 362.285 ;
        RECT 1398.090 362.005 1398.370 362.285 ;
        RECT 1398.710 362.005 1398.990 362.285 ;
        RECT 1389.410 361.385 1389.690 361.665 ;
        RECT 1390.030 361.385 1390.310 361.665 ;
        RECT 1390.650 361.385 1390.930 361.665 ;
        RECT 1391.270 361.385 1391.550 361.665 ;
        RECT 1391.890 361.385 1392.170 361.665 ;
        RECT 1392.510 361.385 1392.790 361.665 ;
        RECT 1393.130 361.385 1393.410 361.665 ;
        RECT 1393.750 361.385 1394.030 361.665 ;
        RECT 1394.370 361.385 1394.650 361.665 ;
        RECT 1394.990 361.385 1395.270 361.665 ;
        RECT 1395.610 361.385 1395.890 361.665 ;
        RECT 1396.230 361.385 1396.510 361.665 ;
        RECT 1396.850 361.385 1397.130 361.665 ;
        RECT 1397.470 361.385 1397.750 361.665 ;
        RECT 1398.090 361.385 1398.370 361.665 ;
        RECT 1398.710 361.385 1398.990 361.665 ;
        RECT 1389.410 360.765 1389.690 361.045 ;
        RECT 1390.030 360.765 1390.310 361.045 ;
        RECT 1390.650 360.765 1390.930 361.045 ;
        RECT 1391.270 360.765 1391.550 361.045 ;
        RECT 1391.890 360.765 1392.170 361.045 ;
        RECT 1392.510 360.765 1392.790 361.045 ;
        RECT 1393.130 360.765 1393.410 361.045 ;
        RECT 1393.750 360.765 1394.030 361.045 ;
        RECT 1394.370 360.765 1394.650 361.045 ;
        RECT 1394.990 360.765 1395.270 361.045 ;
        RECT 1395.610 360.765 1395.890 361.045 ;
        RECT 1396.230 360.765 1396.510 361.045 ;
        RECT 1396.850 360.765 1397.130 361.045 ;
        RECT 1397.470 360.765 1397.750 361.045 ;
        RECT 1398.090 360.765 1398.370 361.045 ;
        RECT 1398.710 360.765 1398.990 361.045 ;
        RECT 1401.260 369.445 1401.540 369.725 ;
        RECT 1401.880 369.445 1402.160 369.725 ;
        RECT 1402.500 369.445 1402.780 369.725 ;
        RECT 1403.120 369.445 1403.400 369.725 ;
        RECT 1403.740 369.445 1404.020 369.725 ;
        RECT 1404.360 369.445 1404.640 369.725 ;
        RECT 1404.980 369.445 1405.260 369.725 ;
        RECT 1405.600 369.445 1405.880 369.725 ;
        RECT 1406.220 369.445 1406.500 369.725 ;
        RECT 1406.840 369.445 1407.120 369.725 ;
        RECT 1407.460 369.445 1407.740 369.725 ;
        RECT 1408.080 369.445 1408.360 369.725 ;
        RECT 1408.700 369.445 1408.980 369.725 ;
        RECT 1409.320 369.445 1409.600 369.725 ;
        RECT 1409.940 369.445 1410.220 369.725 ;
        RECT 1410.560 369.445 1410.840 369.725 ;
        RECT 1401.260 368.825 1401.540 369.105 ;
        RECT 1401.880 368.825 1402.160 369.105 ;
        RECT 1402.500 368.825 1402.780 369.105 ;
        RECT 1403.120 368.825 1403.400 369.105 ;
        RECT 1403.740 368.825 1404.020 369.105 ;
        RECT 1404.360 368.825 1404.640 369.105 ;
        RECT 1404.980 368.825 1405.260 369.105 ;
        RECT 1405.600 368.825 1405.880 369.105 ;
        RECT 1406.220 368.825 1406.500 369.105 ;
        RECT 1406.840 368.825 1407.120 369.105 ;
        RECT 1407.460 368.825 1407.740 369.105 ;
        RECT 1408.080 368.825 1408.360 369.105 ;
        RECT 1408.700 368.825 1408.980 369.105 ;
        RECT 1409.320 368.825 1409.600 369.105 ;
        RECT 1409.940 368.825 1410.220 369.105 ;
        RECT 1410.560 368.825 1410.840 369.105 ;
        RECT 1401.260 368.205 1401.540 368.485 ;
        RECT 1401.880 368.205 1402.160 368.485 ;
        RECT 1402.500 368.205 1402.780 368.485 ;
        RECT 1403.120 368.205 1403.400 368.485 ;
        RECT 1403.740 368.205 1404.020 368.485 ;
        RECT 1404.360 368.205 1404.640 368.485 ;
        RECT 1404.980 368.205 1405.260 368.485 ;
        RECT 1405.600 368.205 1405.880 368.485 ;
        RECT 1406.220 368.205 1406.500 368.485 ;
        RECT 1406.840 368.205 1407.120 368.485 ;
        RECT 1407.460 368.205 1407.740 368.485 ;
        RECT 1408.080 368.205 1408.360 368.485 ;
        RECT 1408.700 368.205 1408.980 368.485 ;
        RECT 1409.320 368.205 1409.600 368.485 ;
        RECT 1409.940 368.205 1410.220 368.485 ;
        RECT 1410.560 368.205 1410.840 368.485 ;
        RECT 1401.260 367.585 1401.540 367.865 ;
        RECT 1401.880 367.585 1402.160 367.865 ;
        RECT 1402.500 367.585 1402.780 367.865 ;
        RECT 1403.120 367.585 1403.400 367.865 ;
        RECT 1403.740 367.585 1404.020 367.865 ;
        RECT 1404.360 367.585 1404.640 367.865 ;
        RECT 1404.980 367.585 1405.260 367.865 ;
        RECT 1405.600 367.585 1405.880 367.865 ;
        RECT 1406.220 367.585 1406.500 367.865 ;
        RECT 1406.840 367.585 1407.120 367.865 ;
        RECT 1407.460 367.585 1407.740 367.865 ;
        RECT 1408.080 367.585 1408.360 367.865 ;
        RECT 1408.700 367.585 1408.980 367.865 ;
        RECT 1409.320 367.585 1409.600 367.865 ;
        RECT 1409.940 367.585 1410.220 367.865 ;
        RECT 1410.560 367.585 1410.840 367.865 ;
        RECT 1401.260 366.965 1401.540 367.245 ;
        RECT 1401.880 366.965 1402.160 367.245 ;
        RECT 1402.500 366.965 1402.780 367.245 ;
        RECT 1403.120 366.965 1403.400 367.245 ;
        RECT 1403.740 366.965 1404.020 367.245 ;
        RECT 1404.360 366.965 1404.640 367.245 ;
        RECT 1404.980 366.965 1405.260 367.245 ;
        RECT 1405.600 366.965 1405.880 367.245 ;
        RECT 1406.220 366.965 1406.500 367.245 ;
        RECT 1406.840 366.965 1407.120 367.245 ;
        RECT 1407.460 366.965 1407.740 367.245 ;
        RECT 1408.080 366.965 1408.360 367.245 ;
        RECT 1408.700 366.965 1408.980 367.245 ;
        RECT 1409.320 366.965 1409.600 367.245 ;
        RECT 1409.940 366.965 1410.220 367.245 ;
        RECT 1410.560 366.965 1410.840 367.245 ;
        RECT 1401.260 366.345 1401.540 366.625 ;
        RECT 1401.880 366.345 1402.160 366.625 ;
        RECT 1402.500 366.345 1402.780 366.625 ;
        RECT 1403.120 366.345 1403.400 366.625 ;
        RECT 1403.740 366.345 1404.020 366.625 ;
        RECT 1404.360 366.345 1404.640 366.625 ;
        RECT 1404.980 366.345 1405.260 366.625 ;
        RECT 1405.600 366.345 1405.880 366.625 ;
        RECT 1406.220 366.345 1406.500 366.625 ;
        RECT 1406.840 366.345 1407.120 366.625 ;
        RECT 1407.460 366.345 1407.740 366.625 ;
        RECT 1408.080 366.345 1408.360 366.625 ;
        RECT 1408.700 366.345 1408.980 366.625 ;
        RECT 1409.320 366.345 1409.600 366.625 ;
        RECT 1409.940 366.345 1410.220 366.625 ;
        RECT 1410.560 366.345 1410.840 366.625 ;
        RECT 1401.260 365.725 1401.540 366.005 ;
        RECT 1401.880 365.725 1402.160 366.005 ;
        RECT 1402.500 365.725 1402.780 366.005 ;
        RECT 1403.120 365.725 1403.400 366.005 ;
        RECT 1403.740 365.725 1404.020 366.005 ;
        RECT 1404.360 365.725 1404.640 366.005 ;
        RECT 1404.980 365.725 1405.260 366.005 ;
        RECT 1405.600 365.725 1405.880 366.005 ;
        RECT 1406.220 365.725 1406.500 366.005 ;
        RECT 1406.840 365.725 1407.120 366.005 ;
        RECT 1407.460 365.725 1407.740 366.005 ;
        RECT 1408.080 365.725 1408.360 366.005 ;
        RECT 1408.700 365.725 1408.980 366.005 ;
        RECT 1409.320 365.725 1409.600 366.005 ;
        RECT 1409.940 365.725 1410.220 366.005 ;
        RECT 1410.560 365.725 1410.840 366.005 ;
        RECT 1401.260 365.105 1401.540 365.385 ;
        RECT 1401.880 365.105 1402.160 365.385 ;
        RECT 1402.500 365.105 1402.780 365.385 ;
        RECT 1403.120 365.105 1403.400 365.385 ;
        RECT 1403.740 365.105 1404.020 365.385 ;
        RECT 1404.360 365.105 1404.640 365.385 ;
        RECT 1404.980 365.105 1405.260 365.385 ;
        RECT 1405.600 365.105 1405.880 365.385 ;
        RECT 1406.220 365.105 1406.500 365.385 ;
        RECT 1406.840 365.105 1407.120 365.385 ;
        RECT 1407.460 365.105 1407.740 365.385 ;
        RECT 1408.080 365.105 1408.360 365.385 ;
        RECT 1408.700 365.105 1408.980 365.385 ;
        RECT 1409.320 365.105 1409.600 365.385 ;
        RECT 1409.940 365.105 1410.220 365.385 ;
        RECT 1410.560 365.105 1410.840 365.385 ;
        RECT 1401.260 364.485 1401.540 364.765 ;
        RECT 1401.880 364.485 1402.160 364.765 ;
        RECT 1402.500 364.485 1402.780 364.765 ;
        RECT 1403.120 364.485 1403.400 364.765 ;
        RECT 1403.740 364.485 1404.020 364.765 ;
        RECT 1404.360 364.485 1404.640 364.765 ;
        RECT 1404.980 364.485 1405.260 364.765 ;
        RECT 1405.600 364.485 1405.880 364.765 ;
        RECT 1406.220 364.485 1406.500 364.765 ;
        RECT 1406.840 364.485 1407.120 364.765 ;
        RECT 1407.460 364.485 1407.740 364.765 ;
        RECT 1408.080 364.485 1408.360 364.765 ;
        RECT 1408.700 364.485 1408.980 364.765 ;
        RECT 1409.320 364.485 1409.600 364.765 ;
        RECT 1409.940 364.485 1410.220 364.765 ;
        RECT 1410.560 364.485 1410.840 364.765 ;
        RECT 1401.260 363.865 1401.540 364.145 ;
        RECT 1401.880 363.865 1402.160 364.145 ;
        RECT 1402.500 363.865 1402.780 364.145 ;
        RECT 1403.120 363.865 1403.400 364.145 ;
        RECT 1403.740 363.865 1404.020 364.145 ;
        RECT 1404.360 363.865 1404.640 364.145 ;
        RECT 1404.980 363.865 1405.260 364.145 ;
        RECT 1405.600 363.865 1405.880 364.145 ;
        RECT 1406.220 363.865 1406.500 364.145 ;
        RECT 1406.840 363.865 1407.120 364.145 ;
        RECT 1407.460 363.865 1407.740 364.145 ;
        RECT 1408.080 363.865 1408.360 364.145 ;
        RECT 1408.700 363.865 1408.980 364.145 ;
        RECT 1409.320 363.865 1409.600 364.145 ;
        RECT 1409.940 363.865 1410.220 364.145 ;
        RECT 1410.560 363.865 1410.840 364.145 ;
        RECT 1401.260 363.245 1401.540 363.525 ;
        RECT 1401.880 363.245 1402.160 363.525 ;
        RECT 1402.500 363.245 1402.780 363.525 ;
        RECT 1403.120 363.245 1403.400 363.525 ;
        RECT 1403.740 363.245 1404.020 363.525 ;
        RECT 1404.360 363.245 1404.640 363.525 ;
        RECT 1404.980 363.245 1405.260 363.525 ;
        RECT 1405.600 363.245 1405.880 363.525 ;
        RECT 1406.220 363.245 1406.500 363.525 ;
        RECT 1406.840 363.245 1407.120 363.525 ;
        RECT 1407.460 363.245 1407.740 363.525 ;
        RECT 1408.080 363.245 1408.360 363.525 ;
        RECT 1408.700 363.245 1408.980 363.525 ;
        RECT 1409.320 363.245 1409.600 363.525 ;
        RECT 1409.940 363.245 1410.220 363.525 ;
        RECT 1410.560 363.245 1410.840 363.525 ;
        RECT 1401.260 362.625 1401.540 362.905 ;
        RECT 1401.880 362.625 1402.160 362.905 ;
        RECT 1402.500 362.625 1402.780 362.905 ;
        RECT 1403.120 362.625 1403.400 362.905 ;
        RECT 1403.740 362.625 1404.020 362.905 ;
        RECT 1404.360 362.625 1404.640 362.905 ;
        RECT 1404.980 362.625 1405.260 362.905 ;
        RECT 1405.600 362.625 1405.880 362.905 ;
        RECT 1406.220 362.625 1406.500 362.905 ;
        RECT 1406.840 362.625 1407.120 362.905 ;
        RECT 1407.460 362.625 1407.740 362.905 ;
        RECT 1408.080 362.625 1408.360 362.905 ;
        RECT 1408.700 362.625 1408.980 362.905 ;
        RECT 1409.320 362.625 1409.600 362.905 ;
        RECT 1409.940 362.625 1410.220 362.905 ;
        RECT 1410.560 362.625 1410.840 362.905 ;
        RECT 1401.260 362.005 1401.540 362.285 ;
        RECT 1401.880 362.005 1402.160 362.285 ;
        RECT 1402.500 362.005 1402.780 362.285 ;
        RECT 1403.120 362.005 1403.400 362.285 ;
        RECT 1403.740 362.005 1404.020 362.285 ;
        RECT 1404.360 362.005 1404.640 362.285 ;
        RECT 1404.980 362.005 1405.260 362.285 ;
        RECT 1405.600 362.005 1405.880 362.285 ;
        RECT 1406.220 362.005 1406.500 362.285 ;
        RECT 1406.840 362.005 1407.120 362.285 ;
        RECT 1407.460 362.005 1407.740 362.285 ;
        RECT 1408.080 362.005 1408.360 362.285 ;
        RECT 1408.700 362.005 1408.980 362.285 ;
        RECT 1409.320 362.005 1409.600 362.285 ;
        RECT 1409.940 362.005 1410.220 362.285 ;
        RECT 1410.560 362.005 1410.840 362.285 ;
        RECT 1401.260 361.385 1401.540 361.665 ;
        RECT 1401.880 361.385 1402.160 361.665 ;
        RECT 1402.500 361.385 1402.780 361.665 ;
        RECT 1403.120 361.385 1403.400 361.665 ;
        RECT 1403.740 361.385 1404.020 361.665 ;
        RECT 1404.360 361.385 1404.640 361.665 ;
        RECT 1404.980 361.385 1405.260 361.665 ;
        RECT 1405.600 361.385 1405.880 361.665 ;
        RECT 1406.220 361.385 1406.500 361.665 ;
        RECT 1406.840 361.385 1407.120 361.665 ;
        RECT 1407.460 361.385 1407.740 361.665 ;
        RECT 1408.080 361.385 1408.360 361.665 ;
        RECT 1408.700 361.385 1408.980 361.665 ;
        RECT 1409.320 361.385 1409.600 361.665 ;
        RECT 1409.940 361.385 1410.220 361.665 ;
        RECT 1410.560 361.385 1410.840 361.665 ;
        RECT 1401.260 360.765 1401.540 361.045 ;
        RECT 1401.880 360.765 1402.160 361.045 ;
        RECT 1402.500 360.765 1402.780 361.045 ;
        RECT 1403.120 360.765 1403.400 361.045 ;
        RECT 1403.740 360.765 1404.020 361.045 ;
        RECT 1404.360 360.765 1404.640 361.045 ;
        RECT 1404.980 360.765 1405.260 361.045 ;
        RECT 1405.600 360.765 1405.880 361.045 ;
        RECT 1406.220 360.765 1406.500 361.045 ;
        RECT 1406.840 360.765 1407.120 361.045 ;
        RECT 1407.460 360.765 1407.740 361.045 ;
        RECT 1408.080 360.765 1408.360 361.045 ;
        RECT 1408.700 360.765 1408.980 361.045 ;
        RECT 1409.320 360.765 1409.600 361.045 ;
        RECT 1409.940 360.765 1410.220 361.045 ;
        RECT 1410.560 360.765 1410.840 361.045 ;
        RECT 1414.410 369.445 1414.690 369.725 ;
        RECT 1415.030 369.445 1415.310 369.725 ;
        RECT 1415.650 369.445 1415.930 369.725 ;
        RECT 1416.270 369.445 1416.550 369.725 ;
        RECT 1416.890 369.445 1417.170 369.725 ;
        RECT 1417.510 369.445 1417.790 369.725 ;
        RECT 1418.130 369.445 1418.410 369.725 ;
        RECT 1418.750 369.445 1419.030 369.725 ;
        RECT 1419.370 369.445 1419.650 369.725 ;
        RECT 1414.410 368.825 1414.690 369.105 ;
        RECT 1415.030 368.825 1415.310 369.105 ;
        RECT 1415.650 368.825 1415.930 369.105 ;
        RECT 1416.270 368.825 1416.550 369.105 ;
        RECT 1416.890 368.825 1417.170 369.105 ;
        RECT 1417.510 368.825 1417.790 369.105 ;
        RECT 1418.130 368.825 1418.410 369.105 ;
        RECT 1418.750 368.825 1419.030 369.105 ;
        RECT 1419.370 368.825 1419.650 369.105 ;
        RECT 1414.410 368.205 1414.690 368.485 ;
        RECT 1415.030 368.205 1415.310 368.485 ;
        RECT 1415.650 368.205 1415.930 368.485 ;
        RECT 1416.270 368.205 1416.550 368.485 ;
        RECT 1416.890 368.205 1417.170 368.485 ;
        RECT 1417.510 368.205 1417.790 368.485 ;
        RECT 1418.130 368.205 1418.410 368.485 ;
        RECT 1418.750 368.205 1419.030 368.485 ;
        RECT 1419.370 368.205 1419.650 368.485 ;
        RECT 1414.410 367.585 1414.690 367.865 ;
        RECT 1415.030 367.585 1415.310 367.865 ;
        RECT 1415.650 367.585 1415.930 367.865 ;
        RECT 1416.270 367.585 1416.550 367.865 ;
        RECT 1416.890 367.585 1417.170 367.865 ;
        RECT 1417.510 367.585 1417.790 367.865 ;
        RECT 1418.130 367.585 1418.410 367.865 ;
        RECT 1418.750 367.585 1419.030 367.865 ;
        RECT 1419.370 367.585 1419.650 367.865 ;
        RECT 1414.410 366.965 1414.690 367.245 ;
        RECT 1415.030 366.965 1415.310 367.245 ;
        RECT 1415.650 366.965 1415.930 367.245 ;
        RECT 1416.270 366.965 1416.550 367.245 ;
        RECT 1416.890 366.965 1417.170 367.245 ;
        RECT 1417.510 366.965 1417.790 367.245 ;
        RECT 1418.130 366.965 1418.410 367.245 ;
        RECT 1418.750 366.965 1419.030 367.245 ;
        RECT 1419.370 366.965 1419.650 367.245 ;
        RECT 1414.410 366.345 1414.690 366.625 ;
        RECT 1415.030 366.345 1415.310 366.625 ;
        RECT 1415.650 366.345 1415.930 366.625 ;
        RECT 1416.270 366.345 1416.550 366.625 ;
        RECT 1416.890 366.345 1417.170 366.625 ;
        RECT 1417.510 366.345 1417.790 366.625 ;
        RECT 1418.130 366.345 1418.410 366.625 ;
        RECT 1418.750 366.345 1419.030 366.625 ;
        RECT 1419.370 366.345 1419.650 366.625 ;
        RECT 1414.410 365.725 1414.690 366.005 ;
        RECT 1415.030 365.725 1415.310 366.005 ;
        RECT 1415.650 365.725 1415.930 366.005 ;
        RECT 1416.270 365.725 1416.550 366.005 ;
        RECT 1416.890 365.725 1417.170 366.005 ;
        RECT 1417.510 365.725 1417.790 366.005 ;
        RECT 1418.130 365.725 1418.410 366.005 ;
        RECT 1418.750 365.725 1419.030 366.005 ;
        RECT 1419.370 365.725 1419.650 366.005 ;
        RECT 1414.410 365.105 1414.690 365.385 ;
        RECT 1415.030 365.105 1415.310 365.385 ;
        RECT 1415.650 365.105 1415.930 365.385 ;
        RECT 1416.270 365.105 1416.550 365.385 ;
        RECT 1416.890 365.105 1417.170 365.385 ;
        RECT 1417.510 365.105 1417.790 365.385 ;
        RECT 1418.130 365.105 1418.410 365.385 ;
        RECT 1418.750 365.105 1419.030 365.385 ;
        RECT 1419.370 365.105 1419.650 365.385 ;
        RECT 1414.410 364.485 1414.690 364.765 ;
        RECT 1415.030 364.485 1415.310 364.765 ;
        RECT 1415.650 364.485 1415.930 364.765 ;
        RECT 1416.270 364.485 1416.550 364.765 ;
        RECT 1416.890 364.485 1417.170 364.765 ;
        RECT 1417.510 364.485 1417.790 364.765 ;
        RECT 1418.130 364.485 1418.410 364.765 ;
        RECT 1418.750 364.485 1419.030 364.765 ;
        RECT 1419.370 364.485 1419.650 364.765 ;
        RECT 1414.410 363.865 1414.690 364.145 ;
        RECT 1415.030 363.865 1415.310 364.145 ;
        RECT 1415.650 363.865 1415.930 364.145 ;
        RECT 1416.270 363.865 1416.550 364.145 ;
        RECT 1416.890 363.865 1417.170 364.145 ;
        RECT 1417.510 363.865 1417.790 364.145 ;
        RECT 1418.130 363.865 1418.410 364.145 ;
        RECT 1418.750 363.865 1419.030 364.145 ;
        RECT 1419.370 363.865 1419.650 364.145 ;
        RECT 1414.410 363.245 1414.690 363.525 ;
        RECT 1415.030 363.245 1415.310 363.525 ;
        RECT 1415.650 363.245 1415.930 363.525 ;
        RECT 1416.270 363.245 1416.550 363.525 ;
        RECT 1416.890 363.245 1417.170 363.525 ;
        RECT 1417.510 363.245 1417.790 363.525 ;
        RECT 1418.130 363.245 1418.410 363.525 ;
        RECT 1418.750 363.245 1419.030 363.525 ;
        RECT 1419.370 363.245 1419.650 363.525 ;
        RECT 1414.410 362.625 1414.690 362.905 ;
        RECT 1415.030 362.625 1415.310 362.905 ;
        RECT 1415.650 362.625 1415.930 362.905 ;
        RECT 1416.270 362.625 1416.550 362.905 ;
        RECT 1416.890 362.625 1417.170 362.905 ;
        RECT 1417.510 362.625 1417.790 362.905 ;
        RECT 1418.130 362.625 1418.410 362.905 ;
        RECT 1418.750 362.625 1419.030 362.905 ;
        RECT 1419.370 362.625 1419.650 362.905 ;
        RECT 1414.410 362.005 1414.690 362.285 ;
        RECT 1415.030 362.005 1415.310 362.285 ;
        RECT 1415.650 362.005 1415.930 362.285 ;
        RECT 1416.270 362.005 1416.550 362.285 ;
        RECT 1416.890 362.005 1417.170 362.285 ;
        RECT 1417.510 362.005 1417.790 362.285 ;
        RECT 1418.130 362.005 1418.410 362.285 ;
        RECT 1418.750 362.005 1419.030 362.285 ;
        RECT 1419.370 362.005 1419.650 362.285 ;
        RECT 1414.410 361.385 1414.690 361.665 ;
        RECT 1415.030 361.385 1415.310 361.665 ;
        RECT 1415.650 361.385 1415.930 361.665 ;
        RECT 1416.270 361.385 1416.550 361.665 ;
        RECT 1416.890 361.385 1417.170 361.665 ;
        RECT 1417.510 361.385 1417.790 361.665 ;
        RECT 1418.130 361.385 1418.410 361.665 ;
        RECT 1418.750 361.385 1419.030 361.665 ;
        RECT 1419.370 361.385 1419.650 361.665 ;
        RECT 1414.410 360.765 1414.690 361.045 ;
        RECT 1415.030 360.765 1415.310 361.045 ;
        RECT 1415.650 360.765 1415.930 361.045 ;
        RECT 1416.270 360.765 1416.550 361.045 ;
        RECT 1416.890 360.765 1417.170 361.045 ;
        RECT 1417.510 360.765 1417.790 361.045 ;
        RECT 1418.130 360.765 1418.410 361.045 ;
        RECT 1418.750 360.765 1419.030 361.045 ;
        RECT 1419.370 360.765 1419.650 361.045 ;
        RECT 3001.630 369.445 3001.910 369.725 ;
        RECT 3002.250 369.445 3002.530 369.725 ;
        RECT 3002.870 369.445 3003.150 369.725 ;
        RECT 3003.490 369.445 3003.770 369.725 ;
        RECT 3004.110 369.445 3004.390 369.725 ;
        RECT 3004.730 369.445 3005.010 369.725 ;
        RECT 3005.350 369.445 3005.630 369.725 ;
        RECT 3005.970 369.445 3006.250 369.725 ;
        RECT 3006.590 369.445 3006.870 369.725 ;
        RECT 3007.210 369.445 3007.490 369.725 ;
        RECT 3007.830 369.445 3008.110 369.725 ;
        RECT 3008.450 369.445 3008.730 369.725 ;
        RECT 3009.070 369.445 3009.350 369.725 ;
        RECT 3009.690 369.445 3009.970 369.725 ;
        RECT 3010.310 369.445 3010.590 369.725 ;
        RECT 3001.630 368.825 3001.910 369.105 ;
        RECT 3002.250 368.825 3002.530 369.105 ;
        RECT 3002.870 368.825 3003.150 369.105 ;
        RECT 3003.490 368.825 3003.770 369.105 ;
        RECT 3004.110 368.825 3004.390 369.105 ;
        RECT 3004.730 368.825 3005.010 369.105 ;
        RECT 3005.350 368.825 3005.630 369.105 ;
        RECT 3005.970 368.825 3006.250 369.105 ;
        RECT 3006.590 368.825 3006.870 369.105 ;
        RECT 3007.210 368.825 3007.490 369.105 ;
        RECT 3007.830 368.825 3008.110 369.105 ;
        RECT 3008.450 368.825 3008.730 369.105 ;
        RECT 3009.070 368.825 3009.350 369.105 ;
        RECT 3009.690 368.825 3009.970 369.105 ;
        RECT 3010.310 368.825 3010.590 369.105 ;
        RECT 3001.630 368.205 3001.910 368.485 ;
        RECT 3002.250 368.205 3002.530 368.485 ;
        RECT 3002.870 368.205 3003.150 368.485 ;
        RECT 3003.490 368.205 3003.770 368.485 ;
        RECT 3004.110 368.205 3004.390 368.485 ;
        RECT 3004.730 368.205 3005.010 368.485 ;
        RECT 3005.350 368.205 3005.630 368.485 ;
        RECT 3005.970 368.205 3006.250 368.485 ;
        RECT 3006.590 368.205 3006.870 368.485 ;
        RECT 3007.210 368.205 3007.490 368.485 ;
        RECT 3007.830 368.205 3008.110 368.485 ;
        RECT 3008.450 368.205 3008.730 368.485 ;
        RECT 3009.070 368.205 3009.350 368.485 ;
        RECT 3009.690 368.205 3009.970 368.485 ;
        RECT 3010.310 368.205 3010.590 368.485 ;
        RECT 3001.630 367.585 3001.910 367.865 ;
        RECT 3002.250 367.585 3002.530 367.865 ;
        RECT 3002.870 367.585 3003.150 367.865 ;
        RECT 3003.490 367.585 3003.770 367.865 ;
        RECT 3004.110 367.585 3004.390 367.865 ;
        RECT 3004.730 367.585 3005.010 367.865 ;
        RECT 3005.350 367.585 3005.630 367.865 ;
        RECT 3005.970 367.585 3006.250 367.865 ;
        RECT 3006.590 367.585 3006.870 367.865 ;
        RECT 3007.210 367.585 3007.490 367.865 ;
        RECT 3007.830 367.585 3008.110 367.865 ;
        RECT 3008.450 367.585 3008.730 367.865 ;
        RECT 3009.070 367.585 3009.350 367.865 ;
        RECT 3009.690 367.585 3009.970 367.865 ;
        RECT 3010.310 367.585 3010.590 367.865 ;
        RECT 3001.630 366.965 3001.910 367.245 ;
        RECT 3002.250 366.965 3002.530 367.245 ;
        RECT 3002.870 366.965 3003.150 367.245 ;
        RECT 3003.490 366.965 3003.770 367.245 ;
        RECT 3004.110 366.965 3004.390 367.245 ;
        RECT 3004.730 366.965 3005.010 367.245 ;
        RECT 3005.350 366.965 3005.630 367.245 ;
        RECT 3005.970 366.965 3006.250 367.245 ;
        RECT 3006.590 366.965 3006.870 367.245 ;
        RECT 3007.210 366.965 3007.490 367.245 ;
        RECT 3007.830 366.965 3008.110 367.245 ;
        RECT 3008.450 366.965 3008.730 367.245 ;
        RECT 3009.070 366.965 3009.350 367.245 ;
        RECT 3009.690 366.965 3009.970 367.245 ;
        RECT 3010.310 366.965 3010.590 367.245 ;
        RECT 3001.630 366.345 3001.910 366.625 ;
        RECT 3002.250 366.345 3002.530 366.625 ;
        RECT 3002.870 366.345 3003.150 366.625 ;
        RECT 3003.490 366.345 3003.770 366.625 ;
        RECT 3004.110 366.345 3004.390 366.625 ;
        RECT 3004.730 366.345 3005.010 366.625 ;
        RECT 3005.350 366.345 3005.630 366.625 ;
        RECT 3005.970 366.345 3006.250 366.625 ;
        RECT 3006.590 366.345 3006.870 366.625 ;
        RECT 3007.210 366.345 3007.490 366.625 ;
        RECT 3007.830 366.345 3008.110 366.625 ;
        RECT 3008.450 366.345 3008.730 366.625 ;
        RECT 3009.070 366.345 3009.350 366.625 ;
        RECT 3009.690 366.345 3009.970 366.625 ;
        RECT 3010.310 366.345 3010.590 366.625 ;
        RECT 3001.630 365.725 3001.910 366.005 ;
        RECT 3002.250 365.725 3002.530 366.005 ;
        RECT 3002.870 365.725 3003.150 366.005 ;
        RECT 3003.490 365.725 3003.770 366.005 ;
        RECT 3004.110 365.725 3004.390 366.005 ;
        RECT 3004.730 365.725 3005.010 366.005 ;
        RECT 3005.350 365.725 3005.630 366.005 ;
        RECT 3005.970 365.725 3006.250 366.005 ;
        RECT 3006.590 365.725 3006.870 366.005 ;
        RECT 3007.210 365.725 3007.490 366.005 ;
        RECT 3007.830 365.725 3008.110 366.005 ;
        RECT 3008.450 365.725 3008.730 366.005 ;
        RECT 3009.070 365.725 3009.350 366.005 ;
        RECT 3009.690 365.725 3009.970 366.005 ;
        RECT 3010.310 365.725 3010.590 366.005 ;
        RECT 3001.630 365.105 3001.910 365.385 ;
        RECT 3002.250 365.105 3002.530 365.385 ;
        RECT 3002.870 365.105 3003.150 365.385 ;
        RECT 3003.490 365.105 3003.770 365.385 ;
        RECT 3004.110 365.105 3004.390 365.385 ;
        RECT 3004.730 365.105 3005.010 365.385 ;
        RECT 3005.350 365.105 3005.630 365.385 ;
        RECT 3005.970 365.105 3006.250 365.385 ;
        RECT 3006.590 365.105 3006.870 365.385 ;
        RECT 3007.210 365.105 3007.490 365.385 ;
        RECT 3007.830 365.105 3008.110 365.385 ;
        RECT 3008.450 365.105 3008.730 365.385 ;
        RECT 3009.070 365.105 3009.350 365.385 ;
        RECT 3009.690 365.105 3009.970 365.385 ;
        RECT 3010.310 365.105 3010.590 365.385 ;
        RECT 3001.630 364.485 3001.910 364.765 ;
        RECT 3002.250 364.485 3002.530 364.765 ;
        RECT 3002.870 364.485 3003.150 364.765 ;
        RECT 3003.490 364.485 3003.770 364.765 ;
        RECT 3004.110 364.485 3004.390 364.765 ;
        RECT 3004.730 364.485 3005.010 364.765 ;
        RECT 3005.350 364.485 3005.630 364.765 ;
        RECT 3005.970 364.485 3006.250 364.765 ;
        RECT 3006.590 364.485 3006.870 364.765 ;
        RECT 3007.210 364.485 3007.490 364.765 ;
        RECT 3007.830 364.485 3008.110 364.765 ;
        RECT 3008.450 364.485 3008.730 364.765 ;
        RECT 3009.070 364.485 3009.350 364.765 ;
        RECT 3009.690 364.485 3009.970 364.765 ;
        RECT 3010.310 364.485 3010.590 364.765 ;
        RECT 3001.630 363.865 3001.910 364.145 ;
        RECT 3002.250 363.865 3002.530 364.145 ;
        RECT 3002.870 363.865 3003.150 364.145 ;
        RECT 3003.490 363.865 3003.770 364.145 ;
        RECT 3004.110 363.865 3004.390 364.145 ;
        RECT 3004.730 363.865 3005.010 364.145 ;
        RECT 3005.350 363.865 3005.630 364.145 ;
        RECT 3005.970 363.865 3006.250 364.145 ;
        RECT 3006.590 363.865 3006.870 364.145 ;
        RECT 3007.210 363.865 3007.490 364.145 ;
        RECT 3007.830 363.865 3008.110 364.145 ;
        RECT 3008.450 363.865 3008.730 364.145 ;
        RECT 3009.070 363.865 3009.350 364.145 ;
        RECT 3009.690 363.865 3009.970 364.145 ;
        RECT 3010.310 363.865 3010.590 364.145 ;
        RECT 3001.630 363.245 3001.910 363.525 ;
        RECT 3002.250 363.245 3002.530 363.525 ;
        RECT 3002.870 363.245 3003.150 363.525 ;
        RECT 3003.490 363.245 3003.770 363.525 ;
        RECT 3004.110 363.245 3004.390 363.525 ;
        RECT 3004.730 363.245 3005.010 363.525 ;
        RECT 3005.350 363.245 3005.630 363.525 ;
        RECT 3005.970 363.245 3006.250 363.525 ;
        RECT 3006.590 363.245 3006.870 363.525 ;
        RECT 3007.210 363.245 3007.490 363.525 ;
        RECT 3007.830 363.245 3008.110 363.525 ;
        RECT 3008.450 363.245 3008.730 363.525 ;
        RECT 3009.070 363.245 3009.350 363.525 ;
        RECT 3009.690 363.245 3009.970 363.525 ;
        RECT 3010.310 363.245 3010.590 363.525 ;
        RECT 3001.630 362.625 3001.910 362.905 ;
        RECT 3002.250 362.625 3002.530 362.905 ;
        RECT 3002.870 362.625 3003.150 362.905 ;
        RECT 3003.490 362.625 3003.770 362.905 ;
        RECT 3004.110 362.625 3004.390 362.905 ;
        RECT 3004.730 362.625 3005.010 362.905 ;
        RECT 3005.350 362.625 3005.630 362.905 ;
        RECT 3005.970 362.625 3006.250 362.905 ;
        RECT 3006.590 362.625 3006.870 362.905 ;
        RECT 3007.210 362.625 3007.490 362.905 ;
        RECT 3007.830 362.625 3008.110 362.905 ;
        RECT 3008.450 362.625 3008.730 362.905 ;
        RECT 3009.070 362.625 3009.350 362.905 ;
        RECT 3009.690 362.625 3009.970 362.905 ;
        RECT 3010.310 362.625 3010.590 362.905 ;
        RECT 3001.630 362.005 3001.910 362.285 ;
        RECT 3002.250 362.005 3002.530 362.285 ;
        RECT 3002.870 362.005 3003.150 362.285 ;
        RECT 3003.490 362.005 3003.770 362.285 ;
        RECT 3004.110 362.005 3004.390 362.285 ;
        RECT 3004.730 362.005 3005.010 362.285 ;
        RECT 3005.350 362.005 3005.630 362.285 ;
        RECT 3005.970 362.005 3006.250 362.285 ;
        RECT 3006.590 362.005 3006.870 362.285 ;
        RECT 3007.210 362.005 3007.490 362.285 ;
        RECT 3007.830 362.005 3008.110 362.285 ;
        RECT 3008.450 362.005 3008.730 362.285 ;
        RECT 3009.070 362.005 3009.350 362.285 ;
        RECT 3009.690 362.005 3009.970 362.285 ;
        RECT 3010.310 362.005 3010.590 362.285 ;
        RECT 3001.630 361.385 3001.910 361.665 ;
        RECT 3002.250 361.385 3002.530 361.665 ;
        RECT 3002.870 361.385 3003.150 361.665 ;
        RECT 3003.490 361.385 3003.770 361.665 ;
        RECT 3004.110 361.385 3004.390 361.665 ;
        RECT 3004.730 361.385 3005.010 361.665 ;
        RECT 3005.350 361.385 3005.630 361.665 ;
        RECT 3005.970 361.385 3006.250 361.665 ;
        RECT 3006.590 361.385 3006.870 361.665 ;
        RECT 3007.210 361.385 3007.490 361.665 ;
        RECT 3007.830 361.385 3008.110 361.665 ;
        RECT 3008.450 361.385 3008.730 361.665 ;
        RECT 3009.070 361.385 3009.350 361.665 ;
        RECT 3009.690 361.385 3009.970 361.665 ;
        RECT 3010.310 361.385 3010.590 361.665 ;
        RECT 3001.630 360.765 3001.910 361.045 ;
        RECT 3002.250 360.765 3002.530 361.045 ;
        RECT 3002.870 360.765 3003.150 361.045 ;
        RECT 3003.490 360.765 3003.770 361.045 ;
        RECT 3004.110 360.765 3004.390 361.045 ;
        RECT 3004.730 360.765 3005.010 361.045 ;
        RECT 3005.350 360.765 3005.630 361.045 ;
        RECT 3005.970 360.765 3006.250 361.045 ;
        RECT 3006.590 360.765 3006.870 361.045 ;
        RECT 3007.210 360.765 3007.490 361.045 ;
        RECT 3007.830 360.765 3008.110 361.045 ;
        RECT 3008.450 360.765 3008.730 361.045 ;
        RECT 3009.070 360.765 3009.350 361.045 ;
        RECT 3009.690 360.765 3009.970 361.045 ;
        RECT 3010.310 360.765 3010.590 361.045 ;
        RECT 3014.030 369.445 3014.310 369.725 ;
        RECT 3014.650 369.445 3014.930 369.725 ;
        RECT 3015.270 369.445 3015.550 369.725 ;
        RECT 3015.890 369.445 3016.170 369.725 ;
        RECT 3016.510 369.445 3016.790 369.725 ;
        RECT 3017.130 369.445 3017.410 369.725 ;
        RECT 3017.750 369.445 3018.030 369.725 ;
        RECT 3018.370 369.445 3018.650 369.725 ;
        RECT 3018.990 369.445 3019.270 369.725 ;
        RECT 3019.610 369.445 3019.890 369.725 ;
        RECT 3014.030 368.825 3014.310 369.105 ;
        RECT 3014.650 368.825 3014.930 369.105 ;
        RECT 3015.270 368.825 3015.550 369.105 ;
        RECT 3015.890 368.825 3016.170 369.105 ;
        RECT 3016.510 368.825 3016.790 369.105 ;
        RECT 3017.130 368.825 3017.410 369.105 ;
        RECT 3017.750 368.825 3018.030 369.105 ;
        RECT 3018.370 368.825 3018.650 369.105 ;
        RECT 3018.990 368.825 3019.270 369.105 ;
        RECT 3019.610 368.825 3019.890 369.105 ;
        RECT 3014.030 368.205 3014.310 368.485 ;
        RECT 3014.650 368.205 3014.930 368.485 ;
        RECT 3015.270 368.205 3015.550 368.485 ;
        RECT 3015.890 368.205 3016.170 368.485 ;
        RECT 3016.510 368.205 3016.790 368.485 ;
        RECT 3017.130 368.205 3017.410 368.485 ;
        RECT 3017.750 368.205 3018.030 368.485 ;
        RECT 3018.370 368.205 3018.650 368.485 ;
        RECT 3018.990 368.205 3019.270 368.485 ;
        RECT 3019.610 368.205 3019.890 368.485 ;
        RECT 3014.030 367.585 3014.310 367.865 ;
        RECT 3014.650 367.585 3014.930 367.865 ;
        RECT 3015.270 367.585 3015.550 367.865 ;
        RECT 3015.890 367.585 3016.170 367.865 ;
        RECT 3016.510 367.585 3016.790 367.865 ;
        RECT 3017.130 367.585 3017.410 367.865 ;
        RECT 3017.750 367.585 3018.030 367.865 ;
        RECT 3018.370 367.585 3018.650 367.865 ;
        RECT 3018.990 367.585 3019.270 367.865 ;
        RECT 3019.610 367.585 3019.890 367.865 ;
        RECT 3014.030 366.965 3014.310 367.245 ;
        RECT 3014.650 366.965 3014.930 367.245 ;
        RECT 3015.270 366.965 3015.550 367.245 ;
        RECT 3015.890 366.965 3016.170 367.245 ;
        RECT 3016.510 366.965 3016.790 367.245 ;
        RECT 3017.130 366.965 3017.410 367.245 ;
        RECT 3017.750 366.965 3018.030 367.245 ;
        RECT 3018.370 366.965 3018.650 367.245 ;
        RECT 3018.990 366.965 3019.270 367.245 ;
        RECT 3019.610 366.965 3019.890 367.245 ;
        RECT 3014.030 366.345 3014.310 366.625 ;
        RECT 3014.650 366.345 3014.930 366.625 ;
        RECT 3015.270 366.345 3015.550 366.625 ;
        RECT 3015.890 366.345 3016.170 366.625 ;
        RECT 3016.510 366.345 3016.790 366.625 ;
        RECT 3017.130 366.345 3017.410 366.625 ;
        RECT 3017.750 366.345 3018.030 366.625 ;
        RECT 3018.370 366.345 3018.650 366.625 ;
        RECT 3018.990 366.345 3019.270 366.625 ;
        RECT 3019.610 366.345 3019.890 366.625 ;
        RECT 3014.030 365.725 3014.310 366.005 ;
        RECT 3014.650 365.725 3014.930 366.005 ;
        RECT 3015.270 365.725 3015.550 366.005 ;
        RECT 3015.890 365.725 3016.170 366.005 ;
        RECT 3016.510 365.725 3016.790 366.005 ;
        RECT 3017.130 365.725 3017.410 366.005 ;
        RECT 3017.750 365.725 3018.030 366.005 ;
        RECT 3018.370 365.725 3018.650 366.005 ;
        RECT 3018.990 365.725 3019.270 366.005 ;
        RECT 3019.610 365.725 3019.890 366.005 ;
        RECT 3014.030 365.105 3014.310 365.385 ;
        RECT 3014.650 365.105 3014.930 365.385 ;
        RECT 3015.270 365.105 3015.550 365.385 ;
        RECT 3015.890 365.105 3016.170 365.385 ;
        RECT 3016.510 365.105 3016.790 365.385 ;
        RECT 3017.130 365.105 3017.410 365.385 ;
        RECT 3017.750 365.105 3018.030 365.385 ;
        RECT 3018.370 365.105 3018.650 365.385 ;
        RECT 3018.990 365.105 3019.270 365.385 ;
        RECT 3019.610 365.105 3019.890 365.385 ;
        RECT 3014.030 364.485 3014.310 364.765 ;
        RECT 3014.650 364.485 3014.930 364.765 ;
        RECT 3015.270 364.485 3015.550 364.765 ;
        RECT 3015.890 364.485 3016.170 364.765 ;
        RECT 3016.510 364.485 3016.790 364.765 ;
        RECT 3017.130 364.485 3017.410 364.765 ;
        RECT 3017.750 364.485 3018.030 364.765 ;
        RECT 3018.370 364.485 3018.650 364.765 ;
        RECT 3018.990 364.485 3019.270 364.765 ;
        RECT 3019.610 364.485 3019.890 364.765 ;
        RECT 3014.030 363.865 3014.310 364.145 ;
        RECT 3014.650 363.865 3014.930 364.145 ;
        RECT 3015.270 363.865 3015.550 364.145 ;
        RECT 3015.890 363.865 3016.170 364.145 ;
        RECT 3016.510 363.865 3016.790 364.145 ;
        RECT 3017.130 363.865 3017.410 364.145 ;
        RECT 3017.750 363.865 3018.030 364.145 ;
        RECT 3018.370 363.865 3018.650 364.145 ;
        RECT 3018.990 363.865 3019.270 364.145 ;
        RECT 3019.610 363.865 3019.890 364.145 ;
        RECT 3014.030 363.245 3014.310 363.525 ;
        RECT 3014.650 363.245 3014.930 363.525 ;
        RECT 3015.270 363.245 3015.550 363.525 ;
        RECT 3015.890 363.245 3016.170 363.525 ;
        RECT 3016.510 363.245 3016.790 363.525 ;
        RECT 3017.130 363.245 3017.410 363.525 ;
        RECT 3017.750 363.245 3018.030 363.525 ;
        RECT 3018.370 363.245 3018.650 363.525 ;
        RECT 3018.990 363.245 3019.270 363.525 ;
        RECT 3019.610 363.245 3019.890 363.525 ;
        RECT 3014.030 362.625 3014.310 362.905 ;
        RECT 3014.650 362.625 3014.930 362.905 ;
        RECT 3015.270 362.625 3015.550 362.905 ;
        RECT 3015.890 362.625 3016.170 362.905 ;
        RECT 3016.510 362.625 3016.790 362.905 ;
        RECT 3017.130 362.625 3017.410 362.905 ;
        RECT 3017.750 362.625 3018.030 362.905 ;
        RECT 3018.370 362.625 3018.650 362.905 ;
        RECT 3018.990 362.625 3019.270 362.905 ;
        RECT 3019.610 362.625 3019.890 362.905 ;
        RECT 3014.030 362.005 3014.310 362.285 ;
        RECT 3014.650 362.005 3014.930 362.285 ;
        RECT 3015.270 362.005 3015.550 362.285 ;
        RECT 3015.890 362.005 3016.170 362.285 ;
        RECT 3016.510 362.005 3016.790 362.285 ;
        RECT 3017.130 362.005 3017.410 362.285 ;
        RECT 3017.750 362.005 3018.030 362.285 ;
        RECT 3018.370 362.005 3018.650 362.285 ;
        RECT 3018.990 362.005 3019.270 362.285 ;
        RECT 3019.610 362.005 3019.890 362.285 ;
        RECT 3014.030 361.385 3014.310 361.665 ;
        RECT 3014.650 361.385 3014.930 361.665 ;
        RECT 3015.270 361.385 3015.550 361.665 ;
        RECT 3015.890 361.385 3016.170 361.665 ;
        RECT 3016.510 361.385 3016.790 361.665 ;
        RECT 3017.130 361.385 3017.410 361.665 ;
        RECT 3017.750 361.385 3018.030 361.665 ;
        RECT 3018.370 361.385 3018.650 361.665 ;
        RECT 3018.990 361.385 3019.270 361.665 ;
        RECT 3019.610 361.385 3019.890 361.665 ;
        RECT 3014.030 360.765 3014.310 361.045 ;
        RECT 3014.650 360.765 3014.930 361.045 ;
        RECT 3015.270 360.765 3015.550 361.045 ;
        RECT 3015.890 360.765 3016.170 361.045 ;
        RECT 3016.510 360.765 3016.790 361.045 ;
        RECT 3017.130 360.765 3017.410 361.045 ;
        RECT 3017.750 360.765 3018.030 361.045 ;
        RECT 3018.370 360.765 3018.650 361.045 ;
        RECT 3018.990 360.765 3019.270 361.045 ;
        RECT 3019.610 360.765 3019.890 361.045 ;
        RECT 3025.880 369.445 3026.160 369.725 ;
        RECT 3026.500 369.445 3026.780 369.725 ;
        RECT 3027.120 369.445 3027.400 369.725 ;
        RECT 3027.740 369.445 3028.020 369.725 ;
        RECT 3028.360 369.445 3028.640 369.725 ;
        RECT 3028.980 369.445 3029.260 369.725 ;
        RECT 3029.600 369.445 3029.880 369.725 ;
        RECT 3030.220 369.445 3030.500 369.725 ;
        RECT 3030.840 369.445 3031.120 369.725 ;
        RECT 3031.460 369.445 3031.740 369.725 ;
        RECT 3032.080 369.445 3032.360 369.725 ;
        RECT 3032.700 369.445 3032.980 369.725 ;
        RECT 3033.320 369.445 3033.600 369.725 ;
        RECT 3033.940 369.445 3034.220 369.725 ;
        RECT 3034.560 369.445 3034.840 369.725 ;
        RECT 3035.180 369.445 3035.460 369.725 ;
        RECT 3025.880 368.825 3026.160 369.105 ;
        RECT 3026.500 368.825 3026.780 369.105 ;
        RECT 3027.120 368.825 3027.400 369.105 ;
        RECT 3027.740 368.825 3028.020 369.105 ;
        RECT 3028.360 368.825 3028.640 369.105 ;
        RECT 3028.980 368.825 3029.260 369.105 ;
        RECT 3029.600 368.825 3029.880 369.105 ;
        RECT 3030.220 368.825 3030.500 369.105 ;
        RECT 3030.840 368.825 3031.120 369.105 ;
        RECT 3031.460 368.825 3031.740 369.105 ;
        RECT 3032.080 368.825 3032.360 369.105 ;
        RECT 3032.700 368.825 3032.980 369.105 ;
        RECT 3033.320 368.825 3033.600 369.105 ;
        RECT 3033.940 368.825 3034.220 369.105 ;
        RECT 3034.560 368.825 3034.840 369.105 ;
        RECT 3035.180 368.825 3035.460 369.105 ;
        RECT 3025.880 368.205 3026.160 368.485 ;
        RECT 3026.500 368.205 3026.780 368.485 ;
        RECT 3027.120 368.205 3027.400 368.485 ;
        RECT 3027.740 368.205 3028.020 368.485 ;
        RECT 3028.360 368.205 3028.640 368.485 ;
        RECT 3028.980 368.205 3029.260 368.485 ;
        RECT 3029.600 368.205 3029.880 368.485 ;
        RECT 3030.220 368.205 3030.500 368.485 ;
        RECT 3030.840 368.205 3031.120 368.485 ;
        RECT 3031.460 368.205 3031.740 368.485 ;
        RECT 3032.080 368.205 3032.360 368.485 ;
        RECT 3032.700 368.205 3032.980 368.485 ;
        RECT 3033.320 368.205 3033.600 368.485 ;
        RECT 3033.940 368.205 3034.220 368.485 ;
        RECT 3034.560 368.205 3034.840 368.485 ;
        RECT 3035.180 368.205 3035.460 368.485 ;
        RECT 3025.880 367.585 3026.160 367.865 ;
        RECT 3026.500 367.585 3026.780 367.865 ;
        RECT 3027.120 367.585 3027.400 367.865 ;
        RECT 3027.740 367.585 3028.020 367.865 ;
        RECT 3028.360 367.585 3028.640 367.865 ;
        RECT 3028.980 367.585 3029.260 367.865 ;
        RECT 3029.600 367.585 3029.880 367.865 ;
        RECT 3030.220 367.585 3030.500 367.865 ;
        RECT 3030.840 367.585 3031.120 367.865 ;
        RECT 3031.460 367.585 3031.740 367.865 ;
        RECT 3032.080 367.585 3032.360 367.865 ;
        RECT 3032.700 367.585 3032.980 367.865 ;
        RECT 3033.320 367.585 3033.600 367.865 ;
        RECT 3033.940 367.585 3034.220 367.865 ;
        RECT 3034.560 367.585 3034.840 367.865 ;
        RECT 3035.180 367.585 3035.460 367.865 ;
        RECT 3025.880 366.965 3026.160 367.245 ;
        RECT 3026.500 366.965 3026.780 367.245 ;
        RECT 3027.120 366.965 3027.400 367.245 ;
        RECT 3027.740 366.965 3028.020 367.245 ;
        RECT 3028.360 366.965 3028.640 367.245 ;
        RECT 3028.980 366.965 3029.260 367.245 ;
        RECT 3029.600 366.965 3029.880 367.245 ;
        RECT 3030.220 366.965 3030.500 367.245 ;
        RECT 3030.840 366.965 3031.120 367.245 ;
        RECT 3031.460 366.965 3031.740 367.245 ;
        RECT 3032.080 366.965 3032.360 367.245 ;
        RECT 3032.700 366.965 3032.980 367.245 ;
        RECT 3033.320 366.965 3033.600 367.245 ;
        RECT 3033.940 366.965 3034.220 367.245 ;
        RECT 3034.560 366.965 3034.840 367.245 ;
        RECT 3035.180 366.965 3035.460 367.245 ;
        RECT 3025.880 366.345 3026.160 366.625 ;
        RECT 3026.500 366.345 3026.780 366.625 ;
        RECT 3027.120 366.345 3027.400 366.625 ;
        RECT 3027.740 366.345 3028.020 366.625 ;
        RECT 3028.360 366.345 3028.640 366.625 ;
        RECT 3028.980 366.345 3029.260 366.625 ;
        RECT 3029.600 366.345 3029.880 366.625 ;
        RECT 3030.220 366.345 3030.500 366.625 ;
        RECT 3030.840 366.345 3031.120 366.625 ;
        RECT 3031.460 366.345 3031.740 366.625 ;
        RECT 3032.080 366.345 3032.360 366.625 ;
        RECT 3032.700 366.345 3032.980 366.625 ;
        RECT 3033.320 366.345 3033.600 366.625 ;
        RECT 3033.940 366.345 3034.220 366.625 ;
        RECT 3034.560 366.345 3034.840 366.625 ;
        RECT 3035.180 366.345 3035.460 366.625 ;
        RECT 3025.880 365.725 3026.160 366.005 ;
        RECT 3026.500 365.725 3026.780 366.005 ;
        RECT 3027.120 365.725 3027.400 366.005 ;
        RECT 3027.740 365.725 3028.020 366.005 ;
        RECT 3028.360 365.725 3028.640 366.005 ;
        RECT 3028.980 365.725 3029.260 366.005 ;
        RECT 3029.600 365.725 3029.880 366.005 ;
        RECT 3030.220 365.725 3030.500 366.005 ;
        RECT 3030.840 365.725 3031.120 366.005 ;
        RECT 3031.460 365.725 3031.740 366.005 ;
        RECT 3032.080 365.725 3032.360 366.005 ;
        RECT 3032.700 365.725 3032.980 366.005 ;
        RECT 3033.320 365.725 3033.600 366.005 ;
        RECT 3033.940 365.725 3034.220 366.005 ;
        RECT 3034.560 365.725 3034.840 366.005 ;
        RECT 3035.180 365.725 3035.460 366.005 ;
        RECT 3025.880 365.105 3026.160 365.385 ;
        RECT 3026.500 365.105 3026.780 365.385 ;
        RECT 3027.120 365.105 3027.400 365.385 ;
        RECT 3027.740 365.105 3028.020 365.385 ;
        RECT 3028.360 365.105 3028.640 365.385 ;
        RECT 3028.980 365.105 3029.260 365.385 ;
        RECT 3029.600 365.105 3029.880 365.385 ;
        RECT 3030.220 365.105 3030.500 365.385 ;
        RECT 3030.840 365.105 3031.120 365.385 ;
        RECT 3031.460 365.105 3031.740 365.385 ;
        RECT 3032.080 365.105 3032.360 365.385 ;
        RECT 3032.700 365.105 3032.980 365.385 ;
        RECT 3033.320 365.105 3033.600 365.385 ;
        RECT 3033.940 365.105 3034.220 365.385 ;
        RECT 3034.560 365.105 3034.840 365.385 ;
        RECT 3035.180 365.105 3035.460 365.385 ;
        RECT 3025.880 364.485 3026.160 364.765 ;
        RECT 3026.500 364.485 3026.780 364.765 ;
        RECT 3027.120 364.485 3027.400 364.765 ;
        RECT 3027.740 364.485 3028.020 364.765 ;
        RECT 3028.360 364.485 3028.640 364.765 ;
        RECT 3028.980 364.485 3029.260 364.765 ;
        RECT 3029.600 364.485 3029.880 364.765 ;
        RECT 3030.220 364.485 3030.500 364.765 ;
        RECT 3030.840 364.485 3031.120 364.765 ;
        RECT 3031.460 364.485 3031.740 364.765 ;
        RECT 3032.080 364.485 3032.360 364.765 ;
        RECT 3032.700 364.485 3032.980 364.765 ;
        RECT 3033.320 364.485 3033.600 364.765 ;
        RECT 3033.940 364.485 3034.220 364.765 ;
        RECT 3034.560 364.485 3034.840 364.765 ;
        RECT 3035.180 364.485 3035.460 364.765 ;
        RECT 3025.880 363.865 3026.160 364.145 ;
        RECT 3026.500 363.865 3026.780 364.145 ;
        RECT 3027.120 363.865 3027.400 364.145 ;
        RECT 3027.740 363.865 3028.020 364.145 ;
        RECT 3028.360 363.865 3028.640 364.145 ;
        RECT 3028.980 363.865 3029.260 364.145 ;
        RECT 3029.600 363.865 3029.880 364.145 ;
        RECT 3030.220 363.865 3030.500 364.145 ;
        RECT 3030.840 363.865 3031.120 364.145 ;
        RECT 3031.460 363.865 3031.740 364.145 ;
        RECT 3032.080 363.865 3032.360 364.145 ;
        RECT 3032.700 363.865 3032.980 364.145 ;
        RECT 3033.320 363.865 3033.600 364.145 ;
        RECT 3033.940 363.865 3034.220 364.145 ;
        RECT 3034.560 363.865 3034.840 364.145 ;
        RECT 3035.180 363.865 3035.460 364.145 ;
        RECT 3025.880 363.245 3026.160 363.525 ;
        RECT 3026.500 363.245 3026.780 363.525 ;
        RECT 3027.120 363.245 3027.400 363.525 ;
        RECT 3027.740 363.245 3028.020 363.525 ;
        RECT 3028.360 363.245 3028.640 363.525 ;
        RECT 3028.980 363.245 3029.260 363.525 ;
        RECT 3029.600 363.245 3029.880 363.525 ;
        RECT 3030.220 363.245 3030.500 363.525 ;
        RECT 3030.840 363.245 3031.120 363.525 ;
        RECT 3031.460 363.245 3031.740 363.525 ;
        RECT 3032.080 363.245 3032.360 363.525 ;
        RECT 3032.700 363.245 3032.980 363.525 ;
        RECT 3033.320 363.245 3033.600 363.525 ;
        RECT 3033.940 363.245 3034.220 363.525 ;
        RECT 3034.560 363.245 3034.840 363.525 ;
        RECT 3035.180 363.245 3035.460 363.525 ;
        RECT 3025.880 362.625 3026.160 362.905 ;
        RECT 3026.500 362.625 3026.780 362.905 ;
        RECT 3027.120 362.625 3027.400 362.905 ;
        RECT 3027.740 362.625 3028.020 362.905 ;
        RECT 3028.360 362.625 3028.640 362.905 ;
        RECT 3028.980 362.625 3029.260 362.905 ;
        RECT 3029.600 362.625 3029.880 362.905 ;
        RECT 3030.220 362.625 3030.500 362.905 ;
        RECT 3030.840 362.625 3031.120 362.905 ;
        RECT 3031.460 362.625 3031.740 362.905 ;
        RECT 3032.080 362.625 3032.360 362.905 ;
        RECT 3032.700 362.625 3032.980 362.905 ;
        RECT 3033.320 362.625 3033.600 362.905 ;
        RECT 3033.940 362.625 3034.220 362.905 ;
        RECT 3034.560 362.625 3034.840 362.905 ;
        RECT 3035.180 362.625 3035.460 362.905 ;
        RECT 3025.880 362.005 3026.160 362.285 ;
        RECT 3026.500 362.005 3026.780 362.285 ;
        RECT 3027.120 362.005 3027.400 362.285 ;
        RECT 3027.740 362.005 3028.020 362.285 ;
        RECT 3028.360 362.005 3028.640 362.285 ;
        RECT 3028.980 362.005 3029.260 362.285 ;
        RECT 3029.600 362.005 3029.880 362.285 ;
        RECT 3030.220 362.005 3030.500 362.285 ;
        RECT 3030.840 362.005 3031.120 362.285 ;
        RECT 3031.460 362.005 3031.740 362.285 ;
        RECT 3032.080 362.005 3032.360 362.285 ;
        RECT 3032.700 362.005 3032.980 362.285 ;
        RECT 3033.320 362.005 3033.600 362.285 ;
        RECT 3033.940 362.005 3034.220 362.285 ;
        RECT 3034.560 362.005 3034.840 362.285 ;
        RECT 3035.180 362.005 3035.460 362.285 ;
        RECT 3025.880 361.385 3026.160 361.665 ;
        RECT 3026.500 361.385 3026.780 361.665 ;
        RECT 3027.120 361.385 3027.400 361.665 ;
        RECT 3027.740 361.385 3028.020 361.665 ;
        RECT 3028.360 361.385 3028.640 361.665 ;
        RECT 3028.980 361.385 3029.260 361.665 ;
        RECT 3029.600 361.385 3029.880 361.665 ;
        RECT 3030.220 361.385 3030.500 361.665 ;
        RECT 3030.840 361.385 3031.120 361.665 ;
        RECT 3031.460 361.385 3031.740 361.665 ;
        RECT 3032.080 361.385 3032.360 361.665 ;
        RECT 3032.700 361.385 3032.980 361.665 ;
        RECT 3033.320 361.385 3033.600 361.665 ;
        RECT 3033.940 361.385 3034.220 361.665 ;
        RECT 3034.560 361.385 3034.840 361.665 ;
        RECT 3035.180 361.385 3035.460 361.665 ;
        RECT 3025.880 360.765 3026.160 361.045 ;
        RECT 3026.500 360.765 3026.780 361.045 ;
        RECT 3027.120 360.765 3027.400 361.045 ;
        RECT 3027.740 360.765 3028.020 361.045 ;
        RECT 3028.360 360.765 3028.640 361.045 ;
        RECT 3028.980 360.765 3029.260 361.045 ;
        RECT 3029.600 360.765 3029.880 361.045 ;
        RECT 3030.220 360.765 3030.500 361.045 ;
        RECT 3030.840 360.765 3031.120 361.045 ;
        RECT 3031.460 360.765 3031.740 361.045 ;
        RECT 3032.080 360.765 3032.360 361.045 ;
        RECT 3032.700 360.765 3032.980 361.045 ;
        RECT 3033.320 360.765 3033.600 361.045 ;
        RECT 3033.940 360.765 3034.220 361.045 ;
        RECT 3034.560 360.765 3034.840 361.045 ;
        RECT 3035.180 360.765 3035.460 361.045 ;
        RECT 3039.410 369.445 3039.690 369.725 ;
        RECT 3040.030 369.445 3040.310 369.725 ;
        RECT 3040.650 369.445 3040.930 369.725 ;
        RECT 3041.270 369.445 3041.550 369.725 ;
        RECT 3041.890 369.445 3042.170 369.725 ;
        RECT 3042.510 369.445 3042.790 369.725 ;
        RECT 3043.130 369.445 3043.410 369.725 ;
        RECT 3043.750 369.445 3044.030 369.725 ;
        RECT 3044.370 369.445 3044.650 369.725 ;
        RECT 3044.990 369.445 3045.270 369.725 ;
        RECT 3045.610 369.445 3045.890 369.725 ;
        RECT 3046.230 369.445 3046.510 369.725 ;
        RECT 3046.850 369.445 3047.130 369.725 ;
        RECT 3047.470 369.445 3047.750 369.725 ;
        RECT 3048.090 369.445 3048.370 369.725 ;
        RECT 3048.710 369.445 3048.990 369.725 ;
        RECT 3039.410 368.825 3039.690 369.105 ;
        RECT 3040.030 368.825 3040.310 369.105 ;
        RECT 3040.650 368.825 3040.930 369.105 ;
        RECT 3041.270 368.825 3041.550 369.105 ;
        RECT 3041.890 368.825 3042.170 369.105 ;
        RECT 3042.510 368.825 3042.790 369.105 ;
        RECT 3043.130 368.825 3043.410 369.105 ;
        RECT 3043.750 368.825 3044.030 369.105 ;
        RECT 3044.370 368.825 3044.650 369.105 ;
        RECT 3044.990 368.825 3045.270 369.105 ;
        RECT 3045.610 368.825 3045.890 369.105 ;
        RECT 3046.230 368.825 3046.510 369.105 ;
        RECT 3046.850 368.825 3047.130 369.105 ;
        RECT 3047.470 368.825 3047.750 369.105 ;
        RECT 3048.090 368.825 3048.370 369.105 ;
        RECT 3048.710 368.825 3048.990 369.105 ;
        RECT 3039.410 368.205 3039.690 368.485 ;
        RECT 3040.030 368.205 3040.310 368.485 ;
        RECT 3040.650 368.205 3040.930 368.485 ;
        RECT 3041.270 368.205 3041.550 368.485 ;
        RECT 3041.890 368.205 3042.170 368.485 ;
        RECT 3042.510 368.205 3042.790 368.485 ;
        RECT 3043.130 368.205 3043.410 368.485 ;
        RECT 3043.750 368.205 3044.030 368.485 ;
        RECT 3044.370 368.205 3044.650 368.485 ;
        RECT 3044.990 368.205 3045.270 368.485 ;
        RECT 3045.610 368.205 3045.890 368.485 ;
        RECT 3046.230 368.205 3046.510 368.485 ;
        RECT 3046.850 368.205 3047.130 368.485 ;
        RECT 3047.470 368.205 3047.750 368.485 ;
        RECT 3048.090 368.205 3048.370 368.485 ;
        RECT 3048.710 368.205 3048.990 368.485 ;
        RECT 3039.410 367.585 3039.690 367.865 ;
        RECT 3040.030 367.585 3040.310 367.865 ;
        RECT 3040.650 367.585 3040.930 367.865 ;
        RECT 3041.270 367.585 3041.550 367.865 ;
        RECT 3041.890 367.585 3042.170 367.865 ;
        RECT 3042.510 367.585 3042.790 367.865 ;
        RECT 3043.130 367.585 3043.410 367.865 ;
        RECT 3043.750 367.585 3044.030 367.865 ;
        RECT 3044.370 367.585 3044.650 367.865 ;
        RECT 3044.990 367.585 3045.270 367.865 ;
        RECT 3045.610 367.585 3045.890 367.865 ;
        RECT 3046.230 367.585 3046.510 367.865 ;
        RECT 3046.850 367.585 3047.130 367.865 ;
        RECT 3047.470 367.585 3047.750 367.865 ;
        RECT 3048.090 367.585 3048.370 367.865 ;
        RECT 3048.710 367.585 3048.990 367.865 ;
        RECT 3039.410 366.965 3039.690 367.245 ;
        RECT 3040.030 366.965 3040.310 367.245 ;
        RECT 3040.650 366.965 3040.930 367.245 ;
        RECT 3041.270 366.965 3041.550 367.245 ;
        RECT 3041.890 366.965 3042.170 367.245 ;
        RECT 3042.510 366.965 3042.790 367.245 ;
        RECT 3043.130 366.965 3043.410 367.245 ;
        RECT 3043.750 366.965 3044.030 367.245 ;
        RECT 3044.370 366.965 3044.650 367.245 ;
        RECT 3044.990 366.965 3045.270 367.245 ;
        RECT 3045.610 366.965 3045.890 367.245 ;
        RECT 3046.230 366.965 3046.510 367.245 ;
        RECT 3046.850 366.965 3047.130 367.245 ;
        RECT 3047.470 366.965 3047.750 367.245 ;
        RECT 3048.090 366.965 3048.370 367.245 ;
        RECT 3048.710 366.965 3048.990 367.245 ;
        RECT 3039.410 366.345 3039.690 366.625 ;
        RECT 3040.030 366.345 3040.310 366.625 ;
        RECT 3040.650 366.345 3040.930 366.625 ;
        RECT 3041.270 366.345 3041.550 366.625 ;
        RECT 3041.890 366.345 3042.170 366.625 ;
        RECT 3042.510 366.345 3042.790 366.625 ;
        RECT 3043.130 366.345 3043.410 366.625 ;
        RECT 3043.750 366.345 3044.030 366.625 ;
        RECT 3044.370 366.345 3044.650 366.625 ;
        RECT 3044.990 366.345 3045.270 366.625 ;
        RECT 3045.610 366.345 3045.890 366.625 ;
        RECT 3046.230 366.345 3046.510 366.625 ;
        RECT 3046.850 366.345 3047.130 366.625 ;
        RECT 3047.470 366.345 3047.750 366.625 ;
        RECT 3048.090 366.345 3048.370 366.625 ;
        RECT 3048.710 366.345 3048.990 366.625 ;
        RECT 3039.410 365.725 3039.690 366.005 ;
        RECT 3040.030 365.725 3040.310 366.005 ;
        RECT 3040.650 365.725 3040.930 366.005 ;
        RECT 3041.270 365.725 3041.550 366.005 ;
        RECT 3041.890 365.725 3042.170 366.005 ;
        RECT 3042.510 365.725 3042.790 366.005 ;
        RECT 3043.130 365.725 3043.410 366.005 ;
        RECT 3043.750 365.725 3044.030 366.005 ;
        RECT 3044.370 365.725 3044.650 366.005 ;
        RECT 3044.990 365.725 3045.270 366.005 ;
        RECT 3045.610 365.725 3045.890 366.005 ;
        RECT 3046.230 365.725 3046.510 366.005 ;
        RECT 3046.850 365.725 3047.130 366.005 ;
        RECT 3047.470 365.725 3047.750 366.005 ;
        RECT 3048.090 365.725 3048.370 366.005 ;
        RECT 3048.710 365.725 3048.990 366.005 ;
        RECT 3039.410 365.105 3039.690 365.385 ;
        RECT 3040.030 365.105 3040.310 365.385 ;
        RECT 3040.650 365.105 3040.930 365.385 ;
        RECT 3041.270 365.105 3041.550 365.385 ;
        RECT 3041.890 365.105 3042.170 365.385 ;
        RECT 3042.510 365.105 3042.790 365.385 ;
        RECT 3043.130 365.105 3043.410 365.385 ;
        RECT 3043.750 365.105 3044.030 365.385 ;
        RECT 3044.370 365.105 3044.650 365.385 ;
        RECT 3044.990 365.105 3045.270 365.385 ;
        RECT 3045.610 365.105 3045.890 365.385 ;
        RECT 3046.230 365.105 3046.510 365.385 ;
        RECT 3046.850 365.105 3047.130 365.385 ;
        RECT 3047.470 365.105 3047.750 365.385 ;
        RECT 3048.090 365.105 3048.370 365.385 ;
        RECT 3048.710 365.105 3048.990 365.385 ;
        RECT 3039.410 364.485 3039.690 364.765 ;
        RECT 3040.030 364.485 3040.310 364.765 ;
        RECT 3040.650 364.485 3040.930 364.765 ;
        RECT 3041.270 364.485 3041.550 364.765 ;
        RECT 3041.890 364.485 3042.170 364.765 ;
        RECT 3042.510 364.485 3042.790 364.765 ;
        RECT 3043.130 364.485 3043.410 364.765 ;
        RECT 3043.750 364.485 3044.030 364.765 ;
        RECT 3044.370 364.485 3044.650 364.765 ;
        RECT 3044.990 364.485 3045.270 364.765 ;
        RECT 3045.610 364.485 3045.890 364.765 ;
        RECT 3046.230 364.485 3046.510 364.765 ;
        RECT 3046.850 364.485 3047.130 364.765 ;
        RECT 3047.470 364.485 3047.750 364.765 ;
        RECT 3048.090 364.485 3048.370 364.765 ;
        RECT 3048.710 364.485 3048.990 364.765 ;
        RECT 3039.410 363.865 3039.690 364.145 ;
        RECT 3040.030 363.865 3040.310 364.145 ;
        RECT 3040.650 363.865 3040.930 364.145 ;
        RECT 3041.270 363.865 3041.550 364.145 ;
        RECT 3041.890 363.865 3042.170 364.145 ;
        RECT 3042.510 363.865 3042.790 364.145 ;
        RECT 3043.130 363.865 3043.410 364.145 ;
        RECT 3043.750 363.865 3044.030 364.145 ;
        RECT 3044.370 363.865 3044.650 364.145 ;
        RECT 3044.990 363.865 3045.270 364.145 ;
        RECT 3045.610 363.865 3045.890 364.145 ;
        RECT 3046.230 363.865 3046.510 364.145 ;
        RECT 3046.850 363.865 3047.130 364.145 ;
        RECT 3047.470 363.865 3047.750 364.145 ;
        RECT 3048.090 363.865 3048.370 364.145 ;
        RECT 3048.710 363.865 3048.990 364.145 ;
        RECT 3039.410 363.245 3039.690 363.525 ;
        RECT 3040.030 363.245 3040.310 363.525 ;
        RECT 3040.650 363.245 3040.930 363.525 ;
        RECT 3041.270 363.245 3041.550 363.525 ;
        RECT 3041.890 363.245 3042.170 363.525 ;
        RECT 3042.510 363.245 3042.790 363.525 ;
        RECT 3043.130 363.245 3043.410 363.525 ;
        RECT 3043.750 363.245 3044.030 363.525 ;
        RECT 3044.370 363.245 3044.650 363.525 ;
        RECT 3044.990 363.245 3045.270 363.525 ;
        RECT 3045.610 363.245 3045.890 363.525 ;
        RECT 3046.230 363.245 3046.510 363.525 ;
        RECT 3046.850 363.245 3047.130 363.525 ;
        RECT 3047.470 363.245 3047.750 363.525 ;
        RECT 3048.090 363.245 3048.370 363.525 ;
        RECT 3048.710 363.245 3048.990 363.525 ;
        RECT 3039.410 362.625 3039.690 362.905 ;
        RECT 3040.030 362.625 3040.310 362.905 ;
        RECT 3040.650 362.625 3040.930 362.905 ;
        RECT 3041.270 362.625 3041.550 362.905 ;
        RECT 3041.890 362.625 3042.170 362.905 ;
        RECT 3042.510 362.625 3042.790 362.905 ;
        RECT 3043.130 362.625 3043.410 362.905 ;
        RECT 3043.750 362.625 3044.030 362.905 ;
        RECT 3044.370 362.625 3044.650 362.905 ;
        RECT 3044.990 362.625 3045.270 362.905 ;
        RECT 3045.610 362.625 3045.890 362.905 ;
        RECT 3046.230 362.625 3046.510 362.905 ;
        RECT 3046.850 362.625 3047.130 362.905 ;
        RECT 3047.470 362.625 3047.750 362.905 ;
        RECT 3048.090 362.625 3048.370 362.905 ;
        RECT 3048.710 362.625 3048.990 362.905 ;
        RECT 3039.410 362.005 3039.690 362.285 ;
        RECT 3040.030 362.005 3040.310 362.285 ;
        RECT 3040.650 362.005 3040.930 362.285 ;
        RECT 3041.270 362.005 3041.550 362.285 ;
        RECT 3041.890 362.005 3042.170 362.285 ;
        RECT 3042.510 362.005 3042.790 362.285 ;
        RECT 3043.130 362.005 3043.410 362.285 ;
        RECT 3043.750 362.005 3044.030 362.285 ;
        RECT 3044.370 362.005 3044.650 362.285 ;
        RECT 3044.990 362.005 3045.270 362.285 ;
        RECT 3045.610 362.005 3045.890 362.285 ;
        RECT 3046.230 362.005 3046.510 362.285 ;
        RECT 3046.850 362.005 3047.130 362.285 ;
        RECT 3047.470 362.005 3047.750 362.285 ;
        RECT 3048.090 362.005 3048.370 362.285 ;
        RECT 3048.710 362.005 3048.990 362.285 ;
        RECT 3039.410 361.385 3039.690 361.665 ;
        RECT 3040.030 361.385 3040.310 361.665 ;
        RECT 3040.650 361.385 3040.930 361.665 ;
        RECT 3041.270 361.385 3041.550 361.665 ;
        RECT 3041.890 361.385 3042.170 361.665 ;
        RECT 3042.510 361.385 3042.790 361.665 ;
        RECT 3043.130 361.385 3043.410 361.665 ;
        RECT 3043.750 361.385 3044.030 361.665 ;
        RECT 3044.370 361.385 3044.650 361.665 ;
        RECT 3044.990 361.385 3045.270 361.665 ;
        RECT 3045.610 361.385 3045.890 361.665 ;
        RECT 3046.230 361.385 3046.510 361.665 ;
        RECT 3046.850 361.385 3047.130 361.665 ;
        RECT 3047.470 361.385 3047.750 361.665 ;
        RECT 3048.090 361.385 3048.370 361.665 ;
        RECT 3048.710 361.385 3048.990 361.665 ;
        RECT 3039.410 360.765 3039.690 361.045 ;
        RECT 3040.030 360.765 3040.310 361.045 ;
        RECT 3040.650 360.765 3040.930 361.045 ;
        RECT 3041.270 360.765 3041.550 361.045 ;
        RECT 3041.890 360.765 3042.170 361.045 ;
        RECT 3042.510 360.765 3042.790 361.045 ;
        RECT 3043.130 360.765 3043.410 361.045 ;
        RECT 3043.750 360.765 3044.030 361.045 ;
        RECT 3044.370 360.765 3044.650 361.045 ;
        RECT 3044.990 360.765 3045.270 361.045 ;
        RECT 3045.610 360.765 3045.890 361.045 ;
        RECT 3046.230 360.765 3046.510 361.045 ;
        RECT 3046.850 360.765 3047.130 361.045 ;
        RECT 3047.470 360.765 3047.750 361.045 ;
        RECT 3048.090 360.765 3048.370 361.045 ;
        RECT 3048.710 360.765 3048.990 361.045 ;
        RECT 3051.260 369.445 3051.540 369.725 ;
        RECT 3051.880 369.445 3052.160 369.725 ;
        RECT 3052.500 369.445 3052.780 369.725 ;
        RECT 3053.120 369.445 3053.400 369.725 ;
        RECT 3053.740 369.445 3054.020 369.725 ;
        RECT 3054.360 369.445 3054.640 369.725 ;
        RECT 3054.980 369.445 3055.260 369.725 ;
        RECT 3055.600 369.445 3055.880 369.725 ;
        RECT 3056.220 369.445 3056.500 369.725 ;
        RECT 3056.840 369.445 3057.120 369.725 ;
        RECT 3057.460 369.445 3057.740 369.725 ;
        RECT 3058.080 369.445 3058.360 369.725 ;
        RECT 3058.700 369.445 3058.980 369.725 ;
        RECT 3059.320 369.445 3059.600 369.725 ;
        RECT 3059.940 369.445 3060.220 369.725 ;
        RECT 3060.560 369.445 3060.840 369.725 ;
        RECT 3051.260 368.825 3051.540 369.105 ;
        RECT 3051.880 368.825 3052.160 369.105 ;
        RECT 3052.500 368.825 3052.780 369.105 ;
        RECT 3053.120 368.825 3053.400 369.105 ;
        RECT 3053.740 368.825 3054.020 369.105 ;
        RECT 3054.360 368.825 3054.640 369.105 ;
        RECT 3054.980 368.825 3055.260 369.105 ;
        RECT 3055.600 368.825 3055.880 369.105 ;
        RECT 3056.220 368.825 3056.500 369.105 ;
        RECT 3056.840 368.825 3057.120 369.105 ;
        RECT 3057.460 368.825 3057.740 369.105 ;
        RECT 3058.080 368.825 3058.360 369.105 ;
        RECT 3058.700 368.825 3058.980 369.105 ;
        RECT 3059.320 368.825 3059.600 369.105 ;
        RECT 3059.940 368.825 3060.220 369.105 ;
        RECT 3060.560 368.825 3060.840 369.105 ;
        RECT 3051.260 368.205 3051.540 368.485 ;
        RECT 3051.880 368.205 3052.160 368.485 ;
        RECT 3052.500 368.205 3052.780 368.485 ;
        RECT 3053.120 368.205 3053.400 368.485 ;
        RECT 3053.740 368.205 3054.020 368.485 ;
        RECT 3054.360 368.205 3054.640 368.485 ;
        RECT 3054.980 368.205 3055.260 368.485 ;
        RECT 3055.600 368.205 3055.880 368.485 ;
        RECT 3056.220 368.205 3056.500 368.485 ;
        RECT 3056.840 368.205 3057.120 368.485 ;
        RECT 3057.460 368.205 3057.740 368.485 ;
        RECT 3058.080 368.205 3058.360 368.485 ;
        RECT 3058.700 368.205 3058.980 368.485 ;
        RECT 3059.320 368.205 3059.600 368.485 ;
        RECT 3059.940 368.205 3060.220 368.485 ;
        RECT 3060.560 368.205 3060.840 368.485 ;
        RECT 3051.260 367.585 3051.540 367.865 ;
        RECT 3051.880 367.585 3052.160 367.865 ;
        RECT 3052.500 367.585 3052.780 367.865 ;
        RECT 3053.120 367.585 3053.400 367.865 ;
        RECT 3053.740 367.585 3054.020 367.865 ;
        RECT 3054.360 367.585 3054.640 367.865 ;
        RECT 3054.980 367.585 3055.260 367.865 ;
        RECT 3055.600 367.585 3055.880 367.865 ;
        RECT 3056.220 367.585 3056.500 367.865 ;
        RECT 3056.840 367.585 3057.120 367.865 ;
        RECT 3057.460 367.585 3057.740 367.865 ;
        RECT 3058.080 367.585 3058.360 367.865 ;
        RECT 3058.700 367.585 3058.980 367.865 ;
        RECT 3059.320 367.585 3059.600 367.865 ;
        RECT 3059.940 367.585 3060.220 367.865 ;
        RECT 3060.560 367.585 3060.840 367.865 ;
        RECT 3051.260 366.965 3051.540 367.245 ;
        RECT 3051.880 366.965 3052.160 367.245 ;
        RECT 3052.500 366.965 3052.780 367.245 ;
        RECT 3053.120 366.965 3053.400 367.245 ;
        RECT 3053.740 366.965 3054.020 367.245 ;
        RECT 3054.360 366.965 3054.640 367.245 ;
        RECT 3054.980 366.965 3055.260 367.245 ;
        RECT 3055.600 366.965 3055.880 367.245 ;
        RECT 3056.220 366.965 3056.500 367.245 ;
        RECT 3056.840 366.965 3057.120 367.245 ;
        RECT 3057.460 366.965 3057.740 367.245 ;
        RECT 3058.080 366.965 3058.360 367.245 ;
        RECT 3058.700 366.965 3058.980 367.245 ;
        RECT 3059.320 366.965 3059.600 367.245 ;
        RECT 3059.940 366.965 3060.220 367.245 ;
        RECT 3060.560 366.965 3060.840 367.245 ;
        RECT 3051.260 366.345 3051.540 366.625 ;
        RECT 3051.880 366.345 3052.160 366.625 ;
        RECT 3052.500 366.345 3052.780 366.625 ;
        RECT 3053.120 366.345 3053.400 366.625 ;
        RECT 3053.740 366.345 3054.020 366.625 ;
        RECT 3054.360 366.345 3054.640 366.625 ;
        RECT 3054.980 366.345 3055.260 366.625 ;
        RECT 3055.600 366.345 3055.880 366.625 ;
        RECT 3056.220 366.345 3056.500 366.625 ;
        RECT 3056.840 366.345 3057.120 366.625 ;
        RECT 3057.460 366.345 3057.740 366.625 ;
        RECT 3058.080 366.345 3058.360 366.625 ;
        RECT 3058.700 366.345 3058.980 366.625 ;
        RECT 3059.320 366.345 3059.600 366.625 ;
        RECT 3059.940 366.345 3060.220 366.625 ;
        RECT 3060.560 366.345 3060.840 366.625 ;
        RECT 3051.260 365.725 3051.540 366.005 ;
        RECT 3051.880 365.725 3052.160 366.005 ;
        RECT 3052.500 365.725 3052.780 366.005 ;
        RECT 3053.120 365.725 3053.400 366.005 ;
        RECT 3053.740 365.725 3054.020 366.005 ;
        RECT 3054.360 365.725 3054.640 366.005 ;
        RECT 3054.980 365.725 3055.260 366.005 ;
        RECT 3055.600 365.725 3055.880 366.005 ;
        RECT 3056.220 365.725 3056.500 366.005 ;
        RECT 3056.840 365.725 3057.120 366.005 ;
        RECT 3057.460 365.725 3057.740 366.005 ;
        RECT 3058.080 365.725 3058.360 366.005 ;
        RECT 3058.700 365.725 3058.980 366.005 ;
        RECT 3059.320 365.725 3059.600 366.005 ;
        RECT 3059.940 365.725 3060.220 366.005 ;
        RECT 3060.560 365.725 3060.840 366.005 ;
        RECT 3051.260 365.105 3051.540 365.385 ;
        RECT 3051.880 365.105 3052.160 365.385 ;
        RECT 3052.500 365.105 3052.780 365.385 ;
        RECT 3053.120 365.105 3053.400 365.385 ;
        RECT 3053.740 365.105 3054.020 365.385 ;
        RECT 3054.360 365.105 3054.640 365.385 ;
        RECT 3054.980 365.105 3055.260 365.385 ;
        RECT 3055.600 365.105 3055.880 365.385 ;
        RECT 3056.220 365.105 3056.500 365.385 ;
        RECT 3056.840 365.105 3057.120 365.385 ;
        RECT 3057.460 365.105 3057.740 365.385 ;
        RECT 3058.080 365.105 3058.360 365.385 ;
        RECT 3058.700 365.105 3058.980 365.385 ;
        RECT 3059.320 365.105 3059.600 365.385 ;
        RECT 3059.940 365.105 3060.220 365.385 ;
        RECT 3060.560 365.105 3060.840 365.385 ;
        RECT 3051.260 364.485 3051.540 364.765 ;
        RECT 3051.880 364.485 3052.160 364.765 ;
        RECT 3052.500 364.485 3052.780 364.765 ;
        RECT 3053.120 364.485 3053.400 364.765 ;
        RECT 3053.740 364.485 3054.020 364.765 ;
        RECT 3054.360 364.485 3054.640 364.765 ;
        RECT 3054.980 364.485 3055.260 364.765 ;
        RECT 3055.600 364.485 3055.880 364.765 ;
        RECT 3056.220 364.485 3056.500 364.765 ;
        RECT 3056.840 364.485 3057.120 364.765 ;
        RECT 3057.460 364.485 3057.740 364.765 ;
        RECT 3058.080 364.485 3058.360 364.765 ;
        RECT 3058.700 364.485 3058.980 364.765 ;
        RECT 3059.320 364.485 3059.600 364.765 ;
        RECT 3059.940 364.485 3060.220 364.765 ;
        RECT 3060.560 364.485 3060.840 364.765 ;
        RECT 3051.260 363.865 3051.540 364.145 ;
        RECT 3051.880 363.865 3052.160 364.145 ;
        RECT 3052.500 363.865 3052.780 364.145 ;
        RECT 3053.120 363.865 3053.400 364.145 ;
        RECT 3053.740 363.865 3054.020 364.145 ;
        RECT 3054.360 363.865 3054.640 364.145 ;
        RECT 3054.980 363.865 3055.260 364.145 ;
        RECT 3055.600 363.865 3055.880 364.145 ;
        RECT 3056.220 363.865 3056.500 364.145 ;
        RECT 3056.840 363.865 3057.120 364.145 ;
        RECT 3057.460 363.865 3057.740 364.145 ;
        RECT 3058.080 363.865 3058.360 364.145 ;
        RECT 3058.700 363.865 3058.980 364.145 ;
        RECT 3059.320 363.865 3059.600 364.145 ;
        RECT 3059.940 363.865 3060.220 364.145 ;
        RECT 3060.560 363.865 3060.840 364.145 ;
        RECT 3051.260 363.245 3051.540 363.525 ;
        RECT 3051.880 363.245 3052.160 363.525 ;
        RECT 3052.500 363.245 3052.780 363.525 ;
        RECT 3053.120 363.245 3053.400 363.525 ;
        RECT 3053.740 363.245 3054.020 363.525 ;
        RECT 3054.360 363.245 3054.640 363.525 ;
        RECT 3054.980 363.245 3055.260 363.525 ;
        RECT 3055.600 363.245 3055.880 363.525 ;
        RECT 3056.220 363.245 3056.500 363.525 ;
        RECT 3056.840 363.245 3057.120 363.525 ;
        RECT 3057.460 363.245 3057.740 363.525 ;
        RECT 3058.080 363.245 3058.360 363.525 ;
        RECT 3058.700 363.245 3058.980 363.525 ;
        RECT 3059.320 363.245 3059.600 363.525 ;
        RECT 3059.940 363.245 3060.220 363.525 ;
        RECT 3060.560 363.245 3060.840 363.525 ;
        RECT 3051.260 362.625 3051.540 362.905 ;
        RECT 3051.880 362.625 3052.160 362.905 ;
        RECT 3052.500 362.625 3052.780 362.905 ;
        RECT 3053.120 362.625 3053.400 362.905 ;
        RECT 3053.740 362.625 3054.020 362.905 ;
        RECT 3054.360 362.625 3054.640 362.905 ;
        RECT 3054.980 362.625 3055.260 362.905 ;
        RECT 3055.600 362.625 3055.880 362.905 ;
        RECT 3056.220 362.625 3056.500 362.905 ;
        RECT 3056.840 362.625 3057.120 362.905 ;
        RECT 3057.460 362.625 3057.740 362.905 ;
        RECT 3058.080 362.625 3058.360 362.905 ;
        RECT 3058.700 362.625 3058.980 362.905 ;
        RECT 3059.320 362.625 3059.600 362.905 ;
        RECT 3059.940 362.625 3060.220 362.905 ;
        RECT 3060.560 362.625 3060.840 362.905 ;
        RECT 3051.260 362.005 3051.540 362.285 ;
        RECT 3051.880 362.005 3052.160 362.285 ;
        RECT 3052.500 362.005 3052.780 362.285 ;
        RECT 3053.120 362.005 3053.400 362.285 ;
        RECT 3053.740 362.005 3054.020 362.285 ;
        RECT 3054.360 362.005 3054.640 362.285 ;
        RECT 3054.980 362.005 3055.260 362.285 ;
        RECT 3055.600 362.005 3055.880 362.285 ;
        RECT 3056.220 362.005 3056.500 362.285 ;
        RECT 3056.840 362.005 3057.120 362.285 ;
        RECT 3057.460 362.005 3057.740 362.285 ;
        RECT 3058.080 362.005 3058.360 362.285 ;
        RECT 3058.700 362.005 3058.980 362.285 ;
        RECT 3059.320 362.005 3059.600 362.285 ;
        RECT 3059.940 362.005 3060.220 362.285 ;
        RECT 3060.560 362.005 3060.840 362.285 ;
        RECT 3051.260 361.385 3051.540 361.665 ;
        RECT 3051.880 361.385 3052.160 361.665 ;
        RECT 3052.500 361.385 3052.780 361.665 ;
        RECT 3053.120 361.385 3053.400 361.665 ;
        RECT 3053.740 361.385 3054.020 361.665 ;
        RECT 3054.360 361.385 3054.640 361.665 ;
        RECT 3054.980 361.385 3055.260 361.665 ;
        RECT 3055.600 361.385 3055.880 361.665 ;
        RECT 3056.220 361.385 3056.500 361.665 ;
        RECT 3056.840 361.385 3057.120 361.665 ;
        RECT 3057.460 361.385 3057.740 361.665 ;
        RECT 3058.080 361.385 3058.360 361.665 ;
        RECT 3058.700 361.385 3058.980 361.665 ;
        RECT 3059.320 361.385 3059.600 361.665 ;
        RECT 3059.940 361.385 3060.220 361.665 ;
        RECT 3060.560 361.385 3060.840 361.665 ;
        RECT 3051.260 360.765 3051.540 361.045 ;
        RECT 3051.880 360.765 3052.160 361.045 ;
        RECT 3052.500 360.765 3052.780 361.045 ;
        RECT 3053.120 360.765 3053.400 361.045 ;
        RECT 3053.740 360.765 3054.020 361.045 ;
        RECT 3054.360 360.765 3054.640 361.045 ;
        RECT 3054.980 360.765 3055.260 361.045 ;
        RECT 3055.600 360.765 3055.880 361.045 ;
        RECT 3056.220 360.765 3056.500 361.045 ;
        RECT 3056.840 360.765 3057.120 361.045 ;
        RECT 3057.460 360.765 3057.740 361.045 ;
        RECT 3058.080 360.765 3058.360 361.045 ;
        RECT 3058.700 360.765 3058.980 361.045 ;
        RECT 3059.320 360.765 3059.600 361.045 ;
        RECT 3059.940 360.765 3060.220 361.045 ;
        RECT 3060.560 360.765 3060.840 361.045 ;
        RECT 3064.410 369.445 3064.690 369.725 ;
        RECT 3065.030 369.445 3065.310 369.725 ;
        RECT 3065.650 369.445 3065.930 369.725 ;
        RECT 3066.270 369.445 3066.550 369.725 ;
        RECT 3066.890 369.445 3067.170 369.725 ;
        RECT 3067.510 369.445 3067.790 369.725 ;
        RECT 3068.130 369.445 3068.410 369.725 ;
        RECT 3068.750 369.445 3069.030 369.725 ;
        RECT 3069.370 369.445 3069.650 369.725 ;
        RECT 3069.990 369.445 3070.270 369.725 ;
        RECT 3070.610 369.445 3070.890 369.725 ;
        RECT 3071.230 369.445 3071.510 369.725 ;
        RECT 3071.850 369.445 3072.130 369.725 ;
        RECT 3072.470 369.445 3072.750 369.725 ;
        RECT 3073.090 369.445 3073.370 369.725 ;
        RECT 3064.410 368.825 3064.690 369.105 ;
        RECT 3065.030 368.825 3065.310 369.105 ;
        RECT 3065.650 368.825 3065.930 369.105 ;
        RECT 3066.270 368.825 3066.550 369.105 ;
        RECT 3066.890 368.825 3067.170 369.105 ;
        RECT 3067.510 368.825 3067.790 369.105 ;
        RECT 3068.130 368.825 3068.410 369.105 ;
        RECT 3068.750 368.825 3069.030 369.105 ;
        RECT 3069.370 368.825 3069.650 369.105 ;
        RECT 3069.990 368.825 3070.270 369.105 ;
        RECT 3070.610 368.825 3070.890 369.105 ;
        RECT 3071.230 368.825 3071.510 369.105 ;
        RECT 3071.850 368.825 3072.130 369.105 ;
        RECT 3072.470 368.825 3072.750 369.105 ;
        RECT 3073.090 368.825 3073.370 369.105 ;
        RECT 3064.410 368.205 3064.690 368.485 ;
        RECT 3065.030 368.205 3065.310 368.485 ;
        RECT 3065.650 368.205 3065.930 368.485 ;
        RECT 3066.270 368.205 3066.550 368.485 ;
        RECT 3066.890 368.205 3067.170 368.485 ;
        RECT 3067.510 368.205 3067.790 368.485 ;
        RECT 3068.130 368.205 3068.410 368.485 ;
        RECT 3068.750 368.205 3069.030 368.485 ;
        RECT 3069.370 368.205 3069.650 368.485 ;
        RECT 3069.990 368.205 3070.270 368.485 ;
        RECT 3070.610 368.205 3070.890 368.485 ;
        RECT 3071.230 368.205 3071.510 368.485 ;
        RECT 3071.850 368.205 3072.130 368.485 ;
        RECT 3072.470 368.205 3072.750 368.485 ;
        RECT 3073.090 368.205 3073.370 368.485 ;
        RECT 3064.410 367.585 3064.690 367.865 ;
        RECT 3065.030 367.585 3065.310 367.865 ;
        RECT 3065.650 367.585 3065.930 367.865 ;
        RECT 3066.270 367.585 3066.550 367.865 ;
        RECT 3066.890 367.585 3067.170 367.865 ;
        RECT 3067.510 367.585 3067.790 367.865 ;
        RECT 3068.130 367.585 3068.410 367.865 ;
        RECT 3068.750 367.585 3069.030 367.865 ;
        RECT 3069.370 367.585 3069.650 367.865 ;
        RECT 3069.990 367.585 3070.270 367.865 ;
        RECT 3070.610 367.585 3070.890 367.865 ;
        RECT 3071.230 367.585 3071.510 367.865 ;
        RECT 3071.850 367.585 3072.130 367.865 ;
        RECT 3072.470 367.585 3072.750 367.865 ;
        RECT 3073.090 367.585 3073.370 367.865 ;
        RECT 3064.410 366.965 3064.690 367.245 ;
        RECT 3065.030 366.965 3065.310 367.245 ;
        RECT 3065.650 366.965 3065.930 367.245 ;
        RECT 3066.270 366.965 3066.550 367.245 ;
        RECT 3066.890 366.965 3067.170 367.245 ;
        RECT 3067.510 366.965 3067.790 367.245 ;
        RECT 3068.130 366.965 3068.410 367.245 ;
        RECT 3068.750 366.965 3069.030 367.245 ;
        RECT 3069.370 366.965 3069.650 367.245 ;
        RECT 3069.990 366.965 3070.270 367.245 ;
        RECT 3070.610 366.965 3070.890 367.245 ;
        RECT 3071.230 366.965 3071.510 367.245 ;
        RECT 3071.850 366.965 3072.130 367.245 ;
        RECT 3072.470 366.965 3072.750 367.245 ;
        RECT 3073.090 366.965 3073.370 367.245 ;
        RECT 3064.410 366.345 3064.690 366.625 ;
        RECT 3065.030 366.345 3065.310 366.625 ;
        RECT 3065.650 366.345 3065.930 366.625 ;
        RECT 3066.270 366.345 3066.550 366.625 ;
        RECT 3066.890 366.345 3067.170 366.625 ;
        RECT 3067.510 366.345 3067.790 366.625 ;
        RECT 3068.130 366.345 3068.410 366.625 ;
        RECT 3068.750 366.345 3069.030 366.625 ;
        RECT 3069.370 366.345 3069.650 366.625 ;
        RECT 3069.990 366.345 3070.270 366.625 ;
        RECT 3070.610 366.345 3070.890 366.625 ;
        RECT 3071.230 366.345 3071.510 366.625 ;
        RECT 3071.850 366.345 3072.130 366.625 ;
        RECT 3072.470 366.345 3072.750 366.625 ;
        RECT 3073.090 366.345 3073.370 366.625 ;
        RECT 3064.410 365.725 3064.690 366.005 ;
        RECT 3065.030 365.725 3065.310 366.005 ;
        RECT 3065.650 365.725 3065.930 366.005 ;
        RECT 3066.270 365.725 3066.550 366.005 ;
        RECT 3066.890 365.725 3067.170 366.005 ;
        RECT 3067.510 365.725 3067.790 366.005 ;
        RECT 3068.130 365.725 3068.410 366.005 ;
        RECT 3068.750 365.725 3069.030 366.005 ;
        RECT 3069.370 365.725 3069.650 366.005 ;
        RECT 3069.990 365.725 3070.270 366.005 ;
        RECT 3070.610 365.725 3070.890 366.005 ;
        RECT 3071.230 365.725 3071.510 366.005 ;
        RECT 3071.850 365.725 3072.130 366.005 ;
        RECT 3072.470 365.725 3072.750 366.005 ;
        RECT 3073.090 365.725 3073.370 366.005 ;
        RECT 3064.410 365.105 3064.690 365.385 ;
        RECT 3065.030 365.105 3065.310 365.385 ;
        RECT 3065.650 365.105 3065.930 365.385 ;
        RECT 3066.270 365.105 3066.550 365.385 ;
        RECT 3066.890 365.105 3067.170 365.385 ;
        RECT 3067.510 365.105 3067.790 365.385 ;
        RECT 3068.130 365.105 3068.410 365.385 ;
        RECT 3068.750 365.105 3069.030 365.385 ;
        RECT 3069.370 365.105 3069.650 365.385 ;
        RECT 3069.990 365.105 3070.270 365.385 ;
        RECT 3070.610 365.105 3070.890 365.385 ;
        RECT 3071.230 365.105 3071.510 365.385 ;
        RECT 3071.850 365.105 3072.130 365.385 ;
        RECT 3072.470 365.105 3072.750 365.385 ;
        RECT 3073.090 365.105 3073.370 365.385 ;
        RECT 3064.410 364.485 3064.690 364.765 ;
        RECT 3065.030 364.485 3065.310 364.765 ;
        RECT 3065.650 364.485 3065.930 364.765 ;
        RECT 3066.270 364.485 3066.550 364.765 ;
        RECT 3066.890 364.485 3067.170 364.765 ;
        RECT 3067.510 364.485 3067.790 364.765 ;
        RECT 3068.130 364.485 3068.410 364.765 ;
        RECT 3068.750 364.485 3069.030 364.765 ;
        RECT 3069.370 364.485 3069.650 364.765 ;
        RECT 3069.990 364.485 3070.270 364.765 ;
        RECT 3070.610 364.485 3070.890 364.765 ;
        RECT 3071.230 364.485 3071.510 364.765 ;
        RECT 3071.850 364.485 3072.130 364.765 ;
        RECT 3072.470 364.485 3072.750 364.765 ;
        RECT 3073.090 364.485 3073.370 364.765 ;
        RECT 3064.410 363.865 3064.690 364.145 ;
        RECT 3065.030 363.865 3065.310 364.145 ;
        RECT 3065.650 363.865 3065.930 364.145 ;
        RECT 3066.270 363.865 3066.550 364.145 ;
        RECT 3066.890 363.865 3067.170 364.145 ;
        RECT 3067.510 363.865 3067.790 364.145 ;
        RECT 3068.130 363.865 3068.410 364.145 ;
        RECT 3068.750 363.865 3069.030 364.145 ;
        RECT 3069.370 363.865 3069.650 364.145 ;
        RECT 3069.990 363.865 3070.270 364.145 ;
        RECT 3070.610 363.865 3070.890 364.145 ;
        RECT 3071.230 363.865 3071.510 364.145 ;
        RECT 3071.850 363.865 3072.130 364.145 ;
        RECT 3072.470 363.865 3072.750 364.145 ;
        RECT 3073.090 363.865 3073.370 364.145 ;
        RECT 3064.410 363.245 3064.690 363.525 ;
        RECT 3065.030 363.245 3065.310 363.525 ;
        RECT 3065.650 363.245 3065.930 363.525 ;
        RECT 3066.270 363.245 3066.550 363.525 ;
        RECT 3066.890 363.245 3067.170 363.525 ;
        RECT 3067.510 363.245 3067.790 363.525 ;
        RECT 3068.130 363.245 3068.410 363.525 ;
        RECT 3068.750 363.245 3069.030 363.525 ;
        RECT 3069.370 363.245 3069.650 363.525 ;
        RECT 3069.990 363.245 3070.270 363.525 ;
        RECT 3070.610 363.245 3070.890 363.525 ;
        RECT 3071.230 363.245 3071.510 363.525 ;
        RECT 3071.850 363.245 3072.130 363.525 ;
        RECT 3072.470 363.245 3072.750 363.525 ;
        RECT 3073.090 363.245 3073.370 363.525 ;
        RECT 3064.410 362.625 3064.690 362.905 ;
        RECT 3065.030 362.625 3065.310 362.905 ;
        RECT 3065.650 362.625 3065.930 362.905 ;
        RECT 3066.270 362.625 3066.550 362.905 ;
        RECT 3066.890 362.625 3067.170 362.905 ;
        RECT 3067.510 362.625 3067.790 362.905 ;
        RECT 3068.130 362.625 3068.410 362.905 ;
        RECT 3068.750 362.625 3069.030 362.905 ;
        RECT 3069.370 362.625 3069.650 362.905 ;
        RECT 3069.990 362.625 3070.270 362.905 ;
        RECT 3070.610 362.625 3070.890 362.905 ;
        RECT 3071.230 362.625 3071.510 362.905 ;
        RECT 3071.850 362.625 3072.130 362.905 ;
        RECT 3072.470 362.625 3072.750 362.905 ;
        RECT 3073.090 362.625 3073.370 362.905 ;
        RECT 3064.410 362.005 3064.690 362.285 ;
        RECT 3065.030 362.005 3065.310 362.285 ;
        RECT 3065.650 362.005 3065.930 362.285 ;
        RECT 3066.270 362.005 3066.550 362.285 ;
        RECT 3066.890 362.005 3067.170 362.285 ;
        RECT 3067.510 362.005 3067.790 362.285 ;
        RECT 3068.130 362.005 3068.410 362.285 ;
        RECT 3068.750 362.005 3069.030 362.285 ;
        RECT 3069.370 362.005 3069.650 362.285 ;
        RECT 3069.990 362.005 3070.270 362.285 ;
        RECT 3070.610 362.005 3070.890 362.285 ;
        RECT 3071.230 362.005 3071.510 362.285 ;
        RECT 3071.850 362.005 3072.130 362.285 ;
        RECT 3072.470 362.005 3072.750 362.285 ;
        RECT 3073.090 362.005 3073.370 362.285 ;
        RECT 3064.410 361.385 3064.690 361.665 ;
        RECT 3065.030 361.385 3065.310 361.665 ;
        RECT 3065.650 361.385 3065.930 361.665 ;
        RECT 3066.270 361.385 3066.550 361.665 ;
        RECT 3066.890 361.385 3067.170 361.665 ;
        RECT 3067.510 361.385 3067.790 361.665 ;
        RECT 3068.130 361.385 3068.410 361.665 ;
        RECT 3068.750 361.385 3069.030 361.665 ;
        RECT 3069.370 361.385 3069.650 361.665 ;
        RECT 3069.990 361.385 3070.270 361.665 ;
        RECT 3070.610 361.385 3070.890 361.665 ;
        RECT 3071.230 361.385 3071.510 361.665 ;
        RECT 3071.850 361.385 3072.130 361.665 ;
        RECT 3072.470 361.385 3072.750 361.665 ;
        RECT 3073.090 361.385 3073.370 361.665 ;
        RECT 3064.410 360.765 3064.690 361.045 ;
        RECT 3065.030 360.765 3065.310 361.045 ;
        RECT 3065.650 360.765 3065.930 361.045 ;
        RECT 3066.270 360.765 3066.550 361.045 ;
        RECT 3066.890 360.765 3067.170 361.045 ;
        RECT 3067.510 360.765 3067.790 361.045 ;
        RECT 3068.130 360.765 3068.410 361.045 ;
        RECT 3068.750 360.765 3069.030 361.045 ;
        RECT 3069.370 360.765 3069.650 361.045 ;
        RECT 3069.990 360.765 3070.270 361.045 ;
        RECT 3070.610 360.765 3070.890 361.045 ;
        RECT 3071.230 360.765 3071.510 361.045 ;
        RECT 3071.850 360.765 3072.130 361.045 ;
        RECT 3072.470 360.765 3072.750 361.045 ;
        RECT 3073.090 360.765 3073.370 361.045 ;
        RECT 3289.030 379.445 3289.310 379.725 ;
        RECT 3289.650 379.445 3289.930 379.725 ;
        RECT 3290.270 379.445 3290.550 379.725 ;
        RECT 3290.890 379.445 3291.170 379.725 ;
        RECT 3291.510 379.445 3291.790 379.725 ;
        RECT 3292.130 379.445 3292.410 379.725 ;
        RECT 3292.750 379.445 3293.030 379.725 ;
        RECT 3293.370 379.445 3293.650 379.725 ;
        RECT 3293.990 379.445 3294.270 379.725 ;
        RECT 3294.610 379.445 3294.890 379.725 ;
        RECT 3295.230 379.445 3295.510 379.725 ;
        RECT 3295.850 379.445 3296.130 379.725 ;
        RECT 3296.470 379.445 3296.750 379.725 ;
        RECT 3297.090 379.445 3297.370 379.725 ;
        RECT 3297.710 379.445 3297.990 379.725 ;
        RECT 3298.330 379.445 3298.610 379.725 ;
        RECT 3289.030 378.825 3289.310 379.105 ;
        RECT 3289.650 378.825 3289.930 379.105 ;
        RECT 3290.270 378.825 3290.550 379.105 ;
        RECT 3290.890 378.825 3291.170 379.105 ;
        RECT 3291.510 378.825 3291.790 379.105 ;
        RECT 3292.130 378.825 3292.410 379.105 ;
        RECT 3292.750 378.825 3293.030 379.105 ;
        RECT 3293.370 378.825 3293.650 379.105 ;
        RECT 3293.990 378.825 3294.270 379.105 ;
        RECT 3294.610 378.825 3294.890 379.105 ;
        RECT 3295.230 378.825 3295.510 379.105 ;
        RECT 3295.850 378.825 3296.130 379.105 ;
        RECT 3296.470 378.825 3296.750 379.105 ;
        RECT 3297.090 378.825 3297.370 379.105 ;
        RECT 3297.710 378.825 3297.990 379.105 ;
        RECT 3298.330 378.825 3298.610 379.105 ;
        RECT 3289.030 378.205 3289.310 378.485 ;
        RECT 3289.650 378.205 3289.930 378.485 ;
        RECT 3290.270 378.205 3290.550 378.485 ;
        RECT 3290.890 378.205 3291.170 378.485 ;
        RECT 3291.510 378.205 3291.790 378.485 ;
        RECT 3292.130 378.205 3292.410 378.485 ;
        RECT 3292.750 378.205 3293.030 378.485 ;
        RECT 3293.370 378.205 3293.650 378.485 ;
        RECT 3293.990 378.205 3294.270 378.485 ;
        RECT 3294.610 378.205 3294.890 378.485 ;
        RECT 3295.230 378.205 3295.510 378.485 ;
        RECT 3295.850 378.205 3296.130 378.485 ;
        RECT 3296.470 378.205 3296.750 378.485 ;
        RECT 3297.090 378.205 3297.370 378.485 ;
        RECT 3297.710 378.205 3297.990 378.485 ;
        RECT 3298.330 378.205 3298.610 378.485 ;
        RECT 3289.030 377.585 3289.310 377.865 ;
        RECT 3289.650 377.585 3289.930 377.865 ;
        RECT 3290.270 377.585 3290.550 377.865 ;
        RECT 3290.890 377.585 3291.170 377.865 ;
        RECT 3291.510 377.585 3291.790 377.865 ;
        RECT 3292.130 377.585 3292.410 377.865 ;
        RECT 3292.750 377.585 3293.030 377.865 ;
        RECT 3293.370 377.585 3293.650 377.865 ;
        RECT 3293.990 377.585 3294.270 377.865 ;
        RECT 3294.610 377.585 3294.890 377.865 ;
        RECT 3295.230 377.585 3295.510 377.865 ;
        RECT 3295.850 377.585 3296.130 377.865 ;
        RECT 3296.470 377.585 3296.750 377.865 ;
        RECT 3297.090 377.585 3297.370 377.865 ;
        RECT 3297.710 377.585 3297.990 377.865 ;
        RECT 3298.330 377.585 3298.610 377.865 ;
        RECT 3289.030 376.965 3289.310 377.245 ;
        RECT 3289.650 376.965 3289.930 377.245 ;
        RECT 3290.270 376.965 3290.550 377.245 ;
        RECT 3290.890 376.965 3291.170 377.245 ;
        RECT 3291.510 376.965 3291.790 377.245 ;
        RECT 3292.130 376.965 3292.410 377.245 ;
        RECT 3292.750 376.965 3293.030 377.245 ;
        RECT 3293.370 376.965 3293.650 377.245 ;
        RECT 3293.990 376.965 3294.270 377.245 ;
        RECT 3294.610 376.965 3294.890 377.245 ;
        RECT 3295.230 376.965 3295.510 377.245 ;
        RECT 3295.850 376.965 3296.130 377.245 ;
        RECT 3296.470 376.965 3296.750 377.245 ;
        RECT 3297.090 376.965 3297.370 377.245 ;
        RECT 3297.710 376.965 3297.990 377.245 ;
        RECT 3298.330 376.965 3298.610 377.245 ;
        RECT 3289.030 376.345 3289.310 376.625 ;
        RECT 3289.650 376.345 3289.930 376.625 ;
        RECT 3290.270 376.345 3290.550 376.625 ;
        RECT 3290.890 376.345 3291.170 376.625 ;
        RECT 3291.510 376.345 3291.790 376.625 ;
        RECT 3292.130 376.345 3292.410 376.625 ;
        RECT 3292.750 376.345 3293.030 376.625 ;
        RECT 3293.370 376.345 3293.650 376.625 ;
        RECT 3293.990 376.345 3294.270 376.625 ;
        RECT 3294.610 376.345 3294.890 376.625 ;
        RECT 3295.230 376.345 3295.510 376.625 ;
        RECT 3295.850 376.345 3296.130 376.625 ;
        RECT 3296.470 376.345 3296.750 376.625 ;
        RECT 3297.090 376.345 3297.370 376.625 ;
        RECT 3297.710 376.345 3297.990 376.625 ;
        RECT 3298.330 376.345 3298.610 376.625 ;
        RECT 3289.030 375.725 3289.310 376.005 ;
        RECT 3289.650 375.725 3289.930 376.005 ;
        RECT 3290.270 375.725 3290.550 376.005 ;
        RECT 3290.890 375.725 3291.170 376.005 ;
        RECT 3291.510 375.725 3291.790 376.005 ;
        RECT 3292.130 375.725 3292.410 376.005 ;
        RECT 3292.750 375.725 3293.030 376.005 ;
        RECT 3293.370 375.725 3293.650 376.005 ;
        RECT 3293.990 375.725 3294.270 376.005 ;
        RECT 3294.610 375.725 3294.890 376.005 ;
        RECT 3295.230 375.725 3295.510 376.005 ;
        RECT 3295.850 375.725 3296.130 376.005 ;
        RECT 3296.470 375.725 3296.750 376.005 ;
        RECT 3297.090 375.725 3297.370 376.005 ;
        RECT 3297.710 375.725 3297.990 376.005 ;
        RECT 3298.330 375.725 3298.610 376.005 ;
        RECT 3289.030 375.105 3289.310 375.385 ;
        RECT 3289.650 375.105 3289.930 375.385 ;
        RECT 3290.270 375.105 3290.550 375.385 ;
        RECT 3290.890 375.105 3291.170 375.385 ;
        RECT 3291.510 375.105 3291.790 375.385 ;
        RECT 3292.130 375.105 3292.410 375.385 ;
        RECT 3292.750 375.105 3293.030 375.385 ;
        RECT 3293.370 375.105 3293.650 375.385 ;
        RECT 3293.990 375.105 3294.270 375.385 ;
        RECT 3294.610 375.105 3294.890 375.385 ;
        RECT 3295.230 375.105 3295.510 375.385 ;
        RECT 3295.850 375.105 3296.130 375.385 ;
        RECT 3296.470 375.105 3296.750 375.385 ;
        RECT 3297.090 375.105 3297.370 375.385 ;
        RECT 3297.710 375.105 3297.990 375.385 ;
        RECT 3298.330 375.105 3298.610 375.385 ;
        RECT 3289.030 374.485 3289.310 374.765 ;
        RECT 3289.650 374.485 3289.930 374.765 ;
        RECT 3290.270 374.485 3290.550 374.765 ;
        RECT 3290.890 374.485 3291.170 374.765 ;
        RECT 3291.510 374.485 3291.790 374.765 ;
        RECT 3292.130 374.485 3292.410 374.765 ;
        RECT 3292.750 374.485 3293.030 374.765 ;
        RECT 3293.370 374.485 3293.650 374.765 ;
        RECT 3293.990 374.485 3294.270 374.765 ;
        RECT 3294.610 374.485 3294.890 374.765 ;
        RECT 3295.230 374.485 3295.510 374.765 ;
        RECT 3295.850 374.485 3296.130 374.765 ;
        RECT 3296.470 374.485 3296.750 374.765 ;
        RECT 3297.090 374.485 3297.370 374.765 ;
        RECT 3297.710 374.485 3297.990 374.765 ;
        RECT 3298.330 374.485 3298.610 374.765 ;
        RECT 3289.030 373.865 3289.310 374.145 ;
        RECT 3289.650 373.865 3289.930 374.145 ;
        RECT 3290.270 373.865 3290.550 374.145 ;
        RECT 3290.890 373.865 3291.170 374.145 ;
        RECT 3291.510 373.865 3291.790 374.145 ;
        RECT 3292.130 373.865 3292.410 374.145 ;
        RECT 3292.750 373.865 3293.030 374.145 ;
        RECT 3293.370 373.865 3293.650 374.145 ;
        RECT 3293.990 373.865 3294.270 374.145 ;
        RECT 3294.610 373.865 3294.890 374.145 ;
        RECT 3295.230 373.865 3295.510 374.145 ;
        RECT 3295.850 373.865 3296.130 374.145 ;
        RECT 3296.470 373.865 3296.750 374.145 ;
        RECT 3297.090 373.865 3297.370 374.145 ;
        RECT 3297.710 373.865 3297.990 374.145 ;
        RECT 3298.330 373.865 3298.610 374.145 ;
        RECT 3289.030 373.245 3289.310 373.525 ;
        RECT 3289.650 373.245 3289.930 373.525 ;
        RECT 3290.270 373.245 3290.550 373.525 ;
        RECT 3290.890 373.245 3291.170 373.525 ;
        RECT 3291.510 373.245 3291.790 373.525 ;
        RECT 3292.130 373.245 3292.410 373.525 ;
        RECT 3292.750 373.245 3293.030 373.525 ;
        RECT 3293.370 373.245 3293.650 373.525 ;
        RECT 3293.990 373.245 3294.270 373.525 ;
        RECT 3294.610 373.245 3294.890 373.525 ;
        RECT 3295.230 373.245 3295.510 373.525 ;
        RECT 3295.850 373.245 3296.130 373.525 ;
        RECT 3296.470 373.245 3296.750 373.525 ;
        RECT 3297.090 373.245 3297.370 373.525 ;
        RECT 3297.710 373.245 3297.990 373.525 ;
        RECT 3298.330 373.245 3298.610 373.525 ;
        RECT 3289.030 372.625 3289.310 372.905 ;
        RECT 3289.650 372.625 3289.930 372.905 ;
        RECT 3290.270 372.625 3290.550 372.905 ;
        RECT 3290.890 372.625 3291.170 372.905 ;
        RECT 3291.510 372.625 3291.790 372.905 ;
        RECT 3292.130 372.625 3292.410 372.905 ;
        RECT 3292.750 372.625 3293.030 372.905 ;
        RECT 3293.370 372.625 3293.650 372.905 ;
        RECT 3293.990 372.625 3294.270 372.905 ;
        RECT 3294.610 372.625 3294.890 372.905 ;
        RECT 3295.230 372.625 3295.510 372.905 ;
        RECT 3295.850 372.625 3296.130 372.905 ;
        RECT 3296.470 372.625 3296.750 372.905 ;
        RECT 3297.090 372.625 3297.370 372.905 ;
        RECT 3297.710 372.625 3297.990 372.905 ;
        RECT 3298.330 372.625 3298.610 372.905 ;
        RECT 3300.880 379.445 3301.160 379.725 ;
        RECT 3301.500 379.445 3301.780 379.725 ;
        RECT 3302.120 379.445 3302.400 379.725 ;
        RECT 3302.740 379.445 3303.020 379.725 ;
        RECT 3303.360 379.445 3303.640 379.725 ;
        RECT 3303.980 379.445 3304.260 379.725 ;
        RECT 3304.600 379.445 3304.880 379.725 ;
        RECT 3305.220 379.445 3305.500 379.725 ;
        RECT 3305.840 379.445 3306.120 379.725 ;
        RECT 3306.460 379.445 3306.740 379.725 ;
        RECT 3307.080 379.445 3307.360 379.725 ;
        RECT 3307.700 379.445 3307.980 379.725 ;
        RECT 3308.320 379.445 3308.600 379.725 ;
        RECT 3308.940 379.445 3309.220 379.725 ;
        RECT 3309.560 379.445 3309.840 379.725 ;
        RECT 3310.180 379.445 3310.460 379.725 ;
        RECT 3300.880 378.825 3301.160 379.105 ;
        RECT 3301.500 378.825 3301.780 379.105 ;
        RECT 3302.120 378.825 3302.400 379.105 ;
        RECT 3302.740 378.825 3303.020 379.105 ;
        RECT 3303.360 378.825 3303.640 379.105 ;
        RECT 3303.980 378.825 3304.260 379.105 ;
        RECT 3304.600 378.825 3304.880 379.105 ;
        RECT 3305.220 378.825 3305.500 379.105 ;
        RECT 3305.840 378.825 3306.120 379.105 ;
        RECT 3306.460 378.825 3306.740 379.105 ;
        RECT 3307.080 378.825 3307.360 379.105 ;
        RECT 3307.700 378.825 3307.980 379.105 ;
        RECT 3308.320 378.825 3308.600 379.105 ;
        RECT 3308.940 378.825 3309.220 379.105 ;
        RECT 3309.560 378.825 3309.840 379.105 ;
        RECT 3310.180 378.825 3310.460 379.105 ;
        RECT 3300.880 378.205 3301.160 378.485 ;
        RECT 3301.500 378.205 3301.780 378.485 ;
        RECT 3302.120 378.205 3302.400 378.485 ;
        RECT 3302.740 378.205 3303.020 378.485 ;
        RECT 3303.360 378.205 3303.640 378.485 ;
        RECT 3303.980 378.205 3304.260 378.485 ;
        RECT 3304.600 378.205 3304.880 378.485 ;
        RECT 3305.220 378.205 3305.500 378.485 ;
        RECT 3305.840 378.205 3306.120 378.485 ;
        RECT 3306.460 378.205 3306.740 378.485 ;
        RECT 3307.080 378.205 3307.360 378.485 ;
        RECT 3307.700 378.205 3307.980 378.485 ;
        RECT 3308.320 378.205 3308.600 378.485 ;
        RECT 3308.940 378.205 3309.220 378.485 ;
        RECT 3309.560 378.205 3309.840 378.485 ;
        RECT 3310.180 378.205 3310.460 378.485 ;
        RECT 3300.880 377.585 3301.160 377.865 ;
        RECT 3301.500 377.585 3301.780 377.865 ;
        RECT 3302.120 377.585 3302.400 377.865 ;
        RECT 3302.740 377.585 3303.020 377.865 ;
        RECT 3303.360 377.585 3303.640 377.865 ;
        RECT 3303.980 377.585 3304.260 377.865 ;
        RECT 3304.600 377.585 3304.880 377.865 ;
        RECT 3305.220 377.585 3305.500 377.865 ;
        RECT 3305.840 377.585 3306.120 377.865 ;
        RECT 3306.460 377.585 3306.740 377.865 ;
        RECT 3307.080 377.585 3307.360 377.865 ;
        RECT 3307.700 377.585 3307.980 377.865 ;
        RECT 3308.320 377.585 3308.600 377.865 ;
        RECT 3308.940 377.585 3309.220 377.865 ;
        RECT 3309.560 377.585 3309.840 377.865 ;
        RECT 3310.180 377.585 3310.460 377.865 ;
        RECT 3300.880 376.965 3301.160 377.245 ;
        RECT 3301.500 376.965 3301.780 377.245 ;
        RECT 3302.120 376.965 3302.400 377.245 ;
        RECT 3302.740 376.965 3303.020 377.245 ;
        RECT 3303.360 376.965 3303.640 377.245 ;
        RECT 3303.980 376.965 3304.260 377.245 ;
        RECT 3304.600 376.965 3304.880 377.245 ;
        RECT 3305.220 376.965 3305.500 377.245 ;
        RECT 3305.840 376.965 3306.120 377.245 ;
        RECT 3306.460 376.965 3306.740 377.245 ;
        RECT 3307.080 376.965 3307.360 377.245 ;
        RECT 3307.700 376.965 3307.980 377.245 ;
        RECT 3308.320 376.965 3308.600 377.245 ;
        RECT 3308.940 376.965 3309.220 377.245 ;
        RECT 3309.560 376.965 3309.840 377.245 ;
        RECT 3310.180 376.965 3310.460 377.245 ;
        RECT 3300.880 376.345 3301.160 376.625 ;
        RECT 3301.500 376.345 3301.780 376.625 ;
        RECT 3302.120 376.345 3302.400 376.625 ;
        RECT 3302.740 376.345 3303.020 376.625 ;
        RECT 3303.360 376.345 3303.640 376.625 ;
        RECT 3303.980 376.345 3304.260 376.625 ;
        RECT 3304.600 376.345 3304.880 376.625 ;
        RECT 3305.220 376.345 3305.500 376.625 ;
        RECT 3305.840 376.345 3306.120 376.625 ;
        RECT 3306.460 376.345 3306.740 376.625 ;
        RECT 3307.080 376.345 3307.360 376.625 ;
        RECT 3307.700 376.345 3307.980 376.625 ;
        RECT 3308.320 376.345 3308.600 376.625 ;
        RECT 3308.940 376.345 3309.220 376.625 ;
        RECT 3309.560 376.345 3309.840 376.625 ;
        RECT 3310.180 376.345 3310.460 376.625 ;
        RECT 3300.880 375.725 3301.160 376.005 ;
        RECT 3301.500 375.725 3301.780 376.005 ;
        RECT 3302.120 375.725 3302.400 376.005 ;
        RECT 3302.740 375.725 3303.020 376.005 ;
        RECT 3303.360 375.725 3303.640 376.005 ;
        RECT 3303.980 375.725 3304.260 376.005 ;
        RECT 3304.600 375.725 3304.880 376.005 ;
        RECT 3305.220 375.725 3305.500 376.005 ;
        RECT 3305.840 375.725 3306.120 376.005 ;
        RECT 3306.460 375.725 3306.740 376.005 ;
        RECT 3307.080 375.725 3307.360 376.005 ;
        RECT 3307.700 375.725 3307.980 376.005 ;
        RECT 3308.320 375.725 3308.600 376.005 ;
        RECT 3308.940 375.725 3309.220 376.005 ;
        RECT 3309.560 375.725 3309.840 376.005 ;
        RECT 3310.180 375.725 3310.460 376.005 ;
        RECT 3300.880 375.105 3301.160 375.385 ;
        RECT 3301.500 375.105 3301.780 375.385 ;
        RECT 3302.120 375.105 3302.400 375.385 ;
        RECT 3302.740 375.105 3303.020 375.385 ;
        RECT 3303.360 375.105 3303.640 375.385 ;
        RECT 3303.980 375.105 3304.260 375.385 ;
        RECT 3304.600 375.105 3304.880 375.385 ;
        RECT 3305.220 375.105 3305.500 375.385 ;
        RECT 3305.840 375.105 3306.120 375.385 ;
        RECT 3306.460 375.105 3306.740 375.385 ;
        RECT 3307.080 375.105 3307.360 375.385 ;
        RECT 3307.700 375.105 3307.980 375.385 ;
        RECT 3308.320 375.105 3308.600 375.385 ;
        RECT 3308.940 375.105 3309.220 375.385 ;
        RECT 3309.560 375.105 3309.840 375.385 ;
        RECT 3310.180 375.105 3310.460 375.385 ;
        RECT 3300.880 374.485 3301.160 374.765 ;
        RECT 3301.500 374.485 3301.780 374.765 ;
        RECT 3302.120 374.485 3302.400 374.765 ;
        RECT 3302.740 374.485 3303.020 374.765 ;
        RECT 3303.360 374.485 3303.640 374.765 ;
        RECT 3303.980 374.485 3304.260 374.765 ;
        RECT 3304.600 374.485 3304.880 374.765 ;
        RECT 3305.220 374.485 3305.500 374.765 ;
        RECT 3305.840 374.485 3306.120 374.765 ;
        RECT 3306.460 374.485 3306.740 374.765 ;
        RECT 3307.080 374.485 3307.360 374.765 ;
        RECT 3307.700 374.485 3307.980 374.765 ;
        RECT 3308.320 374.485 3308.600 374.765 ;
        RECT 3308.940 374.485 3309.220 374.765 ;
        RECT 3309.560 374.485 3309.840 374.765 ;
        RECT 3310.180 374.485 3310.460 374.765 ;
        RECT 3300.880 373.865 3301.160 374.145 ;
        RECT 3301.500 373.865 3301.780 374.145 ;
        RECT 3302.120 373.865 3302.400 374.145 ;
        RECT 3302.740 373.865 3303.020 374.145 ;
        RECT 3303.360 373.865 3303.640 374.145 ;
        RECT 3303.980 373.865 3304.260 374.145 ;
        RECT 3304.600 373.865 3304.880 374.145 ;
        RECT 3305.220 373.865 3305.500 374.145 ;
        RECT 3305.840 373.865 3306.120 374.145 ;
        RECT 3306.460 373.865 3306.740 374.145 ;
        RECT 3307.080 373.865 3307.360 374.145 ;
        RECT 3307.700 373.865 3307.980 374.145 ;
        RECT 3308.320 373.865 3308.600 374.145 ;
        RECT 3308.940 373.865 3309.220 374.145 ;
        RECT 3309.560 373.865 3309.840 374.145 ;
        RECT 3310.180 373.865 3310.460 374.145 ;
        RECT 3300.880 373.245 3301.160 373.525 ;
        RECT 3301.500 373.245 3301.780 373.525 ;
        RECT 3302.120 373.245 3302.400 373.525 ;
        RECT 3302.740 373.245 3303.020 373.525 ;
        RECT 3303.360 373.245 3303.640 373.525 ;
        RECT 3303.980 373.245 3304.260 373.525 ;
        RECT 3304.600 373.245 3304.880 373.525 ;
        RECT 3305.220 373.245 3305.500 373.525 ;
        RECT 3305.840 373.245 3306.120 373.525 ;
        RECT 3306.460 373.245 3306.740 373.525 ;
        RECT 3307.080 373.245 3307.360 373.525 ;
        RECT 3307.700 373.245 3307.980 373.525 ;
        RECT 3308.320 373.245 3308.600 373.525 ;
        RECT 3308.940 373.245 3309.220 373.525 ;
        RECT 3309.560 373.245 3309.840 373.525 ;
        RECT 3310.180 373.245 3310.460 373.525 ;
        RECT 3300.880 372.625 3301.160 372.905 ;
        RECT 3301.500 372.625 3301.780 372.905 ;
        RECT 3302.120 372.625 3302.400 372.905 ;
        RECT 3302.740 372.625 3303.020 372.905 ;
        RECT 3303.360 372.625 3303.640 372.905 ;
        RECT 3303.980 372.625 3304.260 372.905 ;
        RECT 3304.600 372.625 3304.880 372.905 ;
        RECT 3305.220 372.625 3305.500 372.905 ;
        RECT 3305.840 372.625 3306.120 372.905 ;
        RECT 3306.460 372.625 3306.740 372.905 ;
        RECT 3307.080 372.625 3307.360 372.905 ;
        RECT 3307.700 372.625 3307.980 372.905 ;
        RECT 3308.320 372.625 3308.600 372.905 ;
        RECT 3308.940 372.625 3309.220 372.905 ;
        RECT 3309.560 372.625 3309.840 372.905 ;
        RECT 3310.180 372.625 3310.460 372.905 ;
        RECT 3314.410 379.445 3314.690 379.725 ;
        RECT 3315.030 379.445 3315.310 379.725 ;
        RECT 3315.650 379.445 3315.930 379.725 ;
        RECT 3316.270 379.445 3316.550 379.725 ;
        RECT 3316.890 379.445 3317.170 379.725 ;
        RECT 3317.510 379.445 3317.790 379.725 ;
        RECT 3318.130 379.445 3318.410 379.725 ;
        RECT 3318.750 379.445 3319.030 379.725 ;
        RECT 3319.370 379.445 3319.650 379.725 ;
        RECT 3319.990 379.445 3320.270 379.725 ;
        RECT 3320.610 379.445 3320.890 379.725 ;
        RECT 3321.230 379.445 3321.510 379.725 ;
        RECT 3321.850 379.445 3322.130 379.725 ;
        RECT 3322.470 379.445 3322.750 379.725 ;
        RECT 3323.090 379.445 3323.370 379.725 ;
        RECT 3323.710 379.445 3323.990 379.725 ;
        RECT 3314.410 378.825 3314.690 379.105 ;
        RECT 3315.030 378.825 3315.310 379.105 ;
        RECT 3315.650 378.825 3315.930 379.105 ;
        RECT 3316.270 378.825 3316.550 379.105 ;
        RECT 3316.890 378.825 3317.170 379.105 ;
        RECT 3317.510 378.825 3317.790 379.105 ;
        RECT 3318.130 378.825 3318.410 379.105 ;
        RECT 3318.750 378.825 3319.030 379.105 ;
        RECT 3319.370 378.825 3319.650 379.105 ;
        RECT 3319.990 378.825 3320.270 379.105 ;
        RECT 3320.610 378.825 3320.890 379.105 ;
        RECT 3321.230 378.825 3321.510 379.105 ;
        RECT 3321.850 378.825 3322.130 379.105 ;
        RECT 3322.470 378.825 3322.750 379.105 ;
        RECT 3323.090 378.825 3323.370 379.105 ;
        RECT 3323.710 378.825 3323.990 379.105 ;
        RECT 3314.410 378.205 3314.690 378.485 ;
        RECT 3315.030 378.205 3315.310 378.485 ;
        RECT 3315.650 378.205 3315.930 378.485 ;
        RECT 3316.270 378.205 3316.550 378.485 ;
        RECT 3316.890 378.205 3317.170 378.485 ;
        RECT 3317.510 378.205 3317.790 378.485 ;
        RECT 3318.130 378.205 3318.410 378.485 ;
        RECT 3318.750 378.205 3319.030 378.485 ;
        RECT 3319.370 378.205 3319.650 378.485 ;
        RECT 3319.990 378.205 3320.270 378.485 ;
        RECT 3320.610 378.205 3320.890 378.485 ;
        RECT 3321.230 378.205 3321.510 378.485 ;
        RECT 3321.850 378.205 3322.130 378.485 ;
        RECT 3322.470 378.205 3322.750 378.485 ;
        RECT 3323.090 378.205 3323.370 378.485 ;
        RECT 3323.710 378.205 3323.990 378.485 ;
        RECT 3314.410 377.585 3314.690 377.865 ;
        RECT 3315.030 377.585 3315.310 377.865 ;
        RECT 3315.650 377.585 3315.930 377.865 ;
        RECT 3316.270 377.585 3316.550 377.865 ;
        RECT 3316.890 377.585 3317.170 377.865 ;
        RECT 3317.510 377.585 3317.790 377.865 ;
        RECT 3318.130 377.585 3318.410 377.865 ;
        RECT 3318.750 377.585 3319.030 377.865 ;
        RECT 3319.370 377.585 3319.650 377.865 ;
        RECT 3319.990 377.585 3320.270 377.865 ;
        RECT 3320.610 377.585 3320.890 377.865 ;
        RECT 3321.230 377.585 3321.510 377.865 ;
        RECT 3321.850 377.585 3322.130 377.865 ;
        RECT 3322.470 377.585 3322.750 377.865 ;
        RECT 3323.090 377.585 3323.370 377.865 ;
        RECT 3323.710 377.585 3323.990 377.865 ;
        RECT 3314.410 376.965 3314.690 377.245 ;
        RECT 3315.030 376.965 3315.310 377.245 ;
        RECT 3315.650 376.965 3315.930 377.245 ;
        RECT 3316.270 376.965 3316.550 377.245 ;
        RECT 3316.890 376.965 3317.170 377.245 ;
        RECT 3317.510 376.965 3317.790 377.245 ;
        RECT 3318.130 376.965 3318.410 377.245 ;
        RECT 3318.750 376.965 3319.030 377.245 ;
        RECT 3319.370 376.965 3319.650 377.245 ;
        RECT 3319.990 376.965 3320.270 377.245 ;
        RECT 3320.610 376.965 3320.890 377.245 ;
        RECT 3321.230 376.965 3321.510 377.245 ;
        RECT 3321.850 376.965 3322.130 377.245 ;
        RECT 3322.470 376.965 3322.750 377.245 ;
        RECT 3323.090 376.965 3323.370 377.245 ;
        RECT 3323.710 376.965 3323.990 377.245 ;
        RECT 3314.410 376.345 3314.690 376.625 ;
        RECT 3315.030 376.345 3315.310 376.625 ;
        RECT 3315.650 376.345 3315.930 376.625 ;
        RECT 3316.270 376.345 3316.550 376.625 ;
        RECT 3316.890 376.345 3317.170 376.625 ;
        RECT 3317.510 376.345 3317.790 376.625 ;
        RECT 3318.130 376.345 3318.410 376.625 ;
        RECT 3318.750 376.345 3319.030 376.625 ;
        RECT 3319.370 376.345 3319.650 376.625 ;
        RECT 3319.990 376.345 3320.270 376.625 ;
        RECT 3320.610 376.345 3320.890 376.625 ;
        RECT 3321.230 376.345 3321.510 376.625 ;
        RECT 3321.850 376.345 3322.130 376.625 ;
        RECT 3322.470 376.345 3322.750 376.625 ;
        RECT 3323.090 376.345 3323.370 376.625 ;
        RECT 3323.710 376.345 3323.990 376.625 ;
        RECT 3314.410 375.725 3314.690 376.005 ;
        RECT 3315.030 375.725 3315.310 376.005 ;
        RECT 3315.650 375.725 3315.930 376.005 ;
        RECT 3316.270 375.725 3316.550 376.005 ;
        RECT 3316.890 375.725 3317.170 376.005 ;
        RECT 3317.510 375.725 3317.790 376.005 ;
        RECT 3318.130 375.725 3318.410 376.005 ;
        RECT 3318.750 375.725 3319.030 376.005 ;
        RECT 3319.370 375.725 3319.650 376.005 ;
        RECT 3319.990 375.725 3320.270 376.005 ;
        RECT 3320.610 375.725 3320.890 376.005 ;
        RECT 3321.230 375.725 3321.510 376.005 ;
        RECT 3321.850 375.725 3322.130 376.005 ;
        RECT 3322.470 375.725 3322.750 376.005 ;
        RECT 3323.090 375.725 3323.370 376.005 ;
        RECT 3323.710 375.725 3323.990 376.005 ;
        RECT 3314.410 375.105 3314.690 375.385 ;
        RECT 3315.030 375.105 3315.310 375.385 ;
        RECT 3315.650 375.105 3315.930 375.385 ;
        RECT 3316.270 375.105 3316.550 375.385 ;
        RECT 3316.890 375.105 3317.170 375.385 ;
        RECT 3317.510 375.105 3317.790 375.385 ;
        RECT 3318.130 375.105 3318.410 375.385 ;
        RECT 3318.750 375.105 3319.030 375.385 ;
        RECT 3319.370 375.105 3319.650 375.385 ;
        RECT 3319.990 375.105 3320.270 375.385 ;
        RECT 3320.610 375.105 3320.890 375.385 ;
        RECT 3321.230 375.105 3321.510 375.385 ;
        RECT 3321.850 375.105 3322.130 375.385 ;
        RECT 3322.470 375.105 3322.750 375.385 ;
        RECT 3323.090 375.105 3323.370 375.385 ;
        RECT 3323.710 375.105 3323.990 375.385 ;
        RECT 3314.410 374.485 3314.690 374.765 ;
        RECT 3315.030 374.485 3315.310 374.765 ;
        RECT 3315.650 374.485 3315.930 374.765 ;
        RECT 3316.270 374.485 3316.550 374.765 ;
        RECT 3316.890 374.485 3317.170 374.765 ;
        RECT 3317.510 374.485 3317.790 374.765 ;
        RECT 3318.130 374.485 3318.410 374.765 ;
        RECT 3318.750 374.485 3319.030 374.765 ;
        RECT 3319.370 374.485 3319.650 374.765 ;
        RECT 3319.990 374.485 3320.270 374.765 ;
        RECT 3320.610 374.485 3320.890 374.765 ;
        RECT 3321.230 374.485 3321.510 374.765 ;
        RECT 3321.850 374.485 3322.130 374.765 ;
        RECT 3322.470 374.485 3322.750 374.765 ;
        RECT 3323.090 374.485 3323.370 374.765 ;
        RECT 3323.710 374.485 3323.990 374.765 ;
        RECT 3314.410 373.865 3314.690 374.145 ;
        RECT 3315.030 373.865 3315.310 374.145 ;
        RECT 3315.650 373.865 3315.930 374.145 ;
        RECT 3316.270 373.865 3316.550 374.145 ;
        RECT 3316.890 373.865 3317.170 374.145 ;
        RECT 3317.510 373.865 3317.790 374.145 ;
        RECT 3318.130 373.865 3318.410 374.145 ;
        RECT 3318.750 373.865 3319.030 374.145 ;
        RECT 3319.370 373.865 3319.650 374.145 ;
        RECT 3319.990 373.865 3320.270 374.145 ;
        RECT 3320.610 373.865 3320.890 374.145 ;
        RECT 3321.230 373.865 3321.510 374.145 ;
        RECT 3321.850 373.865 3322.130 374.145 ;
        RECT 3322.470 373.865 3322.750 374.145 ;
        RECT 3323.090 373.865 3323.370 374.145 ;
        RECT 3323.710 373.865 3323.990 374.145 ;
        RECT 3314.410 373.245 3314.690 373.525 ;
        RECT 3315.030 373.245 3315.310 373.525 ;
        RECT 3315.650 373.245 3315.930 373.525 ;
        RECT 3316.270 373.245 3316.550 373.525 ;
        RECT 3316.890 373.245 3317.170 373.525 ;
        RECT 3317.510 373.245 3317.790 373.525 ;
        RECT 3318.130 373.245 3318.410 373.525 ;
        RECT 3318.750 373.245 3319.030 373.525 ;
        RECT 3319.370 373.245 3319.650 373.525 ;
        RECT 3319.990 373.245 3320.270 373.525 ;
        RECT 3320.610 373.245 3320.890 373.525 ;
        RECT 3321.230 373.245 3321.510 373.525 ;
        RECT 3321.850 373.245 3322.130 373.525 ;
        RECT 3322.470 373.245 3322.750 373.525 ;
        RECT 3323.090 373.245 3323.370 373.525 ;
        RECT 3323.710 373.245 3323.990 373.525 ;
        RECT 3314.410 372.625 3314.690 372.905 ;
        RECT 3315.030 372.625 3315.310 372.905 ;
        RECT 3315.650 372.625 3315.930 372.905 ;
        RECT 3316.270 372.625 3316.550 372.905 ;
        RECT 3316.890 372.625 3317.170 372.905 ;
        RECT 3317.510 372.625 3317.790 372.905 ;
        RECT 3318.130 372.625 3318.410 372.905 ;
        RECT 3318.750 372.625 3319.030 372.905 ;
        RECT 3319.370 372.625 3319.650 372.905 ;
        RECT 3319.990 372.625 3320.270 372.905 ;
        RECT 3320.610 372.625 3320.890 372.905 ;
        RECT 3321.230 372.625 3321.510 372.905 ;
        RECT 3321.850 372.625 3322.130 372.905 ;
        RECT 3322.470 372.625 3322.750 372.905 ;
        RECT 3323.090 372.625 3323.370 372.905 ;
        RECT 3323.710 372.625 3323.990 372.905 ;
        RECT 3326.260 379.445 3326.540 379.725 ;
        RECT 3326.880 379.445 3327.160 379.725 ;
        RECT 3327.500 379.445 3327.780 379.725 ;
        RECT 3328.120 379.445 3328.400 379.725 ;
        RECT 3328.740 379.445 3329.020 379.725 ;
        RECT 3329.360 379.445 3329.640 379.725 ;
        RECT 3329.980 379.445 3330.260 379.725 ;
        RECT 3330.600 379.445 3330.880 379.725 ;
        RECT 3331.220 379.445 3331.500 379.725 ;
        RECT 3331.840 379.445 3332.120 379.725 ;
        RECT 3332.460 379.445 3332.740 379.725 ;
        RECT 3333.080 379.445 3333.360 379.725 ;
        RECT 3333.700 379.445 3333.980 379.725 ;
        RECT 3334.320 379.445 3334.600 379.725 ;
        RECT 3334.940 379.445 3335.220 379.725 ;
        RECT 3335.560 379.445 3335.840 379.725 ;
        RECT 3326.260 378.825 3326.540 379.105 ;
        RECT 3326.880 378.825 3327.160 379.105 ;
        RECT 3327.500 378.825 3327.780 379.105 ;
        RECT 3328.120 378.825 3328.400 379.105 ;
        RECT 3328.740 378.825 3329.020 379.105 ;
        RECT 3329.360 378.825 3329.640 379.105 ;
        RECT 3329.980 378.825 3330.260 379.105 ;
        RECT 3330.600 378.825 3330.880 379.105 ;
        RECT 3331.220 378.825 3331.500 379.105 ;
        RECT 3331.840 378.825 3332.120 379.105 ;
        RECT 3332.460 378.825 3332.740 379.105 ;
        RECT 3333.080 378.825 3333.360 379.105 ;
        RECT 3333.700 378.825 3333.980 379.105 ;
        RECT 3334.320 378.825 3334.600 379.105 ;
        RECT 3334.940 378.825 3335.220 379.105 ;
        RECT 3335.560 378.825 3335.840 379.105 ;
        RECT 3326.260 378.205 3326.540 378.485 ;
        RECT 3326.880 378.205 3327.160 378.485 ;
        RECT 3327.500 378.205 3327.780 378.485 ;
        RECT 3328.120 378.205 3328.400 378.485 ;
        RECT 3328.740 378.205 3329.020 378.485 ;
        RECT 3329.360 378.205 3329.640 378.485 ;
        RECT 3329.980 378.205 3330.260 378.485 ;
        RECT 3330.600 378.205 3330.880 378.485 ;
        RECT 3331.220 378.205 3331.500 378.485 ;
        RECT 3331.840 378.205 3332.120 378.485 ;
        RECT 3332.460 378.205 3332.740 378.485 ;
        RECT 3333.080 378.205 3333.360 378.485 ;
        RECT 3333.700 378.205 3333.980 378.485 ;
        RECT 3334.320 378.205 3334.600 378.485 ;
        RECT 3334.940 378.205 3335.220 378.485 ;
        RECT 3335.560 378.205 3335.840 378.485 ;
        RECT 3326.260 377.585 3326.540 377.865 ;
        RECT 3326.880 377.585 3327.160 377.865 ;
        RECT 3327.500 377.585 3327.780 377.865 ;
        RECT 3328.120 377.585 3328.400 377.865 ;
        RECT 3328.740 377.585 3329.020 377.865 ;
        RECT 3329.360 377.585 3329.640 377.865 ;
        RECT 3329.980 377.585 3330.260 377.865 ;
        RECT 3330.600 377.585 3330.880 377.865 ;
        RECT 3331.220 377.585 3331.500 377.865 ;
        RECT 3331.840 377.585 3332.120 377.865 ;
        RECT 3332.460 377.585 3332.740 377.865 ;
        RECT 3333.080 377.585 3333.360 377.865 ;
        RECT 3333.700 377.585 3333.980 377.865 ;
        RECT 3334.320 377.585 3334.600 377.865 ;
        RECT 3334.940 377.585 3335.220 377.865 ;
        RECT 3335.560 377.585 3335.840 377.865 ;
        RECT 3326.260 376.965 3326.540 377.245 ;
        RECT 3326.880 376.965 3327.160 377.245 ;
        RECT 3327.500 376.965 3327.780 377.245 ;
        RECT 3328.120 376.965 3328.400 377.245 ;
        RECT 3328.740 376.965 3329.020 377.245 ;
        RECT 3329.360 376.965 3329.640 377.245 ;
        RECT 3329.980 376.965 3330.260 377.245 ;
        RECT 3330.600 376.965 3330.880 377.245 ;
        RECT 3331.220 376.965 3331.500 377.245 ;
        RECT 3331.840 376.965 3332.120 377.245 ;
        RECT 3332.460 376.965 3332.740 377.245 ;
        RECT 3333.080 376.965 3333.360 377.245 ;
        RECT 3333.700 376.965 3333.980 377.245 ;
        RECT 3334.320 376.965 3334.600 377.245 ;
        RECT 3334.940 376.965 3335.220 377.245 ;
        RECT 3335.560 376.965 3335.840 377.245 ;
        RECT 3326.260 376.345 3326.540 376.625 ;
        RECT 3326.880 376.345 3327.160 376.625 ;
        RECT 3327.500 376.345 3327.780 376.625 ;
        RECT 3328.120 376.345 3328.400 376.625 ;
        RECT 3328.740 376.345 3329.020 376.625 ;
        RECT 3329.360 376.345 3329.640 376.625 ;
        RECT 3329.980 376.345 3330.260 376.625 ;
        RECT 3330.600 376.345 3330.880 376.625 ;
        RECT 3331.220 376.345 3331.500 376.625 ;
        RECT 3331.840 376.345 3332.120 376.625 ;
        RECT 3332.460 376.345 3332.740 376.625 ;
        RECT 3333.080 376.345 3333.360 376.625 ;
        RECT 3333.700 376.345 3333.980 376.625 ;
        RECT 3334.320 376.345 3334.600 376.625 ;
        RECT 3334.940 376.345 3335.220 376.625 ;
        RECT 3335.560 376.345 3335.840 376.625 ;
        RECT 3326.260 375.725 3326.540 376.005 ;
        RECT 3326.880 375.725 3327.160 376.005 ;
        RECT 3327.500 375.725 3327.780 376.005 ;
        RECT 3328.120 375.725 3328.400 376.005 ;
        RECT 3328.740 375.725 3329.020 376.005 ;
        RECT 3329.360 375.725 3329.640 376.005 ;
        RECT 3329.980 375.725 3330.260 376.005 ;
        RECT 3330.600 375.725 3330.880 376.005 ;
        RECT 3331.220 375.725 3331.500 376.005 ;
        RECT 3331.840 375.725 3332.120 376.005 ;
        RECT 3332.460 375.725 3332.740 376.005 ;
        RECT 3333.080 375.725 3333.360 376.005 ;
        RECT 3333.700 375.725 3333.980 376.005 ;
        RECT 3334.320 375.725 3334.600 376.005 ;
        RECT 3334.940 375.725 3335.220 376.005 ;
        RECT 3335.560 375.725 3335.840 376.005 ;
        RECT 3326.260 375.105 3326.540 375.385 ;
        RECT 3326.880 375.105 3327.160 375.385 ;
        RECT 3327.500 375.105 3327.780 375.385 ;
        RECT 3328.120 375.105 3328.400 375.385 ;
        RECT 3328.740 375.105 3329.020 375.385 ;
        RECT 3329.360 375.105 3329.640 375.385 ;
        RECT 3329.980 375.105 3330.260 375.385 ;
        RECT 3330.600 375.105 3330.880 375.385 ;
        RECT 3331.220 375.105 3331.500 375.385 ;
        RECT 3331.840 375.105 3332.120 375.385 ;
        RECT 3332.460 375.105 3332.740 375.385 ;
        RECT 3333.080 375.105 3333.360 375.385 ;
        RECT 3333.700 375.105 3333.980 375.385 ;
        RECT 3334.320 375.105 3334.600 375.385 ;
        RECT 3334.940 375.105 3335.220 375.385 ;
        RECT 3335.560 375.105 3335.840 375.385 ;
        RECT 3326.260 374.485 3326.540 374.765 ;
        RECT 3326.880 374.485 3327.160 374.765 ;
        RECT 3327.500 374.485 3327.780 374.765 ;
        RECT 3328.120 374.485 3328.400 374.765 ;
        RECT 3328.740 374.485 3329.020 374.765 ;
        RECT 3329.360 374.485 3329.640 374.765 ;
        RECT 3329.980 374.485 3330.260 374.765 ;
        RECT 3330.600 374.485 3330.880 374.765 ;
        RECT 3331.220 374.485 3331.500 374.765 ;
        RECT 3331.840 374.485 3332.120 374.765 ;
        RECT 3332.460 374.485 3332.740 374.765 ;
        RECT 3333.080 374.485 3333.360 374.765 ;
        RECT 3333.700 374.485 3333.980 374.765 ;
        RECT 3334.320 374.485 3334.600 374.765 ;
        RECT 3334.940 374.485 3335.220 374.765 ;
        RECT 3335.560 374.485 3335.840 374.765 ;
        RECT 3326.260 373.865 3326.540 374.145 ;
        RECT 3326.880 373.865 3327.160 374.145 ;
        RECT 3327.500 373.865 3327.780 374.145 ;
        RECT 3328.120 373.865 3328.400 374.145 ;
        RECT 3328.740 373.865 3329.020 374.145 ;
        RECT 3329.360 373.865 3329.640 374.145 ;
        RECT 3329.980 373.865 3330.260 374.145 ;
        RECT 3330.600 373.865 3330.880 374.145 ;
        RECT 3331.220 373.865 3331.500 374.145 ;
        RECT 3331.840 373.865 3332.120 374.145 ;
        RECT 3332.460 373.865 3332.740 374.145 ;
        RECT 3333.080 373.865 3333.360 374.145 ;
        RECT 3333.700 373.865 3333.980 374.145 ;
        RECT 3334.320 373.865 3334.600 374.145 ;
        RECT 3334.940 373.865 3335.220 374.145 ;
        RECT 3335.560 373.865 3335.840 374.145 ;
        RECT 3326.260 373.245 3326.540 373.525 ;
        RECT 3326.880 373.245 3327.160 373.525 ;
        RECT 3327.500 373.245 3327.780 373.525 ;
        RECT 3328.120 373.245 3328.400 373.525 ;
        RECT 3328.740 373.245 3329.020 373.525 ;
        RECT 3329.360 373.245 3329.640 373.525 ;
        RECT 3329.980 373.245 3330.260 373.525 ;
        RECT 3330.600 373.245 3330.880 373.525 ;
        RECT 3331.220 373.245 3331.500 373.525 ;
        RECT 3331.840 373.245 3332.120 373.525 ;
        RECT 3332.460 373.245 3332.740 373.525 ;
        RECT 3333.080 373.245 3333.360 373.525 ;
        RECT 3333.700 373.245 3333.980 373.525 ;
        RECT 3334.320 373.245 3334.600 373.525 ;
        RECT 3334.940 373.245 3335.220 373.525 ;
        RECT 3335.560 373.245 3335.840 373.525 ;
        RECT 3326.260 372.625 3326.540 372.905 ;
        RECT 3326.880 372.625 3327.160 372.905 ;
        RECT 3327.500 372.625 3327.780 372.905 ;
        RECT 3328.120 372.625 3328.400 372.905 ;
        RECT 3328.740 372.625 3329.020 372.905 ;
        RECT 3329.360 372.625 3329.640 372.905 ;
        RECT 3329.980 372.625 3330.260 372.905 ;
        RECT 3330.600 372.625 3330.880 372.905 ;
        RECT 3331.220 372.625 3331.500 372.905 ;
        RECT 3331.840 372.625 3332.120 372.905 ;
        RECT 3332.460 372.625 3332.740 372.905 ;
        RECT 3333.080 372.625 3333.360 372.905 ;
        RECT 3333.700 372.625 3333.980 372.905 ;
        RECT 3334.320 372.625 3334.600 372.905 ;
        RECT 3334.940 372.625 3335.220 372.905 ;
        RECT 3335.560 372.625 3335.840 372.905 ;
        RECT 3339.410 379.445 3339.690 379.725 ;
        RECT 3340.030 379.445 3340.310 379.725 ;
        RECT 3340.650 379.445 3340.930 379.725 ;
        RECT 3341.270 379.445 3341.550 379.725 ;
        RECT 3341.890 379.445 3342.170 379.725 ;
        RECT 3342.510 379.445 3342.790 379.725 ;
        RECT 3343.130 379.445 3343.410 379.725 ;
        RECT 3343.750 379.445 3344.030 379.725 ;
        RECT 3344.370 379.445 3344.650 379.725 ;
        RECT 3344.990 379.445 3345.270 379.725 ;
        RECT 3345.610 379.445 3345.890 379.725 ;
        RECT 3346.230 379.445 3346.510 379.725 ;
        RECT 3346.850 379.445 3347.130 379.725 ;
        RECT 3347.470 379.445 3347.750 379.725 ;
        RECT 3348.090 379.445 3348.370 379.725 ;
        RECT 3339.410 378.825 3339.690 379.105 ;
        RECT 3340.030 378.825 3340.310 379.105 ;
        RECT 3340.650 378.825 3340.930 379.105 ;
        RECT 3341.270 378.825 3341.550 379.105 ;
        RECT 3341.890 378.825 3342.170 379.105 ;
        RECT 3342.510 378.825 3342.790 379.105 ;
        RECT 3343.130 378.825 3343.410 379.105 ;
        RECT 3343.750 378.825 3344.030 379.105 ;
        RECT 3344.370 378.825 3344.650 379.105 ;
        RECT 3344.990 378.825 3345.270 379.105 ;
        RECT 3345.610 378.825 3345.890 379.105 ;
        RECT 3346.230 378.825 3346.510 379.105 ;
        RECT 3346.850 378.825 3347.130 379.105 ;
        RECT 3347.470 378.825 3347.750 379.105 ;
        RECT 3348.090 378.825 3348.370 379.105 ;
        RECT 3339.410 378.205 3339.690 378.485 ;
        RECT 3340.030 378.205 3340.310 378.485 ;
        RECT 3340.650 378.205 3340.930 378.485 ;
        RECT 3341.270 378.205 3341.550 378.485 ;
        RECT 3341.890 378.205 3342.170 378.485 ;
        RECT 3342.510 378.205 3342.790 378.485 ;
        RECT 3343.130 378.205 3343.410 378.485 ;
        RECT 3343.750 378.205 3344.030 378.485 ;
        RECT 3344.370 378.205 3344.650 378.485 ;
        RECT 3344.990 378.205 3345.270 378.485 ;
        RECT 3345.610 378.205 3345.890 378.485 ;
        RECT 3346.230 378.205 3346.510 378.485 ;
        RECT 3346.850 378.205 3347.130 378.485 ;
        RECT 3347.470 378.205 3347.750 378.485 ;
        RECT 3348.090 378.205 3348.370 378.485 ;
        RECT 3339.410 377.585 3339.690 377.865 ;
        RECT 3340.030 377.585 3340.310 377.865 ;
        RECT 3340.650 377.585 3340.930 377.865 ;
        RECT 3341.270 377.585 3341.550 377.865 ;
        RECT 3341.890 377.585 3342.170 377.865 ;
        RECT 3342.510 377.585 3342.790 377.865 ;
        RECT 3343.130 377.585 3343.410 377.865 ;
        RECT 3343.750 377.585 3344.030 377.865 ;
        RECT 3344.370 377.585 3344.650 377.865 ;
        RECT 3344.990 377.585 3345.270 377.865 ;
        RECT 3345.610 377.585 3345.890 377.865 ;
        RECT 3346.230 377.585 3346.510 377.865 ;
        RECT 3346.850 377.585 3347.130 377.865 ;
        RECT 3347.470 377.585 3347.750 377.865 ;
        RECT 3348.090 377.585 3348.370 377.865 ;
        RECT 3339.410 376.965 3339.690 377.245 ;
        RECT 3340.030 376.965 3340.310 377.245 ;
        RECT 3340.650 376.965 3340.930 377.245 ;
        RECT 3341.270 376.965 3341.550 377.245 ;
        RECT 3341.890 376.965 3342.170 377.245 ;
        RECT 3342.510 376.965 3342.790 377.245 ;
        RECT 3343.130 376.965 3343.410 377.245 ;
        RECT 3343.750 376.965 3344.030 377.245 ;
        RECT 3344.370 376.965 3344.650 377.245 ;
        RECT 3344.990 376.965 3345.270 377.245 ;
        RECT 3345.610 376.965 3345.890 377.245 ;
        RECT 3346.230 376.965 3346.510 377.245 ;
        RECT 3346.850 376.965 3347.130 377.245 ;
        RECT 3347.470 376.965 3347.750 377.245 ;
        RECT 3348.090 376.965 3348.370 377.245 ;
        RECT 3339.410 376.345 3339.690 376.625 ;
        RECT 3340.030 376.345 3340.310 376.625 ;
        RECT 3340.650 376.345 3340.930 376.625 ;
        RECT 3341.270 376.345 3341.550 376.625 ;
        RECT 3341.890 376.345 3342.170 376.625 ;
        RECT 3342.510 376.345 3342.790 376.625 ;
        RECT 3343.130 376.345 3343.410 376.625 ;
        RECT 3343.750 376.345 3344.030 376.625 ;
        RECT 3344.370 376.345 3344.650 376.625 ;
        RECT 3344.990 376.345 3345.270 376.625 ;
        RECT 3345.610 376.345 3345.890 376.625 ;
        RECT 3346.230 376.345 3346.510 376.625 ;
        RECT 3346.850 376.345 3347.130 376.625 ;
        RECT 3347.470 376.345 3347.750 376.625 ;
        RECT 3348.090 376.345 3348.370 376.625 ;
        RECT 3339.410 375.725 3339.690 376.005 ;
        RECT 3340.030 375.725 3340.310 376.005 ;
        RECT 3340.650 375.725 3340.930 376.005 ;
        RECT 3341.270 375.725 3341.550 376.005 ;
        RECT 3341.890 375.725 3342.170 376.005 ;
        RECT 3342.510 375.725 3342.790 376.005 ;
        RECT 3343.130 375.725 3343.410 376.005 ;
        RECT 3343.750 375.725 3344.030 376.005 ;
        RECT 3344.370 375.725 3344.650 376.005 ;
        RECT 3344.990 375.725 3345.270 376.005 ;
        RECT 3345.610 375.725 3345.890 376.005 ;
        RECT 3346.230 375.725 3346.510 376.005 ;
        RECT 3346.850 375.725 3347.130 376.005 ;
        RECT 3347.470 375.725 3347.750 376.005 ;
        RECT 3348.090 375.725 3348.370 376.005 ;
        RECT 3339.410 375.105 3339.690 375.385 ;
        RECT 3340.030 375.105 3340.310 375.385 ;
        RECT 3340.650 375.105 3340.930 375.385 ;
        RECT 3341.270 375.105 3341.550 375.385 ;
        RECT 3341.890 375.105 3342.170 375.385 ;
        RECT 3342.510 375.105 3342.790 375.385 ;
        RECT 3343.130 375.105 3343.410 375.385 ;
        RECT 3343.750 375.105 3344.030 375.385 ;
        RECT 3344.370 375.105 3344.650 375.385 ;
        RECT 3344.990 375.105 3345.270 375.385 ;
        RECT 3345.610 375.105 3345.890 375.385 ;
        RECT 3346.230 375.105 3346.510 375.385 ;
        RECT 3346.850 375.105 3347.130 375.385 ;
        RECT 3347.470 375.105 3347.750 375.385 ;
        RECT 3348.090 375.105 3348.370 375.385 ;
        RECT 3339.410 374.485 3339.690 374.765 ;
        RECT 3340.030 374.485 3340.310 374.765 ;
        RECT 3340.650 374.485 3340.930 374.765 ;
        RECT 3341.270 374.485 3341.550 374.765 ;
        RECT 3341.890 374.485 3342.170 374.765 ;
        RECT 3342.510 374.485 3342.790 374.765 ;
        RECT 3343.130 374.485 3343.410 374.765 ;
        RECT 3343.750 374.485 3344.030 374.765 ;
        RECT 3344.370 374.485 3344.650 374.765 ;
        RECT 3344.990 374.485 3345.270 374.765 ;
        RECT 3345.610 374.485 3345.890 374.765 ;
        RECT 3346.230 374.485 3346.510 374.765 ;
        RECT 3346.850 374.485 3347.130 374.765 ;
        RECT 3347.470 374.485 3347.750 374.765 ;
        RECT 3348.090 374.485 3348.370 374.765 ;
        RECT 3339.410 373.865 3339.690 374.145 ;
        RECT 3340.030 373.865 3340.310 374.145 ;
        RECT 3340.650 373.865 3340.930 374.145 ;
        RECT 3341.270 373.865 3341.550 374.145 ;
        RECT 3341.890 373.865 3342.170 374.145 ;
        RECT 3342.510 373.865 3342.790 374.145 ;
        RECT 3343.130 373.865 3343.410 374.145 ;
        RECT 3343.750 373.865 3344.030 374.145 ;
        RECT 3344.370 373.865 3344.650 374.145 ;
        RECT 3344.990 373.865 3345.270 374.145 ;
        RECT 3345.610 373.865 3345.890 374.145 ;
        RECT 3346.230 373.865 3346.510 374.145 ;
        RECT 3346.850 373.865 3347.130 374.145 ;
        RECT 3347.470 373.865 3347.750 374.145 ;
        RECT 3348.090 373.865 3348.370 374.145 ;
        RECT 3339.410 373.245 3339.690 373.525 ;
        RECT 3340.030 373.245 3340.310 373.525 ;
        RECT 3340.650 373.245 3340.930 373.525 ;
        RECT 3341.270 373.245 3341.550 373.525 ;
        RECT 3341.890 373.245 3342.170 373.525 ;
        RECT 3342.510 373.245 3342.790 373.525 ;
        RECT 3343.130 373.245 3343.410 373.525 ;
        RECT 3343.750 373.245 3344.030 373.525 ;
        RECT 3344.370 373.245 3344.650 373.525 ;
        RECT 3344.990 373.245 3345.270 373.525 ;
        RECT 3345.610 373.245 3345.890 373.525 ;
        RECT 3346.230 373.245 3346.510 373.525 ;
        RECT 3346.850 373.245 3347.130 373.525 ;
        RECT 3347.470 373.245 3347.750 373.525 ;
        RECT 3348.090 373.245 3348.370 373.525 ;
        RECT 3339.410 372.625 3339.690 372.905 ;
        RECT 3340.030 372.625 3340.310 372.905 ;
        RECT 3340.650 372.625 3340.930 372.905 ;
        RECT 3341.270 372.625 3341.550 372.905 ;
        RECT 3341.890 372.625 3342.170 372.905 ;
        RECT 3342.510 372.625 3342.790 372.905 ;
        RECT 3343.130 372.625 3343.410 372.905 ;
        RECT 3343.750 372.625 3344.030 372.905 ;
        RECT 3344.370 372.625 3344.650 372.905 ;
        RECT 3344.990 372.625 3345.270 372.905 ;
        RECT 3345.610 372.625 3345.890 372.905 ;
        RECT 3346.230 372.625 3346.510 372.905 ;
        RECT 3346.850 372.625 3347.130 372.905 ;
        RECT 3347.470 372.625 3347.750 372.905 ;
        RECT 3348.090 372.625 3348.370 372.905 ;
      LAYER Metal3 ;
        RECT 1896.360 4698.600 1905.860 4708.600 ;
        RECT 1908.760 4698.600 1919.010 4708.600 ;
        RECT 1920.610 4698.600 1930.860 4708.600 ;
        RECT 1934.140 4698.600 1944.390 4708.600 ;
        RECT 1945.990 4698.600 1956.240 4708.600 ;
        RECT 1959.140 4698.600 1968.640 4708.600 ;
        RECT 2996.360 4698.600 3005.860 4708.600 ;
        RECT 3008.760 4698.600 3019.010 4708.600 ;
        RECT 3020.610 4698.600 3030.860 4708.600 ;
        RECT 3034.140 4698.600 3044.390 4708.600 ;
        RECT 3045.990 4698.600 3056.240 4708.600 ;
        RECT 3059.140 4698.600 3068.640 4708.600 ;
        RECT 350.000 4384.140 379.080 4393.640 ;
        RECT 350.000 4370.990 379.080 4381.240 ;
        RECT 3499.960 4379.140 3530.000 4388.640 ;
        RECT 350.000 4359.140 379.080 4369.390 ;
        RECT 3499.960 4365.990 3530.000 4376.240 ;
        RECT 350.000 4345.610 379.080 4355.860 ;
        RECT 3499.960 4354.140 3530.000 4364.390 ;
        RECT 350.000 4333.760 379.080 4344.010 ;
        RECT 3499.960 4340.610 3530.000 4350.860 ;
        RECT 350.000 4321.360 379.080 4330.860 ;
        RECT 3499.960 4328.760 3530.000 4339.010 ;
        RECT 3499.960 4316.360 3530.000 4325.860 ;
        RECT 350.000 4179.140 377.080 4188.640 ;
        RECT 350.000 4165.990 377.080 4176.240 ;
        RECT 350.000 4154.140 377.080 4164.390 ;
        RECT 350.000 4140.610 377.080 4150.860 ;
        RECT 350.000 4128.760 377.080 4139.010 ;
        RECT 350.000 4116.360 377.080 4125.860 ;
        RECT 350.000 3974.140 367.080 3983.640 ;
        RECT 350.000 3960.990 367.080 3971.240 ;
        RECT 350.000 3949.140 367.080 3959.390 ;
        RECT 3499.960 3949.140 3530.000 3958.640 ;
        RECT 350.000 3935.610 367.080 3945.860 ;
        RECT 3499.960 3935.990 3530.000 3946.240 ;
        RECT 350.000 3923.760 367.080 3934.010 ;
        RECT 3499.960 3924.140 3530.000 3934.390 ;
        RECT 350.000 3911.360 367.080 3920.860 ;
        RECT 3499.960 3910.610 3530.000 3920.860 ;
        RECT 3499.960 3898.760 3530.000 3909.010 ;
        RECT 3499.960 3886.360 3530.000 3895.860 ;
        RECT 3499.960 2444.140 3530.000 2453.640 ;
        RECT 3499.960 2430.990 3530.000 2441.240 ;
        RECT 3499.960 2419.140 3530.000 2429.390 ;
        RECT 3499.960 2405.610 3530.000 2415.860 ;
        RECT 3499.960 2393.760 3530.000 2404.010 ;
        RECT 3499.960 2381.360 3530.000 2390.860 ;
        RECT 350.000 2334.140 377.080 2343.640 ;
        RECT 350.000 2320.990 377.080 2331.240 ;
        RECT 350.000 2309.140 377.080 2319.390 ;
        RECT 350.000 2295.610 377.080 2305.860 ;
        RECT 350.000 2283.760 377.080 2294.010 ;
        RECT 350.000 2271.360 377.080 2280.860 ;
        RECT 3511.960 2229.140 3530.000 2238.640 ;
        RECT 3511.960 2215.990 3530.000 2226.240 ;
        RECT 3511.960 2204.140 3530.000 2214.390 ;
        RECT 3511.960 2190.610 3530.000 2200.860 ;
        RECT 3511.960 2180.400 3530.000 2189.010 ;
        RECT 3511.960 2166.360 3530.000 2175.860 ;
        RECT 350.000 2129.140 367.080 2138.640 ;
        RECT 350.000 2115.990 367.080 2126.240 ;
        RECT 350.000 2104.140 367.080 2114.390 ;
        RECT 350.000 2090.610 367.080 2100.860 ;
        RECT 350.000 2078.760 367.080 2089.010 ;
        RECT 350.000 2066.360 367.080 2075.860 ;
        RECT 3511.960 2014.140 3530.000 2023.640 ;
        RECT 3511.960 2000.990 3530.000 2011.240 ;
        RECT 3511.960 1989.140 3530.000 1999.390 ;
        RECT 3511.960 1975.610 3530.000 1985.860 ;
        RECT 3511.960 1963.760 3530.000 1974.010 ;
        RECT 3511.960 1951.360 3530.000 1960.860 ;
        RECT 350.000 694.140 377.080 703.640 ;
        RECT 350.000 680.990 377.080 691.240 ;
        RECT 350.000 669.140 377.080 679.390 ;
        RECT 350.000 655.610 377.080 665.860 ;
        RECT 350.000 643.760 377.080 654.010 ;
        RECT 350.000 631.360 377.080 640.860 ;
        RECT 350.000 489.140 377.080 498.640 ;
        RECT 350.000 475.990 377.080 486.240 ;
        RECT 350.000 464.140 377.080 474.390 ;
        RECT 350.000 450.610 377.080 460.860 ;
        RECT 350.000 438.760 377.080 449.010 ;
        RECT 350.000 426.360 377.080 435.860 ;
        RECT 3276.360 372.440 3285.860 380.440 ;
        RECT 3288.760 372.440 3299.010 380.440 ;
        RECT 3300.610 372.440 3310.860 380.440 ;
        RECT 3314.140 372.440 3324.390 380.440 ;
        RECT 3325.990 372.440 3336.240 380.440 ;
        RECT 3339.140 372.440 3348.640 380.440 ;
        RECT 526.360 360.440 535.860 370.440 ;
        RECT 538.760 360.440 549.010 370.440 ;
        RECT 550.610 360.440 560.860 370.440 ;
        RECT 564.140 360.440 574.390 370.440 ;
        RECT 575.990 360.440 586.240 370.440 ;
        RECT 589.140 360.440 598.640 370.440 ;
        RECT 1351.360 360.440 1360.860 370.440 ;
        RECT 1363.760 360.440 1374.010 370.440 ;
        RECT 1375.610 360.440 1385.860 370.440 ;
        RECT 1389.140 360.440 1399.390 370.440 ;
        RECT 1400.990 360.440 1411.240 370.440 ;
        RECT 1414.140 360.440 1423.640 370.440 ;
        RECT 3001.360 360.440 3010.860 370.440 ;
        RECT 3013.760 360.440 3024.010 370.440 ;
        RECT 3025.610 360.440 3035.860 370.440 ;
        RECT 3039.140 360.440 3049.390 370.440 ;
        RECT 3050.990 360.440 3061.240 370.440 ;
        RECT 3064.140 360.440 3073.640 370.440 ;
      LAYER Via3 ;
        RECT 1896.705 4708.095 1896.985 4708.375 ;
        RECT 1897.415 4708.095 1897.695 4708.375 ;
        RECT 1898.125 4708.095 1898.405 4708.375 ;
        RECT 1898.835 4708.095 1899.115 4708.375 ;
        RECT 1899.545 4708.095 1899.825 4708.375 ;
        RECT 1896.705 4707.385 1896.985 4707.665 ;
        RECT 1897.415 4707.385 1897.695 4707.665 ;
        RECT 1898.125 4707.385 1898.405 4707.665 ;
        RECT 1898.835 4707.385 1899.115 4707.665 ;
        RECT 1899.545 4707.385 1899.825 4707.665 ;
        RECT 1896.705 4706.675 1896.985 4706.955 ;
        RECT 1897.415 4706.675 1897.695 4706.955 ;
        RECT 1898.125 4706.675 1898.405 4706.955 ;
        RECT 1898.835 4706.675 1899.115 4706.955 ;
        RECT 1899.545 4706.675 1899.825 4706.955 ;
        RECT 1896.705 4705.965 1896.985 4706.245 ;
        RECT 1897.415 4705.965 1897.695 4706.245 ;
        RECT 1898.125 4705.965 1898.405 4706.245 ;
        RECT 1898.835 4705.965 1899.115 4706.245 ;
        RECT 1899.545 4705.965 1899.825 4706.245 ;
        RECT 1896.705 4705.255 1896.985 4705.535 ;
        RECT 1897.415 4705.255 1897.695 4705.535 ;
        RECT 1898.125 4705.255 1898.405 4705.535 ;
        RECT 1898.835 4705.255 1899.115 4705.535 ;
        RECT 1899.545 4705.255 1899.825 4705.535 ;
        RECT 1896.705 4704.545 1896.985 4704.825 ;
        RECT 1897.415 4704.545 1897.695 4704.825 ;
        RECT 1898.125 4704.545 1898.405 4704.825 ;
        RECT 1898.835 4704.545 1899.115 4704.825 ;
        RECT 1899.545 4704.545 1899.825 4704.825 ;
        RECT 1896.705 4703.835 1896.985 4704.115 ;
        RECT 1897.415 4703.835 1897.695 4704.115 ;
        RECT 1898.125 4703.835 1898.405 4704.115 ;
        RECT 1898.835 4703.835 1899.115 4704.115 ;
        RECT 1899.545 4703.835 1899.825 4704.115 ;
        RECT 1896.705 4703.125 1896.985 4703.405 ;
        RECT 1897.415 4703.125 1897.695 4703.405 ;
        RECT 1898.125 4703.125 1898.405 4703.405 ;
        RECT 1898.835 4703.125 1899.115 4703.405 ;
        RECT 1899.545 4703.125 1899.825 4703.405 ;
        RECT 1896.705 4702.415 1896.985 4702.695 ;
        RECT 1897.415 4702.415 1897.695 4702.695 ;
        RECT 1898.125 4702.415 1898.405 4702.695 ;
        RECT 1898.835 4702.415 1899.115 4702.695 ;
        RECT 1899.545 4702.415 1899.825 4702.695 ;
        RECT 1896.705 4701.705 1896.985 4701.985 ;
        RECT 1897.415 4701.705 1897.695 4701.985 ;
        RECT 1898.125 4701.705 1898.405 4701.985 ;
        RECT 1898.835 4701.705 1899.115 4701.985 ;
        RECT 1899.545 4701.705 1899.825 4701.985 ;
        RECT 1896.705 4700.995 1896.985 4701.275 ;
        RECT 1897.415 4700.995 1897.695 4701.275 ;
        RECT 1898.125 4700.995 1898.405 4701.275 ;
        RECT 1898.835 4700.995 1899.115 4701.275 ;
        RECT 1899.545 4700.995 1899.825 4701.275 ;
        RECT 1896.705 4700.285 1896.985 4700.565 ;
        RECT 1897.415 4700.285 1897.695 4700.565 ;
        RECT 1898.125 4700.285 1898.405 4700.565 ;
        RECT 1898.835 4700.285 1899.115 4700.565 ;
        RECT 1899.545 4700.285 1899.825 4700.565 ;
        RECT 1896.705 4699.575 1896.985 4699.855 ;
        RECT 1897.415 4699.575 1897.695 4699.855 ;
        RECT 1898.125 4699.575 1898.405 4699.855 ;
        RECT 1898.835 4699.575 1899.115 4699.855 ;
        RECT 1899.545 4699.575 1899.825 4699.855 ;
        RECT 1896.705 4698.865 1896.985 4699.145 ;
        RECT 1897.415 4698.865 1897.695 4699.145 ;
        RECT 1898.125 4698.865 1898.405 4699.145 ;
        RECT 1898.835 4698.865 1899.115 4699.145 ;
        RECT 1899.545 4698.865 1899.825 4699.145 ;
        RECT 1909.145 4708.095 1909.425 4708.375 ;
        RECT 1909.855 4708.095 1910.135 4708.375 ;
        RECT 1910.565 4708.095 1910.845 4708.375 ;
        RECT 1911.275 4708.095 1911.555 4708.375 ;
        RECT 1911.985 4708.095 1912.265 4708.375 ;
        RECT 1912.695 4708.095 1912.975 4708.375 ;
        RECT 1913.405 4708.095 1913.685 4708.375 ;
        RECT 1914.115 4708.095 1914.395 4708.375 ;
        RECT 1914.825 4708.095 1915.105 4708.375 ;
        RECT 1915.535 4708.095 1915.815 4708.375 ;
        RECT 1916.245 4708.095 1916.525 4708.375 ;
        RECT 1916.955 4708.095 1917.235 4708.375 ;
        RECT 1917.665 4708.095 1917.945 4708.375 ;
        RECT 1918.375 4708.095 1918.655 4708.375 ;
        RECT 1909.145 4707.385 1909.425 4707.665 ;
        RECT 1909.855 4707.385 1910.135 4707.665 ;
        RECT 1910.565 4707.385 1910.845 4707.665 ;
        RECT 1911.275 4707.385 1911.555 4707.665 ;
        RECT 1911.985 4707.385 1912.265 4707.665 ;
        RECT 1912.695 4707.385 1912.975 4707.665 ;
        RECT 1913.405 4707.385 1913.685 4707.665 ;
        RECT 1914.115 4707.385 1914.395 4707.665 ;
        RECT 1914.825 4707.385 1915.105 4707.665 ;
        RECT 1915.535 4707.385 1915.815 4707.665 ;
        RECT 1916.245 4707.385 1916.525 4707.665 ;
        RECT 1916.955 4707.385 1917.235 4707.665 ;
        RECT 1917.665 4707.385 1917.945 4707.665 ;
        RECT 1918.375 4707.385 1918.655 4707.665 ;
        RECT 1909.145 4706.675 1909.425 4706.955 ;
        RECT 1909.855 4706.675 1910.135 4706.955 ;
        RECT 1910.565 4706.675 1910.845 4706.955 ;
        RECT 1911.275 4706.675 1911.555 4706.955 ;
        RECT 1911.985 4706.675 1912.265 4706.955 ;
        RECT 1912.695 4706.675 1912.975 4706.955 ;
        RECT 1913.405 4706.675 1913.685 4706.955 ;
        RECT 1914.115 4706.675 1914.395 4706.955 ;
        RECT 1914.825 4706.675 1915.105 4706.955 ;
        RECT 1915.535 4706.675 1915.815 4706.955 ;
        RECT 1916.245 4706.675 1916.525 4706.955 ;
        RECT 1916.955 4706.675 1917.235 4706.955 ;
        RECT 1917.665 4706.675 1917.945 4706.955 ;
        RECT 1918.375 4706.675 1918.655 4706.955 ;
        RECT 1909.145 4705.965 1909.425 4706.245 ;
        RECT 1909.855 4705.965 1910.135 4706.245 ;
        RECT 1910.565 4705.965 1910.845 4706.245 ;
        RECT 1911.275 4705.965 1911.555 4706.245 ;
        RECT 1911.985 4705.965 1912.265 4706.245 ;
        RECT 1912.695 4705.965 1912.975 4706.245 ;
        RECT 1913.405 4705.965 1913.685 4706.245 ;
        RECT 1914.115 4705.965 1914.395 4706.245 ;
        RECT 1914.825 4705.965 1915.105 4706.245 ;
        RECT 1915.535 4705.965 1915.815 4706.245 ;
        RECT 1916.245 4705.965 1916.525 4706.245 ;
        RECT 1916.955 4705.965 1917.235 4706.245 ;
        RECT 1917.665 4705.965 1917.945 4706.245 ;
        RECT 1918.375 4705.965 1918.655 4706.245 ;
        RECT 1909.145 4705.255 1909.425 4705.535 ;
        RECT 1909.855 4705.255 1910.135 4705.535 ;
        RECT 1910.565 4705.255 1910.845 4705.535 ;
        RECT 1911.275 4705.255 1911.555 4705.535 ;
        RECT 1911.985 4705.255 1912.265 4705.535 ;
        RECT 1912.695 4705.255 1912.975 4705.535 ;
        RECT 1913.405 4705.255 1913.685 4705.535 ;
        RECT 1914.115 4705.255 1914.395 4705.535 ;
        RECT 1914.825 4705.255 1915.105 4705.535 ;
        RECT 1915.535 4705.255 1915.815 4705.535 ;
        RECT 1916.245 4705.255 1916.525 4705.535 ;
        RECT 1916.955 4705.255 1917.235 4705.535 ;
        RECT 1917.665 4705.255 1917.945 4705.535 ;
        RECT 1918.375 4705.255 1918.655 4705.535 ;
        RECT 1909.145 4704.545 1909.425 4704.825 ;
        RECT 1909.855 4704.545 1910.135 4704.825 ;
        RECT 1910.565 4704.545 1910.845 4704.825 ;
        RECT 1911.275 4704.545 1911.555 4704.825 ;
        RECT 1911.985 4704.545 1912.265 4704.825 ;
        RECT 1912.695 4704.545 1912.975 4704.825 ;
        RECT 1913.405 4704.545 1913.685 4704.825 ;
        RECT 1914.115 4704.545 1914.395 4704.825 ;
        RECT 1914.825 4704.545 1915.105 4704.825 ;
        RECT 1915.535 4704.545 1915.815 4704.825 ;
        RECT 1916.245 4704.545 1916.525 4704.825 ;
        RECT 1916.955 4704.545 1917.235 4704.825 ;
        RECT 1917.665 4704.545 1917.945 4704.825 ;
        RECT 1918.375 4704.545 1918.655 4704.825 ;
        RECT 1909.145 4703.835 1909.425 4704.115 ;
        RECT 1909.855 4703.835 1910.135 4704.115 ;
        RECT 1910.565 4703.835 1910.845 4704.115 ;
        RECT 1911.275 4703.835 1911.555 4704.115 ;
        RECT 1911.985 4703.835 1912.265 4704.115 ;
        RECT 1912.695 4703.835 1912.975 4704.115 ;
        RECT 1913.405 4703.835 1913.685 4704.115 ;
        RECT 1914.115 4703.835 1914.395 4704.115 ;
        RECT 1914.825 4703.835 1915.105 4704.115 ;
        RECT 1915.535 4703.835 1915.815 4704.115 ;
        RECT 1916.245 4703.835 1916.525 4704.115 ;
        RECT 1916.955 4703.835 1917.235 4704.115 ;
        RECT 1917.665 4703.835 1917.945 4704.115 ;
        RECT 1918.375 4703.835 1918.655 4704.115 ;
        RECT 1909.145 4703.125 1909.425 4703.405 ;
        RECT 1909.855 4703.125 1910.135 4703.405 ;
        RECT 1910.565 4703.125 1910.845 4703.405 ;
        RECT 1911.275 4703.125 1911.555 4703.405 ;
        RECT 1911.985 4703.125 1912.265 4703.405 ;
        RECT 1912.695 4703.125 1912.975 4703.405 ;
        RECT 1913.405 4703.125 1913.685 4703.405 ;
        RECT 1914.115 4703.125 1914.395 4703.405 ;
        RECT 1914.825 4703.125 1915.105 4703.405 ;
        RECT 1915.535 4703.125 1915.815 4703.405 ;
        RECT 1916.245 4703.125 1916.525 4703.405 ;
        RECT 1916.955 4703.125 1917.235 4703.405 ;
        RECT 1917.665 4703.125 1917.945 4703.405 ;
        RECT 1918.375 4703.125 1918.655 4703.405 ;
        RECT 1909.145 4702.415 1909.425 4702.695 ;
        RECT 1909.855 4702.415 1910.135 4702.695 ;
        RECT 1910.565 4702.415 1910.845 4702.695 ;
        RECT 1911.275 4702.415 1911.555 4702.695 ;
        RECT 1911.985 4702.415 1912.265 4702.695 ;
        RECT 1912.695 4702.415 1912.975 4702.695 ;
        RECT 1913.405 4702.415 1913.685 4702.695 ;
        RECT 1914.115 4702.415 1914.395 4702.695 ;
        RECT 1914.825 4702.415 1915.105 4702.695 ;
        RECT 1915.535 4702.415 1915.815 4702.695 ;
        RECT 1916.245 4702.415 1916.525 4702.695 ;
        RECT 1916.955 4702.415 1917.235 4702.695 ;
        RECT 1917.665 4702.415 1917.945 4702.695 ;
        RECT 1918.375 4702.415 1918.655 4702.695 ;
        RECT 1909.145 4701.705 1909.425 4701.985 ;
        RECT 1909.855 4701.705 1910.135 4701.985 ;
        RECT 1910.565 4701.705 1910.845 4701.985 ;
        RECT 1911.275 4701.705 1911.555 4701.985 ;
        RECT 1911.985 4701.705 1912.265 4701.985 ;
        RECT 1912.695 4701.705 1912.975 4701.985 ;
        RECT 1913.405 4701.705 1913.685 4701.985 ;
        RECT 1914.115 4701.705 1914.395 4701.985 ;
        RECT 1914.825 4701.705 1915.105 4701.985 ;
        RECT 1915.535 4701.705 1915.815 4701.985 ;
        RECT 1916.245 4701.705 1916.525 4701.985 ;
        RECT 1916.955 4701.705 1917.235 4701.985 ;
        RECT 1917.665 4701.705 1917.945 4701.985 ;
        RECT 1918.375 4701.705 1918.655 4701.985 ;
        RECT 1909.145 4700.995 1909.425 4701.275 ;
        RECT 1909.855 4700.995 1910.135 4701.275 ;
        RECT 1910.565 4700.995 1910.845 4701.275 ;
        RECT 1911.275 4700.995 1911.555 4701.275 ;
        RECT 1911.985 4700.995 1912.265 4701.275 ;
        RECT 1912.695 4700.995 1912.975 4701.275 ;
        RECT 1913.405 4700.995 1913.685 4701.275 ;
        RECT 1914.115 4700.995 1914.395 4701.275 ;
        RECT 1914.825 4700.995 1915.105 4701.275 ;
        RECT 1915.535 4700.995 1915.815 4701.275 ;
        RECT 1916.245 4700.995 1916.525 4701.275 ;
        RECT 1916.955 4700.995 1917.235 4701.275 ;
        RECT 1917.665 4700.995 1917.945 4701.275 ;
        RECT 1918.375 4700.995 1918.655 4701.275 ;
        RECT 1909.145 4700.285 1909.425 4700.565 ;
        RECT 1909.855 4700.285 1910.135 4700.565 ;
        RECT 1910.565 4700.285 1910.845 4700.565 ;
        RECT 1911.275 4700.285 1911.555 4700.565 ;
        RECT 1911.985 4700.285 1912.265 4700.565 ;
        RECT 1912.695 4700.285 1912.975 4700.565 ;
        RECT 1913.405 4700.285 1913.685 4700.565 ;
        RECT 1914.115 4700.285 1914.395 4700.565 ;
        RECT 1914.825 4700.285 1915.105 4700.565 ;
        RECT 1915.535 4700.285 1915.815 4700.565 ;
        RECT 1916.245 4700.285 1916.525 4700.565 ;
        RECT 1916.955 4700.285 1917.235 4700.565 ;
        RECT 1917.665 4700.285 1917.945 4700.565 ;
        RECT 1918.375 4700.285 1918.655 4700.565 ;
        RECT 1909.145 4699.575 1909.425 4699.855 ;
        RECT 1909.855 4699.575 1910.135 4699.855 ;
        RECT 1910.565 4699.575 1910.845 4699.855 ;
        RECT 1911.275 4699.575 1911.555 4699.855 ;
        RECT 1911.985 4699.575 1912.265 4699.855 ;
        RECT 1912.695 4699.575 1912.975 4699.855 ;
        RECT 1913.405 4699.575 1913.685 4699.855 ;
        RECT 1914.115 4699.575 1914.395 4699.855 ;
        RECT 1914.825 4699.575 1915.105 4699.855 ;
        RECT 1915.535 4699.575 1915.815 4699.855 ;
        RECT 1916.245 4699.575 1916.525 4699.855 ;
        RECT 1916.955 4699.575 1917.235 4699.855 ;
        RECT 1917.665 4699.575 1917.945 4699.855 ;
        RECT 1918.375 4699.575 1918.655 4699.855 ;
        RECT 1909.145 4698.865 1909.425 4699.145 ;
        RECT 1909.855 4698.865 1910.135 4699.145 ;
        RECT 1910.565 4698.865 1910.845 4699.145 ;
        RECT 1911.275 4698.865 1911.555 4699.145 ;
        RECT 1911.985 4698.865 1912.265 4699.145 ;
        RECT 1912.695 4698.865 1912.975 4699.145 ;
        RECT 1913.405 4698.865 1913.685 4699.145 ;
        RECT 1914.115 4698.865 1914.395 4699.145 ;
        RECT 1914.825 4698.865 1915.105 4699.145 ;
        RECT 1915.535 4698.865 1915.815 4699.145 ;
        RECT 1916.245 4698.865 1916.525 4699.145 ;
        RECT 1916.955 4698.865 1917.235 4699.145 ;
        RECT 1917.665 4698.865 1917.945 4699.145 ;
        RECT 1918.375 4698.865 1918.655 4699.145 ;
        RECT 1920.995 4708.095 1921.275 4708.375 ;
        RECT 1921.705 4708.095 1921.985 4708.375 ;
        RECT 1922.415 4708.095 1922.695 4708.375 ;
        RECT 1923.125 4708.095 1923.405 4708.375 ;
        RECT 1923.835 4708.095 1924.115 4708.375 ;
        RECT 1924.545 4708.095 1924.825 4708.375 ;
        RECT 1925.255 4708.095 1925.535 4708.375 ;
        RECT 1925.965 4708.095 1926.245 4708.375 ;
        RECT 1926.675 4708.095 1926.955 4708.375 ;
        RECT 1927.385 4708.095 1927.665 4708.375 ;
        RECT 1928.095 4708.095 1928.375 4708.375 ;
        RECT 1928.805 4708.095 1929.085 4708.375 ;
        RECT 1929.515 4708.095 1929.795 4708.375 ;
        RECT 1930.225 4708.095 1930.505 4708.375 ;
        RECT 1920.995 4707.385 1921.275 4707.665 ;
        RECT 1921.705 4707.385 1921.985 4707.665 ;
        RECT 1922.415 4707.385 1922.695 4707.665 ;
        RECT 1923.125 4707.385 1923.405 4707.665 ;
        RECT 1923.835 4707.385 1924.115 4707.665 ;
        RECT 1924.545 4707.385 1924.825 4707.665 ;
        RECT 1925.255 4707.385 1925.535 4707.665 ;
        RECT 1925.965 4707.385 1926.245 4707.665 ;
        RECT 1926.675 4707.385 1926.955 4707.665 ;
        RECT 1927.385 4707.385 1927.665 4707.665 ;
        RECT 1928.095 4707.385 1928.375 4707.665 ;
        RECT 1928.805 4707.385 1929.085 4707.665 ;
        RECT 1929.515 4707.385 1929.795 4707.665 ;
        RECT 1930.225 4707.385 1930.505 4707.665 ;
        RECT 1920.995 4706.675 1921.275 4706.955 ;
        RECT 1921.705 4706.675 1921.985 4706.955 ;
        RECT 1922.415 4706.675 1922.695 4706.955 ;
        RECT 1923.125 4706.675 1923.405 4706.955 ;
        RECT 1923.835 4706.675 1924.115 4706.955 ;
        RECT 1924.545 4706.675 1924.825 4706.955 ;
        RECT 1925.255 4706.675 1925.535 4706.955 ;
        RECT 1925.965 4706.675 1926.245 4706.955 ;
        RECT 1926.675 4706.675 1926.955 4706.955 ;
        RECT 1927.385 4706.675 1927.665 4706.955 ;
        RECT 1928.095 4706.675 1928.375 4706.955 ;
        RECT 1928.805 4706.675 1929.085 4706.955 ;
        RECT 1929.515 4706.675 1929.795 4706.955 ;
        RECT 1930.225 4706.675 1930.505 4706.955 ;
        RECT 1920.995 4705.965 1921.275 4706.245 ;
        RECT 1921.705 4705.965 1921.985 4706.245 ;
        RECT 1922.415 4705.965 1922.695 4706.245 ;
        RECT 1923.125 4705.965 1923.405 4706.245 ;
        RECT 1923.835 4705.965 1924.115 4706.245 ;
        RECT 1924.545 4705.965 1924.825 4706.245 ;
        RECT 1925.255 4705.965 1925.535 4706.245 ;
        RECT 1925.965 4705.965 1926.245 4706.245 ;
        RECT 1926.675 4705.965 1926.955 4706.245 ;
        RECT 1927.385 4705.965 1927.665 4706.245 ;
        RECT 1928.095 4705.965 1928.375 4706.245 ;
        RECT 1928.805 4705.965 1929.085 4706.245 ;
        RECT 1929.515 4705.965 1929.795 4706.245 ;
        RECT 1930.225 4705.965 1930.505 4706.245 ;
        RECT 1920.995 4705.255 1921.275 4705.535 ;
        RECT 1921.705 4705.255 1921.985 4705.535 ;
        RECT 1922.415 4705.255 1922.695 4705.535 ;
        RECT 1923.125 4705.255 1923.405 4705.535 ;
        RECT 1923.835 4705.255 1924.115 4705.535 ;
        RECT 1924.545 4705.255 1924.825 4705.535 ;
        RECT 1925.255 4705.255 1925.535 4705.535 ;
        RECT 1925.965 4705.255 1926.245 4705.535 ;
        RECT 1926.675 4705.255 1926.955 4705.535 ;
        RECT 1927.385 4705.255 1927.665 4705.535 ;
        RECT 1928.095 4705.255 1928.375 4705.535 ;
        RECT 1928.805 4705.255 1929.085 4705.535 ;
        RECT 1929.515 4705.255 1929.795 4705.535 ;
        RECT 1930.225 4705.255 1930.505 4705.535 ;
        RECT 1920.995 4704.545 1921.275 4704.825 ;
        RECT 1921.705 4704.545 1921.985 4704.825 ;
        RECT 1922.415 4704.545 1922.695 4704.825 ;
        RECT 1923.125 4704.545 1923.405 4704.825 ;
        RECT 1923.835 4704.545 1924.115 4704.825 ;
        RECT 1924.545 4704.545 1924.825 4704.825 ;
        RECT 1925.255 4704.545 1925.535 4704.825 ;
        RECT 1925.965 4704.545 1926.245 4704.825 ;
        RECT 1926.675 4704.545 1926.955 4704.825 ;
        RECT 1927.385 4704.545 1927.665 4704.825 ;
        RECT 1928.095 4704.545 1928.375 4704.825 ;
        RECT 1928.805 4704.545 1929.085 4704.825 ;
        RECT 1929.515 4704.545 1929.795 4704.825 ;
        RECT 1930.225 4704.545 1930.505 4704.825 ;
        RECT 1920.995 4703.835 1921.275 4704.115 ;
        RECT 1921.705 4703.835 1921.985 4704.115 ;
        RECT 1922.415 4703.835 1922.695 4704.115 ;
        RECT 1923.125 4703.835 1923.405 4704.115 ;
        RECT 1923.835 4703.835 1924.115 4704.115 ;
        RECT 1924.545 4703.835 1924.825 4704.115 ;
        RECT 1925.255 4703.835 1925.535 4704.115 ;
        RECT 1925.965 4703.835 1926.245 4704.115 ;
        RECT 1926.675 4703.835 1926.955 4704.115 ;
        RECT 1927.385 4703.835 1927.665 4704.115 ;
        RECT 1928.095 4703.835 1928.375 4704.115 ;
        RECT 1928.805 4703.835 1929.085 4704.115 ;
        RECT 1929.515 4703.835 1929.795 4704.115 ;
        RECT 1930.225 4703.835 1930.505 4704.115 ;
        RECT 1920.995 4703.125 1921.275 4703.405 ;
        RECT 1921.705 4703.125 1921.985 4703.405 ;
        RECT 1922.415 4703.125 1922.695 4703.405 ;
        RECT 1923.125 4703.125 1923.405 4703.405 ;
        RECT 1923.835 4703.125 1924.115 4703.405 ;
        RECT 1924.545 4703.125 1924.825 4703.405 ;
        RECT 1925.255 4703.125 1925.535 4703.405 ;
        RECT 1925.965 4703.125 1926.245 4703.405 ;
        RECT 1926.675 4703.125 1926.955 4703.405 ;
        RECT 1927.385 4703.125 1927.665 4703.405 ;
        RECT 1928.095 4703.125 1928.375 4703.405 ;
        RECT 1928.805 4703.125 1929.085 4703.405 ;
        RECT 1929.515 4703.125 1929.795 4703.405 ;
        RECT 1930.225 4703.125 1930.505 4703.405 ;
        RECT 1920.995 4702.415 1921.275 4702.695 ;
        RECT 1921.705 4702.415 1921.985 4702.695 ;
        RECT 1922.415 4702.415 1922.695 4702.695 ;
        RECT 1923.125 4702.415 1923.405 4702.695 ;
        RECT 1923.835 4702.415 1924.115 4702.695 ;
        RECT 1924.545 4702.415 1924.825 4702.695 ;
        RECT 1925.255 4702.415 1925.535 4702.695 ;
        RECT 1925.965 4702.415 1926.245 4702.695 ;
        RECT 1926.675 4702.415 1926.955 4702.695 ;
        RECT 1927.385 4702.415 1927.665 4702.695 ;
        RECT 1928.095 4702.415 1928.375 4702.695 ;
        RECT 1928.805 4702.415 1929.085 4702.695 ;
        RECT 1929.515 4702.415 1929.795 4702.695 ;
        RECT 1930.225 4702.415 1930.505 4702.695 ;
        RECT 1920.995 4701.705 1921.275 4701.985 ;
        RECT 1921.705 4701.705 1921.985 4701.985 ;
        RECT 1922.415 4701.705 1922.695 4701.985 ;
        RECT 1923.125 4701.705 1923.405 4701.985 ;
        RECT 1923.835 4701.705 1924.115 4701.985 ;
        RECT 1924.545 4701.705 1924.825 4701.985 ;
        RECT 1925.255 4701.705 1925.535 4701.985 ;
        RECT 1925.965 4701.705 1926.245 4701.985 ;
        RECT 1926.675 4701.705 1926.955 4701.985 ;
        RECT 1927.385 4701.705 1927.665 4701.985 ;
        RECT 1928.095 4701.705 1928.375 4701.985 ;
        RECT 1928.805 4701.705 1929.085 4701.985 ;
        RECT 1929.515 4701.705 1929.795 4701.985 ;
        RECT 1930.225 4701.705 1930.505 4701.985 ;
        RECT 1920.995 4700.995 1921.275 4701.275 ;
        RECT 1921.705 4700.995 1921.985 4701.275 ;
        RECT 1922.415 4700.995 1922.695 4701.275 ;
        RECT 1923.125 4700.995 1923.405 4701.275 ;
        RECT 1923.835 4700.995 1924.115 4701.275 ;
        RECT 1924.545 4700.995 1924.825 4701.275 ;
        RECT 1925.255 4700.995 1925.535 4701.275 ;
        RECT 1925.965 4700.995 1926.245 4701.275 ;
        RECT 1926.675 4700.995 1926.955 4701.275 ;
        RECT 1927.385 4700.995 1927.665 4701.275 ;
        RECT 1928.095 4700.995 1928.375 4701.275 ;
        RECT 1928.805 4700.995 1929.085 4701.275 ;
        RECT 1929.515 4700.995 1929.795 4701.275 ;
        RECT 1930.225 4700.995 1930.505 4701.275 ;
        RECT 1920.995 4700.285 1921.275 4700.565 ;
        RECT 1921.705 4700.285 1921.985 4700.565 ;
        RECT 1922.415 4700.285 1922.695 4700.565 ;
        RECT 1923.125 4700.285 1923.405 4700.565 ;
        RECT 1923.835 4700.285 1924.115 4700.565 ;
        RECT 1924.545 4700.285 1924.825 4700.565 ;
        RECT 1925.255 4700.285 1925.535 4700.565 ;
        RECT 1925.965 4700.285 1926.245 4700.565 ;
        RECT 1926.675 4700.285 1926.955 4700.565 ;
        RECT 1927.385 4700.285 1927.665 4700.565 ;
        RECT 1928.095 4700.285 1928.375 4700.565 ;
        RECT 1928.805 4700.285 1929.085 4700.565 ;
        RECT 1929.515 4700.285 1929.795 4700.565 ;
        RECT 1930.225 4700.285 1930.505 4700.565 ;
        RECT 1920.995 4699.575 1921.275 4699.855 ;
        RECT 1921.705 4699.575 1921.985 4699.855 ;
        RECT 1922.415 4699.575 1922.695 4699.855 ;
        RECT 1923.125 4699.575 1923.405 4699.855 ;
        RECT 1923.835 4699.575 1924.115 4699.855 ;
        RECT 1924.545 4699.575 1924.825 4699.855 ;
        RECT 1925.255 4699.575 1925.535 4699.855 ;
        RECT 1925.965 4699.575 1926.245 4699.855 ;
        RECT 1926.675 4699.575 1926.955 4699.855 ;
        RECT 1927.385 4699.575 1927.665 4699.855 ;
        RECT 1928.095 4699.575 1928.375 4699.855 ;
        RECT 1928.805 4699.575 1929.085 4699.855 ;
        RECT 1929.515 4699.575 1929.795 4699.855 ;
        RECT 1930.225 4699.575 1930.505 4699.855 ;
        RECT 1920.995 4698.865 1921.275 4699.145 ;
        RECT 1921.705 4698.865 1921.985 4699.145 ;
        RECT 1922.415 4698.865 1922.695 4699.145 ;
        RECT 1923.125 4698.865 1923.405 4699.145 ;
        RECT 1923.835 4698.865 1924.115 4699.145 ;
        RECT 1924.545 4698.865 1924.825 4699.145 ;
        RECT 1925.255 4698.865 1925.535 4699.145 ;
        RECT 1925.965 4698.865 1926.245 4699.145 ;
        RECT 1926.675 4698.865 1926.955 4699.145 ;
        RECT 1927.385 4698.865 1927.665 4699.145 ;
        RECT 1928.095 4698.865 1928.375 4699.145 ;
        RECT 1928.805 4698.865 1929.085 4699.145 ;
        RECT 1929.515 4698.865 1929.795 4699.145 ;
        RECT 1930.225 4698.865 1930.505 4699.145 ;
        RECT 1934.525 4708.095 1934.805 4708.375 ;
        RECT 1935.235 4708.095 1935.515 4708.375 ;
        RECT 1935.945 4708.095 1936.225 4708.375 ;
        RECT 1936.655 4708.095 1936.935 4708.375 ;
        RECT 1937.365 4708.095 1937.645 4708.375 ;
        RECT 1938.075 4708.095 1938.355 4708.375 ;
        RECT 1938.785 4708.095 1939.065 4708.375 ;
        RECT 1939.495 4708.095 1939.775 4708.375 ;
        RECT 1940.205 4708.095 1940.485 4708.375 ;
        RECT 1940.915 4708.095 1941.195 4708.375 ;
        RECT 1941.625 4708.095 1941.905 4708.375 ;
        RECT 1942.335 4708.095 1942.615 4708.375 ;
        RECT 1943.045 4708.095 1943.325 4708.375 ;
        RECT 1943.755 4708.095 1944.035 4708.375 ;
        RECT 1934.525 4707.385 1934.805 4707.665 ;
        RECT 1935.235 4707.385 1935.515 4707.665 ;
        RECT 1935.945 4707.385 1936.225 4707.665 ;
        RECT 1936.655 4707.385 1936.935 4707.665 ;
        RECT 1937.365 4707.385 1937.645 4707.665 ;
        RECT 1938.075 4707.385 1938.355 4707.665 ;
        RECT 1938.785 4707.385 1939.065 4707.665 ;
        RECT 1939.495 4707.385 1939.775 4707.665 ;
        RECT 1940.205 4707.385 1940.485 4707.665 ;
        RECT 1940.915 4707.385 1941.195 4707.665 ;
        RECT 1941.625 4707.385 1941.905 4707.665 ;
        RECT 1942.335 4707.385 1942.615 4707.665 ;
        RECT 1943.045 4707.385 1943.325 4707.665 ;
        RECT 1943.755 4707.385 1944.035 4707.665 ;
        RECT 1934.525 4706.675 1934.805 4706.955 ;
        RECT 1935.235 4706.675 1935.515 4706.955 ;
        RECT 1935.945 4706.675 1936.225 4706.955 ;
        RECT 1936.655 4706.675 1936.935 4706.955 ;
        RECT 1937.365 4706.675 1937.645 4706.955 ;
        RECT 1938.075 4706.675 1938.355 4706.955 ;
        RECT 1938.785 4706.675 1939.065 4706.955 ;
        RECT 1939.495 4706.675 1939.775 4706.955 ;
        RECT 1940.205 4706.675 1940.485 4706.955 ;
        RECT 1940.915 4706.675 1941.195 4706.955 ;
        RECT 1941.625 4706.675 1941.905 4706.955 ;
        RECT 1942.335 4706.675 1942.615 4706.955 ;
        RECT 1943.045 4706.675 1943.325 4706.955 ;
        RECT 1943.755 4706.675 1944.035 4706.955 ;
        RECT 1934.525 4705.965 1934.805 4706.245 ;
        RECT 1935.235 4705.965 1935.515 4706.245 ;
        RECT 1935.945 4705.965 1936.225 4706.245 ;
        RECT 1936.655 4705.965 1936.935 4706.245 ;
        RECT 1937.365 4705.965 1937.645 4706.245 ;
        RECT 1938.075 4705.965 1938.355 4706.245 ;
        RECT 1938.785 4705.965 1939.065 4706.245 ;
        RECT 1939.495 4705.965 1939.775 4706.245 ;
        RECT 1940.205 4705.965 1940.485 4706.245 ;
        RECT 1940.915 4705.965 1941.195 4706.245 ;
        RECT 1941.625 4705.965 1941.905 4706.245 ;
        RECT 1942.335 4705.965 1942.615 4706.245 ;
        RECT 1943.045 4705.965 1943.325 4706.245 ;
        RECT 1943.755 4705.965 1944.035 4706.245 ;
        RECT 1934.525 4705.255 1934.805 4705.535 ;
        RECT 1935.235 4705.255 1935.515 4705.535 ;
        RECT 1935.945 4705.255 1936.225 4705.535 ;
        RECT 1936.655 4705.255 1936.935 4705.535 ;
        RECT 1937.365 4705.255 1937.645 4705.535 ;
        RECT 1938.075 4705.255 1938.355 4705.535 ;
        RECT 1938.785 4705.255 1939.065 4705.535 ;
        RECT 1939.495 4705.255 1939.775 4705.535 ;
        RECT 1940.205 4705.255 1940.485 4705.535 ;
        RECT 1940.915 4705.255 1941.195 4705.535 ;
        RECT 1941.625 4705.255 1941.905 4705.535 ;
        RECT 1942.335 4705.255 1942.615 4705.535 ;
        RECT 1943.045 4705.255 1943.325 4705.535 ;
        RECT 1943.755 4705.255 1944.035 4705.535 ;
        RECT 1934.525 4704.545 1934.805 4704.825 ;
        RECT 1935.235 4704.545 1935.515 4704.825 ;
        RECT 1935.945 4704.545 1936.225 4704.825 ;
        RECT 1936.655 4704.545 1936.935 4704.825 ;
        RECT 1937.365 4704.545 1937.645 4704.825 ;
        RECT 1938.075 4704.545 1938.355 4704.825 ;
        RECT 1938.785 4704.545 1939.065 4704.825 ;
        RECT 1939.495 4704.545 1939.775 4704.825 ;
        RECT 1940.205 4704.545 1940.485 4704.825 ;
        RECT 1940.915 4704.545 1941.195 4704.825 ;
        RECT 1941.625 4704.545 1941.905 4704.825 ;
        RECT 1942.335 4704.545 1942.615 4704.825 ;
        RECT 1943.045 4704.545 1943.325 4704.825 ;
        RECT 1943.755 4704.545 1944.035 4704.825 ;
        RECT 1934.525 4703.835 1934.805 4704.115 ;
        RECT 1935.235 4703.835 1935.515 4704.115 ;
        RECT 1935.945 4703.835 1936.225 4704.115 ;
        RECT 1936.655 4703.835 1936.935 4704.115 ;
        RECT 1937.365 4703.835 1937.645 4704.115 ;
        RECT 1938.075 4703.835 1938.355 4704.115 ;
        RECT 1938.785 4703.835 1939.065 4704.115 ;
        RECT 1939.495 4703.835 1939.775 4704.115 ;
        RECT 1940.205 4703.835 1940.485 4704.115 ;
        RECT 1940.915 4703.835 1941.195 4704.115 ;
        RECT 1941.625 4703.835 1941.905 4704.115 ;
        RECT 1942.335 4703.835 1942.615 4704.115 ;
        RECT 1943.045 4703.835 1943.325 4704.115 ;
        RECT 1943.755 4703.835 1944.035 4704.115 ;
        RECT 1934.525 4703.125 1934.805 4703.405 ;
        RECT 1935.235 4703.125 1935.515 4703.405 ;
        RECT 1935.945 4703.125 1936.225 4703.405 ;
        RECT 1936.655 4703.125 1936.935 4703.405 ;
        RECT 1937.365 4703.125 1937.645 4703.405 ;
        RECT 1938.075 4703.125 1938.355 4703.405 ;
        RECT 1938.785 4703.125 1939.065 4703.405 ;
        RECT 1939.495 4703.125 1939.775 4703.405 ;
        RECT 1940.205 4703.125 1940.485 4703.405 ;
        RECT 1940.915 4703.125 1941.195 4703.405 ;
        RECT 1941.625 4703.125 1941.905 4703.405 ;
        RECT 1942.335 4703.125 1942.615 4703.405 ;
        RECT 1943.045 4703.125 1943.325 4703.405 ;
        RECT 1943.755 4703.125 1944.035 4703.405 ;
        RECT 1934.525 4702.415 1934.805 4702.695 ;
        RECT 1935.235 4702.415 1935.515 4702.695 ;
        RECT 1935.945 4702.415 1936.225 4702.695 ;
        RECT 1936.655 4702.415 1936.935 4702.695 ;
        RECT 1937.365 4702.415 1937.645 4702.695 ;
        RECT 1938.075 4702.415 1938.355 4702.695 ;
        RECT 1938.785 4702.415 1939.065 4702.695 ;
        RECT 1939.495 4702.415 1939.775 4702.695 ;
        RECT 1940.205 4702.415 1940.485 4702.695 ;
        RECT 1940.915 4702.415 1941.195 4702.695 ;
        RECT 1941.625 4702.415 1941.905 4702.695 ;
        RECT 1942.335 4702.415 1942.615 4702.695 ;
        RECT 1943.045 4702.415 1943.325 4702.695 ;
        RECT 1943.755 4702.415 1944.035 4702.695 ;
        RECT 1934.525 4701.705 1934.805 4701.985 ;
        RECT 1935.235 4701.705 1935.515 4701.985 ;
        RECT 1935.945 4701.705 1936.225 4701.985 ;
        RECT 1936.655 4701.705 1936.935 4701.985 ;
        RECT 1937.365 4701.705 1937.645 4701.985 ;
        RECT 1938.075 4701.705 1938.355 4701.985 ;
        RECT 1938.785 4701.705 1939.065 4701.985 ;
        RECT 1939.495 4701.705 1939.775 4701.985 ;
        RECT 1940.205 4701.705 1940.485 4701.985 ;
        RECT 1940.915 4701.705 1941.195 4701.985 ;
        RECT 1941.625 4701.705 1941.905 4701.985 ;
        RECT 1942.335 4701.705 1942.615 4701.985 ;
        RECT 1943.045 4701.705 1943.325 4701.985 ;
        RECT 1943.755 4701.705 1944.035 4701.985 ;
        RECT 1934.525 4700.995 1934.805 4701.275 ;
        RECT 1935.235 4700.995 1935.515 4701.275 ;
        RECT 1935.945 4700.995 1936.225 4701.275 ;
        RECT 1936.655 4700.995 1936.935 4701.275 ;
        RECT 1937.365 4700.995 1937.645 4701.275 ;
        RECT 1938.075 4700.995 1938.355 4701.275 ;
        RECT 1938.785 4700.995 1939.065 4701.275 ;
        RECT 1939.495 4700.995 1939.775 4701.275 ;
        RECT 1940.205 4700.995 1940.485 4701.275 ;
        RECT 1940.915 4700.995 1941.195 4701.275 ;
        RECT 1941.625 4700.995 1941.905 4701.275 ;
        RECT 1942.335 4700.995 1942.615 4701.275 ;
        RECT 1943.045 4700.995 1943.325 4701.275 ;
        RECT 1943.755 4700.995 1944.035 4701.275 ;
        RECT 1934.525 4700.285 1934.805 4700.565 ;
        RECT 1935.235 4700.285 1935.515 4700.565 ;
        RECT 1935.945 4700.285 1936.225 4700.565 ;
        RECT 1936.655 4700.285 1936.935 4700.565 ;
        RECT 1937.365 4700.285 1937.645 4700.565 ;
        RECT 1938.075 4700.285 1938.355 4700.565 ;
        RECT 1938.785 4700.285 1939.065 4700.565 ;
        RECT 1939.495 4700.285 1939.775 4700.565 ;
        RECT 1940.205 4700.285 1940.485 4700.565 ;
        RECT 1940.915 4700.285 1941.195 4700.565 ;
        RECT 1941.625 4700.285 1941.905 4700.565 ;
        RECT 1942.335 4700.285 1942.615 4700.565 ;
        RECT 1943.045 4700.285 1943.325 4700.565 ;
        RECT 1943.755 4700.285 1944.035 4700.565 ;
        RECT 1934.525 4699.575 1934.805 4699.855 ;
        RECT 1935.235 4699.575 1935.515 4699.855 ;
        RECT 1935.945 4699.575 1936.225 4699.855 ;
        RECT 1936.655 4699.575 1936.935 4699.855 ;
        RECT 1937.365 4699.575 1937.645 4699.855 ;
        RECT 1938.075 4699.575 1938.355 4699.855 ;
        RECT 1938.785 4699.575 1939.065 4699.855 ;
        RECT 1939.495 4699.575 1939.775 4699.855 ;
        RECT 1940.205 4699.575 1940.485 4699.855 ;
        RECT 1940.915 4699.575 1941.195 4699.855 ;
        RECT 1941.625 4699.575 1941.905 4699.855 ;
        RECT 1942.335 4699.575 1942.615 4699.855 ;
        RECT 1943.045 4699.575 1943.325 4699.855 ;
        RECT 1943.755 4699.575 1944.035 4699.855 ;
        RECT 1934.525 4698.865 1934.805 4699.145 ;
        RECT 1935.235 4698.865 1935.515 4699.145 ;
        RECT 1935.945 4698.865 1936.225 4699.145 ;
        RECT 1936.655 4698.865 1936.935 4699.145 ;
        RECT 1937.365 4698.865 1937.645 4699.145 ;
        RECT 1938.075 4698.865 1938.355 4699.145 ;
        RECT 1938.785 4698.865 1939.065 4699.145 ;
        RECT 1939.495 4698.865 1939.775 4699.145 ;
        RECT 1940.205 4698.865 1940.485 4699.145 ;
        RECT 1940.915 4698.865 1941.195 4699.145 ;
        RECT 1941.625 4698.865 1941.905 4699.145 ;
        RECT 1942.335 4698.865 1942.615 4699.145 ;
        RECT 1943.045 4698.865 1943.325 4699.145 ;
        RECT 1943.755 4698.865 1944.035 4699.145 ;
        RECT 1946.375 4708.095 1946.655 4708.375 ;
        RECT 1947.085 4708.095 1947.365 4708.375 ;
        RECT 1947.795 4708.095 1948.075 4708.375 ;
        RECT 1948.505 4708.095 1948.785 4708.375 ;
        RECT 1949.215 4708.095 1949.495 4708.375 ;
        RECT 1949.925 4708.095 1950.205 4708.375 ;
        RECT 1950.635 4708.095 1950.915 4708.375 ;
        RECT 1951.345 4708.095 1951.625 4708.375 ;
        RECT 1952.055 4708.095 1952.335 4708.375 ;
        RECT 1952.765 4708.095 1953.045 4708.375 ;
        RECT 1953.475 4708.095 1953.755 4708.375 ;
        RECT 1954.185 4708.095 1954.465 4708.375 ;
        RECT 1954.895 4708.095 1955.175 4708.375 ;
        RECT 1955.605 4708.095 1955.885 4708.375 ;
        RECT 1946.375 4707.385 1946.655 4707.665 ;
        RECT 1947.085 4707.385 1947.365 4707.665 ;
        RECT 1947.795 4707.385 1948.075 4707.665 ;
        RECT 1948.505 4707.385 1948.785 4707.665 ;
        RECT 1949.215 4707.385 1949.495 4707.665 ;
        RECT 1949.925 4707.385 1950.205 4707.665 ;
        RECT 1950.635 4707.385 1950.915 4707.665 ;
        RECT 1951.345 4707.385 1951.625 4707.665 ;
        RECT 1952.055 4707.385 1952.335 4707.665 ;
        RECT 1952.765 4707.385 1953.045 4707.665 ;
        RECT 1953.475 4707.385 1953.755 4707.665 ;
        RECT 1954.185 4707.385 1954.465 4707.665 ;
        RECT 1954.895 4707.385 1955.175 4707.665 ;
        RECT 1955.605 4707.385 1955.885 4707.665 ;
        RECT 1946.375 4706.675 1946.655 4706.955 ;
        RECT 1947.085 4706.675 1947.365 4706.955 ;
        RECT 1947.795 4706.675 1948.075 4706.955 ;
        RECT 1948.505 4706.675 1948.785 4706.955 ;
        RECT 1949.215 4706.675 1949.495 4706.955 ;
        RECT 1949.925 4706.675 1950.205 4706.955 ;
        RECT 1950.635 4706.675 1950.915 4706.955 ;
        RECT 1951.345 4706.675 1951.625 4706.955 ;
        RECT 1952.055 4706.675 1952.335 4706.955 ;
        RECT 1952.765 4706.675 1953.045 4706.955 ;
        RECT 1953.475 4706.675 1953.755 4706.955 ;
        RECT 1954.185 4706.675 1954.465 4706.955 ;
        RECT 1954.895 4706.675 1955.175 4706.955 ;
        RECT 1955.605 4706.675 1955.885 4706.955 ;
        RECT 1946.375 4705.965 1946.655 4706.245 ;
        RECT 1947.085 4705.965 1947.365 4706.245 ;
        RECT 1947.795 4705.965 1948.075 4706.245 ;
        RECT 1948.505 4705.965 1948.785 4706.245 ;
        RECT 1949.215 4705.965 1949.495 4706.245 ;
        RECT 1949.925 4705.965 1950.205 4706.245 ;
        RECT 1950.635 4705.965 1950.915 4706.245 ;
        RECT 1951.345 4705.965 1951.625 4706.245 ;
        RECT 1952.055 4705.965 1952.335 4706.245 ;
        RECT 1952.765 4705.965 1953.045 4706.245 ;
        RECT 1953.475 4705.965 1953.755 4706.245 ;
        RECT 1954.185 4705.965 1954.465 4706.245 ;
        RECT 1954.895 4705.965 1955.175 4706.245 ;
        RECT 1955.605 4705.965 1955.885 4706.245 ;
        RECT 1946.375 4705.255 1946.655 4705.535 ;
        RECT 1947.085 4705.255 1947.365 4705.535 ;
        RECT 1947.795 4705.255 1948.075 4705.535 ;
        RECT 1948.505 4705.255 1948.785 4705.535 ;
        RECT 1949.215 4705.255 1949.495 4705.535 ;
        RECT 1949.925 4705.255 1950.205 4705.535 ;
        RECT 1950.635 4705.255 1950.915 4705.535 ;
        RECT 1951.345 4705.255 1951.625 4705.535 ;
        RECT 1952.055 4705.255 1952.335 4705.535 ;
        RECT 1952.765 4705.255 1953.045 4705.535 ;
        RECT 1953.475 4705.255 1953.755 4705.535 ;
        RECT 1954.185 4705.255 1954.465 4705.535 ;
        RECT 1954.895 4705.255 1955.175 4705.535 ;
        RECT 1955.605 4705.255 1955.885 4705.535 ;
        RECT 1946.375 4704.545 1946.655 4704.825 ;
        RECT 1947.085 4704.545 1947.365 4704.825 ;
        RECT 1947.795 4704.545 1948.075 4704.825 ;
        RECT 1948.505 4704.545 1948.785 4704.825 ;
        RECT 1949.215 4704.545 1949.495 4704.825 ;
        RECT 1949.925 4704.545 1950.205 4704.825 ;
        RECT 1950.635 4704.545 1950.915 4704.825 ;
        RECT 1951.345 4704.545 1951.625 4704.825 ;
        RECT 1952.055 4704.545 1952.335 4704.825 ;
        RECT 1952.765 4704.545 1953.045 4704.825 ;
        RECT 1953.475 4704.545 1953.755 4704.825 ;
        RECT 1954.185 4704.545 1954.465 4704.825 ;
        RECT 1954.895 4704.545 1955.175 4704.825 ;
        RECT 1955.605 4704.545 1955.885 4704.825 ;
        RECT 1946.375 4703.835 1946.655 4704.115 ;
        RECT 1947.085 4703.835 1947.365 4704.115 ;
        RECT 1947.795 4703.835 1948.075 4704.115 ;
        RECT 1948.505 4703.835 1948.785 4704.115 ;
        RECT 1949.215 4703.835 1949.495 4704.115 ;
        RECT 1949.925 4703.835 1950.205 4704.115 ;
        RECT 1950.635 4703.835 1950.915 4704.115 ;
        RECT 1951.345 4703.835 1951.625 4704.115 ;
        RECT 1952.055 4703.835 1952.335 4704.115 ;
        RECT 1952.765 4703.835 1953.045 4704.115 ;
        RECT 1953.475 4703.835 1953.755 4704.115 ;
        RECT 1954.185 4703.835 1954.465 4704.115 ;
        RECT 1954.895 4703.835 1955.175 4704.115 ;
        RECT 1955.605 4703.835 1955.885 4704.115 ;
        RECT 1946.375 4703.125 1946.655 4703.405 ;
        RECT 1947.085 4703.125 1947.365 4703.405 ;
        RECT 1947.795 4703.125 1948.075 4703.405 ;
        RECT 1948.505 4703.125 1948.785 4703.405 ;
        RECT 1949.215 4703.125 1949.495 4703.405 ;
        RECT 1949.925 4703.125 1950.205 4703.405 ;
        RECT 1950.635 4703.125 1950.915 4703.405 ;
        RECT 1951.345 4703.125 1951.625 4703.405 ;
        RECT 1952.055 4703.125 1952.335 4703.405 ;
        RECT 1952.765 4703.125 1953.045 4703.405 ;
        RECT 1953.475 4703.125 1953.755 4703.405 ;
        RECT 1954.185 4703.125 1954.465 4703.405 ;
        RECT 1954.895 4703.125 1955.175 4703.405 ;
        RECT 1955.605 4703.125 1955.885 4703.405 ;
        RECT 1946.375 4702.415 1946.655 4702.695 ;
        RECT 1947.085 4702.415 1947.365 4702.695 ;
        RECT 1947.795 4702.415 1948.075 4702.695 ;
        RECT 1948.505 4702.415 1948.785 4702.695 ;
        RECT 1949.215 4702.415 1949.495 4702.695 ;
        RECT 1949.925 4702.415 1950.205 4702.695 ;
        RECT 1950.635 4702.415 1950.915 4702.695 ;
        RECT 1951.345 4702.415 1951.625 4702.695 ;
        RECT 1952.055 4702.415 1952.335 4702.695 ;
        RECT 1952.765 4702.415 1953.045 4702.695 ;
        RECT 1953.475 4702.415 1953.755 4702.695 ;
        RECT 1954.185 4702.415 1954.465 4702.695 ;
        RECT 1954.895 4702.415 1955.175 4702.695 ;
        RECT 1955.605 4702.415 1955.885 4702.695 ;
        RECT 1946.375 4701.705 1946.655 4701.985 ;
        RECT 1947.085 4701.705 1947.365 4701.985 ;
        RECT 1947.795 4701.705 1948.075 4701.985 ;
        RECT 1948.505 4701.705 1948.785 4701.985 ;
        RECT 1949.215 4701.705 1949.495 4701.985 ;
        RECT 1949.925 4701.705 1950.205 4701.985 ;
        RECT 1950.635 4701.705 1950.915 4701.985 ;
        RECT 1951.345 4701.705 1951.625 4701.985 ;
        RECT 1952.055 4701.705 1952.335 4701.985 ;
        RECT 1952.765 4701.705 1953.045 4701.985 ;
        RECT 1953.475 4701.705 1953.755 4701.985 ;
        RECT 1954.185 4701.705 1954.465 4701.985 ;
        RECT 1954.895 4701.705 1955.175 4701.985 ;
        RECT 1955.605 4701.705 1955.885 4701.985 ;
        RECT 1946.375 4700.995 1946.655 4701.275 ;
        RECT 1947.085 4700.995 1947.365 4701.275 ;
        RECT 1947.795 4700.995 1948.075 4701.275 ;
        RECT 1948.505 4700.995 1948.785 4701.275 ;
        RECT 1949.215 4700.995 1949.495 4701.275 ;
        RECT 1949.925 4700.995 1950.205 4701.275 ;
        RECT 1950.635 4700.995 1950.915 4701.275 ;
        RECT 1951.345 4700.995 1951.625 4701.275 ;
        RECT 1952.055 4700.995 1952.335 4701.275 ;
        RECT 1952.765 4700.995 1953.045 4701.275 ;
        RECT 1953.475 4700.995 1953.755 4701.275 ;
        RECT 1954.185 4700.995 1954.465 4701.275 ;
        RECT 1954.895 4700.995 1955.175 4701.275 ;
        RECT 1955.605 4700.995 1955.885 4701.275 ;
        RECT 1946.375 4700.285 1946.655 4700.565 ;
        RECT 1947.085 4700.285 1947.365 4700.565 ;
        RECT 1947.795 4700.285 1948.075 4700.565 ;
        RECT 1948.505 4700.285 1948.785 4700.565 ;
        RECT 1949.215 4700.285 1949.495 4700.565 ;
        RECT 1949.925 4700.285 1950.205 4700.565 ;
        RECT 1950.635 4700.285 1950.915 4700.565 ;
        RECT 1951.345 4700.285 1951.625 4700.565 ;
        RECT 1952.055 4700.285 1952.335 4700.565 ;
        RECT 1952.765 4700.285 1953.045 4700.565 ;
        RECT 1953.475 4700.285 1953.755 4700.565 ;
        RECT 1954.185 4700.285 1954.465 4700.565 ;
        RECT 1954.895 4700.285 1955.175 4700.565 ;
        RECT 1955.605 4700.285 1955.885 4700.565 ;
        RECT 1946.375 4699.575 1946.655 4699.855 ;
        RECT 1947.085 4699.575 1947.365 4699.855 ;
        RECT 1947.795 4699.575 1948.075 4699.855 ;
        RECT 1948.505 4699.575 1948.785 4699.855 ;
        RECT 1949.215 4699.575 1949.495 4699.855 ;
        RECT 1949.925 4699.575 1950.205 4699.855 ;
        RECT 1950.635 4699.575 1950.915 4699.855 ;
        RECT 1951.345 4699.575 1951.625 4699.855 ;
        RECT 1952.055 4699.575 1952.335 4699.855 ;
        RECT 1952.765 4699.575 1953.045 4699.855 ;
        RECT 1953.475 4699.575 1953.755 4699.855 ;
        RECT 1954.185 4699.575 1954.465 4699.855 ;
        RECT 1954.895 4699.575 1955.175 4699.855 ;
        RECT 1955.605 4699.575 1955.885 4699.855 ;
        RECT 1946.375 4698.865 1946.655 4699.145 ;
        RECT 1947.085 4698.865 1947.365 4699.145 ;
        RECT 1947.795 4698.865 1948.075 4699.145 ;
        RECT 1948.505 4698.865 1948.785 4699.145 ;
        RECT 1949.215 4698.865 1949.495 4699.145 ;
        RECT 1949.925 4698.865 1950.205 4699.145 ;
        RECT 1950.635 4698.865 1950.915 4699.145 ;
        RECT 1951.345 4698.865 1951.625 4699.145 ;
        RECT 1952.055 4698.865 1952.335 4699.145 ;
        RECT 1952.765 4698.865 1953.045 4699.145 ;
        RECT 1953.475 4698.865 1953.755 4699.145 ;
        RECT 1954.185 4698.865 1954.465 4699.145 ;
        RECT 1954.895 4698.865 1955.175 4699.145 ;
        RECT 1955.605 4698.865 1955.885 4699.145 ;
        RECT 1959.485 4708.095 1959.765 4708.375 ;
        RECT 1960.195 4708.095 1960.475 4708.375 ;
        RECT 1960.905 4708.095 1961.185 4708.375 ;
        RECT 1961.615 4708.095 1961.895 4708.375 ;
        RECT 1962.325 4708.095 1962.605 4708.375 ;
        RECT 1963.035 4708.095 1963.315 4708.375 ;
        RECT 1963.745 4708.095 1964.025 4708.375 ;
        RECT 1964.455 4708.095 1964.735 4708.375 ;
        RECT 1965.165 4708.095 1965.445 4708.375 ;
        RECT 1965.875 4708.095 1966.155 4708.375 ;
        RECT 1966.585 4708.095 1966.865 4708.375 ;
        RECT 1967.295 4708.095 1967.575 4708.375 ;
        RECT 1968.005 4708.095 1968.285 4708.375 ;
        RECT 1959.485 4707.385 1959.765 4707.665 ;
        RECT 1960.195 4707.385 1960.475 4707.665 ;
        RECT 1960.905 4707.385 1961.185 4707.665 ;
        RECT 1961.615 4707.385 1961.895 4707.665 ;
        RECT 1962.325 4707.385 1962.605 4707.665 ;
        RECT 1963.035 4707.385 1963.315 4707.665 ;
        RECT 1963.745 4707.385 1964.025 4707.665 ;
        RECT 1964.455 4707.385 1964.735 4707.665 ;
        RECT 1965.165 4707.385 1965.445 4707.665 ;
        RECT 1965.875 4707.385 1966.155 4707.665 ;
        RECT 1966.585 4707.385 1966.865 4707.665 ;
        RECT 1967.295 4707.385 1967.575 4707.665 ;
        RECT 1968.005 4707.385 1968.285 4707.665 ;
        RECT 1959.485 4706.675 1959.765 4706.955 ;
        RECT 1960.195 4706.675 1960.475 4706.955 ;
        RECT 1960.905 4706.675 1961.185 4706.955 ;
        RECT 1961.615 4706.675 1961.895 4706.955 ;
        RECT 1962.325 4706.675 1962.605 4706.955 ;
        RECT 1963.035 4706.675 1963.315 4706.955 ;
        RECT 1963.745 4706.675 1964.025 4706.955 ;
        RECT 1964.455 4706.675 1964.735 4706.955 ;
        RECT 1965.165 4706.675 1965.445 4706.955 ;
        RECT 1965.875 4706.675 1966.155 4706.955 ;
        RECT 1966.585 4706.675 1966.865 4706.955 ;
        RECT 1967.295 4706.675 1967.575 4706.955 ;
        RECT 1968.005 4706.675 1968.285 4706.955 ;
        RECT 1959.485 4705.965 1959.765 4706.245 ;
        RECT 1960.195 4705.965 1960.475 4706.245 ;
        RECT 1960.905 4705.965 1961.185 4706.245 ;
        RECT 1961.615 4705.965 1961.895 4706.245 ;
        RECT 1962.325 4705.965 1962.605 4706.245 ;
        RECT 1963.035 4705.965 1963.315 4706.245 ;
        RECT 1963.745 4705.965 1964.025 4706.245 ;
        RECT 1964.455 4705.965 1964.735 4706.245 ;
        RECT 1965.165 4705.965 1965.445 4706.245 ;
        RECT 1965.875 4705.965 1966.155 4706.245 ;
        RECT 1966.585 4705.965 1966.865 4706.245 ;
        RECT 1967.295 4705.965 1967.575 4706.245 ;
        RECT 1968.005 4705.965 1968.285 4706.245 ;
        RECT 1959.485 4705.255 1959.765 4705.535 ;
        RECT 1960.195 4705.255 1960.475 4705.535 ;
        RECT 1960.905 4705.255 1961.185 4705.535 ;
        RECT 1961.615 4705.255 1961.895 4705.535 ;
        RECT 1962.325 4705.255 1962.605 4705.535 ;
        RECT 1963.035 4705.255 1963.315 4705.535 ;
        RECT 1963.745 4705.255 1964.025 4705.535 ;
        RECT 1964.455 4705.255 1964.735 4705.535 ;
        RECT 1965.165 4705.255 1965.445 4705.535 ;
        RECT 1965.875 4705.255 1966.155 4705.535 ;
        RECT 1966.585 4705.255 1966.865 4705.535 ;
        RECT 1967.295 4705.255 1967.575 4705.535 ;
        RECT 1968.005 4705.255 1968.285 4705.535 ;
        RECT 1959.485 4704.545 1959.765 4704.825 ;
        RECT 1960.195 4704.545 1960.475 4704.825 ;
        RECT 1960.905 4704.545 1961.185 4704.825 ;
        RECT 1961.615 4704.545 1961.895 4704.825 ;
        RECT 1962.325 4704.545 1962.605 4704.825 ;
        RECT 1963.035 4704.545 1963.315 4704.825 ;
        RECT 1963.745 4704.545 1964.025 4704.825 ;
        RECT 1964.455 4704.545 1964.735 4704.825 ;
        RECT 1965.165 4704.545 1965.445 4704.825 ;
        RECT 1965.875 4704.545 1966.155 4704.825 ;
        RECT 1966.585 4704.545 1966.865 4704.825 ;
        RECT 1967.295 4704.545 1967.575 4704.825 ;
        RECT 1968.005 4704.545 1968.285 4704.825 ;
        RECT 1959.485 4703.835 1959.765 4704.115 ;
        RECT 1960.195 4703.835 1960.475 4704.115 ;
        RECT 1960.905 4703.835 1961.185 4704.115 ;
        RECT 1961.615 4703.835 1961.895 4704.115 ;
        RECT 1962.325 4703.835 1962.605 4704.115 ;
        RECT 1963.035 4703.835 1963.315 4704.115 ;
        RECT 1963.745 4703.835 1964.025 4704.115 ;
        RECT 1964.455 4703.835 1964.735 4704.115 ;
        RECT 1965.165 4703.835 1965.445 4704.115 ;
        RECT 1965.875 4703.835 1966.155 4704.115 ;
        RECT 1966.585 4703.835 1966.865 4704.115 ;
        RECT 1967.295 4703.835 1967.575 4704.115 ;
        RECT 1968.005 4703.835 1968.285 4704.115 ;
        RECT 1959.485 4703.125 1959.765 4703.405 ;
        RECT 1960.195 4703.125 1960.475 4703.405 ;
        RECT 1960.905 4703.125 1961.185 4703.405 ;
        RECT 1961.615 4703.125 1961.895 4703.405 ;
        RECT 1962.325 4703.125 1962.605 4703.405 ;
        RECT 1963.035 4703.125 1963.315 4703.405 ;
        RECT 1963.745 4703.125 1964.025 4703.405 ;
        RECT 1964.455 4703.125 1964.735 4703.405 ;
        RECT 1965.165 4703.125 1965.445 4703.405 ;
        RECT 1965.875 4703.125 1966.155 4703.405 ;
        RECT 1966.585 4703.125 1966.865 4703.405 ;
        RECT 1967.295 4703.125 1967.575 4703.405 ;
        RECT 1968.005 4703.125 1968.285 4703.405 ;
        RECT 1959.485 4702.415 1959.765 4702.695 ;
        RECT 1960.195 4702.415 1960.475 4702.695 ;
        RECT 1960.905 4702.415 1961.185 4702.695 ;
        RECT 1961.615 4702.415 1961.895 4702.695 ;
        RECT 1962.325 4702.415 1962.605 4702.695 ;
        RECT 1963.035 4702.415 1963.315 4702.695 ;
        RECT 1963.745 4702.415 1964.025 4702.695 ;
        RECT 1964.455 4702.415 1964.735 4702.695 ;
        RECT 1965.165 4702.415 1965.445 4702.695 ;
        RECT 1965.875 4702.415 1966.155 4702.695 ;
        RECT 1966.585 4702.415 1966.865 4702.695 ;
        RECT 1967.295 4702.415 1967.575 4702.695 ;
        RECT 1968.005 4702.415 1968.285 4702.695 ;
        RECT 1959.485 4701.705 1959.765 4701.985 ;
        RECT 1960.195 4701.705 1960.475 4701.985 ;
        RECT 1960.905 4701.705 1961.185 4701.985 ;
        RECT 1961.615 4701.705 1961.895 4701.985 ;
        RECT 1962.325 4701.705 1962.605 4701.985 ;
        RECT 1963.035 4701.705 1963.315 4701.985 ;
        RECT 1963.745 4701.705 1964.025 4701.985 ;
        RECT 1964.455 4701.705 1964.735 4701.985 ;
        RECT 1965.165 4701.705 1965.445 4701.985 ;
        RECT 1965.875 4701.705 1966.155 4701.985 ;
        RECT 1966.585 4701.705 1966.865 4701.985 ;
        RECT 1967.295 4701.705 1967.575 4701.985 ;
        RECT 1968.005 4701.705 1968.285 4701.985 ;
        RECT 1959.485 4700.995 1959.765 4701.275 ;
        RECT 1960.195 4700.995 1960.475 4701.275 ;
        RECT 1960.905 4700.995 1961.185 4701.275 ;
        RECT 1961.615 4700.995 1961.895 4701.275 ;
        RECT 1962.325 4700.995 1962.605 4701.275 ;
        RECT 1963.035 4700.995 1963.315 4701.275 ;
        RECT 1963.745 4700.995 1964.025 4701.275 ;
        RECT 1964.455 4700.995 1964.735 4701.275 ;
        RECT 1965.165 4700.995 1965.445 4701.275 ;
        RECT 1965.875 4700.995 1966.155 4701.275 ;
        RECT 1966.585 4700.995 1966.865 4701.275 ;
        RECT 1967.295 4700.995 1967.575 4701.275 ;
        RECT 1968.005 4700.995 1968.285 4701.275 ;
        RECT 1959.485 4700.285 1959.765 4700.565 ;
        RECT 1960.195 4700.285 1960.475 4700.565 ;
        RECT 1960.905 4700.285 1961.185 4700.565 ;
        RECT 1961.615 4700.285 1961.895 4700.565 ;
        RECT 1962.325 4700.285 1962.605 4700.565 ;
        RECT 1963.035 4700.285 1963.315 4700.565 ;
        RECT 1963.745 4700.285 1964.025 4700.565 ;
        RECT 1964.455 4700.285 1964.735 4700.565 ;
        RECT 1965.165 4700.285 1965.445 4700.565 ;
        RECT 1965.875 4700.285 1966.155 4700.565 ;
        RECT 1966.585 4700.285 1966.865 4700.565 ;
        RECT 1967.295 4700.285 1967.575 4700.565 ;
        RECT 1968.005 4700.285 1968.285 4700.565 ;
        RECT 1959.485 4699.575 1959.765 4699.855 ;
        RECT 1960.195 4699.575 1960.475 4699.855 ;
        RECT 1960.905 4699.575 1961.185 4699.855 ;
        RECT 1961.615 4699.575 1961.895 4699.855 ;
        RECT 1962.325 4699.575 1962.605 4699.855 ;
        RECT 1963.035 4699.575 1963.315 4699.855 ;
        RECT 1963.745 4699.575 1964.025 4699.855 ;
        RECT 1964.455 4699.575 1964.735 4699.855 ;
        RECT 1965.165 4699.575 1965.445 4699.855 ;
        RECT 1965.875 4699.575 1966.155 4699.855 ;
        RECT 1966.585 4699.575 1966.865 4699.855 ;
        RECT 1967.295 4699.575 1967.575 4699.855 ;
        RECT 1968.005 4699.575 1968.285 4699.855 ;
        RECT 1959.485 4698.865 1959.765 4699.145 ;
        RECT 1960.195 4698.865 1960.475 4699.145 ;
        RECT 1960.905 4698.865 1961.185 4699.145 ;
        RECT 1961.615 4698.865 1961.895 4699.145 ;
        RECT 1962.325 4698.865 1962.605 4699.145 ;
        RECT 1963.035 4698.865 1963.315 4699.145 ;
        RECT 1963.745 4698.865 1964.025 4699.145 ;
        RECT 1964.455 4698.865 1964.735 4699.145 ;
        RECT 1965.165 4698.865 1965.445 4699.145 ;
        RECT 1965.875 4698.865 1966.155 4699.145 ;
        RECT 1966.585 4698.865 1966.865 4699.145 ;
        RECT 1967.295 4698.865 1967.575 4699.145 ;
        RECT 1968.005 4698.865 1968.285 4699.145 ;
        RECT 2996.705 4708.095 2996.985 4708.375 ;
        RECT 2997.415 4708.095 2997.695 4708.375 ;
        RECT 2998.125 4708.095 2998.405 4708.375 ;
        RECT 2998.835 4708.095 2999.115 4708.375 ;
        RECT 2999.545 4708.095 2999.825 4708.375 ;
        RECT 3000.255 4708.095 3000.535 4708.375 ;
        RECT 3000.965 4708.095 3001.245 4708.375 ;
        RECT 3001.675 4708.095 3001.955 4708.375 ;
        RECT 3002.385 4708.095 3002.665 4708.375 ;
        RECT 3003.095 4708.095 3003.375 4708.375 ;
        RECT 3003.805 4708.095 3004.085 4708.375 ;
        RECT 3004.515 4708.095 3004.795 4708.375 ;
        RECT 3005.225 4708.095 3005.505 4708.375 ;
        RECT 2996.705 4707.385 2996.985 4707.665 ;
        RECT 2997.415 4707.385 2997.695 4707.665 ;
        RECT 2998.125 4707.385 2998.405 4707.665 ;
        RECT 2998.835 4707.385 2999.115 4707.665 ;
        RECT 2999.545 4707.385 2999.825 4707.665 ;
        RECT 3000.255 4707.385 3000.535 4707.665 ;
        RECT 3000.965 4707.385 3001.245 4707.665 ;
        RECT 3001.675 4707.385 3001.955 4707.665 ;
        RECT 3002.385 4707.385 3002.665 4707.665 ;
        RECT 3003.095 4707.385 3003.375 4707.665 ;
        RECT 3003.805 4707.385 3004.085 4707.665 ;
        RECT 3004.515 4707.385 3004.795 4707.665 ;
        RECT 3005.225 4707.385 3005.505 4707.665 ;
        RECT 2996.705 4706.675 2996.985 4706.955 ;
        RECT 2997.415 4706.675 2997.695 4706.955 ;
        RECT 2998.125 4706.675 2998.405 4706.955 ;
        RECT 2998.835 4706.675 2999.115 4706.955 ;
        RECT 2999.545 4706.675 2999.825 4706.955 ;
        RECT 3000.255 4706.675 3000.535 4706.955 ;
        RECT 3000.965 4706.675 3001.245 4706.955 ;
        RECT 3001.675 4706.675 3001.955 4706.955 ;
        RECT 3002.385 4706.675 3002.665 4706.955 ;
        RECT 3003.095 4706.675 3003.375 4706.955 ;
        RECT 3003.805 4706.675 3004.085 4706.955 ;
        RECT 3004.515 4706.675 3004.795 4706.955 ;
        RECT 3005.225 4706.675 3005.505 4706.955 ;
        RECT 2996.705 4705.965 2996.985 4706.245 ;
        RECT 2997.415 4705.965 2997.695 4706.245 ;
        RECT 2998.125 4705.965 2998.405 4706.245 ;
        RECT 2998.835 4705.965 2999.115 4706.245 ;
        RECT 2999.545 4705.965 2999.825 4706.245 ;
        RECT 3000.255 4705.965 3000.535 4706.245 ;
        RECT 3000.965 4705.965 3001.245 4706.245 ;
        RECT 3001.675 4705.965 3001.955 4706.245 ;
        RECT 3002.385 4705.965 3002.665 4706.245 ;
        RECT 3003.095 4705.965 3003.375 4706.245 ;
        RECT 3003.805 4705.965 3004.085 4706.245 ;
        RECT 3004.515 4705.965 3004.795 4706.245 ;
        RECT 3005.225 4705.965 3005.505 4706.245 ;
        RECT 2996.705 4705.255 2996.985 4705.535 ;
        RECT 2997.415 4705.255 2997.695 4705.535 ;
        RECT 2998.125 4705.255 2998.405 4705.535 ;
        RECT 2998.835 4705.255 2999.115 4705.535 ;
        RECT 2999.545 4705.255 2999.825 4705.535 ;
        RECT 3000.255 4705.255 3000.535 4705.535 ;
        RECT 3000.965 4705.255 3001.245 4705.535 ;
        RECT 3001.675 4705.255 3001.955 4705.535 ;
        RECT 3002.385 4705.255 3002.665 4705.535 ;
        RECT 3003.095 4705.255 3003.375 4705.535 ;
        RECT 3003.805 4705.255 3004.085 4705.535 ;
        RECT 3004.515 4705.255 3004.795 4705.535 ;
        RECT 3005.225 4705.255 3005.505 4705.535 ;
        RECT 2996.705 4704.545 2996.985 4704.825 ;
        RECT 2997.415 4704.545 2997.695 4704.825 ;
        RECT 2998.125 4704.545 2998.405 4704.825 ;
        RECT 2998.835 4704.545 2999.115 4704.825 ;
        RECT 2999.545 4704.545 2999.825 4704.825 ;
        RECT 3000.255 4704.545 3000.535 4704.825 ;
        RECT 3000.965 4704.545 3001.245 4704.825 ;
        RECT 3001.675 4704.545 3001.955 4704.825 ;
        RECT 3002.385 4704.545 3002.665 4704.825 ;
        RECT 3003.095 4704.545 3003.375 4704.825 ;
        RECT 3003.805 4704.545 3004.085 4704.825 ;
        RECT 3004.515 4704.545 3004.795 4704.825 ;
        RECT 3005.225 4704.545 3005.505 4704.825 ;
        RECT 2996.705 4703.835 2996.985 4704.115 ;
        RECT 2997.415 4703.835 2997.695 4704.115 ;
        RECT 2998.125 4703.835 2998.405 4704.115 ;
        RECT 2998.835 4703.835 2999.115 4704.115 ;
        RECT 2999.545 4703.835 2999.825 4704.115 ;
        RECT 3000.255 4703.835 3000.535 4704.115 ;
        RECT 3000.965 4703.835 3001.245 4704.115 ;
        RECT 3001.675 4703.835 3001.955 4704.115 ;
        RECT 3002.385 4703.835 3002.665 4704.115 ;
        RECT 3003.095 4703.835 3003.375 4704.115 ;
        RECT 3003.805 4703.835 3004.085 4704.115 ;
        RECT 3004.515 4703.835 3004.795 4704.115 ;
        RECT 3005.225 4703.835 3005.505 4704.115 ;
        RECT 2996.705 4703.125 2996.985 4703.405 ;
        RECT 2997.415 4703.125 2997.695 4703.405 ;
        RECT 2998.125 4703.125 2998.405 4703.405 ;
        RECT 2998.835 4703.125 2999.115 4703.405 ;
        RECT 2999.545 4703.125 2999.825 4703.405 ;
        RECT 3000.255 4703.125 3000.535 4703.405 ;
        RECT 3000.965 4703.125 3001.245 4703.405 ;
        RECT 3001.675 4703.125 3001.955 4703.405 ;
        RECT 3002.385 4703.125 3002.665 4703.405 ;
        RECT 3003.095 4703.125 3003.375 4703.405 ;
        RECT 3003.805 4703.125 3004.085 4703.405 ;
        RECT 3004.515 4703.125 3004.795 4703.405 ;
        RECT 3005.225 4703.125 3005.505 4703.405 ;
        RECT 2996.705 4702.415 2996.985 4702.695 ;
        RECT 2997.415 4702.415 2997.695 4702.695 ;
        RECT 2998.125 4702.415 2998.405 4702.695 ;
        RECT 2998.835 4702.415 2999.115 4702.695 ;
        RECT 2999.545 4702.415 2999.825 4702.695 ;
        RECT 3000.255 4702.415 3000.535 4702.695 ;
        RECT 3000.965 4702.415 3001.245 4702.695 ;
        RECT 3001.675 4702.415 3001.955 4702.695 ;
        RECT 3002.385 4702.415 3002.665 4702.695 ;
        RECT 3003.095 4702.415 3003.375 4702.695 ;
        RECT 3003.805 4702.415 3004.085 4702.695 ;
        RECT 3004.515 4702.415 3004.795 4702.695 ;
        RECT 3005.225 4702.415 3005.505 4702.695 ;
        RECT 2996.705 4701.705 2996.985 4701.985 ;
        RECT 2997.415 4701.705 2997.695 4701.985 ;
        RECT 2998.125 4701.705 2998.405 4701.985 ;
        RECT 2998.835 4701.705 2999.115 4701.985 ;
        RECT 2999.545 4701.705 2999.825 4701.985 ;
        RECT 3000.255 4701.705 3000.535 4701.985 ;
        RECT 3000.965 4701.705 3001.245 4701.985 ;
        RECT 3001.675 4701.705 3001.955 4701.985 ;
        RECT 3002.385 4701.705 3002.665 4701.985 ;
        RECT 3003.095 4701.705 3003.375 4701.985 ;
        RECT 3003.805 4701.705 3004.085 4701.985 ;
        RECT 3004.515 4701.705 3004.795 4701.985 ;
        RECT 3005.225 4701.705 3005.505 4701.985 ;
        RECT 2996.705 4700.995 2996.985 4701.275 ;
        RECT 2997.415 4700.995 2997.695 4701.275 ;
        RECT 2998.125 4700.995 2998.405 4701.275 ;
        RECT 2998.835 4700.995 2999.115 4701.275 ;
        RECT 2999.545 4700.995 2999.825 4701.275 ;
        RECT 3000.255 4700.995 3000.535 4701.275 ;
        RECT 3000.965 4700.995 3001.245 4701.275 ;
        RECT 3001.675 4700.995 3001.955 4701.275 ;
        RECT 3002.385 4700.995 3002.665 4701.275 ;
        RECT 3003.095 4700.995 3003.375 4701.275 ;
        RECT 3003.805 4700.995 3004.085 4701.275 ;
        RECT 3004.515 4700.995 3004.795 4701.275 ;
        RECT 3005.225 4700.995 3005.505 4701.275 ;
        RECT 2996.705 4700.285 2996.985 4700.565 ;
        RECT 2997.415 4700.285 2997.695 4700.565 ;
        RECT 2998.125 4700.285 2998.405 4700.565 ;
        RECT 2998.835 4700.285 2999.115 4700.565 ;
        RECT 2999.545 4700.285 2999.825 4700.565 ;
        RECT 3000.255 4700.285 3000.535 4700.565 ;
        RECT 3000.965 4700.285 3001.245 4700.565 ;
        RECT 3001.675 4700.285 3001.955 4700.565 ;
        RECT 3002.385 4700.285 3002.665 4700.565 ;
        RECT 3003.095 4700.285 3003.375 4700.565 ;
        RECT 3003.805 4700.285 3004.085 4700.565 ;
        RECT 3004.515 4700.285 3004.795 4700.565 ;
        RECT 3005.225 4700.285 3005.505 4700.565 ;
        RECT 2996.705 4699.575 2996.985 4699.855 ;
        RECT 2997.415 4699.575 2997.695 4699.855 ;
        RECT 2998.125 4699.575 2998.405 4699.855 ;
        RECT 2998.835 4699.575 2999.115 4699.855 ;
        RECT 2999.545 4699.575 2999.825 4699.855 ;
        RECT 3000.255 4699.575 3000.535 4699.855 ;
        RECT 3000.965 4699.575 3001.245 4699.855 ;
        RECT 3001.675 4699.575 3001.955 4699.855 ;
        RECT 3002.385 4699.575 3002.665 4699.855 ;
        RECT 3003.095 4699.575 3003.375 4699.855 ;
        RECT 3003.805 4699.575 3004.085 4699.855 ;
        RECT 3004.515 4699.575 3004.795 4699.855 ;
        RECT 3005.225 4699.575 3005.505 4699.855 ;
        RECT 2996.705 4698.865 2996.985 4699.145 ;
        RECT 2997.415 4698.865 2997.695 4699.145 ;
        RECT 2998.125 4698.865 2998.405 4699.145 ;
        RECT 2998.835 4698.865 2999.115 4699.145 ;
        RECT 2999.545 4698.865 2999.825 4699.145 ;
        RECT 3000.255 4698.865 3000.535 4699.145 ;
        RECT 3000.965 4698.865 3001.245 4699.145 ;
        RECT 3001.675 4698.865 3001.955 4699.145 ;
        RECT 3002.385 4698.865 3002.665 4699.145 ;
        RECT 3003.095 4698.865 3003.375 4699.145 ;
        RECT 3003.805 4698.865 3004.085 4699.145 ;
        RECT 3004.515 4698.865 3004.795 4699.145 ;
        RECT 3005.225 4698.865 3005.505 4699.145 ;
        RECT 3009.145 4708.095 3009.425 4708.375 ;
        RECT 3009.855 4708.095 3010.135 4708.375 ;
        RECT 3010.565 4708.095 3010.845 4708.375 ;
        RECT 3011.275 4708.095 3011.555 4708.375 ;
        RECT 3011.985 4708.095 3012.265 4708.375 ;
        RECT 3012.695 4708.095 3012.975 4708.375 ;
        RECT 3013.405 4708.095 3013.685 4708.375 ;
        RECT 3014.115 4708.095 3014.395 4708.375 ;
        RECT 3014.825 4708.095 3015.105 4708.375 ;
        RECT 3015.535 4708.095 3015.815 4708.375 ;
        RECT 3016.245 4708.095 3016.525 4708.375 ;
        RECT 3016.955 4708.095 3017.235 4708.375 ;
        RECT 3017.665 4708.095 3017.945 4708.375 ;
        RECT 3018.375 4708.095 3018.655 4708.375 ;
        RECT 3009.145 4707.385 3009.425 4707.665 ;
        RECT 3009.855 4707.385 3010.135 4707.665 ;
        RECT 3010.565 4707.385 3010.845 4707.665 ;
        RECT 3011.275 4707.385 3011.555 4707.665 ;
        RECT 3011.985 4707.385 3012.265 4707.665 ;
        RECT 3012.695 4707.385 3012.975 4707.665 ;
        RECT 3013.405 4707.385 3013.685 4707.665 ;
        RECT 3014.115 4707.385 3014.395 4707.665 ;
        RECT 3014.825 4707.385 3015.105 4707.665 ;
        RECT 3015.535 4707.385 3015.815 4707.665 ;
        RECT 3016.245 4707.385 3016.525 4707.665 ;
        RECT 3016.955 4707.385 3017.235 4707.665 ;
        RECT 3017.665 4707.385 3017.945 4707.665 ;
        RECT 3018.375 4707.385 3018.655 4707.665 ;
        RECT 3009.145 4706.675 3009.425 4706.955 ;
        RECT 3009.855 4706.675 3010.135 4706.955 ;
        RECT 3010.565 4706.675 3010.845 4706.955 ;
        RECT 3011.275 4706.675 3011.555 4706.955 ;
        RECT 3011.985 4706.675 3012.265 4706.955 ;
        RECT 3012.695 4706.675 3012.975 4706.955 ;
        RECT 3013.405 4706.675 3013.685 4706.955 ;
        RECT 3014.115 4706.675 3014.395 4706.955 ;
        RECT 3014.825 4706.675 3015.105 4706.955 ;
        RECT 3015.535 4706.675 3015.815 4706.955 ;
        RECT 3016.245 4706.675 3016.525 4706.955 ;
        RECT 3016.955 4706.675 3017.235 4706.955 ;
        RECT 3017.665 4706.675 3017.945 4706.955 ;
        RECT 3018.375 4706.675 3018.655 4706.955 ;
        RECT 3009.145 4705.965 3009.425 4706.245 ;
        RECT 3009.855 4705.965 3010.135 4706.245 ;
        RECT 3010.565 4705.965 3010.845 4706.245 ;
        RECT 3011.275 4705.965 3011.555 4706.245 ;
        RECT 3011.985 4705.965 3012.265 4706.245 ;
        RECT 3012.695 4705.965 3012.975 4706.245 ;
        RECT 3013.405 4705.965 3013.685 4706.245 ;
        RECT 3014.115 4705.965 3014.395 4706.245 ;
        RECT 3014.825 4705.965 3015.105 4706.245 ;
        RECT 3015.535 4705.965 3015.815 4706.245 ;
        RECT 3016.245 4705.965 3016.525 4706.245 ;
        RECT 3016.955 4705.965 3017.235 4706.245 ;
        RECT 3017.665 4705.965 3017.945 4706.245 ;
        RECT 3018.375 4705.965 3018.655 4706.245 ;
        RECT 3009.145 4705.255 3009.425 4705.535 ;
        RECT 3009.855 4705.255 3010.135 4705.535 ;
        RECT 3010.565 4705.255 3010.845 4705.535 ;
        RECT 3011.275 4705.255 3011.555 4705.535 ;
        RECT 3011.985 4705.255 3012.265 4705.535 ;
        RECT 3012.695 4705.255 3012.975 4705.535 ;
        RECT 3013.405 4705.255 3013.685 4705.535 ;
        RECT 3014.115 4705.255 3014.395 4705.535 ;
        RECT 3014.825 4705.255 3015.105 4705.535 ;
        RECT 3015.535 4705.255 3015.815 4705.535 ;
        RECT 3016.245 4705.255 3016.525 4705.535 ;
        RECT 3016.955 4705.255 3017.235 4705.535 ;
        RECT 3017.665 4705.255 3017.945 4705.535 ;
        RECT 3018.375 4705.255 3018.655 4705.535 ;
        RECT 3009.145 4704.545 3009.425 4704.825 ;
        RECT 3009.855 4704.545 3010.135 4704.825 ;
        RECT 3010.565 4704.545 3010.845 4704.825 ;
        RECT 3011.275 4704.545 3011.555 4704.825 ;
        RECT 3011.985 4704.545 3012.265 4704.825 ;
        RECT 3012.695 4704.545 3012.975 4704.825 ;
        RECT 3013.405 4704.545 3013.685 4704.825 ;
        RECT 3014.115 4704.545 3014.395 4704.825 ;
        RECT 3014.825 4704.545 3015.105 4704.825 ;
        RECT 3015.535 4704.545 3015.815 4704.825 ;
        RECT 3016.245 4704.545 3016.525 4704.825 ;
        RECT 3016.955 4704.545 3017.235 4704.825 ;
        RECT 3017.665 4704.545 3017.945 4704.825 ;
        RECT 3018.375 4704.545 3018.655 4704.825 ;
        RECT 3009.145 4703.835 3009.425 4704.115 ;
        RECT 3009.855 4703.835 3010.135 4704.115 ;
        RECT 3010.565 4703.835 3010.845 4704.115 ;
        RECT 3011.275 4703.835 3011.555 4704.115 ;
        RECT 3011.985 4703.835 3012.265 4704.115 ;
        RECT 3012.695 4703.835 3012.975 4704.115 ;
        RECT 3013.405 4703.835 3013.685 4704.115 ;
        RECT 3014.115 4703.835 3014.395 4704.115 ;
        RECT 3014.825 4703.835 3015.105 4704.115 ;
        RECT 3015.535 4703.835 3015.815 4704.115 ;
        RECT 3016.245 4703.835 3016.525 4704.115 ;
        RECT 3016.955 4703.835 3017.235 4704.115 ;
        RECT 3017.665 4703.835 3017.945 4704.115 ;
        RECT 3018.375 4703.835 3018.655 4704.115 ;
        RECT 3009.145 4703.125 3009.425 4703.405 ;
        RECT 3009.855 4703.125 3010.135 4703.405 ;
        RECT 3010.565 4703.125 3010.845 4703.405 ;
        RECT 3011.275 4703.125 3011.555 4703.405 ;
        RECT 3011.985 4703.125 3012.265 4703.405 ;
        RECT 3012.695 4703.125 3012.975 4703.405 ;
        RECT 3013.405 4703.125 3013.685 4703.405 ;
        RECT 3014.115 4703.125 3014.395 4703.405 ;
        RECT 3014.825 4703.125 3015.105 4703.405 ;
        RECT 3015.535 4703.125 3015.815 4703.405 ;
        RECT 3016.245 4703.125 3016.525 4703.405 ;
        RECT 3016.955 4703.125 3017.235 4703.405 ;
        RECT 3017.665 4703.125 3017.945 4703.405 ;
        RECT 3018.375 4703.125 3018.655 4703.405 ;
        RECT 3009.145 4702.415 3009.425 4702.695 ;
        RECT 3009.855 4702.415 3010.135 4702.695 ;
        RECT 3010.565 4702.415 3010.845 4702.695 ;
        RECT 3011.275 4702.415 3011.555 4702.695 ;
        RECT 3011.985 4702.415 3012.265 4702.695 ;
        RECT 3012.695 4702.415 3012.975 4702.695 ;
        RECT 3013.405 4702.415 3013.685 4702.695 ;
        RECT 3014.115 4702.415 3014.395 4702.695 ;
        RECT 3014.825 4702.415 3015.105 4702.695 ;
        RECT 3015.535 4702.415 3015.815 4702.695 ;
        RECT 3016.245 4702.415 3016.525 4702.695 ;
        RECT 3016.955 4702.415 3017.235 4702.695 ;
        RECT 3017.665 4702.415 3017.945 4702.695 ;
        RECT 3018.375 4702.415 3018.655 4702.695 ;
        RECT 3009.145 4701.705 3009.425 4701.985 ;
        RECT 3009.855 4701.705 3010.135 4701.985 ;
        RECT 3010.565 4701.705 3010.845 4701.985 ;
        RECT 3011.275 4701.705 3011.555 4701.985 ;
        RECT 3011.985 4701.705 3012.265 4701.985 ;
        RECT 3012.695 4701.705 3012.975 4701.985 ;
        RECT 3013.405 4701.705 3013.685 4701.985 ;
        RECT 3014.115 4701.705 3014.395 4701.985 ;
        RECT 3014.825 4701.705 3015.105 4701.985 ;
        RECT 3015.535 4701.705 3015.815 4701.985 ;
        RECT 3016.245 4701.705 3016.525 4701.985 ;
        RECT 3016.955 4701.705 3017.235 4701.985 ;
        RECT 3017.665 4701.705 3017.945 4701.985 ;
        RECT 3018.375 4701.705 3018.655 4701.985 ;
        RECT 3009.145 4700.995 3009.425 4701.275 ;
        RECT 3009.855 4700.995 3010.135 4701.275 ;
        RECT 3010.565 4700.995 3010.845 4701.275 ;
        RECT 3011.275 4700.995 3011.555 4701.275 ;
        RECT 3011.985 4700.995 3012.265 4701.275 ;
        RECT 3012.695 4700.995 3012.975 4701.275 ;
        RECT 3013.405 4700.995 3013.685 4701.275 ;
        RECT 3014.115 4700.995 3014.395 4701.275 ;
        RECT 3014.825 4700.995 3015.105 4701.275 ;
        RECT 3015.535 4700.995 3015.815 4701.275 ;
        RECT 3016.245 4700.995 3016.525 4701.275 ;
        RECT 3016.955 4700.995 3017.235 4701.275 ;
        RECT 3017.665 4700.995 3017.945 4701.275 ;
        RECT 3018.375 4700.995 3018.655 4701.275 ;
        RECT 3009.145 4700.285 3009.425 4700.565 ;
        RECT 3009.855 4700.285 3010.135 4700.565 ;
        RECT 3010.565 4700.285 3010.845 4700.565 ;
        RECT 3011.275 4700.285 3011.555 4700.565 ;
        RECT 3011.985 4700.285 3012.265 4700.565 ;
        RECT 3012.695 4700.285 3012.975 4700.565 ;
        RECT 3013.405 4700.285 3013.685 4700.565 ;
        RECT 3014.115 4700.285 3014.395 4700.565 ;
        RECT 3014.825 4700.285 3015.105 4700.565 ;
        RECT 3015.535 4700.285 3015.815 4700.565 ;
        RECT 3016.245 4700.285 3016.525 4700.565 ;
        RECT 3016.955 4700.285 3017.235 4700.565 ;
        RECT 3017.665 4700.285 3017.945 4700.565 ;
        RECT 3018.375 4700.285 3018.655 4700.565 ;
        RECT 3009.145 4699.575 3009.425 4699.855 ;
        RECT 3009.855 4699.575 3010.135 4699.855 ;
        RECT 3010.565 4699.575 3010.845 4699.855 ;
        RECT 3011.275 4699.575 3011.555 4699.855 ;
        RECT 3011.985 4699.575 3012.265 4699.855 ;
        RECT 3012.695 4699.575 3012.975 4699.855 ;
        RECT 3013.405 4699.575 3013.685 4699.855 ;
        RECT 3014.115 4699.575 3014.395 4699.855 ;
        RECT 3014.825 4699.575 3015.105 4699.855 ;
        RECT 3015.535 4699.575 3015.815 4699.855 ;
        RECT 3016.245 4699.575 3016.525 4699.855 ;
        RECT 3016.955 4699.575 3017.235 4699.855 ;
        RECT 3017.665 4699.575 3017.945 4699.855 ;
        RECT 3018.375 4699.575 3018.655 4699.855 ;
        RECT 3009.145 4698.865 3009.425 4699.145 ;
        RECT 3009.855 4698.865 3010.135 4699.145 ;
        RECT 3010.565 4698.865 3010.845 4699.145 ;
        RECT 3011.275 4698.865 3011.555 4699.145 ;
        RECT 3011.985 4698.865 3012.265 4699.145 ;
        RECT 3012.695 4698.865 3012.975 4699.145 ;
        RECT 3013.405 4698.865 3013.685 4699.145 ;
        RECT 3014.115 4698.865 3014.395 4699.145 ;
        RECT 3014.825 4698.865 3015.105 4699.145 ;
        RECT 3015.535 4698.865 3015.815 4699.145 ;
        RECT 3016.245 4698.865 3016.525 4699.145 ;
        RECT 3016.955 4698.865 3017.235 4699.145 ;
        RECT 3017.665 4698.865 3017.945 4699.145 ;
        RECT 3018.375 4698.865 3018.655 4699.145 ;
        RECT 3025.255 4708.095 3025.535 4708.375 ;
        RECT 3025.965 4708.095 3026.245 4708.375 ;
        RECT 3026.675 4708.095 3026.955 4708.375 ;
        RECT 3027.385 4708.095 3027.665 4708.375 ;
        RECT 3028.095 4708.095 3028.375 4708.375 ;
        RECT 3028.805 4708.095 3029.085 4708.375 ;
        RECT 3029.515 4708.095 3029.795 4708.375 ;
        RECT 3030.225 4708.095 3030.505 4708.375 ;
        RECT 3025.255 4707.385 3025.535 4707.665 ;
        RECT 3025.965 4707.385 3026.245 4707.665 ;
        RECT 3026.675 4707.385 3026.955 4707.665 ;
        RECT 3027.385 4707.385 3027.665 4707.665 ;
        RECT 3028.095 4707.385 3028.375 4707.665 ;
        RECT 3028.805 4707.385 3029.085 4707.665 ;
        RECT 3029.515 4707.385 3029.795 4707.665 ;
        RECT 3030.225 4707.385 3030.505 4707.665 ;
        RECT 3025.255 4706.675 3025.535 4706.955 ;
        RECT 3025.965 4706.675 3026.245 4706.955 ;
        RECT 3026.675 4706.675 3026.955 4706.955 ;
        RECT 3027.385 4706.675 3027.665 4706.955 ;
        RECT 3028.095 4706.675 3028.375 4706.955 ;
        RECT 3028.805 4706.675 3029.085 4706.955 ;
        RECT 3029.515 4706.675 3029.795 4706.955 ;
        RECT 3030.225 4706.675 3030.505 4706.955 ;
        RECT 3025.255 4705.965 3025.535 4706.245 ;
        RECT 3025.965 4705.965 3026.245 4706.245 ;
        RECT 3026.675 4705.965 3026.955 4706.245 ;
        RECT 3027.385 4705.965 3027.665 4706.245 ;
        RECT 3028.095 4705.965 3028.375 4706.245 ;
        RECT 3028.805 4705.965 3029.085 4706.245 ;
        RECT 3029.515 4705.965 3029.795 4706.245 ;
        RECT 3030.225 4705.965 3030.505 4706.245 ;
        RECT 3025.255 4705.255 3025.535 4705.535 ;
        RECT 3025.965 4705.255 3026.245 4705.535 ;
        RECT 3026.675 4705.255 3026.955 4705.535 ;
        RECT 3027.385 4705.255 3027.665 4705.535 ;
        RECT 3028.095 4705.255 3028.375 4705.535 ;
        RECT 3028.805 4705.255 3029.085 4705.535 ;
        RECT 3029.515 4705.255 3029.795 4705.535 ;
        RECT 3030.225 4705.255 3030.505 4705.535 ;
        RECT 3025.255 4704.545 3025.535 4704.825 ;
        RECT 3025.965 4704.545 3026.245 4704.825 ;
        RECT 3026.675 4704.545 3026.955 4704.825 ;
        RECT 3027.385 4704.545 3027.665 4704.825 ;
        RECT 3028.095 4704.545 3028.375 4704.825 ;
        RECT 3028.805 4704.545 3029.085 4704.825 ;
        RECT 3029.515 4704.545 3029.795 4704.825 ;
        RECT 3030.225 4704.545 3030.505 4704.825 ;
        RECT 3025.255 4703.835 3025.535 4704.115 ;
        RECT 3025.965 4703.835 3026.245 4704.115 ;
        RECT 3026.675 4703.835 3026.955 4704.115 ;
        RECT 3027.385 4703.835 3027.665 4704.115 ;
        RECT 3028.095 4703.835 3028.375 4704.115 ;
        RECT 3028.805 4703.835 3029.085 4704.115 ;
        RECT 3029.515 4703.835 3029.795 4704.115 ;
        RECT 3030.225 4703.835 3030.505 4704.115 ;
        RECT 3025.255 4703.125 3025.535 4703.405 ;
        RECT 3025.965 4703.125 3026.245 4703.405 ;
        RECT 3026.675 4703.125 3026.955 4703.405 ;
        RECT 3027.385 4703.125 3027.665 4703.405 ;
        RECT 3028.095 4703.125 3028.375 4703.405 ;
        RECT 3028.805 4703.125 3029.085 4703.405 ;
        RECT 3029.515 4703.125 3029.795 4703.405 ;
        RECT 3030.225 4703.125 3030.505 4703.405 ;
        RECT 3025.255 4702.415 3025.535 4702.695 ;
        RECT 3025.965 4702.415 3026.245 4702.695 ;
        RECT 3026.675 4702.415 3026.955 4702.695 ;
        RECT 3027.385 4702.415 3027.665 4702.695 ;
        RECT 3028.095 4702.415 3028.375 4702.695 ;
        RECT 3028.805 4702.415 3029.085 4702.695 ;
        RECT 3029.515 4702.415 3029.795 4702.695 ;
        RECT 3030.225 4702.415 3030.505 4702.695 ;
        RECT 3025.255 4701.705 3025.535 4701.985 ;
        RECT 3025.965 4701.705 3026.245 4701.985 ;
        RECT 3026.675 4701.705 3026.955 4701.985 ;
        RECT 3027.385 4701.705 3027.665 4701.985 ;
        RECT 3028.095 4701.705 3028.375 4701.985 ;
        RECT 3028.805 4701.705 3029.085 4701.985 ;
        RECT 3029.515 4701.705 3029.795 4701.985 ;
        RECT 3030.225 4701.705 3030.505 4701.985 ;
        RECT 3025.255 4700.995 3025.535 4701.275 ;
        RECT 3025.965 4700.995 3026.245 4701.275 ;
        RECT 3026.675 4700.995 3026.955 4701.275 ;
        RECT 3027.385 4700.995 3027.665 4701.275 ;
        RECT 3028.095 4700.995 3028.375 4701.275 ;
        RECT 3028.805 4700.995 3029.085 4701.275 ;
        RECT 3029.515 4700.995 3029.795 4701.275 ;
        RECT 3030.225 4700.995 3030.505 4701.275 ;
        RECT 3025.255 4700.285 3025.535 4700.565 ;
        RECT 3025.965 4700.285 3026.245 4700.565 ;
        RECT 3026.675 4700.285 3026.955 4700.565 ;
        RECT 3027.385 4700.285 3027.665 4700.565 ;
        RECT 3028.095 4700.285 3028.375 4700.565 ;
        RECT 3028.805 4700.285 3029.085 4700.565 ;
        RECT 3029.515 4700.285 3029.795 4700.565 ;
        RECT 3030.225 4700.285 3030.505 4700.565 ;
        RECT 3025.255 4699.575 3025.535 4699.855 ;
        RECT 3025.965 4699.575 3026.245 4699.855 ;
        RECT 3026.675 4699.575 3026.955 4699.855 ;
        RECT 3027.385 4699.575 3027.665 4699.855 ;
        RECT 3028.095 4699.575 3028.375 4699.855 ;
        RECT 3028.805 4699.575 3029.085 4699.855 ;
        RECT 3029.515 4699.575 3029.795 4699.855 ;
        RECT 3030.225 4699.575 3030.505 4699.855 ;
        RECT 3025.255 4698.865 3025.535 4699.145 ;
        RECT 3025.965 4698.865 3026.245 4699.145 ;
        RECT 3026.675 4698.865 3026.955 4699.145 ;
        RECT 3027.385 4698.865 3027.665 4699.145 ;
        RECT 3028.095 4698.865 3028.375 4699.145 ;
        RECT 3028.805 4698.865 3029.085 4699.145 ;
        RECT 3029.515 4698.865 3029.795 4699.145 ;
        RECT 3030.225 4698.865 3030.505 4699.145 ;
        RECT 3034.525 4708.095 3034.805 4708.375 ;
        RECT 3035.235 4708.095 3035.515 4708.375 ;
        RECT 3035.945 4708.095 3036.225 4708.375 ;
        RECT 3036.655 4708.095 3036.935 4708.375 ;
        RECT 3037.365 4708.095 3037.645 4708.375 ;
        RECT 3038.075 4708.095 3038.355 4708.375 ;
        RECT 3038.785 4708.095 3039.065 4708.375 ;
        RECT 3039.495 4708.095 3039.775 4708.375 ;
        RECT 3040.205 4708.095 3040.485 4708.375 ;
        RECT 3040.915 4708.095 3041.195 4708.375 ;
        RECT 3041.625 4708.095 3041.905 4708.375 ;
        RECT 3042.335 4708.095 3042.615 4708.375 ;
        RECT 3043.045 4708.095 3043.325 4708.375 ;
        RECT 3043.755 4708.095 3044.035 4708.375 ;
        RECT 3034.525 4707.385 3034.805 4707.665 ;
        RECT 3035.235 4707.385 3035.515 4707.665 ;
        RECT 3035.945 4707.385 3036.225 4707.665 ;
        RECT 3036.655 4707.385 3036.935 4707.665 ;
        RECT 3037.365 4707.385 3037.645 4707.665 ;
        RECT 3038.075 4707.385 3038.355 4707.665 ;
        RECT 3038.785 4707.385 3039.065 4707.665 ;
        RECT 3039.495 4707.385 3039.775 4707.665 ;
        RECT 3040.205 4707.385 3040.485 4707.665 ;
        RECT 3040.915 4707.385 3041.195 4707.665 ;
        RECT 3041.625 4707.385 3041.905 4707.665 ;
        RECT 3042.335 4707.385 3042.615 4707.665 ;
        RECT 3043.045 4707.385 3043.325 4707.665 ;
        RECT 3043.755 4707.385 3044.035 4707.665 ;
        RECT 3034.525 4706.675 3034.805 4706.955 ;
        RECT 3035.235 4706.675 3035.515 4706.955 ;
        RECT 3035.945 4706.675 3036.225 4706.955 ;
        RECT 3036.655 4706.675 3036.935 4706.955 ;
        RECT 3037.365 4706.675 3037.645 4706.955 ;
        RECT 3038.075 4706.675 3038.355 4706.955 ;
        RECT 3038.785 4706.675 3039.065 4706.955 ;
        RECT 3039.495 4706.675 3039.775 4706.955 ;
        RECT 3040.205 4706.675 3040.485 4706.955 ;
        RECT 3040.915 4706.675 3041.195 4706.955 ;
        RECT 3041.625 4706.675 3041.905 4706.955 ;
        RECT 3042.335 4706.675 3042.615 4706.955 ;
        RECT 3043.045 4706.675 3043.325 4706.955 ;
        RECT 3043.755 4706.675 3044.035 4706.955 ;
        RECT 3034.525 4705.965 3034.805 4706.245 ;
        RECT 3035.235 4705.965 3035.515 4706.245 ;
        RECT 3035.945 4705.965 3036.225 4706.245 ;
        RECT 3036.655 4705.965 3036.935 4706.245 ;
        RECT 3037.365 4705.965 3037.645 4706.245 ;
        RECT 3038.075 4705.965 3038.355 4706.245 ;
        RECT 3038.785 4705.965 3039.065 4706.245 ;
        RECT 3039.495 4705.965 3039.775 4706.245 ;
        RECT 3040.205 4705.965 3040.485 4706.245 ;
        RECT 3040.915 4705.965 3041.195 4706.245 ;
        RECT 3041.625 4705.965 3041.905 4706.245 ;
        RECT 3042.335 4705.965 3042.615 4706.245 ;
        RECT 3043.045 4705.965 3043.325 4706.245 ;
        RECT 3043.755 4705.965 3044.035 4706.245 ;
        RECT 3034.525 4705.255 3034.805 4705.535 ;
        RECT 3035.235 4705.255 3035.515 4705.535 ;
        RECT 3035.945 4705.255 3036.225 4705.535 ;
        RECT 3036.655 4705.255 3036.935 4705.535 ;
        RECT 3037.365 4705.255 3037.645 4705.535 ;
        RECT 3038.075 4705.255 3038.355 4705.535 ;
        RECT 3038.785 4705.255 3039.065 4705.535 ;
        RECT 3039.495 4705.255 3039.775 4705.535 ;
        RECT 3040.205 4705.255 3040.485 4705.535 ;
        RECT 3040.915 4705.255 3041.195 4705.535 ;
        RECT 3041.625 4705.255 3041.905 4705.535 ;
        RECT 3042.335 4705.255 3042.615 4705.535 ;
        RECT 3043.045 4705.255 3043.325 4705.535 ;
        RECT 3043.755 4705.255 3044.035 4705.535 ;
        RECT 3034.525 4704.545 3034.805 4704.825 ;
        RECT 3035.235 4704.545 3035.515 4704.825 ;
        RECT 3035.945 4704.545 3036.225 4704.825 ;
        RECT 3036.655 4704.545 3036.935 4704.825 ;
        RECT 3037.365 4704.545 3037.645 4704.825 ;
        RECT 3038.075 4704.545 3038.355 4704.825 ;
        RECT 3038.785 4704.545 3039.065 4704.825 ;
        RECT 3039.495 4704.545 3039.775 4704.825 ;
        RECT 3040.205 4704.545 3040.485 4704.825 ;
        RECT 3040.915 4704.545 3041.195 4704.825 ;
        RECT 3041.625 4704.545 3041.905 4704.825 ;
        RECT 3042.335 4704.545 3042.615 4704.825 ;
        RECT 3043.045 4704.545 3043.325 4704.825 ;
        RECT 3043.755 4704.545 3044.035 4704.825 ;
        RECT 3034.525 4703.835 3034.805 4704.115 ;
        RECT 3035.235 4703.835 3035.515 4704.115 ;
        RECT 3035.945 4703.835 3036.225 4704.115 ;
        RECT 3036.655 4703.835 3036.935 4704.115 ;
        RECT 3037.365 4703.835 3037.645 4704.115 ;
        RECT 3038.075 4703.835 3038.355 4704.115 ;
        RECT 3038.785 4703.835 3039.065 4704.115 ;
        RECT 3039.495 4703.835 3039.775 4704.115 ;
        RECT 3040.205 4703.835 3040.485 4704.115 ;
        RECT 3040.915 4703.835 3041.195 4704.115 ;
        RECT 3041.625 4703.835 3041.905 4704.115 ;
        RECT 3042.335 4703.835 3042.615 4704.115 ;
        RECT 3043.045 4703.835 3043.325 4704.115 ;
        RECT 3043.755 4703.835 3044.035 4704.115 ;
        RECT 3034.525 4703.125 3034.805 4703.405 ;
        RECT 3035.235 4703.125 3035.515 4703.405 ;
        RECT 3035.945 4703.125 3036.225 4703.405 ;
        RECT 3036.655 4703.125 3036.935 4703.405 ;
        RECT 3037.365 4703.125 3037.645 4703.405 ;
        RECT 3038.075 4703.125 3038.355 4703.405 ;
        RECT 3038.785 4703.125 3039.065 4703.405 ;
        RECT 3039.495 4703.125 3039.775 4703.405 ;
        RECT 3040.205 4703.125 3040.485 4703.405 ;
        RECT 3040.915 4703.125 3041.195 4703.405 ;
        RECT 3041.625 4703.125 3041.905 4703.405 ;
        RECT 3042.335 4703.125 3042.615 4703.405 ;
        RECT 3043.045 4703.125 3043.325 4703.405 ;
        RECT 3043.755 4703.125 3044.035 4703.405 ;
        RECT 3034.525 4702.415 3034.805 4702.695 ;
        RECT 3035.235 4702.415 3035.515 4702.695 ;
        RECT 3035.945 4702.415 3036.225 4702.695 ;
        RECT 3036.655 4702.415 3036.935 4702.695 ;
        RECT 3037.365 4702.415 3037.645 4702.695 ;
        RECT 3038.075 4702.415 3038.355 4702.695 ;
        RECT 3038.785 4702.415 3039.065 4702.695 ;
        RECT 3039.495 4702.415 3039.775 4702.695 ;
        RECT 3040.205 4702.415 3040.485 4702.695 ;
        RECT 3040.915 4702.415 3041.195 4702.695 ;
        RECT 3041.625 4702.415 3041.905 4702.695 ;
        RECT 3042.335 4702.415 3042.615 4702.695 ;
        RECT 3043.045 4702.415 3043.325 4702.695 ;
        RECT 3043.755 4702.415 3044.035 4702.695 ;
        RECT 3034.525 4701.705 3034.805 4701.985 ;
        RECT 3035.235 4701.705 3035.515 4701.985 ;
        RECT 3035.945 4701.705 3036.225 4701.985 ;
        RECT 3036.655 4701.705 3036.935 4701.985 ;
        RECT 3037.365 4701.705 3037.645 4701.985 ;
        RECT 3038.075 4701.705 3038.355 4701.985 ;
        RECT 3038.785 4701.705 3039.065 4701.985 ;
        RECT 3039.495 4701.705 3039.775 4701.985 ;
        RECT 3040.205 4701.705 3040.485 4701.985 ;
        RECT 3040.915 4701.705 3041.195 4701.985 ;
        RECT 3041.625 4701.705 3041.905 4701.985 ;
        RECT 3042.335 4701.705 3042.615 4701.985 ;
        RECT 3043.045 4701.705 3043.325 4701.985 ;
        RECT 3043.755 4701.705 3044.035 4701.985 ;
        RECT 3034.525 4700.995 3034.805 4701.275 ;
        RECT 3035.235 4700.995 3035.515 4701.275 ;
        RECT 3035.945 4700.995 3036.225 4701.275 ;
        RECT 3036.655 4700.995 3036.935 4701.275 ;
        RECT 3037.365 4700.995 3037.645 4701.275 ;
        RECT 3038.075 4700.995 3038.355 4701.275 ;
        RECT 3038.785 4700.995 3039.065 4701.275 ;
        RECT 3039.495 4700.995 3039.775 4701.275 ;
        RECT 3040.205 4700.995 3040.485 4701.275 ;
        RECT 3040.915 4700.995 3041.195 4701.275 ;
        RECT 3041.625 4700.995 3041.905 4701.275 ;
        RECT 3042.335 4700.995 3042.615 4701.275 ;
        RECT 3043.045 4700.995 3043.325 4701.275 ;
        RECT 3043.755 4700.995 3044.035 4701.275 ;
        RECT 3034.525 4700.285 3034.805 4700.565 ;
        RECT 3035.235 4700.285 3035.515 4700.565 ;
        RECT 3035.945 4700.285 3036.225 4700.565 ;
        RECT 3036.655 4700.285 3036.935 4700.565 ;
        RECT 3037.365 4700.285 3037.645 4700.565 ;
        RECT 3038.075 4700.285 3038.355 4700.565 ;
        RECT 3038.785 4700.285 3039.065 4700.565 ;
        RECT 3039.495 4700.285 3039.775 4700.565 ;
        RECT 3040.205 4700.285 3040.485 4700.565 ;
        RECT 3040.915 4700.285 3041.195 4700.565 ;
        RECT 3041.625 4700.285 3041.905 4700.565 ;
        RECT 3042.335 4700.285 3042.615 4700.565 ;
        RECT 3043.045 4700.285 3043.325 4700.565 ;
        RECT 3043.755 4700.285 3044.035 4700.565 ;
        RECT 3034.525 4699.575 3034.805 4699.855 ;
        RECT 3035.235 4699.575 3035.515 4699.855 ;
        RECT 3035.945 4699.575 3036.225 4699.855 ;
        RECT 3036.655 4699.575 3036.935 4699.855 ;
        RECT 3037.365 4699.575 3037.645 4699.855 ;
        RECT 3038.075 4699.575 3038.355 4699.855 ;
        RECT 3038.785 4699.575 3039.065 4699.855 ;
        RECT 3039.495 4699.575 3039.775 4699.855 ;
        RECT 3040.205 4699.575 3040.485 4699.855 ;
        RECT 3040.915 4699.575 3041.195 4699.855 ;
        RECT 3041.625 4699.575 3041.905 4699.855 ;
        RECT 3042.335 4699.575 3042.615 4699.855 ;
        RECT 3043.045 4699.575 3043.325 4699.855 ;
        RECT 3043.755 4699.575 3044.035 4699.855 ;
        RECT 3034.525 4698.865 3034.805 4699.145 ;
        RECT 3035.235 4698.865 3035.515 4699.145 ;
        RECT 3035.945 4698.865 3036.225 4699.145 ;
        RECT 3036.655 4698.865 3036.935 4699.145 ;
        RECT 3037.365 4698.865 3037.645 4699.145 ;
        RECT 3038.075 4698.865 3038.355 4699.145 ;
        RECT 3038.785 4698.865 3039.065 4699.145 ;
        RECT 3039.495 4698.865 3039.775 4699.145 ;
        RECT 3040.205 4698.865 3040.485 4699.145 ;
        RECT 3040.915 4698.865 3041.195 4699.145 ;
        RECT 3041.625 4698.865 3041.905 4699.145 ;
        RECT 3042.335 4698.865 3042.615 4699.145 ;
        RECT 3043.045 4698.865 3043.325 4699.145 ;
        RECT 3043.755 4698.865 3044.035 4699.145 ;
        RECT 3046.375 4708.095 3046.655 4708.375 ;
        RECT 3047.085 4708.095 3047.365 4708.375 ;
        RECT 3047.795 4708.095 3048.075 4708.375 ;
        RECT 3048.505 4708.095 3048.785 4708.375 ;
        RECT 3049.215 4708.095 3049.495 4708.375 ;
        RECT 3049.925 4708.095 3050.205 4708.375 ;
        RECT 3050.635 4708.095 3050.915 4708.375 ;
        RECT 3051.345 4708.095 3051.625 4708.375 ;
        RECT 3052.055 4708.095 3052.335 4708.375 ;
        RECT 3052.765 4708.095 3053.045 4708.375 ;
        RECT 3053.475 4708.095 3053.755 4708.375 ;
        RECT 3054.185 4708.095 3054.465 4708.375 ;
        RECT 3054.895 4708.095 3055.175 4708.375 ;
        RECT 3055.605 4708.095 3055.885 4708.375 ;
        RECT 3046.375 4707.385 3046.655 4707.665 ;
        RECT 3047.085 4707.385 3047.365 4707.665 ;
        RECT 3047.795 4707.385 3048.075 4707.665 ;
        RECT 3048.505 4707.385 3048.785 4707.665 ;
        RECT 3049.215 4707.385 3049.495 4707.665 ;
        RECT 3049.925 4707.385 3050.205 4707.665 ;
        RECT 3050.635 4707.385 3050.915 4707.665 ;
        RECT 3051.345 4707.385 3051.625 4707.665 ;
        RECT 3052.055 4707.385 3052.335 4707.665 ;
        RECT 3052.765 4707.385 3053.045 4707.665 ;
        RECT 3053.475 4707.385 3053.755 4707.665 ;
        RECT 3054.185 4707.385 3054.465 4707.665 ;
        RECT 3054.895 4707.385 3055.175 4707.665 ;
        RECT 3055.605 4707.385 3055.885 4707.665 ;
        RECT 3046.375 4706.675 3046.655 4706.955 ;
        RECT 3047.085 4706.675 3047.365 4706.955 ;
        RECT 3047.795 4706.675 3048.075 4706.955 ;
        RECT 3048.505 4706.675 3048.785 4706.955 ;
        RECT 3049.215 4706.675 3049.495 4706.955 ;
        RECT 3049.925 4706.675 3050.205 4706.955 ;
        RECT 3050.635 4706.675 3050.915 4706.955 ;
        RECT 3051.345 4706.675 3051.625 4706.955 ;
        RECT 3052.055 4706.675 3052.335 4706.955 ;
        RECT 3052.765 4706.675 3053.045 4706.955 ;
        RECT 3053.475 4706.675 3053.755 4706.955 ;
        RECT 3054.185 4706.675 3054.465 4706.955 ;
        RECT 3054.895 4706.675 3055.175 4706.955 ;
        RECT 3055.605 4706.675 3055.885 4706.955 ;
        RECT 3046.375 4705.965 3046.655 4706.245 ;
        RECT 3047.085 4705.965 3047.365 4706.245 ;
        RECT 3047.795 4705.965 3048.075 4706.245 ;
        RECT 3048.505 4705.965 3048.785 4706.245 ;
        RECT 3049.215 4705.965 3049.495 4706.245 ;
        RECT 3049.925 4705.965 3050.205 4706.245 ;
        RECT 3050.635 4705.965 3050.915 4706.245 ;
        RECT 3051.345 4705.965 3051.625 4706.245 ;
        RECT 3052.055 4705.965 3052.335 4706.245 ;
        RECT 3052.765 4705.965 3053.045 4706.245 ;
        RECT 3053.475 4705.965 3053.755 4706.245 ;
        RECT 3054.185 4705.965 3054.465 4706.245 ;
        RECT 3054.895 4705.965 3055.175 4706.245 ;
        RECT 3055.605 4705.965 3055.885 4706.245 ;
        RECT 3046.375 4705.255 3046.655 4705.535 ;
        RECT 3047.085 4705.255 3047.365 4705.535 ;
        RECT 3047.795 4705.255 3048.075 4705.535 ;
        RECT 3048.505 4705.255 3048.785 4705.535 ;
        RECT 3049.215 4705.255 3049.495 4705.535 ;
        RECT 3049.925 4705.255 3050.205 4705.535 ;
        RECT 3050.635 4705.255 3050.915 4705.535 ;
        RECT 3051.345 4705.255 3051.625 4705.535 ;
        RECT 3052.055 4705.255 3052.335 4705.535 ;
        RECT 3052.765 4705.255 3053.045 4705.535 ;
        RECT 3053.475 4705.255 3053.755 4705.535 ;
        RECT 3054.185 4705.255 3054.465 4705.535 ;
        RECT 3054.895 4705.255 3055.175 4705.535 ;
        RECT 3055.605 4705.255 3055.885 4705.535 ;
        RECT 3046.375 4704.545 3046.655 4704.825 ;
        RECT 3047.085 4704.545 3047.365 4704.825 ;
        RECT 3047.795 4704.545 3048.075 4704.825 ;
        RECT 3048.505 4704.545 3048.785 4704.825 ;
        RECT 3049.215 4704.545 3049.495 4704.825 ;
        RECT 3049.925 4704.545 3050.205 4704.825 ;
        RECT 3050.635 4704.545 3050.915 4704.825 ;
        RECT 3051.345 4704.545 3051.625 4704.825 ;
        RECT 3052.055 4704.545 3052.335 4704.825 ;
        RECT 3052.765 4704.545 3053.045 4704.825 ;
        RECT 3053.475 4704.545 3053.755 4704.825 ;
        RECT 3054.185 4704.545 3054.465 4704.825 ;
        RECT 3054.895 4704.545 3055.175 4704.825 ;
        RECT 3055.605 4704.545 3055.885 4704.825 ;
        RECT 3046.375 4703.835 3046.655 4704.115 ;
        RECT 3047.085 4703.835 3047.365 4704.115 ;
        RECT 3047.795 4703.835 3048.075 4704.115 ;
        RECT 3048.505 4703.835 3048.785 4704.115 ;
        RECT 3049.215 4703.835 3049.495 4704.115 ;
        RECT 3049.925 4703.835 3050.205 4704.115 ;
        RECT 3050.635 4703.835 3050.915 4704.115 ;
        RECT 3051.345 4703.835 3051.625 4704.115 ;
        RECT 3052.055 4703.835 3052.335 4704.115 ;
        RECT 3052.765 4703.835 3053.045 4704.115 ;
        RECT 3053.475 4703.835 3053.755 4704.115 ;
        RECT 3054.185 4703.835 3054.465 4704.115 ;
        RECT 3054.895 4703.835 3055.175 4704.115 ;
        RECT 3055.605 4703.835 3055.885 4704.115 ;
        RECT 3046.375 4703.125 3046.655 4703.405 ;
        RECT 3047.085 4703.125 3047.365 4703.405 ;
        RECT 3047.795 4703.125 3048.075 4703.405 ;
        RECT 3048.505 4703.125 3048.785 4703.405 ;
        RECT 3049.215 4703.125 3049.495 4703.405 ;
        RECT 3049.925 4703.125 3050.205 4703.405 ;
        RECT 3050.635 4703.125 3050.915 4703.405 ;
        RECT 3051.345 4703.125 3051.625 4703.405 ;
        RECT 3052.055 4703.125 3052.335 4703.405 ;
        RECT 3052.765 4703.125 3053.045 4703.405 ;
        RECT 3053.475 4703.125 3053.755 4703.405 ;
        RECT 3054.185 4703.125 3054.465 4703.405 ;
        RECT 3054.895 4703.125 3055.175 4703.405 ;
        RECT 3055.605 4703.125 3055.885 4703.405 ;
        RECT 3046.375 4702.415 3046.655 4702.695 ;
        RECT 3047.085 4702.415 3047.365 4702.695 ;
        RECT 3047.795 4702.415 3048.075 4702.695 ;
        RECT 3048.505 4702.415 3048.785 4702.695 ;
        RECT 3049.215 4702.415 3049.495 4702.695 ;
        RECT 3049.925 4702.415 3050.205 4702.695 ;
        RECT 3050.635 4702.415 3050.915 4702.695 ;
        RECT 3051.345 4702.415 3051.625 4702.695 ;
        RECT 3052.055 4702.415 3052.335 4702.695 ;
        RECT 3052.765 4702.415 3053.045 4702.695 ;
        RECT 3053.475 4702.415 3053.755 4702.695 ;
        RECT 3054.185 4702.415 3054.465 4702.695 ;
        RECT 3054.895 4702.415 3055.175 4702.695 ;
        RECT 3055.605 4702.415 3055.885 4702.695 ;
        RECT 3046.375 4701.705 3046.655 4701.985 ;
        RECT 3047.085 4701.705 3047.365 4701.985 ;
        RECT 3047.795 4701.705 3048.075 4701.985 ;
        RECT 3048.505 4701.705 3048.785 4701.985 ;
        RECT 3049.215 4701.705 3049.495 4701.985 ;
        RECT 3049.925 4701.705 3050.205 4701.985 ;
        RECT 3050.635 4701.705 3050.915 4701.985 ;
        RECT 3051.345 4701.705 3051.625 4701.985 ;
        RECT 3052.055 4701.705 3052.335 4701.985 ;
        RECT 3052.765 4701.705 3053.045 4701.985 ;
        RECT 3053.475 4701.705 3053.755 4701.985 ;
        RECT 3054.185 4701.705 3054.465 4701.985 ;
        RECT 3054.895 4701.705 3055.175 4701.985 ;
        RECT 3055.605 4701.705 3055.885 4701.985 ;
        RECT 3046.375 4700.995 3046.655 4701.275 ;
        RECT 3047.085 4700.995 3047.365 4701.275 ;
        RECT 3047.795 4700.995 3048.075 4701.275 ;
        RECT 3048.505 4700.995 3048.785 4701.275 ;
        RECT 3049.215 4700.995 3049.495 4701.275 ;
        RECT 3049.925 4700.995 3050.205 4701.275 ;
        RECT 3050.635 4700.995 3050.915 4701.275 ;
        RECT 3051.345 4700.995 3051.625 4701.275 ;
        RECT 3052.055 4700.995 3052.335 4701.275 ;
        RECT 3052.765 4700.995 3053.045 4701.275 ;
        RECT 3053.475 4700.995 3053.755 4701.275 ;
        RECT 3054.185 4700.995 3054.465 4701.275 ;
        RECT 3054.895 4700.995 3055.175 4701.275 ;
        RECT 3055.605 4700.995 3055.885 4701.275 ;
        RECT 3046.375 4700.285 3046.655 4700.565 ;
        RECT 3047.085 4700.285 3047.365 4700.565 ;
        RECT 3047.795 4700.285 3048.075 4700.565 ;
        RECT 3048.505 4700.285 3048.785 4700.565 ;
        RECT 3049.215 4700.285 3049.495 4700.565 ;
        RECT 3049.925 4700.285 3050.205 4700.565 ;
        RECT 3050.635 4700.285 3050.915 4700.565 ;
        RECT 3051.345 4700.285 3051.625 4700.565 ;
        RECT 3052.055 4700.285 3052.335 4700.565 ;
        RECT 3052.765 4700.285 3053.045 4700.565 ;
        RECT 3053.475 4700.285 3053.755 4700.565 ;
        RECT 3054.185 4700.285 3054.465 4700.565 ;
        RECT 3054.895 4700.285 3055.175 4700.565 ;
        RECT 3055.605 4700.285 3055.885 4700.565 ;
        RECT 3046.375 4699.575 3046.655 4699.855 ;
        RECT 3047.085 4699.575 3047.365 4699.855 ;
        RECT 3047.795 4699.575 3048.075 4699.855 ;
        RECT 3048.505 4699.575 3048.785 4699.855 ;
        RECT 3049.215 4699.575 3049.495 4699.855 ;
        RECT 3049.925 4699.575 3050.205 4699.855 ;
        RECT 3050.635 4699.575 3050.915 4699.855 ;
        RECT 3051.345 4699.575 3051.625 4699.855 ;
        RECT 3052.055 4699.575 3052.335 4699.855 ;
        RECT 3052.765 4699.575 3053.045 4699.855 ;
        RECT 3053.475 4699.575 3053.755 4699.855 ;
        RECT 3054.185 4699.575 3054.465 4699.855 ;
        RECT 3054.895 4699.575 3055.175 4699.855 ;
        RECT 3055.605 4699.575 3055.885 4699.855 ;
        RECT 3046.375 4698.865 3046.655 4699.145 ;
        RECT 3047.085 4698.865 3047.365 4699.145 ;
        RECT 3047.795 4698.865 3048.075 4699.145 ;
        RECT 3048.505 4698.865 3048.785 4699.145 ;
        RECT 3049.215 4698.865 3049.495 4699.145 ;
        RECT 3049.925 4698.865 3050.205 4699.145 ;
        RECT 3050.635 4698.865 3050.915 4699.145 ;
        RECT 3051.345 4698.865 3051.625 4699.145 ;
        RECT 3052.055 4698.865 3052.335 4699.145 ;
        RECT 3052.765 4698.865 3053.045 4699.145 ;
        RECT 3053.475 4698.865 3053.755 4699.145 ;
        RECT 3054.185 4698.865 3054.465 4699.145 ;
        RECT 3054.895 4698.865 3055.175 4699.145 ;
        RECT 3055.605 4698.865 3055.885 4699.145 ;
        RECT 3059.485 4708.095 3059.765 4708.375 ;
        RECT 3060.195 4708.095 3060.475 4708.375 ;
        RECT 3060.905 4708.095 3061.185 4708.375 ;
        RECT 3061.615 4708.095 3061.895 4708.375 ;
        RECT 3062.325 4708.095 3062.605 4708.375 ;
        RECT 3063.035 4708.095 3063.315 4708.375 ;
        RECT 3063.745 4708.095 3064.025 4708.375 ;
        RECT 3064.455 4708.095 3064.735 4708.375 ;
        RECT 3065.165 4708.095 3065.445 4708.375 ;
        RECT 3065.875 4708.095 3066.155 4708.375 ;
        RECT 3066.585 4708.095 3066.865 4708.375 ;
        RECT 3067.295 4708.095 3067.575 4708.375 ;
        RECT 3068.005 4708.095 3068.285 4708.375 ;
        RECT 3059.485 4707.385 3059.765 4707.665 ;
        RECT 3060.195 4707.385 3060.475 4707.665 ;
        RECT 3060.905 4707.385 3061.185 4707.665 ;
        RECT 3061.615 4707.385 3061.895 4707.665 ;
        RECT 3062.325 4707.385 3062.605 4707.665 ;
        RECT 3063.035 4707.385 3063.315 4707.665 ;
        RECT 3063.745 4707.385 3064.025 4707.665 ;
        RECT 3064.455 4707.385 3064.735 4707.665 ;
        RECT 3065.165 4707.385 3065.445 4707.665 ;
        RECT 3065.875 4707.385 3066.155 4707.665 ;
        RECT 3066.585 4707.385 3066.865 4707.665 ;
        RECT 3067.295 4707.385 3067.575 4707.665 ;
        RECT 3068.005 4707.385 3068.285 4707.665 ;
        RECT 3059.485 4706.675 3059.765 4706.955 ;
        RECT 3060.195 4706.675 3060.475 4706.955 ;
        RECT 3060.905 4706.675 3061.185 4706.955 ;
        RECT 3061.615 4706.675 3061.895 4706.955 ;
        RECT 3062.325 4706.675 3062.605 4706.955 ;
        RECT 3063.035 4706.675 3063.315 4706.955 ;
        RECT 3063.745 4706.675 3064.025 4706.955 ;
        RECT 3064.455 4706.675 3064.735 4706.955 ;
        RECT 3065.165 4706.675 3065.445 4706.955 ;
        RECT 3065.875 4706.675 3066.155 4706.955 ;
        RECT 3066.585 4706.675 3066.865 4706.955 ;
        RECT 3067.295 4706.675 3067.575 4706.955 ;
        RECT 3068.005 4706.675 3068.285 4706.955 ;
        RECT 3059.485 4705.965 3059.765 4706.245 ;
        RECT 3060.195 4705.965 3060.475 4706.245 ;
        RECT 3060.905 4705.965 3061.185 4706.245 ;
        RECT 3061.615 4705.965 3061.895 4706.245 ;
        RECT 3062.325 4705.965 3062.605 4706.245 ;
        RECT 3063.035 4705.965 3063.315 4706.245 ;
        RECT 3063.745 4705.965 3064.025 4706.245 ;
        RECT 3064.455 4705.965 3064.735 4706.245 ;
        RECT 3065.165 4705.965 3065.445 4706.245 ;
        RECT 3065.875 4705.965 3066.155 4706.245 ;
        RECT 3066.585 4705.965 3066.865 4706.245 ;
        RECT 3067.295 4705.965 3067.575 4706.245 ;
        RECT 3068.005 4705.965 3068.285 4706.245 ;
        RECT 3059.485 4705.255 3059.765 4705.535 ;
        RECT 3060.195 4705.255 3060.475 4705.535 ;
        RECT 3060.905 4705.255 3061.185 4705.535 ;
        RECT 3061.615 4705.255 3061.895 4705.535 ;
        RECT 3062.325 4705.255 3062.605 4705.535 ;
        RECT 3063.035 4705.255 3063.315 4705.535 ;
        RECT 3063.745 4705.255 3064.025 4705.535 ;
        RECT 3064.455 4705.255 3064.735 4705.535 ;
        RECT 3065.165 4705.255 3065.445 4705.535 ;
        RECT 3065.875 4705.255 3066.155 4705.535 ;
        RECT 3066.585 4705.255 3066.865 4705.535 ;
        RECT 3067.295 4705.255 3067.575 4705.535 ;
        RECT 3068.005 4705.255 3068.285 4705.535 ;
        RECT 3059.485 4704.545 3059.765 4704.825 ;
        RECT 3060.195 4704.545 3060.475 4704.825 ;
        RECT 3060.905 4704.545 3061.185 4704.825 ;
        RECT 3061.615 4704.545 3061.895 4704.825 ;
        RECT 3062.325 4704.545 3062.605 4704.825 ;
        RECT 3063.035 4704.545 3063.315 4704.825 ;
        RECT 3063.745 4704.545 3064.025 4704.825 ;
        RECT 3064.455 4704.545 3064.735 4704.825 ;
        RECT 3065.165 4704.545 3065.445 4704.825 ;
        RECT 3065.875 4704.545 3066.155 4704.825 ;
        RECT 3066.585 4704.545 3066.865 4704.825 ;
        RECT 3067.295 4704.545 3067.575 4704.825 ;
        RECT 3068.005 4704.545 3068.285 4704.825 ;
        RECT 3059.485 4703.835 3059.765 4704.115 ;
        RECT 3060.195 4703.835 3060.475 4704.115 ;
        RECT 3060.905 4703.835 3061.185 4704.115 ;
        RECT 3061.615 4703.835 3061.895 4704.115 ;
        RECT 3062.325 4703.835 3062.605 4704.115 ;
        RECT 3063.035 4703.835 3063.315 4704.115 ;
        RECT 3063.745 4703.835 3064.025 4704.115 ;
        RECT 3064.455 4703.835 3064.735 4704.115 ;
        RECT 3065.165 4703.835 3065.445 4704.115 ;
        RECT 3065.875 4703.835 3066.155 4704.115 ;
        RECT 3066.585 4703.835 3066.865 4704.115 ;
        RECT 3067.295 4703.835 3067.575 4704.115 ;
        RECT 3068.005 4703.835 3068.285 4704.115 ;
        RECT 3059.485 4703.125 3059.765 4703.405 ;
        RECT 3060.195 4703.125 3060.475 4703.405 ;
        RECT 3060.905 4703.125 3061.185 4703.405 ;
        RECT 3061.615 4703.125 3061.895 4703.405 ;
        RECT 3062.325 4703.125 3062.605 4703.405 ;
        RECT 3063.035 4703.125 3063.315 4703.405 ;
        RECT 3063.745 4703.125 3064.025 4703.405 ;
        RECT 3064.455 4703.125 3064.735 4703.405 ;
        RECT 3065.165 4703.125 3065.445 4703.405 ;
        RECT 3065.875 4703.125 3066.155 4703.405 ;
        RECT 3066.585 4703.125 3066.865 4703.405 ;
        RECT 3067.295 4703.125 3067.575 4703.405 ;
        RECT 3068.005 4703.125 3068.285 4703.405 ;
        RECT 3059.485 4702.415 3059.765 4702.695 ;
        RECT 3060.195 4702.415 3060.475 4702.695 ;
        RECT 3060.905 4702.415 3061.185 4702.695 ;
        RECT 3061.615 4702.415 3061.895 4702.695 ;
        RECT 3062.325 4702.415 3062.605 4702.695 ;
        RECT 3063.035 4702.415 3063.315 4702.695 ;
        RECT 3063.745 4702.415 3064.025 4702.695 ;
        RECT 3064.455 4702.415 3064.735 4702.695 ;
        RECT 3065.165 4702.415 3065.445 4702.695 ;
        RECT 3065.875 4702.415 3066.155 4702.695 ;
        RECT 3066.585 4702.415 3066.865 4702.695 ;
        RECT 3067.295 4702.415 3067.575 4702.695 ;
        RECT 3068.005 4702.415 3068.285 4702.695 ;
        RECT 3059.485 4701.705 3059.765 4701.985 ;
        RECT 3060.195 4701.705 3060.475 4701.985 ;
        RECT 3060.905 4701.705 3061.185 4701.985 ;
        RECT 3061.615 4701.705 3061.895 4701.985 ;
        RECT 3062.325 4701.705 3062.605 4701.985 ;
        RECT 3063.035 4701.705 3063.315 4701.985 ;
        RECT 3063.745 4701.705 3064.025 4701.985 ;
        RECT 3064.455 4701.705 3064.735 4701.985 ;
        RECT 3065.165 4701.705 3065.445 4701.985 ;
        RECT 3065.875 4701.705 3066.155 4701.985 ;
        RECT 3066.585 4701.705 3066.865 4701.985 ;
        RECT 3067.295 4701.705 3067.575 4701.985 ;
        RECT 3068.005 4701.705 3068.285 4701.985 ;
        RECT 3059.485 4700.995 3059.765 4701.275 ;
        RECT 3060.195 4700.995 3060.475 4701.275 ;
        RECT 3060.905 4700.995 3061.185 4701.275 ;
        RECT 3061.615 4700.995 3061.895 4701.275 ;
        RECT 3062.325 4700.995 3062.605 4701.275 ;
        RECT 3063.035 4700.995 3063.315 4701.275 ;
        RECT 3063.745 4700.995 3064.025 4701.275 ;
        RECT 3064.455 4700.995 3064.735 4701.275 ;
        RECT 3065.165 4700.995 3065.445 4701.275 ;
        RECT 3065.875 4700.995 3066.155 4701.275 ;
        RECT 3066.585 4700.995 3066.865 4701.275 ;
        RECT 3067.295 4700.995 3067.575 4701.275 ;
        RECT 3068.005 4700.995 3068.285 4701.275 ;
        RECT 3059.485 4700.285 3059.765 4700.565 ;
        RECT 3060.195 4700.285 3060.475 4700.565 ;
        RECT 3060.905 4700.285 3061.185 4700.565 ;
        RECT 3061.615 4700.285 3061.895 4700.565 ;
        RECT 3062.325 4700.285 3062.605 4700.565 ;
        RECT 3063.035 4700.285 3063.315 4700.565 ;
        RECT 3063.745 4700.285 3064.025 4700.565 ;
        RECT 3064.455 4700.285 3064.735 4700.565 ;
        RECT 3065.165 4700.285 3065.445 4700.565 ;
        RECT 3065.875 4700.285 3066.155 4700.565 ;
        RECT 3066.585 4700.285 3066.865 4700.565 ;
        RECT 3067.295 4700.285 3067.575 4700.565 ;
        RECT 3068.005 4700.285 3068.285 4700.565 ;
        RECT 3059.485 4699.575 3059.765 4699.855 ;
        RECT 3060.195 4699.575 3060.475 4699.855 ;
        RECT 3060.905 4699.575 3061.185 4699.855 ;
        RECT 3061.615 4699.575 3061.895 4699.855 ;
        RECT 3062.325 4699.575 3062.605 4699.855 ;
        RECT 3063.035 4699.575 3063.315 4699.855 ;
        RECT 3063.745 4699.575 3064.025 4699.855 ;
        RECT 3064.455 4699.575 3064.735 4699.855 ;
        RECT 3065.165 4699.575 3065.445 4699.855 ;
        RECT 3065.875 4699.575 3066.155 4699.855 ;
        RECT 3066.585 4699.575 3066.865 4699.855 ;
        RECT 3067.295 4699.575 3067.575 4699.855 ;
        RECT 3068.005 4699.575 3068.285 4699.855 ;
        RECT 3059.485 4698.865 3059.765 4699.145 ;
        RECT 3060.195 4698.865 3060.475 4699.145 ;
        RECT 3060.905 4698.865 3061.185 4699.145 ;
        RECT 3061.615 4698.865 3061.895 4699.145 ;
        RECT 3062.325 4698.865 3062.605 4699.145 ;
        RECT 3063.035 4698.865 3063.315 4699.145 ;
        RECT 3063.745 4698.865 3064.025 4699.145 ;
        RECT 3064.455 4698.865 3064.735 4699.145 ;
        RECT 3065.165 4698.865 3065.445 4699.145 ;
        RECT 3065.875 4698.865 3066.155 4699.145 ;
        RECT 3066.585 4698.865 3066.865 4699.145 ;
        RECT 3067.295 4698.865 3067.575 4699.145 ;
        RECT 3068.005 4698.865 3068.285 4699.145 ;
        RECT 369.330 4392.970 369.610 4393.250 ;
        RECT 370.040 4392.970 370.320 4393.250 ;
        RECT 370.750 4392.970 371.030 4393.250 ;
        RECT 371.460 4392.970 371.740 4393.250 ;
        RECT 372.170 4392.970 372.450 4393.250 ;
        RECT 372.880 4392.970 373.160 4393.250 ;
        RECT 373.590 4392.970 373.870 4393.250 ;
        RECT 374.300 4392.970 374.580 4393.250 ;
        RECT 375.010 4392.970 375.290 4393.250 ;
        RECT 375.720 4392.970 376.000 4393.250 ;
        RECT 376.430 4392.970 376.710 4393.250 ;
        RECT 377.140 4392.970 377.420 4393.250 ;
        RECT 377.850 4392.970 378.130 4393.250 ;
        RECT 378.560 4392.970 378.840 4393.250 ;
        RECT 369.330 4392.260 369.610 4392.540 ;
        RECT 370.040 4392.260 370.320 4392.540 ;
        RECT 370.750 4392.260 371.030 4392.540 ;
        RECT 371.460 4392.260 371.740 4392.540 ;
        RECT 372.170 4392.260 372.450 4392.540 ;
        RECT 372.880 4392.260 373.160 4392.540 ;
        RECT 373.590 4392.260 373.870 4392.540 ;
        RECT 374.300 4392.260 374.580 4392.540 ;
        RECT 375.010 4392.260 375.290 4392.540 ;
        RECT 375.720 4392.260 376.000 4392.540 ;
        RECT 376.430 4392.260 376.710 4392.540 ;
        RECT 377.140 4392.260 377.420 4392.540 ;
        RECT 377.850 4392.260 378.130 4392.540 ;
        RECT 378.560 4392.260 378.840 4392.540 ;
        RECT 369.330 4391.550 369.610 4391.830 ;
        RECT 370.040 4391.550 370.320 4391.830 ;
        RECT 370.750 4391.550 371.030 4391.830 ;
        RECT 371.460 4391.550 371.740 4391.830 ;
        RECT 372.170 4391.550 372.450 4391.830 ;
        RECT 372.880 4391.550 373.160 4391.830 ;
        RECT 373.590 4391.550 373.870 4391.830 ;
        RECT 374.300 4391.550 374.580 4391.830 ;
        RECT 375.010 4391.550 375.290 4391.830 ;
        RECT 375.720 4391.550 376.000 4391.830 ;
        RECT 376.430 4391.550 376.710 4391.830 ;
        RECT 377.140 4391.550 377.420 4391.830 ;
        RECT 377.850 4391.550 378.130 4391.830 ;
        RECT 378.560 4391.550 378.840 4391.830 ;
        RECT 369.330 4390.840 369.610 4391.120 ;
        RECT 370.040 4390.840 370.320 4391.120 ;
        RECT 370.750 4390.840 371.030 4391.120 ;
        RECT 371.460 4390.840 371.740 4391.120 ;
        RECT 372.170 4390.840 372.450 4391.120 ;
        RECT 372.880 4390.840 373.160 4391.120 ;
        RECT 373.590 4390.840 373.870 4391.120 ;
        RECT 374.300 4390.840 374.580 4391.120 ;
        RECT 375.010 4390.840 375.290 4391.120 ;
        RECT 375.720 4390.840 376.000 4391.120 ;
        RECT 376.430 4390.840 376.710 4391.120 ;
        RECT 377.140 4390.840 377.420 4391.120 ;
        RECT 377.850 4390.840 378.130 4391.120 ;
        RECT 378.560 4390.840 378.840 4391.120 ;
        RECT 369.330 4390.130 369.610 4390.410 ;
        RECT 370.040 4390.130 370.320 4390.410 ;
        RECT 370.750 4390.130 371.030 4390.410 ;
        RECT 371.460 4390.130 371.740 4390.410 ;
        RECT 372.170 4390.130 372.450 4390.410 ;
        RECT 372.880 4390.130 373.160 4390.410 ;
        RECT 373.590 4390.130 373.870 4390.410 ;
        RECT 374.300 4390.130 374.580 4390.410 ;
        RECT 375.010 4390.130 375.290 4390.410 ;
        RECT 375.720 4390.130 376.000 4390.410 ;
        RECT 376.430 4390.130 376.710 4390.410 ;
        RECT 377.140 4390.130 377.420 4390.410 ;
        RECT 377.850 4390.130 378.130 4390.410 ;
        RECT 378.560 4390.130 378.840 4390.410 ;
        RECT 369.330 4389.420 369.610 4389.700 ;
        RECT 370.040 4389.420 370.320 4389.700 ;
        RECT 370.750 4389.420 371.030 4389.700 ;
        RECT 371.460 4389.420 371.740 4389.700 ;
        RECT 372.170 4389.420 372.450 4389.700 ;
        RECT 372.880 4389.420 373.160 4389.700 ;
        RECT 373.590 4389.420 373.870 4389.700 ;
        RECT 374.300 4389.420 374.580 4389.700 ;
        RECT 375.010 4389.420 375.290 4389.700 ;
        RECT 375.720 4389.420 376.000 4389.700 ;
        RECT 376.430 4389.420 376.710 4389.700 ;
        RECT 377.140 4389.420 377.420 4389.700 ;
        RECT 377.850 4389.420 378.130 4389.700 ;
        RECT 378.560 4389.420 378.840 4389.700 ;
        RECT 369.330 4388.710 369.610 4388.990 ;
        RECT 370.040 4388.710 370.320 4388.990 ;
        RECT 370.750 4388.710 371.030 4388.990 ;
        RECT 371.460 4388.710 371.740 4388.990 ;
        RECT 372.170 4388.710 372.450 4388.990 ;
        RECT 372.880 4388.710 373.160 4388.990 ;
        RECT 373.590 4388.710 373.870 4388.990 ;
        RECT 374.300 4388.710 374.580 4388.990 ;
        RECT 375.010 4388.710 375.290 4388.990 ;
        RECT 375.720 4388.710 376.000 4388.990 ;
        RECT 376.430 4388.710 376.710 4388.990 ;
        RECT 377.140 4388.710 377.420 4388.990 ;
        RECT 377.850 4388.710 378.130 4388.990 ;
        RECT 378.560 4388.710 378.840 4388.990 ;
        RECT 369.330 4388.000 369.610 4388.280 ;
        RECT 370.040 4388.000 370.320 4388.280 ;
        RECT 370.750 4388.000 371.030 4388.280 ;
        RECT 371.460 4388.000 371.740 4388.280 ;
        RECT 372.170 4388.000 372.450 4388.280 ;
        RECT 372.880 4388.000 373.160 4388.280 ;
        RECT 373.590 4388.000 373.870 4388.280 ;
        RECT 374.300 4388.000 374.580 4388.280 ;
        RECT 375.010 4388.000 375.290 4388.280 ;
        RECT 375.720 4388.000 376.000 4388.280 ;
        RECT 376.430 4388.000 376.710 4388.280 ;
        RECT 377.140 4388.000 377.420 4388.280 ;
        RECT 377.850 4388.000 378.130 4388.280 ;
        RECT 378.560 4388.000 378.840 4388.280 ;
        RECT 369.330 4387.290 369.610 4387.570 ;
        RECT 370.040 4387.290 370.320 4387.570 ;
        RECT 370.750 4387.290 371.030 4387.570 ;
        RECT 371.460 4387.290 371.740 4387.570 ;
        RECT 372.170 4387.290 372.450 4387.570 ;
        RECT 372.880 4387.290 373.160 4387.570 ;
        RECT 373.590 4387.290 373.870 4387.570 ;
        RECT 374.300 4387.290 374.580 4387.570 ;
        RECT 375.010 4387.290 375.290 4387.570 ;
        RECT 375.720 4387.290 376.000 4387.570 ;
        RECT 376.430 4387.290 376.710 4387.570 ;
        RECT 377.140 4387.290 377.420 4387.570 ;
        RECT 377.850 4387.290 378.130 4387.570 ;
        RECT 378.560 4387.290 378.840 4387.570 ;
        RECT 369.330 4386.580 369.610 4386.860 ;
        RECT 370.040 4386.580 370.320 4386.860 ;
        RECT 370.750 4386.580 371.030 4386.860 ;
        RECT 371.460 4386.580 371.740 4386.860 ;
        RECT 372.170 4386.580 372.450 4386.860 ;
        RECT 372.880 4386.580 373.160 4386.860 ;
        RECT 373.590 4386.580 373.870 4386.860 ;
        RECT 374.300 4386.580 374.580 4386.860 ;
        RECT 375.010 4386.580 375.290 4386.860 ;
        RECT 375.720 4386.580 376.000 4386.860 ;
        RECT 376.430 4386.580 376.710 4386.860 ;
        RECT 377.140 4386.580 377.420 4386.860 ;
        RECT 377.850 4386.580 378.130 4386.860 ;
        RECT 378.560 4386.580 378.840 4386.860 ;
        RECT 369.330 4385.870 369.610 4386.150 ;
        RECT 370.040 4385.870 370.320 4386.150 ;
        RECT 370.750 4385.870 371.030 4386.150 ;
        RECT 371.460 4385.870 371.740 4386.150 ;
        RECT 372.170 4385.870 372.450 4386.150 ;
        RECT 372.880 4385.870 373.160 4386.150 ;
        RECT 373.590 4385.870 373.870 4386.150 ;
        RECT 374.300 4385.870 374.580 4386.150 ;
        RECT 375.010 4385.870 375.290 4386.150 ;
        RECT 375.720 4385.870 376.000 4386.150 ;
        RECT 376.430 4385.870 376.710 4386.150 ;
        RECT 377.140 4385.870 377.420 4386.150 ;
        RECT 377.850 4385.870 378.130 4386.150 ;
        RECT 378.560 4385.870 378.840 4386.150 ;
        RECT 369.330 4385.160 369.610 4385.440 ;
        RECT 370.040 4385.160 370.320 4385.440 ;
        RECT 370.750 4385.160 371.030 4385.440 ;
        RECT 371.460 4385.160 371.740 4385.440 ;
        RECT 372.170 4385.160 372.450 4385.440 ;
        RECT 372.880 4385.160 373.160 4385.440 ;
        RECT 373.590 4385.160 373.870 4385.440 ;
        RECT 374.300 4385.160 374.580 4385.440 ;
        RECT 375.010 4385.160 375.290 4385.440 ;
        RECT 375.720 4385.160 376.000 4385.440 ;
        RECT 376.430 4385.160 376.710 4385.440 ;
        RECT 377.140 4385.160 377.420 4385.440 ;
        RECT 377.850 4385.160 378.130 4385.440 ;
        RECT 378.560 4385.160 378.840 4385.440 ;
        RECT 369.330 4384.450 369.610 4384.730 ;
        RECT 370.040 4384.450 370.320 4384.730 ;
        RECT 370.750 4384.450 371.030 4384.730 ;
        RECT 371.460 4384.450 371.740 4384.730 ;
        RECT 372.170 4384.450 372.450 4384.730 ;
        RECT 372.880 4384.450 373.160 4384.730 ;
        RECT 373.590 4384.450 373.870 4384.730 ;
        RECT 374.300 4384.450 374.580 4384.730 ;
        RECT 375.010 4384.450 375.290 4384.730 ;
        RECT 375.720 4384.450 376.000 4384.730 ;
        RECT 376.430 4384.450 376.710 4384.730 ;
        RECT 377.140 4384.450 377.420 4384.730 ;
        RECT 377.850 4384.450 378.130 4384.730 ;
        RECT 378.560 4384.450 378.840 4384.730 ;
        RECT 3500.200 4388.050 3500.480 4388.330 ;
        RECT 3500.910 4388.050 3501.190 4388.330 ;
        RECT 3501.620 4388.050 3501.900 4388.330 ;
        RECT 3502.330 4388.050 3502.610 4388.330 ;
        RECT 3503.040 4388.050 3503.320 4388.330 ;
        RECT 3503.750 4388.050 3504.030 4388.330 ;
        RECT 3504.460 4388.050 3504.740 4388.330 ;
        RECT 3505.170 4388.050 3505.450 4388.330 ;
        RECT 3505.880 4388.050 3506.160 4388.330 ;
        RECT 3506.590 4388.050 3506.870 4388.330 ;
        RECT 3507.300 4388.050 3507.580 4388.330 ;
        RECT 3508.010 4388.050 3508.290 4388.330 ;
        RECT 3508.720 4388.050 3509.000 4388.330 ;
        RECT 3509.430 4388.050 3509.710 4388.330 ;
        RECT 3500.200 4387.340 3500.480 4387.620 ;
        RECT 3500.910 4387.340 3501.190 4387.620 ;
        RECT 3501.620 4387.340 3501.900 4387.620 ;
        RECT 3502.330 4387.340 3502.610 4387.620 ;
        RECT 3503.040 4387.340 3503.320 4387.620 ;
        RECT 3503.750 4387.340 3504.030 4387.620 ;
        RECT 3504.460 4387.340 3504.740 4387.620 ;
        RECT 3505.170 4387.340 3505.450 4387.620 ;
        RECT 3505.880 4387.340 3506.160 4387.620 ;
        RECT 3506.590 4387.340 3506.870 4387.620 ;
        RECT 3507.300 4387.340 3507.580 4387.620 ;
        RECT 3508.010 4387.340 3508.290 4387.620 ;
        RECT 3508.720 4387.340 3509.000 4387.620 ;
        RECT 3509.430 4387.340 3509.710 4387.620 ;
        RECT 3500.200 4386.630 3500.480 4386.910 ;
        RECT 3500.910 4386.630 3501.190 4386.910 ;
        RECT 3501.620 4386.630 3501.900 4386.910 ;
        RECT 3502.330 4386.630 3502.610 4386.910 ;
        RECT 3503.040 4386.630 3503.320 4386.910 ;
        RECT 3503.750 4386.630 3504.030 4386.910 ;
        RECT 3504.460 4386.630 3504.740 4386.910 ;
        RECT 3505.170 4386.630 3505.450 4386.910 ;
        RECT 3505.880 4386.630 3506.160 4386.910 ;
        RECT 3506.590 4386.630 3506.870 4386.910 ;
        RECT 3507.300 4386.630 3507.580 4386.910 ;
        RECT 3508.010 4386.630 3508.290 4386.910 ;
        RECT 3508.720 4386.630 3509.000 4386.910 ;
        RECT 3509.430 4386.630 3509.710 4386.910 ;
        RECT 3500.200 4385.920 3500.480 4386.200 ;
        RECT 3500.910 4385.920 3501.190 4386.200 ;
        RECT 3501.620 4385.920 3501.900 4386.200 ;
        RECT 3502.330 4385.920 3502.610 4386.200 ;
        RECT 3503.040 4385.920 3503.320 4386.200 ;
        RECT 3503.750 4385.920 3504.030 4386.200 ;
        RECT 3504.460 4385.920 3504.740 4386.200 ;
        RECT 3505.170 4385.920 3505.450 4386.200 ;
        RECT 3505.880 4385.920 3506.160 4386.200 ;
        RECT 3506.590 4385.920 3506.870 4386.200 ;
        RECT 3507.300 4385.920 3507.580 4386.200 ;
        RECT 3508.010 4385.920 3508.290 4386.200 ;
        RECT 3508.720 4385.920 3509.000 4386.200 ;
        RECT 3509.430 4385.920 3509.710 4386.200 ;
        RECT 3500.200 4385.210 3500.480 4385.490 ;
        RECT 3500.910 4385.210 3501.190 4385.490 ;
        RECT 3501.620 4385.210 3501.900 4385.490 ;
        RECT 3502.330 4385.210 3502.610 4385.490 ;
        RECT 3503.040 4385.210 3503.320 4385.490 ;
        RECT 3503.750 4385.210 3504.030 4385.490 ;
        RECT 3504.460 4385.210 3504.740 4385.490 ;
        RECT 3505.170 4385.210 3505.450 4385.490 ;
        RECT 3505.880 4385.210 3506.160 4385.490 ;
        RECT 3506.590 4385.210 3506.870 4385.490 ;
        RECT 3507.300 4385.210 3507.580 4385.490 ;
        RECT 3508.010 4385.210 3508.290 4385.490 ;
        RECT 3508.720 4385.210 3509.000 4385.490 ;
        RECT 3509.430 4385.210 3509.710 4385.490 ;
        RECT 3500.200 4384.500 3500.480 4384.780 ;
        RECT 3500.910 4384.500 3501.190 4384.780 ;
        RECT 3501.620 4384.500 3501.900 4384.780 ;
        RECT 3502.330 4384.500 3502.610 4384.780 ;
        RECT 3503.040 4384.500 3503.320 4384.780 ;
        RECT 3503.750 4384.500 3504.030 4384.780 ;
        RECT 3504.460 4384.500 3504.740 4384.780 ;
        RECT 3505.170 4384.500 3505.450 4384.780 ;
        RECT 3505.880 4384.500 3506.160 4384.780 ;
        RECT 3506.590 4384.500 3506.870 4384.780 ;
        RECT 3507.300 4384.500 3507.580 4384.780 ;
        RECT 3508.010 4384.500 3508.290 4384.780 ;
        RECT 3508.720 4384.500 3509.000 4384.780 ;
        RECT 3509.430 4384.500 3509.710 4384.780 ;
        RECT 3500.200 4383.790 3500.480 4384.070 ;
        RECT 3500.910 4383.790 3501.190 4384.070 ;
        RECT 3501.620 4383.790 3501.900 4384.070 ;
        RECT 3502.330 4383.790 3502.610 4384.070 ;
        RECT 3503.040 4383.790 3503.320 4384.070 ;
        RECT 3503.750 4383.790 3504.030 4384.070 ;
        RECT 3504.460 4383.790 3504.740 4384.070 ;
        RECT 3505.170 4383.790 3505.450 4384.070 ;
        RECT 3505.880 4383.790 3506.160 4384.070 ;
        RECT 3506.590 4383.790 3506.870 4384.070 ;
        RECT 3507.300 4383.790 3507.580 4384.070 ;
        RECT 3508.010 4383.790 3508.290 4384.070 ;
        RECT 3508.720 4383.790 3509.000 4384.070 ;
        RECT 3509.430 4383.790 3509.710 4384.070 ;
        RECT 3500.200 4383.080 3500.480 4383.360 ;
        RECT 3500.910 4383.080 3501.190 4383.360 ;
        RECT 3501.620 4383.080 3501.900 4383.360 ;
        RECT 3502.330 4383.080 3502.610 4383.360 ;
        RECT 3503.040 4383.080 3503.320 4383.360 ;
        RECT 3503.750 4383.080 3504.030 4383.360 ;
        RECT 3504.460 4383.080 3504.740 4383.360 ;
        RECT 3505.170 4383.080 3505.450 4383.360 ;
        RECT 3505.880 4383.080 3506.160 4383.360 ;
        RECT 3506.590 4383.080 3506.870 4383.360 ;
        RECT 3507.300 4383.080 3507.580 4383.360 ;
        RECT 3508.010 4383.080 3508.290 4383.360 ;
        RECT 3508.720 4383.080 3509.000 4383.360 ;
        RECT 3509.430 4383.080 3509.710 4383.360 ;
        RECT 3500.200 4382.370 3500.480 4382.650 ;
        RECT 3500.910 4382.370 3501.190 4382.650 ;
        RECT 3501.620 4382.370 3501.900 4382.650 ;
        RECT 3502.330 4382.370 3502.610 4382.650 ;
        RECT 3503.040 4382.370 3503.320 4382.650 ;
        RECT 3503.750 4382.370 3504.030 4382.650 ;
        RECT 3504.460 4382.370 3504.740 4382.650 ;
        RECT 3505.170 4382.370 3505.450 4382.650 ;
        RECT 3505.880 4382.370 3506.160 4382.650 ;
        RECT 3506.590 4382.370 3506.870 4382.650 ;
        RECT 3507.300 4382.370 3507.580 4382.650 ;
        RECT 3508.010 4382.370 3508.290 4382.650 ;
        RECT 3508.720 4382.370 3509.000 4382.650 ;
        RECT 3509.430 4382.370 3509.710 4382.650 ;
        RECT 3500.200 4381.660 3500.480 4381.940 ;
        RECT 3500.910 4381.660 3501.190 4381.940 ;
        RECT 3501.620 4381.660 3501.900 4381.940 ;
        RECT 3502.330 4381.660 3502.610 4381.940 ;
        RECT 3503.040 4381.660 3503.320 4381.940 ;
        RECT 3503.750 4381.660 3504.030 4381.940 ;
        RECT 3504.460 4381.660 3504.740 4381.940 ;
        RECT 3505.170 4381.660 3505.450 4381.940 ;
        RECT 3505.880 4381.660 3506.160 4381.940 ;
        RECT 3506.590 4381.660 3506.870 4381.940 ;
        RECT 3507.300 4381.660 3507.580 4381.940 ;
        RECT 3508.010 4381.660 3508.290 4381.940 ;
        RECT 3508.720 4381.660 3509.000 4381.940 ;
        RECT 3509.430 4381.660 3509.710 4381.940 ;
        RECT 369.275 4380.565 369.555 4380.845 ;
        RECT 369.985 4380.565 370.265 4380.845 ;
        RECT 370.695 4380.565 370.975 4380.845 ;
        RECT 371.405 4380.565 371.685 4380.845 ;
        RECT 372.115 4380.565 372.395 4380.845 ;
        RECT 372.825 4380.565 373.105 4380.845 ;
        RECT 373.535 4380.565 373.815 4380.845 ;
        RECT 374.245 4380.565 374.525 4380.845 ;
        RECT 374.955 4380.565 375.235 4380.845 ;
        RECT 375.665 4380.565 375.945 4380.845 ;
        RECT 376.375 4380.565 376.655 4380.845 ;
        RECT 377.085 4380.565 377.365 4380.845 ;
        RECT 377.795 4380.565 378.075 4380.845 ;
        RECT 378.505 4380.565 378.785 4380.845 ;
        RECT 369.275 4379.855 369.555 4380.135 ;
        RECT 369.985 4379.855 370.265 4380.135 ;
        RECT 370.695 4379.855 370.975 4380.135 ;
        RECT 371.405 4379.855 371.685 4380.135 ;
        RECT 372.115 4379.855 372.395 4380.135 ;
        RECT 372.825 4379.855 373.105 4380.135 ;
        RECT 373.535 4379.855 373.815 4380.135 ;
        RECT 374.245 4379.855 374.525 4380.135 ;
        RECT 374.955 4379.855 375.235 4380.135 ;
        RECT 375.665 4379.855 375.945 4380.135 ;
        RECT 376.375 4379.855 376.655 4380.135 ;
        RECT 377.085 4379.855 377.365 4380.135 ;
        RECT 377.795 4379.855 378.075 4380.135 ;
        RECT 378.505 4379.855 378.785 4380.135 ;
        RECT 369.275 4379.145 369.555 4379.425 ;
        RECT 369.985 4379.145 370.265 4379.425 ;
        RECT 370.695 4379.145 370.975 4379.425 ;
        RECT 371.405 4379.145 371.685 4379.425 ;
        RECT 372.115 4379.145 372.395 4379.425 ;
        RECT 372.825 4379.145 373.105 4379.425 ;
        RECT 373.535 4379.145 373.815 4379.425 ;
        RECT 374.245 4379.145 374.525 4379.425 ;
        RECT 374.955 4379.145 375.235 4379.425 ;
        RECT 375.665 4379.145 375.945 4379.425 ;
        RECT 376.375 4379.145 376.655 4379.425 ;
        RECT 377.085 4379.145 377.365 4379.425 ;
        RECT 377.795 4379.145 378.075 4379.425 ;
        RECT 378.505 4379.145 378.785 4379.425 ;
        RECT 3500.200 4380.950 3500.480 4381.230 ;
        RECT 3500.910 4380.950 3501.190 4381.230 ;
        RECT 3501.620 4380.950 3501.900 4381.230 ;
        RECT 3502.330 4380.950 3502.610 4381.230 ;
        RECT 3503.040 4380.950 3503.320 4381.230 ;
        RECT 3503.750 4380.950 3504.030 4381.230 ;
        RECT 3504.460 4380.950 3504.740 4381.230 ;
        RECT 3505.170 4380.950 3505.450 4381.230 ;
        RECT 3505.880 4380.950 3506.160 4381.230 ;
        RECT 3506.590 4380.950 3506.870 4381.230 ;
        RECT 3507.300 4380.950 3507.580 4381.230 ;
        RECT 3508.010 4380.950 3508.290 4381.230 ;
        RECT 3508.720 4380.950 3509.000 4381.230 ;
        RECT 3509.430 4380.950 3509.710 4381.230 ;
        RECT 3500.200 4380.240 3500.480 4380.520 ;
        RECT 3500.910 4380.240 3501.190 4380.520 ;
        RECT 3501.620 4380.240 3501.900 4380.520 ;
        RECT 3502.330 4380.240 3502.610 4380.520 ;
        RECT 3503.040 4380.240 3503.320 4380.520 ;
        RECT 3503.750 4380.240 3504.030 4380.520 ;
        RECT 3504.460 4380.240 3504.740 4380.520 ;
        RECT 3505.170 4380.240 3505.450 4380.520 ;
        RECT 3505.880 4380.240 3506.160 4380.520 ;
        RECT 3506.590 4380.240 3506.870 4380.520 ;
        RECT 3507.300 4380.240 3507.580 4380.520 ;
        RECT 3508.010 4380.240 3508.290 4380.520 ;
        RECT 3508.720 4380.240 3509.000 4380.520 ;
        RECT 3509.430 4380.240 3509.710 4380.520 ;
        RECT 3500.200 4379.530 3500.480 4379.810 ;
        RECT 3500.910 4379.530 3501.190 4379.810 ;
        RECT 3501.620 4379.530 3501.900 4379.810 ;
        RECT 3502.330 4379.530 3502.610 4379.810 ;
        RECT 3503.040 4379.530 3503.320 4379.810 ;
        RECT 3503.750 4379.530 3504.030 4379.810 ;
        RECT 3504.460 4379.530 3504.740 4379.810 ;
        RECT 3505.170 4379.530 3505.450 4379.810 ;
        RECT 3505.880 4379.530 3506.160 4379.810 ;
        RECT 3506.590 4379.530 3506.870 4379.810 ;
        RECT 3507.300 4379.530 3507.580 4379.810 ;
        RECT 3508.010 4379.530 3508.290 4379.810 ;
        RECT 3508.720 4379.530 3509.000 4379.810 ;
        RECT 3509.430 4379.530 3509.710 4379.810 ;
        RECT 369.275 4378.435 369.555 4378.715 ;
        RECT 369.985 4378.435 370.265 4378.715 ;
        RECT 370.695 4378.435 370.975 4378.715 ;
        RECT 371.405 4378.435 371.685 4378.715 ;
        RECT 372.115 4378.435 372.395 4378.715 ;
        RECT 372.825 4378.435 373.105 4378.715 ;
        RECT 373.535 4378.435 373.815 4378.715 ;
        RECT 374.245 4378.435 374.525 4378.715 ;
        RECT 374.955 4378.435 375.235 4378.715 ;
        RECT 375.665 4378.435 375.945 4378.715 ;
        RECT 376.375 4378.435 376.655 4378.715 ;
        RECT 377.085 4378.435 377.365 4378.715 ;
        RECT 377.795 4378.435 378.075 4378.715 ;
        RECT 378.505 4378.435 378.785 4378.715 ;
        RECT 369.275 4377.725 369.555 4378.005 ;
        RECT 369.985 4377.725 370.265 4378.005 ;
        RECT 370.695 4377.725 370.975 4378.005 ;
        RECT 371.405 4377.725 371.685 4378.005 ;
        RECT 372.115 4377.725 372.395 4378.005 ;
        RECT 372.825 4377.725 373.105 4378.005 ;
        RECT 373.535 4377.725 373.815 4378.005 ;
        RECT 374.245 4377.725 374.525 4378.005 ;
        RECT 374.955 4377.725 375.235 4378.005 ;
        RECT 375.665 4377.725 375.945 4378.005 ;
        RECT 376.375 4377.725 376.655 4378.005 ;
        RECT 377.085 4377.725 377.365 4378.005 ;
        RECT 377.795 4377.725 378.075 4378.005 ;
        RECT 378.505 4377.725 378.785 4378.005 ;
        RECT 369.275 4377.015 369.555 4377.295 ;
        RECT 369.985 4377.015 370.265 4377.295 ;
        RECT 370.695 4377.015 370.975 4377.295 ;
        RECT 371.405 4377.015 371.685 4377.295 ;
        RECT 372.115 4377.015 372.395 4377.295 ;
        RECT 372.825 4377.015 373.105 4377.295 ;
        RECT 373.535 4377.015 373.815 4377.295 ;
        RECT 374.245 4377.015 374.525 4377.295 ;
        RECT 374.955 4377.015 375.235 4377.295 ;
        RECT 375.665 4377.015 375.945 4377.295 ;
        RECT 376.375 4377.015 376.655 4377.295 ;
        RECT 377.085 4377.015 377.365 4377.295 ;
        RECT 377.795 4377.015 378.075 4377.295 ;
        RECT 378.505 4377.015 378.785 4377.295 ;
        RECT 369.275 4376.305 369.555 4376.585 ;
        RECT 369.985 4376.305 370.265 4376.585 ;
        RECT 370.695 4376.305 370.975 4376.585 ;
        RECT 371.405 4376.305 371.685 4376.585 ;
        RECT 372.115 4376.305 372.395 4376.585 ;
        RECT 372.825 4376.305 373.105 4376.585 ;
        RECT 373.535 4376.305 373.815 4376.585 ;
        RECT 374.245 4376.305 374.525 4376.585 ;
        RECT 374.955 4376.305 375.235 4376.585 ;
        RECT 375.665 4376.305 375.945 4376.585 ;
        RECT 376.375 4376.305 376.655 4376.585 ;
        RECT 377.085 4376.305 377.365 4376.585 ;
        RECT 377.795 4376.305 378.075 4376.585 ;
        RECT 378.505 4376.305 378.785 4376.585 ;
        RECT 369.275 4375.595 369.555 4375.875 ;
        RECT 369.985 4375.595 370.265 4375.875 ;
        RECT 370.695 4375.595 370.975 4375.875 ;
        RECT 371.405 4375.595 371.685 4375.875 ;
        RECT 372.115 4375.595 372.395 4375.875 ;
        RECT 372.825 4375.595 373.105 4375.875 ;
        RECT 373.535 4375.595 373.815 4375.875 ;
        RECT 374.245 4375.595 374.525 4375.875 ;
        RECT 374.955 4375.595 375.235 4375.875 ;
        RECT 375.665 4375.595 375.945 4375.875 ;
        RECT 376.375 4375.595 376.655 4375.875 ;
        RECT 377.085 4375.595 377.365 4375.875 ;
        RECT 377.795 4375.595 378.075 4375.875 ;
        RECT 378.505 4375.595 378.785 4375.875 ;
        RECT 369.275 4374.885 369.555 4375.165 ;
        RECT 369.985 4374.885 370.265 4375.165 ;
        RECT 370.695 4374.885 370.975 4375.165 ;
        RECT 371.405 4374.885 371.685 4375.165 ;
        RECT 372.115 4374.885 372.395 4375.165 ;
        RECT 372.825 4374.885 373.105 4375.165 ;
        RECT 373.535 4374.885 373.815 4375.165 ;
        RECT 374.245 4374.885 374.525 4375.165 ;
        RECT 374.955 4374.885 375.235 4375.165 ;
        RECT 375.665 4374.885 375.945 4375.165 ;
        RECT 376.375 4374.885 376.655 4375.165 ;
        RECT 377.085 4374.885 377.365 4375.165 ;
        RECT 377.795 4374.885 378.075 4375.165 ;
        RECT 378.505 4374.885 378.785 4375.165 ;
        RECT 369.275 4374.175 369.555 4374.455 ;
        RECT 369.985 4374.175 370.265 4374.455 ;
        RECT 370.695 4374.175 370.975 4374.455 ;
        RECT 371.405 4374.175 371.685 4374.455 ;
        RECT 372.115 4374.175 372.395 4374.455 ;
        RECT 372.825 4374.175 373.105 4374.455 ;
        RECT 373.535 4374.175 373.815 4374.455 ;
        RECT 374.245 4374.175 374.525 4374.455 ;
        RECT 374.955 4374.175 375.235 4374.455 ;
        RECT 375.665 4374.175 375.945 4374.455 ;
        RECT 376.375 4374.175 376.655 4374.455 ;
        RECT 377.085 4374.175 377.365 4374.455 ;
        RECT 377.795 4374.175 378.075 4374.455 ;
        RECT 378.505 4374.175 378.785 4374.455 ;
        RECT 369.275 4373.465 369.555 4373.745 ;
        RECT 369.985 4373.465 370.265 4373.745 ;
        RECT 370.695 4373.465 370.975 4373.745 ;
        RECT 371.405 4373.465 371.685 4373.745 ;
        RECT 372.115 4373.465 372.395 4373.745 ;
        RECT 372.825 4373.465 373.105 4373.745 ;
        RECT 373.535 4373.465 373.815 4373.745 ;
        RECT 374.245 4373.465 374.525 4373.745 ;
        RECT 374.955 4373.465 375.235 4373.745 ;
        RECT 375.665 4373.465 375.945 4373.745 ;
        RECT 376.375 4373.465 376.655 4373.745 ;
        RECT 377.085 4373.465 377.365 4373.745 ;
        RECT 377.795 4373.465 378.075 4373.745 ;
        RECT 378.505 4373.465 378.785 4373.745 ;
        RECT 369.275 4372.755 369.555 4373.035 ;
        RECT 369.985 4372.755 370.265 4373.035 ;
        RECT 370.695 4372.755 370.975 4373.035 ;
        RECT 371.405 4372.755 371.685 4373.035 ;
        RECT 372.115 4372.755 372.395 4373.035 ;
        RECT 372.825 4372.755 373.105 4373.035 ;
        RECT 373.535 4372.755 373.815 4373.035 ;
        RECT 374.245 4372.755 374.525 4373.035 ;
        RECT 374.955 4372.755 375.235 4373.035 ;
        RECT 375.665 4372.755 375.945 4373.035 ;
        RECT 376.375 4372.755 376.655 4373.035 ;
        RECT 377.085 4372.755 377.365 4373.035 ;
        RECT 377.795 4372.755 378.075 4373.035 ;
        RECT 378.505 4372.755 378.785 4373.035 ;
        RECT 369.275 4372.045 369.555 4372.325 ;
        RECT 369.985 4372.045 370.265 4372.325 ;
        RECT 370.695 4372.045 370.975 4372.325 ;
        RECT 371.405 4372.045 371.685 4372.325 ;
        RECT 372.115 4372.045 372.395 4372.325 ;
        RECT 372.825 4372.045 373.105 4372.325 ;
        RECT 373.535 4372.045 373.815 4372.325 ;
        RECT 374.245 4372.045 374.525 4372.325 ;
        RECT 374.955 4372.045 375.235 4372.325 ;
        RECT 375.665 4372.045 375.945 4372.325 ;
        RECT 376.375 4372.045 376.655 4372.325 ;
        RECT 377.085 4372.045 377.365 4372.325 ;
        RECT 377.795 4372.045 378.075 4372.325 ;
        RECT 378.505 4372.045 378.785 4372.325 ;
        RECT 369.275 4371.335 369.555 4371.615 ;
        RECT 369.985 4371.335 370.265 4371.615 ;
        RECT 370.695 4371.335 370.975 4371.615 ;
        RECT 371.405 4371.335 371.685 4371.615 ;
        RECT 372.115 4371.335 372.395 4371.615 ;
        RECT 372.825 4371.335 373.105 4371.615 ;
        RECT 373.535 4371.335 373.815 4371.615 ;
        RECT 374.245 4371.335 374.525 4371.615 ;
        RECT 374.955 4371.335 375.235 4371.615 ;
        RECT 375.665 4371.335 375.945 4371.615 ;
        RECT 376.375 4371.335 376.655 4371.615 ;
        RECT 377.085 4371.335 377.365 4371.615 ;
        RECT 377.795 4371.335 378.075 4371.615 ;
        RECT 378.505 4371.335 378.785 4371.615 ;
        RECT 3500.255 4375.615 3500.535 4375.895 ;
        RECT 3500.965 4375.615 3501.245 4375.895 ;
        RECT 3501.675 4375.615 3501.955 4375.895 ;
        RECT 3502.385 4375.615 3502.665 4375.895 ;
        RECT 3503.095 4375.615 3503.375 4375.895 ;
        RECT 3503.805 4375.615 3504.085 4375.895 ;
        RECT 3504.515 4375.615 3504.795 4375.895 ;
        RECT 3505.225 4375.615 3505.505 4375.895 ;
        RECT 3505.935 4375.615 3506.215 4375.895 ;
        RECT 3506.645 4375.615 3506.925 4375.895 ;
        RECT 3507.355 4375.615 3507.635 4375.895 ;
        RECT 3508.065 4375.615 3508.345 4375.895 ;
        RECT 3508.775 4375.615 3509.055 4375.895 ;
        RECT 3509.485 4375.615 3509.765 4375.895 ;
        RECT 3500.255 4374.905 3500.535 4375.185 ;
        RECT 3500.965 4374.905 3501.245 4375.185 ;
        RECT 3501.675 4374.905 3501.955 4375.185 ;
        RECT 3502.385 4374.905 3502.665 4375.185 ;
        RECT 3503.095 4374.905 3503.375 4375.185 ;
        RECT 3503.805 4374.905 3504.085 4375.185 ;
        RECT 3504.515 4374.905 3504.795 4375.185 ;
        RECT 3505.225 4374.905 3505.505 4375.185 ;
        RECT 3505.935 4374.905 3506.215 4375.185 ;
        RECT 3506.645 4374.905 3506.925 4375.185 ;
        RECT 3507.355 4374.905 3507.635 4375.185 ;
        RECT 3508.065 4374.905 3508.345 4375.185 ;
        RECT 3508.775 4374.905 3509.055 4375.185 ;
        RECT 3509.485 4374.905 3509.765 4375.185 ;
        RECT 3500.255 4374.195 3500.535 4374.475 ;
        RECT 3500.965 4374.195 3501.245 4374.475 ;
        RECT 3501.675 4374.195 3501.955 4374.475 ;
        RECT 3502.385 4374.195 3502.665 4374.475 ;
        RECT 3503.095 4374.195 3503.375 4374.475 ;
        RECT 3503.805 4374.195 3504.085 4374.475 ;
        RECT 3504.515 4374.195 3504.795 4374.475 ;
        RECT 3505.225 4374.195 3505.505 4374.475 ;
        RECT 3505.935 4374.195 3506.215 4374.475 ;
        RECT 3506.645 4374.195 3506.925 4374.475 ;
        RECT 3507.355 4374.195 3507.635 4374.475 ;
        RECT 3508.065 4374.195 3508.345 4374.475 ;
        RECT 3508.775 4374.195 3509.055 4374.475 ;
        RECT 3509.485 4374.195 3509.765 4374.475 ;
        RECT 3500.255 4373.485 3500.535 4373.765 ;
        RECT 3500.965 4373.485 3501.245 4373.765 ;
        RECT 3501.675 4373.485 3501.955 4373.765 ;
        RECT 3502.385 4373.485 3502.665 4373.765 ;
        RECT 3503.095 4373.485 3503.375 4373.765 ;
        RECT 3503.805 4373.485 3504.085 4373.765 ;
        RECT 3504.515 4373.485 3504.795 4373.765 ;
        RECT 3505.225 4373.485 3505.505 4373.765 ;
        RECT 3505.935 4373.485 3506.215 4373.765 ;
        RECT 3506.645 4373.485 3506.925 4373.765 ;
        RECT 3507.355 4373.485 3507.635 4373.765 ;
        RECT 3508.065 4373.485 3508.345 4373.765 ;
        RECT 3508.775 4373.485 3509.055 4373.765 ;
        RECT 3509.485 4373.485 3509.765 4373.765 ;
        RECT 3500.255 4372.775 3500.535 4373.055 ;
        RECT 3500.965 4372.775 3501.245 4373.055 ;
        RECT 3501.675 4372.775 3501.955 4373.055 ;
        RECT 3502.385 4372.775 3502.665 4373.055 ;
        RECT 3503.095 4372.775 3503.375 4373.055 ;
        RECT 3503.805 4372.775 3504.085 4373.055 ;
        RECT 3504.515 4372.775 3504.795 4373.055 ;
        RECT 3505.225 4372.775 3505.505 4373.055 ;
        RECT 3505.935 4372.775 3506.215 4373.055 ;
        RECT 3506.645 4372.775 3506.925 4373.055 ;
        RECT 3507.355 4372.775 3507.635 4373.055 ;
        RECT 3508.065 4372.775 3508.345 4373.055 ;
        RECT 3508.775 4372.775 3509.055 4373.055 ;
        RECT 3509.485 4372.775 3509.765 4373.055 ;
        RECT 3500.255 4372.065 3500.535 4372.345 ;
        RECT 3500.965 4372.065 3501.245 4372.345 ;
        RECT 3501.675 4372.065 3501.955 4372.345 ;
        RECT 3502.385 4372.065 3502.665 4372.345 ;
        RECT 3503.095 4372.065 3503.375 4372.345 ;
        RECT 3503.805 4372.065 3504.085 4372.345 ;
        RECT 3504.515 4372.065 3504.795 4372.345 ;
        RECT 3505.225 4372.065 3505.505 4372.345 ;
        RECT 3505.935 4372.065 3506.215 4372.345 ;
        RECT 3506.645 4372.065 3506.925 4372.345 ;
        RECT 3507.355 4372.065 3507.635 4372.345 ;
        RECT 3508.065 4372.065 3508.345 4372.345 ;
        RECT 3508.775 4372.065 3509.055 4372.345 ;
        RECT 3509.485 4372.065 3509.765 4372.345 ;
        RECT 3500.255 4371.355 3500.535 4371.635 ;
        RECT 3500.965 4371.355 3501.245 4371.635 ;
        RECT 3501.675 4371.355 3501.955 4371.635 ;
        RECT 3502.385 4371.355 3502.665 4371.635 ;
        RECT 3503.095 4371.355 3503.375 4371.635 ;
        RECT 3503.805 4371.355 3504.085 4371.635 ;
        RECT 3504.515 4371.355 3504.795 4371.635 ;
        RECT 3505.225 4371.355 3505.505 4371.635 ;
        RECT 3505.935 4371.355 3506.215 4371.635 ;
        RECT 3506.645 4371.355 3506.925 4371.635 ;
        RECT 3507.355 4371.355 3507.635 4371.635 ;
        RECT 3508.065 4371.355 3508.345 4371.635 ;
        RECT 3508.775 4371.355 3509.055 4371.635 ;
        RECT 3509.485 4371.355 3509.765 4371.635 ;
        RECT 3500.255 4370.645 3500.535 4370.925 ;
        RECT 3500.965 4370.645 3501.245 4370.925 ;
        RECT 3501.675 4370.645 3501.955 4370.925 ;
        RECT 3502.385 4370.645 3502.665 4370.925 ;
        RECT 3503.095 4370.645 3503.375 4370.925 ;
        RECT 3503.805 4370.645 3504.085 4370.925 ;
        RECT 3504.515 4370.645 3504.795 4370.925 ;
        RECT 3505.225 4370.645 3505.505 4370.925 ;
        RECT 3505.935 4370.645 3506.215 4370.925 ;
        RECT 3506.645 4370.645 3506.925 4370.925 ;
        RECT 3507.355 4370.645 3507.635 4370.925 ;
        RECT 3508.065 4370.645 3508.345 4370.925 ;
        RECT 3508.775 4370.645 3509.055 4370.925 ;
        RECT 3509.485 4370.645 3509.765 4370.925 ;
        RECT 3500.255 4369.935 3500.535 4370.215 ;
        RECT 3500.965 4369.935 3501.245 4370.215 ;
        RECT 3501.675 4369.935 3501.955 4370.215 ;
        RECT 3502.385 4369.935 3502.665 4370.215 ;
        RECT 3503.095 4369.935 3503.375 4370.215 ;
        RECT 3503.805 4369.935 3504.085 4370.215 ;
        RECT 3504.515 4369.935 3504.795 4370.215 ;
        RECT 3505.225 4369.935 3505.505 4370.215 ;
        RECT 3505.935 4369.935 3506.215 4370.215 ;
        RECT 3506.645 4369.935 3506.925 4370.215 ;
        RECT 3507.355 4369.935 3507.635 4370.215 ;
        RECT 3508.065 4369.935 3508.345 4370.215 ;
        RECT 3508.775 4369.935 3509.055 4370.215 ;
        RECT 3509.485 4369.935 3509.765 4370.215 ;
        RECT 369.275 4368.715 369.555 4368.995 ;
        RECT 369.985 4368.715 370.265 4368.995 ;
        RECT 370.695 4368.715 370.975 4368.995 ;
        RECT 371.405 4368.715 371.685 4368.995 ;
        RECT 372.115 4368.715 372.395 4368.995 ;
        RECT 372.825 4368.715 373.105 4368.995 ;
        RECT 373.535 4368.715 373.815 4368.995 ;
        RECT 374.245 4368.715 374.525 4368.995 ;
        RECT 374.955 4368.715 375.235 4368.995 ;
        RECT 375.665 4368.715 375.945 4368.995 ;
        RECT 376.375 4368.715 376.655 4368.995 ;
        RECT 377.085 4368.715 377.365 4368.995 ;
        RECT 377.795 4368.715 378.075 4368.995 ;
        RECT 378.505 4368.715 378.785 4368.995 ;
        RECT 369.275 4368.005 369.555 4368.285 ;
        RECT 369.985 4368.005 370.265 4368.285 ;
        RECT 370.695 4368.005 370.975 4368.285 ;
        RECT 371.405 4368.005 371.685 4368.285 ;
        RECT 372.115 4368.005 372.395 4368.285 ;
        RECT 372.825 4368.005 373.105 4368.285 ;
        RECT 373.535 4368.005 373.815 4368.285 ;
        RECT 374.245 4368.005 374.525 4368.285 ;
        RECT 374.955 4368.005 375.235 4368.285 ;
        RECT 375.665 4368.005 375.945 4368.285 ;
        RECT 376.375 4368.005 376.655 4368.285 ;
        RECT 377.085 4368.005 377.365 4368.285 ;
        RECT 377.795 4368.005 378.075 4368.285 ;
        RECT 378.505 4368.005 378.785 4368.285 ;
        RECT 369.275 4367.295 369.555 4367.575 ;
        RECT 369.985 4367.295 370.265 4367.575 ;
        RECT 370.695 4367.295 370.975 4367.575 ;
        RECT 371.405 4367.295 371.685 4367.575 ;
        RECT 372.115 4367.295 372.395 4367.575 ;
        RECT 372.825 4367.295 373.105 4367.575 ;
        RECT 373.535 4367.295 373.815 4367.575 ;
        RECT 374.245 4367.295 374.525 4367.575 ;
        RECT 374.955 4367.295 375.235 4367.575 ;
        RECT 375.665 4367.295 375.945 4367.575 ;
        RECT 376.375 4367.295 376.655 4367.575 ;
        RECT 377.085 4367.295 377.365 4367.575 ;
        RECT 377.795 4367.295 378.075 4367.575 ;
        RECT 378.505 4367.295 378.785 4367.575 ;
        RECT 369.275 4366.585 369.555 4366.865 ;
        RECT 369.985 4366.585 370.265 4366.865 ;
        RECT 370.695 4366.585 370.975 4366.865 ;
        RECT 371.405 4366.585 371.685 4366.865 ;
        RECT 372.115 4366.585 372.395 4366.865 ;
        RECT 372.825 4366.585 373.105 4366.865 ;
        RECT 373.535 4366.585 373.815 4366.865 ;
        RECT 374.245 4366.585 374.525 4366.865 ;
        RECT 374.955 4366.585 375.235 4366.865 ;
        RECT 375.665 4366.585 375.945 4366.865 ;
        RECT 376.375 4366.585 376.655 4366.865 ;
        RECT 377.085 4366.585 377.365 4366.865 ;
        RECT 377.795 4366.585 378.075 4366.865 ;
        RECT 378.505 4366.585 378.785 4366.865 ;
        RECT 369.275 4365.875 369.555 4366.155 ;
        RECT 369.985 4365.875 370.265 4366.155 ;
        RECT 370.695 4365.875 370.975 4366.155 ;
        RECT 371.405 4365.875 371.685 4366.155 ;
        RECT 372.115 4365.875 372.395 4366.155 ;
        RECT 372.825 4365.875 373.105 4366.155 ;
        RECT 373.535 4365.875 373.815 4366.155 ;
        RECT 374.245 4365.875 374.525 4366.155 ;
        RECT 374.955 4365.875 375.235 4366.155 ;
        RECT 375.665 4365.875 375.945 4366.155 ;
        RECT 376.375 4365.875 376.655 4366.155 ;
        RECT 377.085 4365.875 377.365 4366.155 ;
        RECT 377.795 4365.875 378.075 4366.155 ;
        RECT 378.505 4365.875 378.785 4366.155 ;
        RECT 3500.255 4369.225 3500.535 4369.505 ;
        RECT 3500.965 4369.225 3501.245 4369.505 ;
        RECT 3501.675 4369.225 3501.955 4369.505 ;
        RECT 3502.385 4369.225 3502.665 4369.505 ;
        RECT 3503.095 4369.225 3503.375 4369.505 ;
        RECT 3503.805 4369.225 3504.085 4369.505 ;
        RECT 3504.515 4369.225 3504.795 4369.505 ;
        RECT 3505.225 4369.225 3505.505 4369.505 ;
        RECT 3505.935 4369.225 3506.215 4369.505 ;
        RECT 3506.645 4369.225 3506.925 4369.505 ;
        RECT 3507.355 4369.225 3507.635 4369.505 ;
        RECT 3508.065 4369.225 3508.345 4369.505 ;
        RECT 3508.775 4369.225 3509.055 4369.505 ;
        RECT 3509.485 4369.225 3509.765 4369.505 ;
        RECT 3500.255 4368.515 3500.535 4368.795 ;
        RECT 3500.965 4368.515 3501.245 4368.795 ;
        RECT 3501.675 4368.515 3501.955 4368.795 ;
        RECT 3502.385 4368.515 3502.665 4368.795 ;
        RECT 3503.095 4368.515 3503.375 4368.795 ;
        RECT 3503.805 4368.515 3504.085 4368.795 ;
        RECT 3504.515 4368.515 3504.795 4368.795 ;
        RECT 3505.225 4368.515 3505.505 4368.795 ;
        RECT 3505.935 4368.515 3506.215 4368.795 ;
        RECT 3506.645 4368.515 3506.925 4368.795 ;
        RECT 3507.355 4368.515 3507.635 4368.795 ;
        RECT 3508.065 4368.515 3508.345 4368.795 ;
        RECT 3508.775 4368.515 3509.055 4368.795 ;
        RECT 3509.485 4368.515 3509.765 4368.795 ;
        RECT 3500.255 4367.805 3500.535 4368.085 ;
        RECT 3500.965 4367.805 3501.245 4368.085 ;
        RECT 3501.675 4367.805 3501.955 4368.085 ;
        RECT 3502.385 4367.805 3502.665 4368.085 ;
        RECT 3503.095 4367.805 3503.375 4368.085 ;
        RECT 3503.805 4367.805 3504.085 4368.085 ;
        RECT 3504.515 4367.805 3504.795 4368.085 ;
        RECT 3505.225 4367.805 3505.505 4368.085 ;
        RECT 3505.935 4367.805 3506.215 4368.085 ;
        RECT 3506.645 4367.805 3506.925 4368.085 ;
        RECT 3507.355 4367.805 3507.635 4368.085 ;
        RECT 3508.065 4367.805 3508.345 4368.085 ;
        RECT 3508.775 4367.805 3509.055 4368.085 ;
        RECT 3509.485 4367.805 3509.765 4368.085 ;
        RECT 3500.255 4367.095 3500.535 4367.375 ;
        RECT 3500.965 4367.095 3501.245 4367.375 ;
        RECT 3501.675 4367.095 3501.955 4367.375 ;
        RECT 3502.385 4367.095 3502.665 4367.375 ;
        RECT 3503.095 4367.095 3503.375 4367.375 ;
        RECT 3503.805 4367.095 3504.085 4367.375 ;
        RECT 3504.515 4367.095 3504.795 4367.375 ;
        RECT 3505.225 4367.095 3505.505 4367.375 ;
        RECT 3505.935 4367.095 3506.215 4367.375 ;
        RECT 3506.645 4367.095 3506.925 4367.375 ;
        RECT 3507.355 4367.095 3507.635 4367.375 ;
        RECT 3508.065 4367.095 3508.345 4367.375 ;
        RECT 3508.775 4367.095 3509.055 4367.375 ;
        RECT 3509.485 4367.095 3509.765 4367.375 ;
        RECT 3500.255 4366.385 3500.535 4366.665 ;
        RECT 3500.965 4366.385 3501.245 4366.665 ;
        RECT 3501.675 4366.385 3501.955 4366.665 ;
        RECT 3502.385 4366.385 3502.665 4366.665 ;
        RECT 3503.095 4366.385 3503.375 4366.665 ;
        RECT 3503.805 4366.385 3504.085 4366.665 ;
        RECT 3504.515 4366.385 3504.795 4366.665 ;
        RECT 3505.225 4366.385 3505.505 4366.665 ;
        RECT 3505.935 4366.385 3506.215 4366.665 ;
        RECT 3506.645 4366.385 3506.925 4366.665 ;
        RECT 3507.355 4366.385 3507.635 4366.665 ;
        RECT 3508.065 4366.385 3508.345 4366.665 ;
        RECT 3508.775 4366.385 3509.055 4366.665 ;
        RECT 3509.485 4366.385 3509.765 4366.665 ;
        RECT 369.275 4365.165 369.555 4365.445 ;
        RECT 369.985 4365.165 370.265 4365.445 ;
        RECT 370.695 4365.165 370.975 4365.445 ;
        RECT 371.405 4365.165 371.685 4365.445 ;
        RECT 372.115 4365.165 372.395 4365.445 ;
        RECT 372.825 4365.165 373.105 4365.445 ;
        RECT 373.535 4365.165 373.815 4365.445 ;
        RECT 374.245 4365.165 374.525 4365.445 ;
        RECT 374.955 4365.165 375.235 4365.445 ;
        RECT 375.665 4365.165 375.945 4365.445 ;
        RECT 376.375 4365.165 376.655 4365.445 ;
        RECT 377.085 4365.165 377.365 4365.445 ;
        RECT 377.795 4365.165 378.075 4365.445 ;
        RECT 378.505 4365.165 378.785 4365.445 ;
        RECT 369.275 4364.455 369.555 4364.735 ;
        RECT 369.985 4364.455 370.265 4364.735 ;
        RECT 370.695 4364.455 370.975 4364.735 ;
        RECT 371.405 4364.455 371.685 4364.735 ;
        RECT 372.115 4364.455 372.395 4364.735 ;
        RECT 372.825 4364.455 373.105 4364.735 ;
        RECT 373.535 4364.455 373.815 4364.735 ;
        RECT 374.245 4364.455 374.525 4364.735 ;
        RECT 374.955 4364.455 375.235 4364.735 ;
        RECT 375.665 4364.455 375.945 4364.735 ;
        RECT 376.375 4364.455 376.655 4364.735 ;
        RECT 377.085 4364.455 377.365 4364.735 ;
        RECT 377.795 4364.455 378.075 4364.735 ;
        RECT 378.505 4364.455 378.785 4364.735 ;
        RECT 369.275 4363.745 369.555 4364.025 ;
        RECT 369.985 4363.745 370.265 4364.025 ;
        RECT 370.695 4363.745 370.975 4364.025 ;
        RECT 371.405 4363.745 371.685 4364.025 ;
        RECT 372.115 4363.745 372.395 4364.025 ;
        RECT 372.825 4363.745 373.105 4364.025 ;
        RECT 373.535 4363.745 373.815 4364.025 ;
        RECT 374.245 4363.745 374.525 4364.025 ;
        RECT 374.955 4363.745 375.235 4364.025 ;
        RECT 375.665 4363.745 375.945 4364.025 ;
        RECT 376.375 4363.745 376.655 4364.025 ;
        RECT 377.085 4363.745 377.365 4364.025 ;
        RECT 377.795 4363.745 378.075 4364.025 ;
        RECT 378.505 4363.745 378.785 4364.025 ;
        RECT 369.275 4363.035 369.555 4363.315 ;
        RECT 369.985 4363.035 370.265 4363.315 ;
        RECT 370.695 4363.035 370.975 4363.315 ;
        RECT 371.405 4363.035 371.685 4363.315 ;
        RECT 372.115 4363.035 372.395 4363.315 ;
        RECT 372.825 4363.035 373.105 4363.315 ;
        RECT 373.535 4363.035 373.815 4363.315 ;
        RECT 374.245 4363.035 374.525 4363.315 ;
        RECT 374.955 4363.035 375.235 4363.315 ;
        RECT 375.665 4363.035 375.945 4363.315 ;
        RECT 376.375 4363.035 376.655 4363.315 ;
        RECT 377.085 4363.035 377.365 4363.315 ;
        RECT 377.795 4363.035 378.075 4363.315 ;
        RECT 378.505 4363.035 378.785 4363.315 ;
        RECT 369.275 4362.325 369.555 4362.605 ;
        RECT 369.985 4362.325 370.265 4362.605 ;
        RECT 370.695 4362.325 370.975 4362.605 ;
        RECT 371.405 4362.325 371.685 4362.605 ;
        RECT 372.115 4362.325 372.395 4362.605 ;
        RECT 372.825 4362.325 373.105 4362.605 ;
        RECT 373.535 4362.325 373.815 4362.605 ;
        RECT 374.245 4362.325 374.525 4362.605 ;
        RECT 374.955 4362.325 375.235 4362.605 ;
        RECT 375.665 4362.325 375.945 4362.605 ;
        RECT 376.375 4362.325 376.655 4362.605 ;
        RECT 377.085 4362.325 377.365 4362.605 ;
        RECT 377.795 4362.325 378.075 4362.605 ;
        RECT 378.505 4362.325 378.785 4362.605 ;
        RECT 369.275 4361.615 369.555 4361.895 ;
        RECT 369.985 4361.615 370.265 4361.895 ;
        RECT 370.695 4361.615 370.975 4361.895 ;
        RECT 371.405 4361.615 371.685 4361.895 ;
        RECT 372.115 4361.615 372.395 4361.895 ;
        RECT 372.825 4361.615 373.105 4361.895 ;
        RECT 373.535 4361.615 373.815 4361.895 ;
        RECT 374.245 4361.615 374.525 4361.895 ;
        RECT 374.955 4361.615 375.235 4361.895 ;
        RECT 375.665 4361.615 375.945 4361.895 ;
        RECT 376.375 4361.615 376.655 4361.895 ;
        RECT 377.085 4361.615 377.365 4361.895 ;
        RECT 377.795 4361.615 378.075 4361.895 ;
        RECT 378.505 4361.615 378.785 4361.895 ;
        RECT 369.275 4360.905 369.555 4361.185 ;
        RECT 369.985 4360.905 370.265 4361.185 ;
        RECT 370.695 4360.905 370.975 4361.185 ;
        RECT 371.405 4360.905 371.685 4361.185 ;
        RECT 372.115 4360.905 372.395 4361.185 ;
        RECT 372.825 4360.905 373.105 4361.185 ;
        RECT 373.535 4360.905 373.815 4361.185 ;
        RECT 374.245 4360.905 374.525 4361.185 ;
        RECT 374.955 4360.905 375.235 4361.185 ;
        RECT 375.665 4360.905 375.945 4361.185 ;
        RECT 376.375 4360.905 376.655 4361.185 ;
        RECT 377.085 4360.905 377.365 4361.185 ;
        RECT 377.795 4360.905 378.075 4361.185 ;
        RECT 378.505 4360.905 378.785 4361.185 ;
        RECT 369.275 4360.195 369.555 4360.475 ;
        RECT 369.985 4360.195 370.265 4360.475 ;
        RECT 370.695 4360.195 370.975 4360.475 ;
        RECT 371.405 4360.195 371.685 4360.475 ;
        RECT 372.115 4360.195 372.395 4360.475 ;
        RECT 372.825 4360.195 373.105 4360.475 ;
        RECT 373.535 4360.195 373.815 4360.475 ;
        RECT 374.245 4360.195 374.525 4360.475 ;
        RECT 374.955 4360.195 375.235 4360.475 ;
        RECT 375.665 4360.195 375.945 4360.475 ;
        RECT 376.375 4360.195 376.655 4360.475 ;
        RECT 377.085 4360.195 377.365 4360.475 ;
        RECT 377.795 4360.195 378.075 4360.475 ;
        RECT 378.505 4360.195 378.785 4360.475 ;
        RECT 369.275 4359.485 369.555 4359.765 ;
        RECT 369.985 4359.485 370.265 4359.765 ;
        RECT 370.695 4359.485 370.975 4359.765 ;
        RECT 371.405 4359.485 371.685 4359.765 ;
        RECT 372.115 4359.485 372.395 4359.765 ;
        RECT 372.825 4359.485 373.105 4359.765 ;
        RECT 373.535 4359.485 373.815 4359.765 ;
        RECT 374.245 4359.485 374.525 4359.765 ;
        RECT 374.955 4359.485 375.235 4359.765 ;
        RECT 375.665 4359.485 375.945 4359.765 ;
        RECT 376.375 4359.485 376.655 4359.765 ;
        RECT 377.085 4359.485 377.365 4359.765 ;
        RECT 377.795 4359.485 378.075 4359.765 ;
        RECT 378.505 4359.485 378.785 4359.765 ;
        RECT 3500.255 4363.765 3500.535 4364.045 ;
        RECT 3500.965 4363.765 3501.245 4364.045 ;
        RECT 3501.675 4363.765 3501.955 4364.045 ;
        RECT 3502.385 4363.765 3502.665 4364.045 ;
        RECT 3503.095 4363.765 3503.375 4364.045 ;
        RECT 3503.805 4363.765 3504.085 4364.045 ;
        RECT 3504.515 4363.765 3504.795 4364.045 ;
        RECT 3505.225 4363.765 3505.505 4364.045 ;
        RECT 3505.935 4363.765 3506.215 4364.045 ;
        RECT 3506.645 4363.765 3506.925 4364.045 ;
        RECT 3507.355 4363.765 3507.635 4364.045 ;
        RECT 3508.065 4363.765 3508.345 4364.045 ;
        RECT 3508.775 4363.765 3509.055 4364.045 ;
        RECT 3509.485 4363.765 3509.765 4364.045 ;
        RECT 3500.255 4363.055 3500.535 4363.335 ;
        RECT 3500.965 4363.055 3501.245 4363.335 ;
        RECT 3501.675 4363.055 3501.955 4363.335 ;
        RECT 3502.385 4363.055 3502.665 4363.335 ;
        RECT 3503.095 4363.055 3503.375 4363.335 ;
        RECT 3503.805 4363.055 3504.085 4363.335 ;
        RECT 3504.515 4363.055 3504.795 4363.335 ;
        RECT 3505.225 4363.055 3505.505 4363.335 ;
        RECT 3505.935 4363.055 3506.215 4363.335 ;
        RECT 3506.645 4363.055 3506.925 4363.335 ;
        RECT 3507.355 4363.055 3507.635 4363.335 ;
        RECT 3508.065 4363.055 3508.345 4363.335 ;
        RECT 3508.775 4363.055 3509.055 4363.335 ;
        RECT 3509.485 4363.055 3509.765 4363.335 ;
        RECT 3500.255 4362.345 3500.535 4362.625 ;
        RECT 3500.965 4362.345 3501.245 4362.625 ;
        RECT 3501.675 4362.345 3501.955 4362.625 ;
        RECT 3502.385 4362.345 3502.665 4362.625 ;
        RECT 3503.095 4362.345 3503.375 4362.625 ;
        RECT 3503.805 4362.345 3504.085 4362.625 ;
        RECT 3504.515 4362.345 3504.795 4362.625 ;
        RECT 3505.225 4362.345 3505.505 4362.625 ;
        RECT 3505.935 4362.345 3506.215 4362.625 ;
        RECT 3506.645 4362.345 3506.925 4362.625 ;
        RECT 3507.355 4362.345 3507.635 4362.625 ;
        RECT 3508.065 4362.345 3508.345 4362.625 ;
        RECT 3508.775 4362.345 3509.055 4362.625 ;
        RECT 3509.485 4362.345 3509.765 4362.625 ;
        RECT 3500.255 4361.635 3500.535 4361.915 ;
        RECT 3500.965 4361.635 3501.245 4361.915 ;
        RECT 3501.675 4361.635 3501.955 4361.915 ;
        RECT 3502.385 4361.635 3502.665 4361.915 ;
        RECT 3503.095 4361.635 3503.375 4361.915 ;
        RECT 3503.805 4361.635 3504.085 4361.915 ;
        RECT 3504.515 4361.635 3504.795 4361.915 ;
        RECT 3505.225 4361.635 3505.505 4361.915 ;
        RECT 3505.935 4361.635 3506.215 4361.915 ;
        RECT 3506.645 4361.635 3506.925 4361.915 ;
        RECT 3507.355 4361.635 3507.635 4361.915 ;
        RECT 3508.065 4361.635 3508.345 4361.915 ;
        RECT 3508.775 4361.635 3509.055 4361.915 ;
        RECT 3509.485 4361.635 3509.765 4361.915 ;
        RECT 3500.255 4360.925 3500.535 4361.205 ;
        RECT 3500.965 4360.925 3501.245 4361.205 ;
        RECT 3501.675 4360.925 3501.955 4361.205 ;
        RECT 3502.385 4360.925 3502.665 4361.205 ;
        RECT 3503.095 4360.925 3503.375 4361.205 ;
        RECT 3503.805 4360.925 3504.085 4361.205 ;
        RECT 3504.515 4360.925 3504.795 4361.205 ;
        RECT 3505.225 4360.925 3505.505 4361.205 ;
        RECT 3505.935 4360.925 3506.215 4361.205 ;
        RECT 3506.645 4360.925 3506.925 4361.205 ;
        RECT 3507.355 4360.925 3507.635 4361.205 ;
        RECT 3508.065 4360.925 3508.345 4361.205 ;
        RECT 3508.775 4360.925 3509.055 4361.205 ;
        RECT 3509.485 4360.925 3509.765 4361.205 ;
        RECT 3500.255 4360.215 3500.535 4360.495 ;
        RECT 3500.965 4360.215 3501.245 4360.495 ;
        RECT 3501.675 4360.215 3501.955 4360.495 ;
        RECT 3502.385 4360.215 3502.665 4360.495 ;
        RECT 3503.095 4360.215 3503.375 4360.495 ;
        RECT 3503.805 4360.215 3504.085 4360.495 ;
        RECT 3504.515 4360.215 3504.795 4360.495 ;
        RECT 3505.225 4360.215 3505.505 4360.495 ;
        RECT 3505.935 4360.215 3506.215 4360.495 ;
        RECT 3506.645 4360.215 3506.925 4360.495 ;
        RECT 3507.355 4360.215 3507.635 4360.495 ;
        RECT 3508.065 4360.215 3508.345 4360.495 ;
        RECT 3508.775 4360.215 3509.055 4360.495 ;
        RECT 3509.485 4360.215 3509.765 4360.495 ;
        RECT 3500.255 4359.505 3500.535 4359.785 ;
        RECT 3500.965 4359.505 3501.245 4359.785 ;
        RECT 3501.675 4359.505 3501.955 4359.785 ;
        RECT 3502.385 4359.505 3502.665 4359.785 ;
        RECT 3503.095 4359.505 3503.375 4359.785 ;
        RECT 3503.805 4359.505 3504.085 4359.785 ;
        RECT 3504.515 4359.505 3504.795 4359.785 ;
        RECT 3505.225 4359.505 3505.505 4359.785 ;
        RECT 3505.935 4359.505 3506.215 4359.785 ;
        RECT 3506.645 4359.505 3506.925 4359.785 ;
        RECT 3507.355 4359.505 3507.635 4359.785 ;
        RECT 3508.065 4359.505 3508.345 4359.785 ;
        RECT 3508.775 4359.505 3509.055 4359.785 ;
        RECT 3509.485 4359.505 3509.765 4359.785 ;
        RECT 3500.255 4358.795 3500.535 4359.075 ;
        RECT 3500.965 4358.795 3501.245 4359.075 ;
        RECT 3501.675 4358.795 3501.955 4359.075 ;
        RECT 3502.385 4358.795 3502.665 4359.075 ;
        RECT 3503.095 4358.795 3503.375 4359.075 ;
        RECT 3503.805 4358.795 3504.085 4359.075 ;
        RECT 3504.515 4358.795 3504.795 4359.075 ;
        RECT 3505.225 4358.795 3505.505 4359.075 ;
        RECT 3505.935 4358.795 3506.215 4359.075 ;
        RECT 3506.645 4358.795 3506.925 4359.075 ;
        RECT 3507.355 4358.795 3507.635 4359.075 ;
        RECT 3508.065 4358.795 3508.345 4359.075 ;
        RECT 3508.775 4358.795 3509.055 4359.075 ;
        RECT 3509.485 4358.795 3509.765 4359.075 ;
        RECT 3500.255 4358.085 3500.535 4358.365 ;
        RECT 3500.965 4358.085 3501.245 4358.365 ;
        RECT 3501.675 4358.085 3501.955 4358.365 ;
        RECT 3502.385 4358.085 3502.665 4358.365 ;
        RECT 3503.095 4358.085 3503.375 4358.365 ;
        RECT 3503.805 4358.085 3504.085 4358.365 ;
        RECT 3504.515 4358.085 3504.795 4358.365 ;
        RECT 3505.225 4358.085 3505.505 4358.365 ;
        RECT 3505.935 4358.085 3506.215 4358.365 ;
        RECT 3506.645 4358.085 3506.925 4358.365 ;
        RECT 3507.355 4358.085 3507.635 4358.365 ;
        RECT 3508.065 4358.085 3508.345 4358.365 ;
        RECT 3508.775 4358.085 3509.055 4358.365 ;
        RECT 3509.485 4358.085 3509.765 4358.365 ;
        RECT 3500.255 4357.375 3500.535 4357.655 ;
        RECT 3500.965 4357.375 3501.245 4357.655 ;
        RECT 3501.675 4357.375 3501.955 4357.655 ;
        RECT 3502.385 4357.375 3502.665 4357.655 ;
        RECT 3503.095 4357.375 3503.375 4357.655 ;
        RECT 3503.805 4357.375 3504.085 4357.655 ;
        RECT 3504.515 4357.375 3504.795 4357.655 ;
        RECT 3505.225 4357.375 3505.505 4357.655 ;
        RECT 3505.935 4357.375 3506.215 4357.655 ;
        RECT 3506.645 4357.375 3506.925 4357.655 ;
        RECT 3507.355 4357.375 3507.635 4357.655 ;
        RECT 3508.065 4357.375 3508.345 4357.655 ;
        RECT 3508.775 4357.375 3509.055 4357.655 ;
        RECT 3509.485 4357.375 3509.765 4357.655 ;
        RECT 3500.255 4356.665 3500.535 4356.945 ;
        RECT 3500.965 4356.665 3501.245 4356.945 ;
        RECT 3501.675 4356.665 3501.955 4356.945 ;
        RECT 3502.385 4356.665 3502.665 4356.945 ;
        RECT 3503.095 4356.665 3503.375 4356.945 ;
        RECT 3503.805 4356.665 3504.085 4356.945 ;
        RECT 3504.515 4356.665 3504.795 4356.945 ;
        RECT 3505.225 4356.665 3505.505 4356.945 ;
        RECT 3505.935 4356.665 3506.215 4356.945 ;
        RECT 3506.645 4356.665 3506.925 4356.945 ;
        RECT 3507.355 4356.665 3507.635 4356.945 ;
        RECT 3508.065 4356.665 3508.345 4356.945 ;
        RECT 3508.775 4356.665 3509.055 4356.945 ;
        RECT 3509.485 4356.665 3509.765 4356.945 ;
        RECT 3500.255 4355.955 3500.535 4356.235 ;
        RECT 3500.965 4355.955 3501.245 4356.235 ;
        RECT 3501.675 4355.955 3501.955 4356.235 ;
        RECT 3502.385 4355.955 3502.665 4356.235 ;
        RECT 3503.095 4355.955 3503.375 4356.235 ;
        RECT 3503.805 4355.955 3504.085 4356.235 ;
        RECT 3504.515 4355.955 3504.795 4356.235 ;
        RECT 3505.225 4355.955 3505.505 4356.235 ;
        RECT 3505.935 4355.955 3506.215 4356.235 ;
        RECT 3506.645 4355.955 3506.925 4356.235 ;
        RECT 3507.355 4355.955 3507.635 4356.235 ;
        RECT 3508.065 4355.955 3508.345 4356.235 ;
        RECT 3508.775 4355.955 3509.055 4356.235 ;
        RECT 3509.485 4355.955 3509.765 4356.235 ;
        RECT 369.275 4355.185 369.555 4355.465 ;
        RECT 369.985 4355.185 370.265 4355.465 ;
        RECT 370.695 4355.185 370.975 4355.465 ;
        RECT 371.405 4355.185 371.685 4355.465 ;
        RECT 372.115 4355.185 372.395 4355.465 ;
        RECT 372.825 4355.185 373.105 4355.465 ;
        RECT 373.535 4355.185 373.815 4355.465 ;
        RECT 374.245 4355.185 374.525 4355.465 ;
        RECT 374.955 4355.185 375.235 4355.465 ;
        RECT 375.665 4355.185 375.945 4355.465 ;
        RECT 376.375 4355.185 376.655 4355.465 ;
        RECT 377.085 4355.185 377.365 4355.465 ;
        RECT 377.795 4355.185 378.075 4355.465 ;
        RECT 378.505 4355.185 378.785 4355.465 ;
        RECT 369.275 4354.475 369.555 4354.755 ;
        RECT 369.985 4354.475 370.265 4354.755 ;
        RECT 370.695 4354.475 370.975 4354.755 ;
        RECT 371.405 4354.475 371.685 4354.755 ;
        RECT 372.115 4354.475 372.395 4354.755 ;
        RECT 372.825 4354.475 373.105 4354.755 ;
        RECT 373.535 4354.475 373.815 4354.755 ;
        RECT 374.245 4354.475 374.525 4354.755 ;
        RECT 374.955 4354.475 375.235 4354.755 ;
        RECT 375.665 4354.475 375.945 4354.755 ;
        RECT 376.375 4354.475 376.655 4354.755 ;
        RECT 377.085 4354.475 377.365 4354.755 ;
        RECT 377.795 4354.475 378.075 4354.755 ;
        RECT 378.505 4354.475 378.785 4354.755 ;
        RECT 3500.255 4355.245 3500.535 4355.525 ;
        RECT 3500.965 4355.245 3501.245 4355.525 ;
        RECT 3501.675 4355.245 3501.955 4355.525 ;
        RECT 3502.385 4355.245 3502.665 4355.525 ;
        RECT 3503.095 4355.245 3503.375 4355.525 ;
        RECT 3503.805 4355.245 3504.085 4355.525 ;
        RECT 3504.515 4355.245 3504.795 4355.525 ;
        RECT 3505.225 4355.245 3505.505 4355.525 ;
        RECT 3505.935 4355.245 3506.215 4355.525 ;
        RECT 3506.645 4355.245 3506.925 4355.525 ;
        RECT 3507.355 4355.245 3507.635 4355.525 ;
        RECT 3508.065 4355.245 3508.345 4355.525 ;
        RECT 3508.775 4355.245 3509.055 4355.525 ;
        RECT 3509.485 4355.245 3509.765 4355.525 ;
        RECT 3500.255 4354.535 3500.535 4354.815 ;
        RECT 3500.965 4354.535 3501.245 4354.815 ;
        RECT 3501.675 4354.535 3501.955 4354.815 ;
        RECT 3502.385 4354.535 3502.665 4354.815 ;
        RECT 3503.095 4354.535 3503.375 4354.815 ;
        RECT 3503.805 4354.535 3504.085 4354.815 ;
        RECT 3504.515 4354.535 3504.795 4354.815 ;
        RECT 3505.225 4354.535 3505.505 4354.815 ;
        RECT 3505.935 4354.535 3506.215 4354.815 ;
        RECT 3506.645 4354.535 3506.925 4354.815 ;
        RECT 3507.355 4354.535 3507.635 4354.815 ;
        RECT 3508.065 4354.535 3508.345 4354.815 ;
        RECT 3508.775 4354.535 3509.055 4354.815 ;
        RECT 3509.485 4354.535 3509.765 4354.815 ;
        RECT 369.275 4353.765 369.555 4354.045 ;
        RECT 369.985 4353.765 370.265 4354.045 ;
        RECT 370.695 4353.765 370.975 4354.045 ;
        RECT 371.405 4353.765 371.685 4354.045 ;
        RECT 372.115 4353.765 372.395 4354.045 ;
        RECT 372.825 4353.765 373.105 4354.045 ;
        RECT 373.535 4353.765 373.815 4354.045 ;
        RECT 374.245 4353.765 374.525 4354.045 ;
        RECT 374.955 4353.765 375.235 4354.045 ;
        RECT 375.665 4353.765 375.945 4354.045 ;
        RECT 376.375 4353.765 376.655 4354.045 ;
        RECT 377.085 4353.765 377.365 4354.045 ;
        RECT 377.795 4353.765 378.075 4354.045 ;
        RECT 378.505 4353.765 378.785 4354.045 ;
        RECT 369.275 4353.055 369.555 4353.335 ;
        RECT 369.985 4353.055 370.265 4353.335 ;
        RECT 370.695 4353.055 370.975 4353.335 ;
        RECT 371.405 4353.055 371.685 4353.335 ;
        RECT 372.115 4353.055 372.395 4353.335 ;
        RECT 372.825 4353.055 373.105 4353.335 ;
        RECT 373.535 4353.055 373.815 4353.335 ;
        RECT 374.245 4353.055 374.525 4353.335 ;
        RECT 374.955 4353.055 375.235 4353.335 ;
        RECT 375.665 4353.055 375.945 4353.335 ;
        RECT 376.375 4353.055 376.655 4353.335 ;
        RECT 377.085 4353.055 377.365 4353.335 ;
        RECT 377.795 4353.055 378.075 4353.335 ;
        RECT 378.505 4353.055 378.785 4353.335 ;
        RECT 369.275 4352.345 369.555 4352.625 ;
        RECT 369.985 4352.345 370.265 4352.625 ;
        RECT 370.695 4352.345 370.975 4352.625 ;
        RECT 371.405 4352.345 371.685 4352.625 ;
        RECT 372.115 4352.345 372.395 4352.625 ;
        RECT 372.825 4352.345 373.105 4352.625 ;
        RECT 373.535 4352.345 373.815 4352.625 ;
        RECT 374.245 4352.345 374.525 4352.625 ;
        RECT 374.955 4352.345 375.235 4352.625 ;
        RECT 375.665 4352.345 375.945 4352.625 ;
        RECT 376.375 4352.345 376.655 4352.625 ;
        RECT 377.085 4352.345 377.365 4352.625 ;
        RECT 377.795 4352.345 378.075 4352.625 ;
        RECT 378.505 4352.345 378.785 4352.625 ;
        RECT 369.275 4351.635 369.555 4351.915 ;
        RECT 369.985 4351.635 370.265 4351.915 ;
        RECT 370.695 4351.635 370.975 4351.915 ;
        RECT 371.405 4351.635 371.685 4351.915 ;
        RECT 372.115 4351.635 372.395 4351.915 ;
        RECT 372.825 4351.635 373.105 4351.915 ;
        RECT 373.535 4351.635 373.815 4351.915 ;
        RECT 374.245 4351.635 374.525 4351.915 ;
        RECT 374.955 4351.635 375.235 4351.915 ;
        RECT 375.665 4351.635 375.945 4351.915 ;
        RECT 376.375 4351.635 376.655 4351.915 ;
        RECT 377.085 4351.635 377.365 4351.915 ;
        RECT 377.795 4351.635 378.075 4351.915 ;
        RECT 378.505 4351.635 378.785 4351.915 ;
        RECT 369.275 4350.925 369.555 4351.205 ;
        RECT 369.985 4350.925 370.265 4351.205 ;
        RECT 370.695 4350.925 370.975 4351.205 ;
        RECT 371.405 4350.925 371.685 4351.205 ;
        RECT 372.115 4350.925 372.395 4351.205 ;
        RECT 372.825 4350.925 373.105 4351.205 ;
        RECT 373.535 4350.925 373.815 4351.205 ;
        RECT 374.245 4350.925 374.525 4351.205 ;
        RECT 374.955 4350.925 375.235 4351.205 ;
        RECT 375.665 4350.925 375.945 4351.205 ;
        RECT 376.375 4350.925 376.655 4351.205 ;
        RECT 377.085 4350.925 377.365 4351.205 ;
        RECT 377.795 4350.925 378.075 4351.205 ;
        RECT 378.505 4350.925 378.785 4351.205 ;
        RECT 369.275 4350.215 369.555 4350.495 ;
        RECT 369.985 4350.215 370.265 4350.495 ;
        RECT 370.695 4350.215 370.975 4350.495 ;
        RECT 371.405 4350.215 371.685 4350.495 ;
        RECT 372.115 4350.215 372.395 4350.495 ;
        RECT 372.825 4350.215 373.105 4350.495 ;
        RECT 373.535 4350.215 373.815 4350.495 ;
        RECT 374.245 4350.215 374.525 4350.495 ;
        RECT 374.955 4350.215 375.235 4350.495 ;
        RECT 375.665 4350.215 375.945 4350.495 ;
        RECT 376.375 4350.215 376.655 4350.495 ;
        RECT 377.085 4350.215 377.365 4350.495 ;
        RECT 377.795 4350.215 378.075 4350.495 ;
        RECT 378.505 4350.215 378.785 4350.495 ;
        RECT 369.275 4349.505 369.555 4349.785 ;
        RECT 369.985 4349.505 370.265 4349.785 ;
        RECT 370.695 4349.505 370.975 4349.785 ;
        RECT 371.405 4349.505 371.685 4349.785 ;
        RECT 372.115 4349.505 372.395 4349.785 ;
        RECT 372.825 4349.505 373.105 4349.785 ;
        RECT 373.535 4349.505 373.815 4349.785 ;
        RECT 374.245 4349.505 374.525 4349.785 ;
        RECT 374.955 4349.505 375.235 4349.785 ;
        RECT 375.665 4349.505 375.945 4349.785 ;
        RECT 376.375 4349.505 376.655 4349.785 ;
        RECT 377.085 4349.505 377.365 4349.785 ;
        RECT 377.795 4349.505 378.075 4349.785 ;
        RECT 378.505 4349.505 378.785 4349.785 ;
        RECT 369.275 4348.795 369.555 4349.075 ;
        RECT 369.985 4348.795 370.265 4349.075 ;
        RECT 370.695 4348.795 370.975 4349.075 ;
        RECT 371.405 4348.795 371.685 4349.075 ;
        RECT 372.115 4348.795 372.395 4349.075 ;
        RECT 372.825 4348.795 373.105 4349.075 ;
        RECT 373.535 4348.795 373.815 4349.075 ;
        RECT 374.245 4348.795 374.525 4349.075 ;
        RECT 374.955 4348.795 375.235 4349.075 ;
        RECT 375.665 4348.795 375.945 4349.075 ;
        RECT 376.375 4348.795 376.655 4349.075 ;
        RECT 377.085 4348.795 377.365 4349.075 ;
        RECT 377.795 4348.795 378.075 4349.075 ;
        RECT 378.505 4348.795 378.785 4349.075 ;
        RECT 369.275 4348.085 369.555 4348.365 ;
        RECT 369.985 4348.085 370.265 4348.365 ;
        RECT 370.695 4348.085 370.975 4348.365 ;
        RECT 371.405 4348.085 371.685 4348.365 ;
        RECT 372.115 4348.085 372.395 4348.365 ;
        RECT 372.825 4348.085 373.105 4348.365 ;
        RECT 373.535 4348.085 373.815 4348.365 ;
        RECT 374.245 4348.085 374.525 4348.365 ;
        RECT 374.955 4348.085 375.235 4348.365 ;
        RECT 375.665 4348.085 375.945 4348.365 ;
        RECT 376.375 4348.085 376.655 4348.365 ;
        RECT 377.085 4348.085 377.365 4348.365 ;
        RECT 377.795 4348.085 378.075 4348.365 ;
        RECT 378.505 4348.085 378.785 4348.365 ;
        RECT 369.275 4347.375 369.555 4347.655 ;
        RECT 369.985 4347.375 370.265 4347.655 ;
        RECT 370.695 4347.375 370.975 4347.655 ;
        RECT 371.405 4347.375 371.685 4347.655 ;
        RECT 372.115 4347.375 372.395 4347.655 ;
        RECT 372.825 4347.375 373.105 4347.655 ;
        RECT 373.535 4347.375 373.815 4347.655 ;
        RECT 374.245 4347.375 374.525 4347.655 ;
        RECT 374.955 4347.375 375.235 4347.655 ;
        RECT 375.665 4347.375 375.945 4347.655 ;
        RECT 376.375 4347.375 376.655 4347.655 ;
        RECT 377.085 4347.375 377.365 4347.655 ;
        RECT 377.795 4347.375 378.075 4347.655 ;
        RECT 378.505 4347.375 378.785 4347.655 ;
        RECT 369.275 4346.665 369.555 4346.945 ;
        RECT 369.985 4346.665 370.265 4346.945 ;
        RECT 370.695 4346.665 370.975 4346.945 ;
        RECT 371.405 4346.665 371.685 4346.945 ;
        RECT 372.115 4346.665 372.395 4346.945 ;
        RECT 372.825 4346.665 373.105 4346.945 ;
        RECT 373.535 4346.665 373.815 4346.945 ;
        RECT 374.245 4346.665 374.525 4346.945 ;
        RECT 374.955 4346.665 375.235 4346.945 ;
        RECT 375.665 4346.665 375.945 4346.945 ;
        RECT 376.375 4346.665 376.655 4346.945 ;
        RECT 377.085 4346.665 377.365 4346.945 ;
        RECT 377.795 4346.665 378.075 4346.945 ;
        RECT 378.505 4346.665 378.785 4346.945 ;
        RECT 369.275 4345.955 369.555 4346.235 ;
        RECT 369.985 4345.955 370.265 4346.235 ;
        RECT 370.695 4345.955 370.975 4346.235 ;
        RECT 371.405 4345.955 371.685 4346.235 ;
        RECT 372.115 4345.955 372.395 4346.235 ;
        RECT 372.825 4345.955 373.105 4346.235 ;
        RECT 373.535 4345.955 373.815 4346.235 ;
        RECT 374.245 4345.955 374.525 4346.235 ;
        RECT 374.955 4345.955 375.235 4346.235 ;
        RECT 375.665 4345.955 375.945 4346.235 ;
        RECT 376.375 4345.955 376.655 4346.235 ;
        RECT 377.085 4345.955 377.365 4346.235 ;
        RECT 377.795 4345.955 378.075 4346.235 ;
        RECT 378.505 4345.955 378.785 4346.235 ;
        RECT 3500.255 4350.235 3500.535 4350.515 ;
        RECT 3500.965 4350.235 3501.245 4350.515 ;
        RECT 3501.675 4350.235 3501.955 4350.515 ;
        RECT 3502.385 4350.235 3502.665 4350.515 ;
        RECT 3503.095 4350.235 3503.375 4350.515 ;
        RECT 3503.805 4350.235 3504.085 4350.515 ;
        RECT 3504.515 4350.235 3504.795 4350.515 ;
        RECT 3505.225 4350.235 3505.505 4350.515 ;
        RECT 3505.935 4350.235 3506.215 4350.515 ;
        RECT 3506.645 4350.235 3506.925 4350.515 ;
        RECT 3507.355 4350.235 3507.635 4350.515 ;
        RECT 3508.065 4350.235 3508.345 4350.515 ;
        RECT 3508.775 4350.235 3509.055 4350.515 ;
        RECT 3509.485 4350.235 3509.765 4350.515 ;
        RECT 3500.255 4349.525 3500.535 4349.805 ;
        RECT 3500.965 4349.525 3501.245 4349.805 ;
        RECT 3501.675 4349.525 3501.955 4349.805 ;
        RECT 3502.385 4349.525 3502.665 4349.805 ;
        RECT 3503.095 4349.525 3503.375 4349.805 ;
        RECT 3503.805 4349.525 3504.085 4349.805 ;
        RECT 3504.515 4349.525 3504.795 4349.805 ;
        RECT 3505.225 4349.525 3505.505 4349.805 ;
        RECT 3505.935 4349.525 3506.215 4349.805 ;
        RECT 3506.645 4349.525 3506.925 4349.805 ;
        RECT 3507.355 4349.525 3507.635 4349.805 ;
        RECT 3508.065 4349.525 3508.345 4349.805 ;
        RECT 3508.775 4349.525 3509.055 4349.805 ;
        RECT 3509.485 4349.525 3509.765 4349.805 ;
        RECT 3500.255 4348.815 3500.535 4349.095 ;
        RECT 3500.965 4348.815 3501.245 4349.095 ;
        RECT 3501.675 4348.815 3501.955 4349.095 ;
        RECT 3502.385 4348.815 3502.665 4349.095 ;
        RECT 3503.095 4348.815 3503.375 4349.095 ;
        RECT 3503.805 4348.815 3504.085 4349.095 ;
        RECT 3504.515 4348.815 3504.795 4349.095 ;
        RECT 3505.225 4348.815 3505.505 4349.095 ;
        RECT 3505.935 4348.815 3506.215 4349.095 ;
        RECT 3506.645 4348.815 3506.925 4349.095 ;
        RECT 3507.355 4348.815 3507.635 4349.095 ;
        RECT 3508.065 4348.815 3508.345 4349.095 ;
        RECT 3508.775 4348.815 3509.055 4349.095 ;
        RECT 3509.485 4348.815 3509.765 4349.095 ;
        RECT 3500.255 4348.105 3500.535 4348.385 ;
        RECT 3500.965 4348.105 3501.245 4348.385 ;
        RECT 3501.675 4348.105 3501.955 4348.385 ;
        RECT 3502.385 4348.105 3502.665 4348.385 ;
        RECT 3503.095 4348.105 3503.375 4348.385 ;
        RECT 3503.805 4348.105 3504.085 4348.385 ;
        RECT 3504.515 4348.105 3504.795 4348.385 ;
        RECT 3505.225 4348.105 3505.505 4348.385 ;
        RECT 3505.935 4348.105 3506.215 4348.385 ;
        RECT 3506.645 4348.105 3506.925 4348.385 ;
        RECT 3507.355 4348.105 3507.635 4348.385 ;
        RECT 3508.065 4348.105 3508.345 4348.385 ;
        RECT 3508.775 4348.105 3509.055 4348.385 ;
        RECT 3509.485 4348.105 3509.765 4348.385 ;
        RECT 3500.255 4347.395 3500.535 4347.675 ;
        RECT 3500.965 4347.395 3501.245 4347.675 ;
        RECT 3501.675 4347.395 3501.955 4347.675 ;
        RECT 3502.385 4347.395 3502.665 4347.675 ;
        RECT 3503.095 4347.395 3503.375 4347.675 ;
        RECT 3503.805 4347.395 3504.085 4347.675 ;
        RECT 3504.515 4347.395 3504.795 4347.675 ;
        RECT 3505.225 4347.395 3505.505 4347.675 ;
        RECT 3505.935 4347.395 3506.215 4347.675 ;
        RECT 3506.645 4347.395 3506.925 4347.675 ;
        RECT 3507.355 4347.395 3507.635 4347.675 ;
        RECT 3508.065 4347.395 3508.345 4347.675 ;
        RECT 3508.775 4347.395 3509.055 4347.675 ;
        RECT 3509.485 4347.395 3509.765 4347.675 ;
        RECT 3500.255 4346.685 3500.535 4346.965 ;
        RECT 3500.965 4346.685 3501.245 4346.965 ;
        RECT 3501.675 4346.685 3501.955 4346.965 ;
        RECT 3502.385 4346.685 3502.665 4346.965 ;
        RECT 3503.095 4346.685 3503.375 4346.965 ;
        RECT 3503.805 4346.685 3504.085 4346.965 ;
        RECT 3504.515 4346.685 3504.795 4346.965 ;
        RECT 3505.225 4346.685 3505.505 4346.965 ;
        RECT 3505.935 4346.685 3506.215 4346.965 ;
        RECT 3506.645 4346.685 3506.925 4346.965 ;
        RECT 3507.355 4346.685 3507.635 4346.965 ;
        RECT 3508.065 4346.685 3508.345 4346.965 ;
        RECT 3508.775 4346.685 3509.055 4346.965 ;
        RECT 3509.485 4346.685 3509.765 4346.965 ;
        RECT 3500.255 4345.975 3500.535 4346.255 ;
        RECT 3500.965 4345.975 3501.245 4346.255 ;
        RECT 3501.675 4345.975 3501.955 4346.255 ;
        RECT 3502.385 4345.975 3502.665 4346.255 ;
        RECT 3503.095 4345.975 3503.375 4346.255 ;
        RECT 3503.805 4345.975 3504.085 4346.255 ;
        RECT 3504.515 4345.975 3504.795 4346.255 ;
        RECT 3505.225 4345.975 3505.505 4346.255 ;
        RECT 3505.935 4345.975 3506.215 4346.255 ;
        RECT 3506.645 4345.975 3506.925 4346.255 ;
        RECT 3507.355 4345.975 3507.635 4346.255 ;
        RECT 3508.065 4345.975 3508.345 4346.255 ;
        RECT 3508.775 4345.975 3509.055 4346.255 ;
        RECT 3509.485 4345.975 3509.765 4346.255 ;
        RECT 3500.255 4345.265 3500.535 4345.545 ;
        RECT 3500.965 4345.265 3501.245 4345.545 ;
        RECT 3501.675 4345.265 3501.955 4345.545 ;
        RECT 3502.385 4345.265 3502.665 4345.545 ;
        RECT 3503.095 4345.265 3503.375 4345.545 ;
        RECT 3503.805 4345.265 3504.085 4345.545 ;
        RECT 3504.515 4345.265 3504.795 4345.545 ;
        RECT 3505.225 4345.265 3505.505 4345.545 ;
        RECT 3505.935 4345.265 3506.215 4345.545 ;
        RECT 3506.645 4345.265 3506.925 4345.545 ;
        RECT 3507.355 4345.265 3507.635 4345.545 ;
        RECT 3508.065 4345.265 3508.345 4345.545 ;
        RECT 3508.775 4345.265 3509.055 4345.545 ;
        RECT 3509.485 4345.265 3509.765 4345.545 ;
        RECT 3500.255 4344.555 3500.535 4344.835 ;
        RECT 3500.965 4344.555 3501.245 4344.835 ;
        RECT 3501.675 4344.555 3501.955 4344.835 ;
        RECT 3502.385 4344.555 3502.665 4344.835 ;
        RECT 3503.095 4344.555 3503.375 4344.835 ;
        RECT 3503.805 4344.555 3504.085 4344.835 ;
        RECT 3504.515 4344.555 3504.795 4344.835 ;
        RECT 3505.225 4344.555 3505.505 4344.835 ;
        RECT 3505.935 4344.555 3506.215 4344.835 ;
        RECT 3506.645 4344.555 3506.925 4344.835 ;
        RECT 3507.355 4344.555 3507.635 4344.835 ;
        RECT 3508.065 4344.555 3508.345 4344.835 ;
        RECT 3508.775 4344.555 3509.055 4344.835 ;
        RECT 3509.485 4344.555 3509.765 4344.835 ;
        RECT 369.275 4343.335 369.555 4343.615 ;
        RECT 369.985 4343.335 370.265 4343.615 ;
        RECT 370.695 4343.335 370.975 4343.615 ;
        RECT 371.405 4343.335 371.685 4343.615 ;
        RECT 372.115 4343.335 372.395 4343.615 ;
        RECT 372.825 4343.335 373.105 4343.615 ;
        RECT 373.535 4343.335 373.815 4343.615 ;
        RECT 374.245 4343.335 374.525 4343.615 ;
        RECT 374.955 4343.335 375.235 4343.615 ;
        RECT 375.665 4343.335 375.945 4343.615 ;
        RECT 376.375 4343.335 376.655 4343.615 ;
        RECT 377.085 4343.335 377.365 4343.615 ;
        RECT 377.795 4343.335 378.075 4343.615 ;
        RECT 378.505 4343.335 378.785 4343.615 ;
        RECT 369.275 4342.625 369.555 4342.905 ;
        RECT 369.985 4342.625 370.265 4342.905 ;
        RECT 370.695 4342.625 370.975 4342.905 ;
        RECT 371.405 4342.625 371.685 4342.905 ;
        RECT 372.115 4342.625 372.395 4342.905 ;
        RECT 372.825 4342.625 373.105 4342.905 ;
        RECT 373.535 4342.625 373.815 4342.905 ;
        RECT 374.245 4342.625 374.525 4342.905 ;
        RECT 374.955 4342.625 375.235 4342.905 ;
        RECT 375.665 4342.625 375.945 4342.905 ;
        RECT 376.375 4342.625 376.655 4342.905 ;
        RECT 377.085 4342.625 377.365 4342.905 ;
        RECT 377.795 4342.625 378.075 4342.905 ;
        RECT 378.505 4342.625 378.785 4342.905 ;
        RECT 369.275 4341.915 369.555 4342.195 ;
        RECT 369.985 4341.915 370.265 4342.195 ;
        RECT 370.695 4341.915 370.975 4342.195 ;
        RECT 371.405 4341.915 371.685 4342.195 ;
        RECT 372.115 4341.915 372.395 4342.195 ;
        RECT 372.825 4341.915 373.105 4342.195 ;
        RECT 373.535 4341.915 373.815 4342.195 ;
        RECT 374.245 4341.915 374.525 4342.195 ;
        RECT 374.955 4341.915 375.235 4342.195 ;
        RECT 375.665 4341.915 375.945 4342.195 ;
        RECT 376.375 4341.915 376.655 4342.195 ;
        RECT 377.085 4341.915 377.365 4342.195 ;
        RECT 377.795 4341.915 378.075 4342.195 ;
        RECT 378.505 4341.915 378.785 4342.195 ;
        RECT 369.275 4341.205 369.555 4341.485 ;
        RECT 369.985 4341.205 370.265 4341.485 ;
        RECT 370.695 4341.205 370.975 4341.485 ;
        RECT 371.405 4341.205 371.685 4341.485 ;
        RECT 372.115 4341.205 372.395 4341.485 ;
        RECT 372.825 4341.205 373.105 4341.485 ;
        RECT 373.535 4341.205 373.815 4341.485 ;
        RECT 374.245 4341.205 374.525 4341.485 ;
        RECT 374.955 4341.205 375.235 4341.485 ;
        RECT 375.665 4341.205 375.945 4341.485 ;
        RECT 376.375 4341.205 376.655 4341.485 ;
        RECT 377.085 4341.205 377.365 4341.485 ;
        RECT 377.795 4341.205 378.075 4341.485 ;
        RECT 378.505 4341.205 378.785 4341.485 ;
        RECT 369.275 4340.495 369.555 4340.775 ;
        RECT 369.985 4340.495 370.265 4340.775 ;
        RECT 370.695 4340.495 370.975 4340.775 ;
        RECT 371.405 4340.495 371.685 4340.775 ;
        RECT 372.115 4340.495 372.395 4340.775 ;
        RECT 372.825 4340.495 373.105 4340.775 ;
        RECT 373.535 4340.495 373.815 4340.775 ;
        RECT 374.245 4340.495 374.525 4340.775 ;
        RECT 374.955 4340.495 375.235 4340.775 ;
        RECT 375.665 4340.495 375.945 4340.775 ;
        RECT 376.375 4340.495 376.655 4340.775 ;
        RECT 377.085 4340.495 377.365 4340.775 ;
        RECT 377.795 4340.495 378.075 4340.775 ;
        RECT 378.505 4340.495 378.785 4340.775 ;
        RECT 3500.255 4343.845 3500.535 4344.125 ;
        RECT 3500.965 4343.845 3501.245 4344.125 ;
        RECT 3501.675 4343.845 3501.955 4344.125 ;
        RECT 3502.385 4343.845 3502.665 4344.125 ;
        RECT 3503.095 4343.845 3503.375 4344.125 ;
        RECT 3503.805 4343.845 3504.085 4344.125 ;
        RECT 3504.515 4343.845 3504.795 4344.125 ;
        RECT 3505.225 4343.845 3505.505 4344.125 ;
        RECT 3505.935 4343.845 3506.215 4344.125 ;
        RECT 3506.645 4343.845 3506.925 4344.125 ;
        RECT 3507.355 4343.845 3507.635 4344.125 ;
        RECT 3508.065 4343.845 3508.345 4344.125 ;
        RECT 3508.775 4343.845 3509.055 4344.125 ;
        RECT 3509.485 4343.845 3509.765 4344.125 ;
        RECT 3500.255 4343.135 3500.535 4343.415 ;
        RECT 3500.965 4343.135 3501.245 4343.415 ;
        RECT 3501.675 4343.135 3501.955 4343.415 ;
        RECT 3502.385 4343.135 3502.665 4343.415 ;
        RECT 3503.095 4343.135 3503.375 4343.415 ;
        RECT 3503.805 4343.135 3504.085 4343.415 ;
        RECT 3504.515 4343.135 3504.795 4343.415 ;
        RECT 3505.225 4343.135 3505.505 4343.415 ;
        RECT 3505.935 4343.135 3506.215 4343.415 ;
        RECT 3506.645 4343.135 3506.925 4343.415 ;
        RECT 3507.355 4343.135 3507.635 4343.415 ;
        RECT 3508.065 4343.135 3508.345 4343.415 ;
        RECT 3508.775 4343.135 3509.055 4343.415 ;
        RECT 3509.485 4343.135 3509.765 4343.415 ;
        RECT 3500.255 4342.425 3500.535 4342.705 ;
        RECT 3500.965 4342.425 3501.245 4342.705 ;
        RECT 3501.675 4342.425 3501.955 4342.705 ;
        RECT 3502.385 4342.425 3502.665 4342.705 ;
        RECT 3503.095 4342.425 3503.375 4342.705 ;
        RECT 3503.805 4342.425 3504.085 4342.705 ;
        RECT 3504.515 4342.425 3504.795 4342.705 ;
        RECT 3505.225 4342.425 3505.505 4342.705 ;
        RECT 3505.935 4342.425 3506.215 4342.705 ;
        RECT 3506.645 4342.425 3506.925 4342.705 ;
        RECT 3507.355 4342.425 3507.635 4342.705 ;
        RECT 3508.065 4342.425 3508.345 4342.705 ;
        RECT 3508.775 4342.425 3509.055 4342.705 ;
        RECT 3509.485 4342.425 3509.765 4342.705 ;
        RECT 3500.255 4341.715 3500.535 4341.995 ;
        RECT 3500.965 4341.715 3501.245 4341.995 ;
        RECT 3501.675 4341.715 3501.955 4341.995 ;
        RECT 3502.385 4341.715 3502.665 4341.995 ;
        RECT 3503.095 4341.715 3503.375 4341.995 ;
        RECT 3503.805 4341.715 3504.085 4341.995 ;
        RECT 3504.515 4341.715 3504.795 4341.995 ;
        RECT 3505.225 4341.715 3505.505 4341.995 ;
        RECT 3505.935 4341.715 3506.215 4341.995 ;
        RECT 3506.645 4341.715 3506.925 4341.995 ;
        RECT 3507.355 4341.715 3507.635 4341.995 ;
        RECT 3508.065 4341.715 3508.345 4341.995 ;
        RECT 3508.775 4341.715 3509.055 4341.995 ;
        RECT 3509.485 4341.715 3509.765 4341.995 ;
        RECT 3500.255 4341.005 3500.535 4341.285 ;
        RECT 3500.965 4341.005 3501.245 4341.285 ;
        RECT 3501.675 4341.005 3501.955 4341.285 ;
        RECT 3502.385 4341.005 3502.665 4341.285 ;
        RECT 3503.095 4341.005 3503.375 4341.285 ;
        RECT 3503.805 4341.005 3504.085 4341.285 ;
        RECT 3504.515 4341.005 3504.795 4341.285 ;
        RECT 3505.225 4341.005 3505.505 4341.285 ;
        RECT 3505.935 4341.005 3506.215 4341.285 ;
        RECT 3506.645 4341.005 3506.925 4341.285 ;
        RECT 3507.355 4341.005 3507.635 4341.285 ;
        RECT 3508.065 4341.005 3508.345 4341.285 ;
        RECT 3508.775 4341.005 3509.055 4341.285 ;
        RECT 3509.485 4341.005 3509.765 4341.285 ;
        RECT 369.275 4339.785 369.555 4340.065 ;
        RECT 369.985 4339.785 370.265 4340.065 ;
        RECT 370.695 4339.785 370.975 4340.065 ;
        RECT 371.405 4339.785 371.685 4340.065 ;
        RECT 372.115 4339.785 372.395 4340.065 ;
        RECT 372.825 4339.785 373.105 4340.065 ;
        RECT 373.535 4339.785 373.815 4340.065 ;
        RECT 374.245 4339.785 374.525 4340.065 ;
        RECT 374.955 4339.785 375.235 4340.065 ;
        RECT 375.665 4339.785 375.945 4340.065 ;
        RECT 376.375 4339.785 376.655 4340.065 ;
        RECT 377.085 4339.785 377.365 4340.065 ;
        RECT 377.795 4339.785 378.075 4340.065 ;
        RECT 378.505 4339.785 378.785 4340.065 ;
        RECT 369.275 4339.075 369.555 4339.355 ;
        RECT 369.985 4339.075 370.265 4339.355 ;
        RECT 370.695 4339.075 370.975 4339.355 ;
        RECT 371.405 4339.075 371.685 4339.355 ;
        RECT 372.115 4339.075 372.395 4339.355 ;
        RECT 372.825 4339.075 373.105 4339.355 ;
        RECT 373.535 4339.075 373.815 4339.355 ;
        RECT 374.245 4339.075 374.525 4339.355 ;
        RECT 374.955 4339.075 375.235 4339.355 ;
        RECT 375.665 4339.075 375.945 4339.355 ;
        RECT 376.375 4339.075 376.655 4339.355 ;
        RECT 377.085 4339.075 377.365 4339.355 ;
        RECT 377.795 4339.075 378.075 4339.355 ;
        RECT 378.505 4339.075 378.785 4339.355 ;
        RECT 369.275 4338.365 369.555 4338.645 ;
        RECT 369.985 4338.365 370.265 4338.645 ;
        RECT 370.695 4338.365 370.975 4338.645 ;
        RECT 371.405 4338.365 371.685 4338.645 ;
        RECT 372.115 4338.365 372.395 4338.645 ;
        RECT 372.825 4338.365 373.105 4338.645 ;
        RECT 373.535 4338.365 373.815 4338.645 ;
        RECT 374.245 4338.365 374.525 4338.645 ;
        RECT 374.955 4338.365 375.235 4338.645 ;
        RECT 375.665 4338.365 375.945 4338.645 ;
        RECT 376.375 4338.365 376.655 4338.645 ;
        RECT 377.085 4338.365 377.365 4338.645 ;
        RECT 377.795 4338.365 378.075 4338.645 ;
        RECT 378.505 4338.365 378.785 4338.645 ;
        RECT 369.275 4337.655 369.555 4337.935 ;
        RECT 369.985 4337.655 370.265 4337.935 ;
        RECT 370.695 4337.655 370.975 4337.935 ;
        RECT 371.405 4337.655 371.685 4337.935 ;
        RECT 372.115 4337.655 372.395 4337.935 ;
        RECT 372.825 4337.655 373.105 4337.935 ;
        RECT 373.535 4337.655 373.815 4337.935 ;
        RECT 374.245 4337.655 374.525 4337.935 ;
        RECT 374.955 4337.655 375.235 4337.935 ;
        RECT 375.665 4337.655 375.945 4337.935 ;
        RECT 376.375 4337.655 376.655 4337.935 ;
        RECT 377.085 4337.655 377.365 4337.935 ;
        RECT 377.795 4337.655 378.075 4337.935 ;
        RECT 378.505 4337.655 378.785 4337.935 ;
        RECT 369.275 4336.945 369.555 4337.225 ;
        RECT 369.985 4336.945 370.265 4337.225 ;
        RECT 370.695 4336.945 370.975 4337.225 ;
        RECT 371.405 4336.945 371.685 4337.225 ;
        RECT 372.115 4336.945 372.395 4337.225 ;
        RECT 372.825 4336.945 373.105 4337.225 ;
        RECT 373.535 4336.945 373.815 4337.225 ;
        RECT 374.245 4336.945 374.525 4337.225 ;
        RECT 374.955 4336.945 375.235 4337.225 ;
        RECT 375.665 4336.945 375.945 4337.225 ;
        RECT 376.375 4336.945 376.655 4337.225 ;
        RECT 377.085 4336.945 377.365 4337.225 ;
        RECT 377.795 4336.945 378.075 4337.225 ;
        RECT 378.505 4336.945 378.785 4337.225 ;
        RECT 369.275 4336.235 369.555 4336.515 ;
        RECT 369.985 4336.235 370.265 4336.515 ;
        RECT 370.695 4336.235 370.975 4336.515 ;
        RECT 371.405 4336.235 371.685 4336.515 ;
        RECT 372.115 4336.235 372.395 4336.515 ;
        RECT 372.825 4336.235 373.105 4336.515 ;
        RECT 373.535 4336.235 373.815 4336.515 ;
        RECT 374.245 4336.235 374.525 4336.515 ;
        RECT 374.955 4336.235 375.235 4336.515 ;
        RECT 375.665 4336.235 375.945 4336.515 ;
        RECT 376.375 4336.235 376.655 4336.515 ;
        RECT 377.085 4336.235 377.365 4336.515 ;
        RECT 377.795 4336.235 378.075 4336.515 ;
        RECT 378.505 4336.235 378.785 4336.515 ;
        RECT 369.275 4335.525 369.555 4335.805 ;
        RECT 369.985 4335.525 370.265 4335.805 ;
        RECT 370.695 4335.525 370.975 4335.805 ;
        RECT 371.405 4335.525 371.685 4335.805 ;
        RECT 372.115 4335.525 372.395 4335.805 ;
        RECT 372.825 4335.525 373.105 4335.805 ;
        RECT 373.535 4335.525 373.815 4335.805 ;
        RECT 374.245 4335.525 374.525 4335.805 ;
        RECT 374.955 4335.525 375.235 4335.805 ;
        RECT 375.665 4335.525 375.945 4335.805 ;
        RECT 376.375 4335.525 376.655 4335.805 ;
        RECT 377.085 4335.525 377.365 4335.805 ;
        RECT 377.795 4335.525 378.075 4335.805 ;
        RECT 378.505 4335.525 378.785 4335.805 ;
        RECT 369.275 4334.815 369.555 4335.095 ;
        RECT 369.985 4334.815 370.265 4335.095 ;
        RECT 370.695 4334.815 370.975 4335.095 ;
        RECT 371.405 4334.815 371.685 4335.095 ;
        RECT 372.115 4334.815 372.395 4335.095 ;
        RECT 372.825 4334.815 373.105 4335.095 ;
        RECT 373.535 4334.815 373.815 4335.095 ;
        RECT 374.245 4334.815 374.525 4335.095 ;
        RECT 374.955 4334.815 375.235 4335.095 ;
        RECT 375.665 4334.815 375.945 4335.095 ;
        RECT 376.375 4334.815 376.655 4335.095 ;
        RECT 377.085 4334.815 377.365 4335.095 ;
        RECT 377.795 4334.815 378.075 4335.095 ;
        RECT 378.505 4334.815 378.785 4335.095 ;
        RECT 369.275 4334.105 369.555 4334.385 ;
        RECT 369.985 4334.105 370.265 4334.385 ;
        RECT 370.695 4334.105 370.975 4334.385 ;
        RECT 371.405 4334.105 371.685 4334.385 ;
        RECT 372.115 4334.105 372.395 4334.385 ;
        RECT 372.825 4334.105 373.105 4334.385 ;
        RECT 373.535 4334.105 373.815 4334.385 ;
        RECT 374.245 4334.105 374.525 4334.385 ;
        RECT 374.955 4334.105 375.235 4334.385 ;
        RECT 375.665 4334.105 375.945 4334.385 ;
        RECT 376.375 4334.105 376.655 4334.385 ;
        RECT 377.085 4334.105 377.365 4334.385 ;
        RECT 377.795 4334.105 378.075 4334.385 ;
        RECT 378.505 4334.105 378.785 4334.385 ;
        RECT 3500.255 4338.385 3500.535 4338.665 ;
        RECT 3500.965 4338.385 3501.245 4338.665 ;
        RECT 3501.675 4338.385 3501.955 4338.665 ;
        RECT 3502.385 4338.385 3502.665 4338.665 ;
        RECT 3503.095 4338.385 3503.375 4338.665 ;
        RECT 3503.805 4338.385 3504.085 4338.665 ;
        RECT 3504.515 4338.385 3504.795 4338.665 ;
        RECT 3505.225 4338.385 3505.505 4338.665 ;
        RECT 3505.935 4338.385 3506.215 4338.665 ;
        RECT 3506.645 4338.385 3506.925 4338.665 ;
        RECT 3507.355 4338.385 3507.635 4338.665 ;
        RECT 3508.065 4338.385 3508.345 4338.665 ;
        RECT 3508.775 4338.385 3509.055 4338.665 ;
        RECT 3509.485 4338.385 3509.765 4338.665 ;
        RECT 3500.255 4337.675 3500.535 4337.955 ;
        RECT 3500.965 4337.675 3501.245 4337.955 ;
        RECT 3501.675 4337.675 3501.955 4337.955 ;
        RECT 3502.385 4337.675 3502.665 4337.955 ;
        RECT 3503.095 4337.675 3503.375 4337.955 ;
        RECT 3503.805 4337.675 3504.085 4337.955 ;
        RECT 3504.515 4337.675 3504.795 4337.955 ;
        RECT 3505.225 4337.675 3505.505 4337.955 ;
        RECT 3505.935 4337.675 3506.215 4337.955 ;
        RECT 3506.645 4337.675 3506.925 4337.955 ;
        RECT 3507.355 4337.675 3507.635 4337.955 ;
        RECT 3508.065 4337.675 3508.345 4337.955 ;
        RECT 3508.775 4337.675 3509.055 4337.955 ;
        RECT 3509.485 4337.675 3509.765 4337.955 ;
        RECT 3500.255 4336.965 3500.535 4337.245 ;
        RECT 3500.965 4336.965 3501.245 4337.245 ;
        RECT 3501.675 4336.965 3501.955 4337.245 ;
        RECT 3502.385 4336.965 3502.665 4337.245 ;
        RECT 3503.095 4336.965 3503.375 4337.245 ;
        RECT 3503.805 4336.965 3504.085 4337.245 ;
        RECT 3504.515 4336.965 3504.795 4337.245 ;
        RECT 3505.225 4336.965 3505.505 4337.245 ;
        RECT 3505.935 4336.965 3506.215 4337.245 ;
        RECT 3506.645 4336.965 3506.925 4337.245 ;
        RECT 3507.355 4336.965 3507.635 4337.245 ;
        RECT 3508.065 4336.965 3508.345 4337.245 ;
        RECT 3508.775 4336.965 3509.055 4337.245 ;
        RECT 3509.485 4336.965 3509.765 4337.245 ;
        RECT 3500.255 4336.255 3500.535 4336.535 ;
        RECT 3500.965 4336.255 3501.245 4336.535 ;
        RECT 3501.675 4336.255 3501.955 4336.535 ;
        RECT 3502.385 4336.255 3502.665 4336.535 ;
        RECT 3503.095 4336.255 3503.375 4336.535 ;
        RECT 3503.805 4336.255 3504.085 4336.535 ;
        RECT 3504.515 4336.255 3504.795 4336.535 ;
        RECT 3505.225 4336.255 3505.505 4336.535 ;
        RECT 3505.935 4336.255 3506.215 4336.535 ;
        RECT 3506.645 4336.255 3506.925 4336.535 ;
        RECT 3507.355 4336.255 3507.635 4336.535 ;
        RECT 3508.065 4336.255 3508.345 4336.535 ;
        RECT 3508.775 4336.255 3509.055 4336.535 ;
        RECT 3509.485 4336.255 3509.765 4336.535 ;
        RECT 3500.255 4335.545 3500.535 4335.825 ;
        RECT 3500.965 4335.545 3501.245 4335.825 ;
        RECT 3501.675 4335.545 3501.955 4335.825 ;
        RECT 3502.385 4335.545 3502.665 4335.825 ;
        RECT 3503.095 4335.545 3503.375 4335.825 ;
        RECT 3503.805 4335.545 3504.085 4335.825 ;
        RECT 3504.515 4335.545 3504.795 4335.825 ;
        RECT 3505.225 4335.545 3505.505 4335.825 ;
        RECT 3505.935 4335.545 3506.215 4335.825 ;
        RECT 3506.645 4335.545 3506.925 4335.825 ;
        RECT 3507.355 4335.545 3507.635 4335.825 ;
        RECT 3508.065 4335.545 3508.345 4335.825 ;
        RECT 3508.775 4335.545 3509.055 4335.825 ;
        RECT 3509.485 4335.545 3509.765 4335.825 ;
        RECT 3500.255 4334.835 3500.535 4335.115 ;
        RECT 3500.965 4334.835 3501.245 4335.115 ;
        RECT 3501.675 4334.835 3501.955 4335.115 ;
        RECT 3502.385 4334.835 3502.665 4335.115 ;
        RECT 3503.095 4334.835 3503.375 4335.115 ;
        RECT 3503.805 4334.835 3504.085 4335.115 ;
        RECT 3504.515 4334.835 3504.795 4335.115 ;
        RECT 3505.225 4334.835 3505.505 4335.115 ;
        RECT 3505.935 4334.835 3506.215 4335.115 ;
        RECT 3506.645 4334.835 3506.925 4335.115 ;
        RECT 3507.355 4334.835 3507.635 4335.115 ;
        RECT 3508.065 4334.835 3508.345 4335.115 ;
        RECT 3508.775 4334.835 3509.055 4335.115 ;
        RECT 3509.485 4334.835 3509.765 4335.115 ;
        RECT 3500.255 4334.125 3500.535 4334.405 ;
        RECT 3500.965 4334.125 3501.245 4334.405 ;
        RECT 3501.675 4334.125 3501.955 4334.405 ;
        RECT 3502.385 4334.125 3502.665 4334.405 ;
        RECT 3503.095 4334.125 3503.375 4334.405 ;
        RECT 3503.805 4334.125 3504.085 4334.405 ;
        RECT 3504.515 4334.125 3504.795 4334.405 ;
        RECT 3505.225 4334.125 3505.505 4334.405 ;
        RECT 3505.935 4334.125 3506.215 4334.405 ;
        RECT 3506.645 4334.125 3506.925 4334.405 ;
        RECT 3507.355 4334.125 3507.635 4334.405 ;
        RECT 3508.065 4334.125 3508.345 4334.405 ;
        RECT 3508.775 4334.125 3509.055 4334.405 ;
        RECT 3509.485 4334.125 3509.765 4334.405 ;
        RECT 3500.255 4333.415 3500.535 4333.695 ;
        RECT 3500.965 4333.415 3501.245 4333.695 ;
        RECT 3501.675 4333.415 3501.955 4333.695 ;
        RECT 3502.385 4333.415 3502.665 4333.695 ;
        RECT 3503.095 4333.415 3503.375 4333.695 ;
        RECT 3503.805 4333.415 3504.085 4333.695 ;
        RECT 3504.515 4333.415 3504.795 4333.695 ;
        RECT 3505.225 4333.415 3505.505 4333.695 ;
        RECT 3505.935 4333.415 3506.215 4333.695 ;
        RECT 3506.645 4333.415 3506.925 4333.695 ;
        RECT 3507.355 4333.415 3507.635 4333.695 ;
        RECT 3508.065 4333.415 3508.345 4333.695 ;
        RECT 3508.775 4333.415 3509.055 4333.695 ;
        RECT 3509.485 4333.415 3509.765 4333.695 ;
        RECT 3500.255 4332.705 3500.535 4332.985 ;
        RECT 3500.965 4332.705 3501.245 4332.985 ;
        RECT 3501.675 4332.705 3501.955 4332.985 ;
        RECT 3502.385 4332.705 3502.665 4332.985 ;
        RECT 3503.095 4332.705 3503.375 4332.985 ;
        RECT 3503.805 4332.705 3504.085 4332.985 ;
        RECT 3504.515 4332.705 3504.795 4332.985 ;
        RECT 3505.225 4332.705 3505.505 4332.985 ;
        RECT 3505.935 4332.705 3506.215 4332.985 ;
        RECT 3506.645 4332.705 3506.925 4332.985 ;
        RECT 3507.355 4332.705 3507.635 4332.985 ;
        RECT 3508.065 4332.705 3508.345 4332.985 ;
        RECT 3508.775 4332.705 3509.055 4332.985 ;
        RECT 3509.485 4332.705 3509.765 4332.985 ;
        RECT 3500.255 4331.995 3500.535 4332.275 ;
        RECT 3500.965 4331.995 3501.245 4332.275 ;
        RECT 3501.675 4331.995 3501.955 4332.275 ;
        RECT 3502.385 4331.995 3502.665 4332.275 ;
        RECT 3503.095 4331.995 3503.375 4332.275 ;
        RECT 3503.805 4331.995 3504.085 4332.275 ;
        RECT 3504.515 4331.995 3504.795 4332.275 ;
        RECT 3505.225 4331.995 3505.505 4332.275 ;
        RECT 3505.935 4331.995 3506.215 4332.275 ;
        RECT 3506.645 4331.995 3506.925 4332.275 ;
        RECT 3507.355 4331.995 3507.635 4332.275 ;
        RECT 3508.065 4331.995 3508.345 4332.275 ;
        RECT 3508.775 4331.995 3509.055 4332.275 ;
        RECT 3509.485 4331.995 3509.765 4332.275 ;
        RECT 3500.255 4331.285 3500.535 4331.565 ;
        RECT 3500.965 4331.285 3501.245 4331.565 ;
        RECT 3501.675 4331.285 3501.955 4331.565 ;
        RECT 3502.385 4331.285 3502.665 4331.565 ;
        RECT 3503.095 4331.285 3503.375 4331.565 ;
        RECT 3503.805 4331.285 3504.085 4331.565 ;
        RECT 3504.515 4331.285 3504.795 4331.565 ;
        RECT 3505.225 4331.285 3505.505 4331.565 ;
        RECT 3505.935 4331.285 3506.215 4331.565 ;
        RECT 3506.645 4331.285 3506.925 4331.565 ;
        RECT 3507.355 4331.285 3507.635 4331.565 ;
        RECT 3508.065 4331.285 3508.345 4331.565 ;
        RECT 3508.775 4331.285 3509.055 4331.565 ;
        RECT 3509.485 4331.285 3509.765 4331.565 ;
        RECT 369.330 4330.190 369.610 4330.470 ;
        RECT 370.040 4330.190 370.320 4330.470 ;
        RECT 370.750 4330.190 371.030 4330.470 ;
        RECT 371.460 4330.190 371.740 4330.470 ;
        RECT 372.170 4330.190 372.450 4330.470 ;
        RECT 372.880 4330.190 373.160 4330.470 ;
        RECT 373.590 4330.190 373.870 4330.470 ;
        RECT 374.300 4330.190 374.580 4330.470 ;
        RECT 375.010 4330.190 375.290 4330.470 ;
        RECT 375.720 4330.190 376.000 4330.470 ;
        RECT 376.430 4330.190 376.710 4330.470 ;
        RECT 377.140 4330.190 377.420 4330.470 ;
        RECT 377.850 4330.190 378.130 4330.470 ;
        RECT 378.560 4330.190 378.840 4330.470 ;
        RECT 369.330 4329.480 369.610 4329.760 ;
        RECT 370.040 4329.480 370.320 4329.760 ;
        RECT 370.750 4329.480 371.030 4329.760 ;
        RECT 371.460 4329.480 371.740 4329.760 ;
        RECT 372.170 4329.480 372.450 4329.760 ;
        RECT 372.880 4329.480 373.160 4329.760 ;
        RECT 373.590 4329.480 373.870 4329.760 ;
        RECT 374.300 4329.480 374.580 4329.760 ;
        RECT 375.010 4329.480 375.290 4329.760 ;
        RECT 375.720 4329.480 376.000 4329.760 ;
        RECT 376.430 4329.480 376.710 4329.760 ;
        RECT 377.140 4329.480 377.420 4329.760 ;
        RECT 377.850 4329.480 378.130 4329.760 ;
        RECT 378.560 4329.480 378.840 4329.760 ;
        RECT 369.330 4328.770 369.610 4329.050 ;
        RECT 370.040 4328.770 370.320 4329.050 ;
        RECT 370.750 4328.770 371.030 4329.050 ;
        RECT 371.460 4328.770 371.740 4329.050 ;
        RECT 372.170 4328.770 372.450 4329.050 ;
        RECT 372.880 4328.770 373.160 4329.050 ;
        RECT 373.590 4328.770 373.870 4329.050 ;
        RECT 374.300 4328.770 374.580 4329.050 ;
        RECT 375.010 4328.770 375.290 4329.050 ;
        RECT 375.720 4328.770 376.000 4329.050 ;
        RECT 376.430 4328.770 376.710 4329.050 ;
        RECT 377.140 4328.770 377.420 4329.050 ;
        RECT 377.850 4328.770 378.130 4329.050 ;
        RECT 378.560 4328.770 378.840 4329.050 ;
        RECT 3500.255 4330.575 3500.535 4330.855 ;
        RECT 3500.965 4330.575 3501.245 4330.855 ;
        RECT 3501.675 4330.575 3501.955 4330.855 ;
        RECT 3502.385 4330.575 3502.665 4330.855 ;
        RECT 3503.095 4330.575 3503.375 4330.855 ;
        RECT 3503.805 4330.575 3504.085 4330.855 ;
        RECT 3504.515 4330.575 3504.795 4330.855 ;
        RECT 3505.225 4330.575 3505.505 4330.855 ;
        RECT 3505.935 4330.575 3506.215 4330.855 ;
        RECT 3506.645 4330.575 3506.925 4330.855 ;
        RECT 3507.355 4330.575 3507.635 4330.855 ;
        RECT 3508.065 4330.575 3508.345 4330.855 ;
        RECT 3508.775 4330.575 3509.055 4330.855 ;
        RECT 3509.485 4330.575 3509.765 4330.855 ;
        RECT 3500.255 4329.865 3500.535 4330.145 ;
        RECT 3500.965 4329.865 3501.245 4330.145 ;
        RECT 3501.675 4329.865 3501.955 4330.145 ;
        RECT 3502.385 4329.865 3502.665 4330.145 ;
        RECT 3503.095 4329.865 3503.375 4330.145 ;
        RECT 3503.805 4329.865 3504.085 4330.145 ;
        RECT 3504.515 4329.865 3504.795 4330.145 ;
        RECT 3505.225 4329.865 3505.505 4330.145 ;
        RECT 3505.935 4329.865 3506.215 4330.145 ;
        RECT 3506.645 4329.865 3506.925 4330.145 ;
        RECT 3507.355 4329.865 3507.635 4330.145 ;
        RECT 3508.065 4329.865 3508.345 4330.145 ;
        RECT 3508.775 4329.865 3509.055 4330.145 ;
        RECT 3509.485 4329.865 3509.765 4330.145 ;
        RECT 3500.255 4329.155 3500.535 4329.435 ;
        RECT 3500.965 4329.155 3501.245 4329.435 ;
        RECT 3501.675 4329.155 3501.955 4329.435 ;
        RECT 3502.385 4329.155 3502.665 4329.435 ;
        RECT 3503.095 4329.155 3503.375 4329.435 ;
        RECT 3503.805 4329.155 3504.085 4329.435 ;
        RECT 3504.515 4329.155 3504.795 4329.435 ;
        RECT 3505.225 4329.155 3505.505 4329.435 ;
        RECT 3505.935 4329.155 3506.215 4329.435 ;
        RECT 3506.645 4329.155 3506.925 4329.435 ;
        RECT 3507.355 4329.155 3507.635 4329.435 ;
        RECT 3508.065 4329.155 3508.345 4329.435 ;
        RECT 3508.775 4329.155 3509.055 4329.435 ;
        RECT 3509.485 4329.155 3509.765 4329.435 ;
        RECT 369.330 4328.060 369.610 4328.340 ;
        RECT 370.040 4328.060 370.320 4328.340 ;
        RECT 370.750 4328.060 371.030 4328.340 ;
        RECT 371.460 4328.060 371.740 4328.340 ;
        RECT 372.170 4328.060 372.450 4328.340 ;
        RECT 372.880 4328.060 373.160 4328.340 ;
        RECT 373.590 4328.060 373.870 4328.340 ;
        RECT 374.300 4328.060 374.580 4328.340 ;
        RECT 375.010 4328.060 375.290 4328.340 ;
        RECT 375.720 4328.060 376.000 4328.340 ;
        RECT 376.430 4328.060 376.710 4328.340 ;
        RECT 377.140 4328.060 377.420 4328.340 ;
        RECT 377.850 4328.060 378.130 4328.340 ;
        RECT 378.560 4328.060 378.840 4328.340 ;
        RECT 369.330 4327.350 369.610 4327.630 ;
        RECT 370.040 4327.350 370.320 4327.630 ;
        RECT 370.750 4327.350 371.030 4327.630 ;
        RECT 371.460 4327.350 371.740 4327.630 ;
        RECT 372.170 4327.350 372.450 4327.630 ;
        RECT 372.880 4327.350 373.160 4327.630 ;
        RECT 373.590 4327.350 373.870 4327.630 ;
        RECT 374.300 4327.350 374.580 4327.630 ;
        RECT 375.010 4327.350 375.290 4327.630 ;
        RECT 375.720 4327.350 376.000 4327.630 ;
        RECT 376.430 4327.350 376.710 4327.630 ;
        RECT 377.140 4327.350 377.420 4327.630 ;
        RECT 377.850 4327.350 378.130 4327.630 ;
        RECT 378.560 4327.350 378.840 4327.630 ;
        RECT 369.330 4326.640 369.610 4326.920 ;
        RECT 370.040 4326.640 370.320 4326.920 ;
        RECT 370.750 4326.640 371.030 4326.920 ;
        RECT 371.460 4326.640 371.740 4326.920 ;
        RECT 372.170 4326.640 372.450 4326.920 ;
        RECT 372.880 4326.640 373.160 4326.920 ;
        RECT 373.590 4326.640 373.870 4326.920 ;
        RECT 374.300 4326.640 374.580 4326.920 ;
        RECT 375.010 4326.640 375.290 4326.920 ;
        RECT 375.720 4326.640 376.000 4326.920 ;
        RECT 376.430 4326.640 376.710 4326.920 ;
        RECT 377.140 4326.640 377.420 4326.920 ;
        RECT 377.850 4326.640 378.130 4326.920 ;
        RECT 378.560 4326.640 378.840 4326.920 ;
        RECT 369.330 4325.930 369.610 4326.210 ;
        RECT 370.040 4325.930 370.320 4326.210 ;
        RECT 370.750 4325.930 371.030 4326.210 ;
        RECT 371.460 4325.930 371.740 4326.210 ;
        RECT 372.170 4325.930 372.450 4326.210 ;
        RECT 372.880 4325.930 373.160 4326.210 ;
        RECT 373.590 4325.930 373.870 4326.210 ;
        RECT 374.300 4325.930 374.580 4326.210 ;
        RECT 375.010 4325.930 375.290 4326.210 ;
        RECT 375.720 4325.930 376.000 4326.210 ;
        RECT 376.430 4325.930 376.710 4326.210 ;
        RECT 377.140 4325.930 377.420 4326.210 ;
        RECT 377.850 4325.930 378.130 4326.210 ;
        RECT 378.560 4325.930 378.840 4326.210 ;
        RECT 369.330 4325.220 369.610 4325.500 ;
        RECT 370.040 4325.220 370.320 4325.500 ;
        RECT 370.750 4325.220 371.030 4325.500 ;
        RECT 371.460 4325.220 371.740 4325.500 ;
        RECT 372.170 4325.220 372.450 4325.500 ;
        RECT 372.880 4325.220 373.160 4325.500 ;
        RECT 373.590 4325.220 373.870 4325.500 ;
        RECT 374.300 4325.220 374.580 4325.500 ;
        RECT 375.010 4325.220 375.290 4325.500 ;
        RECT 375.720 4325.220 376.000 4325.500 ;
        RECT 376.430 4325.220 376.710 4325.500 ;
        RECT 377.140 4325.220 377.420 4325.500 ;
        RECT 377.850 4325.220 378.130 4325.500 ;
        RECT 378.560 4325.220 378.840 4325.500 ;
        RECT 369.330 4324.510 369.610 4324.790 ;
        RECT 370.040 4324.510 370.320 4324.790 ;
        RECT 370.750 4324.510 371.030 4324.790 ;
        RECT 371.460 4324.510 371.740 4324.790 ;
        RECT 372.170 4324.510 372.450 4324.790 ;
        RECT 372.880 4324.510 373.160 4324.790 ;
        RECT 373.590 4324.510 373.870 4324.790 ;
        RECT 374.300 4324.510 374.580 4324.790 ;
        RECT 375.010 4324.510 375.290 4324.790 ;
        RECT 375.720 4324.510 376.000 4324.790 ;
        RECT 376.430 4324.510 376.710 4324.790 ;
        RECT 377.140 4324.510 377.420 4324.790 ;
        RECT 377.850 4324.510 378.130 4324.790 ;
        RECT 378.560 4324.510 378.840 4324.790 ;
        RECT 369.330 4323.800 369.610 4324.080 ;
        RECT 370.040 4323.800 370.320 4324.080 ;
        RECT 370.750 4323.800 371.030 4324.080 ;
        RECT 371.460 4323.800 371.740 4324.080 ;
        RECT 372.170 4323.800 372.450 4324.080 ;
        RECT 372.880 4323.800 373.160 4324.080 ;
        RECT 373.590 4323.800 373.870 4324.080 ;
        RECT 374.300 4323.800 374.580 4324.080 ;
        RECT 375.010 4323.800 375.290 4324.080 ;
        RECT 375.720 4323.800 376.000 4324.080 ;
        RECT 376.430 4323.800 376.710 4324.080 ;
        RECT 377.140 4323.800 377.420 4324.080 ;
        RECT 377.850 4323.800 378.130 4324.080 ;
        RECT 378.560 4323.800 378.840 4324.080 ;
        RECT 369.330 4323.090 369.610 4323.370 ;
        RECT 370.040 4323.090 370.320 4323.370 ;
        RECT 370.750 4323.090 371.030 4323.370 ;
        RECT 371.460 4323.090 371.740 4323.370 ;
        RECT 372.170 4323.090 372.450 4323.370 ;
        RECT 372.880 4323.090 373.160 4323.370 ;
        RECT 373.590 4323.090 373.870 4323.370 ;
        RECT 374.300 4323.090 374.580 4323.370 ;
        RECT 375.010 4323.090 375.290 4323.370 ;
        RECT 375.720 4323.090 376.000 4323.370 ;
        RECT 376.430 4323.090 376.710 4323.370 ;
        RECT 377.140 4323.090 377.420 4323.370 ;
        RECT 377.850 4323.090 378.130 4323.370 ;
        RECT 378.560 4323.090 378.840 4323.370 ;
        RECT 369.330 4322.380 369.610 4322.660 ;
        RECT 370.040 4322.380 370.320 4322.660 ;
        RECT 370.750 4322.380 371.030 4322.660 ;
        RECT 371.460 4322.380 371.740 4322.660 ;
        RECT 372.170 4322.380 372.450 4322.660 ;
        RECT 372.880 4322.380 373.160 4322.660 ;
        RECT 373.590 4322.380 373.870 4322.660 ;
        RECT 374.300 4322.380 374.580 4322.660 ;
        RECT 375.010 4322.380 375.290 4322.660 ;
        RECT 375.720 4322.380 376.000 4322.660 ;
        RECT 376.430 4322.380 376.710 4322.660 ;
        RECT 377.140 4322.380 377.420 4322.660 ;
        RECT 377.850 4322.380 378.130 4322.660 ;
        RECT 378.560 4322.380 378.840 4322.660 ;
        RECT 369.330 4321.670 369.610 4321.950 ;
        RECT 370.040 4321.670 370.320 4321.950 ;
        RECT 370.750 4321.670 371.030 4321.950 ;
        RECT 371.460 4321.670 371.740 4321.950 ;
        RECT 372.170 4321.670 372.450 4321.950 ;
        RECT 372.880 4321.670 373.160 4321.950 ;
        RECT 373.590 4321.670 373.870 4321.950 ;
        RECT 374.300 4321.670 374.580 4321.950 ;
        RECT 375.010 4321.670 375.290 4321.950 ;
        RECT 375.720 4321.670 376.000 4321.950 ;
        RECT 376.430 4321.670 376.710 4321.950 ;
        RECT 377.140 4321.670 377.420 4321.950 ;
        RECT 377.850 4321.670 378.130 4321.950 ;
        RECT 378.560 4321.670 378.840 4321.950 ;
        RECT 3500.200 4325.270 3500.480 4325.550 ;
        RECT 3500.910 4325.270 3501.190 4325.550 ;
        RECT 3501.620 4325.270 3501.900 4325.550 ;
        RECT 3502.330 4325.270 3502.610 4325.550 ;
        RECT 3503.040 4325.270 3503.320 4325.550 ;
        RECT 3503.750 4325.270 3504.030 4325.550 ;
        RECT 3504.460 4325.270 3504.740 4325.550 ;
        RECT 3505.170 4325.270 3505.450 4325.550 ;
        RECT 3505.880 4325.270 3506.160 4325.550 ;
        RECT 3506.590 4325.270 3506.870 4325.550 ;
        RECT 3507.300 4325.270 3507.580 4325.550 ;
        RECT 3508.010 4325.270 3508.290 4325.550 ;
        RECT 3508.720 4325.270 3509.000 4325.550 ;
        RECT 3509.430 4325.270 3509.710 4325.550 ;
        RECT 3500.200 4324.560 3500.480 4324.840 ;
        RECT 3500.910 4324.560 3501.190 4324.840 ;
        RECT 3501.620 4324.560 3501.900 4324.840 ;
        RECT 3502.330 4324.560 3502.610 4324.840 ;
        RECT 3503.040 4324.560 3503.320 4324.840 ;
        RECT 3503.750 4324.560 3504.030 4324.840 ;
        RECT 3504.460 4324.560 3504.740 4324.840 ;
        RECT 3505.170 4324.560 3505.450 4324.840 ;
        RECT 3505.880 4324.560 3506.160 4324.840 ;
        RECT 3506.590 4324.560 3506.870 4324.840 ;
        RECT 3507.300 4324.560 3507.580 4324.840 ;
        RECT 3508.010 4324.560 3508.290 4324.840 ;
        RECT 3508.720 4324.560 3509.000 4324.840 ;
        RECT 3509.430 4324.560 3509.710 4324.840 ;
        RECT 3500.200 4323.850 3500.480 4324.130 ;
        RECT 3500.910 4323.850 3501.190 4324.130 ;
        RECT 3501.620 4323.850 3501.900 4324.130 ;
        RECT 3502.330 4323.850 3502.610 4324.130 ;
        RECT 3503.040 4323.850 3503.320 4324.130 ;
        RECT 3503.750 4323.850 3504.030 4324.130 ;
        RECT 3504.460 4323.850 3504.740 4324.130 ;
        RECT 3505.170 4323.850 3505.450 4324.130 ;
        RECT 3505.880 4323.850 3506.160 4324.130 ;
        RECT 3506.590 4323.850 3506.870 4324.130 ;
        RECT 3507.300 4323.850 3507.580 4324.130 ;
        RECT 3508.010 4323.850 3508.290 4324.130 ;
        RECT 3508.720 4323.850 3509.000 4324.130 ;
        RECT 3509.430 4323.850 3509.710 4324.130 ;
        RECT 3500.200 4323.140 3500.480 4323.420 ;
        RECT 3500.910 4323.140 3501.190 4323.420 ;
        RECT 3501.620 4323.140 3501.900 4323.420 ;
        RECT 3502.330 4323.140 3502.610 4323.420 ;
        RECT 3503.040 4323.140 3503.320 4323.420 ;
        RECT 3503.750 4323.140 3504.030 4323.420 ;
        RECT 3504.460 4323.140 3504.740 4323.420 ;
        RECT 3505.170 4323.140 3505.450 4323.420 ;
        RECT 3505.880 4323.140 3506.160 4323.420 ;
        RECT 3506.590 4323.140 3506.870 4323.420 ;
        RECT 3507.300 4323.140 3507.580 4323.420 ;
        RECT 3508.010 4323.140 3508.290 4323.420 ;
        RECT 3508.720 4323.140 3509.000 4323.420 ;
        RECT 3509.430 4323.140 3509.710 4323.420 ;
        RECT 3500.200 4322.430 3500.480 4322.710 ;
        RECT 3500.910 4322.430 3501.190 4322.710 ;
        RECT 3501.620 4322.430 3501.900 4322.710 ;
        RECT 3502.330 4322.430 3502.610 4322.710 ;
        RECT 3503.040 4322.430 3503.320 4322.710 ;
        RECT 3503.750 4322.430 3504.030 4322.710 ;
        RECT 3504.460 4322.430 3504.740 4322.710 ;
        RECT 3505.170 4322.430 3505.450 4322.710 ;
        RECT 3505.880 4322.430 3506.160 4322.710 ;
        RECT 3506.590 4322.430 3506.870 4322.710 ;
        RECT 3507.300 4322.430 3507.580 4322.710 ;
        RECT 3508.010 4322.430 3508.290 4322.710 ;
        RECT 3508.720 4322.430 3509.000 4322.710 ;
        RECT 3509.430 4322.430 3509.710 4322.710 ;
        RECT 3500.200 4321.720 3500.480 4322.000 ;
        RECT 3500.910 4321.720 3501.190 4322.000 ;
        RECT 3501.620 4321.720 3501.900 4322.000 ;
        RECT 3502.330 4321.720 3502.610 4322.000 ;
        RECT 3503.040 4321.720 3503.320 4322.000 ;
        RECT 3503.750 4321.720 3504.030 4322.000 ;
        RECT 3504.460 4321.720 3504.740 4322.000 ;
        RECT 3505.170 4321.720 3505.450 4322.000 ;
        RECT 3505.880 4321.720 3506.160 4322.000 ;
        RECT 3506.590 4321.720 3506.870 4322.000 ;
        RECT 3507.300 4321.720 3507.580 4322.000 ;
        RECT 3508.010 4321.720 3508.290 4322.000 ;
        RECT 3508.720 4321.720 3509.000 4322.000 ;
        RECT 3509.430 4321.720 3509.710 4322.000 ;
        RECT 3500.200 4321.010 3500.480 4321.290 ;
        RECT 3500.910 4321.010 3501.190 4321.290 ;
        RECT 3501.620 4321.010 3501.900 4321.290 ;
        RECT 3502.330 4321.010 3502.610 4321.290 ;
        RECT 3503.040 4321.010 3503.320 4321.290 ;
        RECT 3503.750 4321.010 3504.030 4321.290 ;
        RECT 3504.460 4321.010 3504.740 4321.290 ;
        RECT 3505.170 4321.010 3505.450 4321.290 ;
        RECT 3505.880 4321.010 3506.160 4321.290 ;
        RECT 3506.590 4321.010 3506.870 4321.290 ;
        RECT 3507.300 4321.010 3507.580 4321.290 ;
        RECT 3508.010 4321.010 3508.290 4321.290 ;
        RECT 3508.720 4321.010 3509.000 4321.290 ;
        RECT 3509.430 4321.010 3509.710 4321.290 ;
        RECT 3500.200 4320.300 3500.480 4320.580 ;
        RECT 3500.910 4320.300 3501.190 4320.580 ;
        RECT 3501.620 4320.300 3501.900 4320.580 ;
        RECT 3502.330 4320.300 3502.610 4320.580 ;
        RECT 3503.040 4320.300 3503.320 4320.580 ;
        RECT 3503.750 4320.300 3504.030 4320.580 ;
        RECT 3504.460 4320.300 3504.740 4320.580 ;
        RECT 3505.170 4320.300 3505.450 4320.580 ;
        RECT 3505.880 4320.300 3506.160 4320.580 ;
        RECT 3506.590 4320.300 3506.870 4320.580 ;
        RECT 3507.300 4320.300 3507.580 4320.580 ;
        RECT 3508.010 4320.300 3508.290 4320.580 ;
        RECT 3508.720 4320.300 3509.000 4320.580 ;
        RECT 3509.430 4320.300 3509.710 4320.580 ;
        RECT 3500.200 4319.590 3500.480 4319.870 ;
        RECT 3500.910 4319.590 3501.190 4319.870 ;
        RECT 3501.620 4319.590 3501.900 4319.870 ;
        RECT 3502.330 4319.590 3502.610 4319.870 ;
        RECT 3503.040 4319.590 3503.320 4319.870 ;
        RECT 3503.750 4319.590 3504.030 4319.870 ;
        RECT 3504.460 4319.590 3504.740 4319.870 ;
        RECT 3505.170 4319.590 3505.450 4319.870 ;
        RECT 3505.880 4319.590 3506.160 4319.870 ;
        RECT 3506.590 4319.590 3506.870 4319.870 ;
        RECT 3507.300 4319.590 3507.580 4319.870 ;
        RECT 3508.010 4319.590 3508.290 4319.870 ;
        RECT 3508.720 4319.590 3509.000 4319.870 ;
        RECT 3509.430 4319.590 3509.710 4319.870 ;
        RECT 3500.200 4318.880 3500.480 4319.160 ;
        RECT 3500.910 4318.880 3501.190 4319.160 ;
        RECT 3501.620 4318.880 3501.900 4319.160 ;
        RECT 3502.330 4318.880 3502.610 4319.160 ;
        RECT 3503.040 4318.880 3503.320 4319.160 ;
        RECT 3503.750 4318.880 3504.030 4319.160 ;
        RECT 3504.460 4318.880 3504.740 4319.160 ;
        RECT 3505.170 4318.880 3505.450 4319.160 ;
        RECT 3505.880 4318.880 3506.160 4319.160 ;
        RECT 3506.590 4318.880 3506.870 4319.160 ;
        RECT 3507.300 4318.880 3507.580 4319.160 ;
        RECT 3508.010 4318.880 3508.290 4319.160 ;
        RECT 3508.720 4318.880 3509.000 4319.160 ;
        RECT 3509.430 4318.880 3509.710 4319.160 ;
        RECT 3500.200 4318.170 3500.480 4318.450 ;
        RECT 3500.910 4318.170 3501.190 4318.450 ;
        RECT 3501.620 4318.170 3501.900 4318.450 ;
        RECT 3502.330 4318.170 3502.610 4318.450 ;
        RECT 3503.040 4318.170 3503.320 4318.450 ;
        RECT 3503.750 4318.170 3504.030 4318.450 ;
        RECT 3504.460 4318.170 3504.740 4318.450 ;
        RECT 3505.170 4318.170 3505.450 4318.450 ;
        RECT 3505.880 4318.170 3506.160 4318.450 ;
        RECT 3506.590 4318.170 3506.870 4318.450 ;
        RECT 3507.300 4318.170 3507.580 4318.450 ;
        RECT 3508.010 4318.170 3508.290 4318.450 ;
        RECT 3508.720 4318.170 3509.000 4318.450 ;
        RECT 3509.430 4318.170 3509.710 4318.450 ;
        RECT 3500.200 4317.460 3500.480 4317.740 ;
        RECT 3500.910 4317.460 3501.190 4317.740 ;
        RECT 3501.620 4317.460 3501.900 4317.740 ;
        RECT 3502.330 4317.460 3502.610 4317.740 ;
        RECT 3503.040 4317.460 3503.320 4317.740 ;
        RECT 3503.750 4317.460 3504.030 4317.740 ;
        RECT 3504.460 4317.460 3504.740 4317.740 ;
        RECT 3505.170 4317.460 3505.450 4317.740 ;
        RECT 3505.880 4317.460 3506.160 4317.740 ;
        RECT 3506.590 4317.460 3506.870 4317.740 ;
        RECT 3507.300 4317.460 3507.580 4317.740 ;
        RECT 3508.010 4317.460 3508.290 4317.740 ;
        RECT 3508.720 4317.460 3509.000 4317.740 ;
        RECT 3509.430 4317.460 3509.710 4317.740 ;
        RECT 3500.200 4316.750 3500.480 4317.030 ;
        RECT 3500.910 4316.750 3501.190 4317.030 ;
        RECT 3501.620 4316.750 3501.900 4317.030 ;
        RECT 3502.330 4316.750 3502.610 4317.030 ;
        RECT 3503.040 4316.750 3503.320 4317.030 ;
        RECT 3503.750 4316.750 3504.030 4317.030 ;
        RECT 3504.460 4316.750 3504.740 4317.030 ;
        RECT 3505.170 4316.750 3505.450 4317.030 ;
        RECT 3505.880 4316.750 3506.160 4317.030 ;
        RECT 3506.590 4316.750 3506.870 4317.030 ;
        RECT 3507.300 4316.750 3507.580 4317.030 ;
        RECT 3508.010 4316.750 3508.290 4317.030 ;
        RECT 3508.720 4316.750 3509.000 4317.030 ;
        RECT 3509.430 4316.750 3509.710 4317.030 ;
        RECT 369.330 4187.970 369.610 4188.250 ;
        RECT 370.040 4187.970 370.320 4188.250 ;
        RECT 370.750 4187.970 371.030 4188.250 ;
        RECT 371.460 4187.970 371.740 4188.250 ;
        RECT 372.170 4187.970 372.450 4188.250 ;
        RECT 372.880 4187.970 373.160 4188.250 ;
        RECT 373.590 4187.970 373.870 4188.250 ;
        RECT 374.300 4187.970 374.580 4188.250 ;
        RECT 375.010 4187.970 375.290 4188.250 ;
        RECT 375.720 4187.970 376.000 4188.250 ;
        RECT 376.430 4187.970 376.710 4188.250 ;
        RECT 369.330 4187.260 369.610 4187.540 ;
        RECT 370.040 4187.260 370.320 4187.540 ;
        RECT 370.750 4187.260 371.030 4187.540 ;
        RECT 371.460 4187.260 371.740 4187.540 ;
        RECT 372.170 4187.260 372.450 4187.540 ;
        RECT 372.880 4187.260 373.160 4187.540 ;
        RECT 373.590 4187.260 373.870 4187.540 ;
        RECT 374.300 4187.260 374.580 4187.540 ;
        RECT 375.010 4187.260 375.290 4187.540 ;
        RECT 375.720 4187.260 376.000 4187.540 ;
        RECT 376.430 4187.260 376.710 4187.540 ;
        RECT 369.330 4186.550 369.610 4186.830 ;
        RECT 370.040 4186.550 370.320 4186.830 ;
        RECT 370.750 4186.550 371.030 4186.830 ;
        RECT 371.460 4186.550 371.740 4186.830 ;
        RECT 372.170 4186.550 372.450 4186.830 ;
        RECT 372.880 4186.550 373.160 4186.830 ;
        RECT 373.590 4186.550 373.870 4186.830 ;
        RECT 374.300 4186.550 374.580 4186.830 ;
        RECT 375.010 4186.550 375.290 4186.830 ;
        RECT 375.720 4186.550 376.000 4186.830 ;
        RECT 376.430 4186.550 376.710 4186.830 ;
        RECT 369.330 4185.840 369.610 4186.120 ;
        RECT 370.040 4185.840 370.320 4186.120 ;
        RECT 370.750 4185.840 371.030 4186.120 ;
        RECT 371.460 4185.840 371.740 4186.120 ;
        RECT 372.170 4185.840 372.450 4186.120 ;
        RECT 372.880 4185.840 373.160 4186.120 ;
        RECT 373.590 4185.840 373.870 4186.120 ;
        RECT 374.300 4185.840 374.580 4186.120 ;
        RECT 375.010 4185.840 375.290 4186.120 ;
        RECT 375.720 4185.840 376.000 4186.120 ;
        RECT 376.430 4185.840 376.710 4186.120 ;
        RECT 369.330 4185.130 369.610 4185.410 ;
        RECT 370.040 4185.130 370.320 4185.410 ;
        RECT 370.750 4185.130 371.030 4185.410 ;
        RECT 371.460 4185.130 371.740 4185.410 ;
        RECT 372.170 4185.130 372.450 4185.410 ;
        RECT 372.880 4185.130 373.160 4185.410 ;
        RECT 373.590 4185.130 373.870 4185.410 ;
        RECT 374.300 4185.130 374.580 4185.410 ;
        RECT 375.010 4185.130 375.290 4185.410 ;
        RECT 375.720 4185.130 376.000 4185.410 ;
        RECT 376.430 4185.130 376.710 4185.410 ;
        RECT 369.330 4184.420 369.610 4184.700 ;
        RECT 370.040 4184.420 370.320 4184.700 ;
        RECT 370.750 4184.420 371.030 4184.700 ;
        RECT 371.460 4184.420 371.740 4184.700 ;
        RECT 372.170 4184.420 372.450 4184.700 ;
        RECT 372.880 4184.420 373.160 4184.700 ;
        RECT 373.590 4184.420 373.870 4184.700 ;
        RECT 374.300 4184.420 374.580 4184.700 ;
        RECT 375.010 4184.420 375.290 4184.700 ;
        RECT 375.720 4184.420 376.000 4184.700 ;
        RECT 376.430 4184.420 376.710 4184.700 ;
        RECT 369.330 4183.710 369.610 4183.990 ;
        RECT 370.040 4183.710 370.320 4183.990 ;
        RECT 370.750 4183.710 371.030 4183.990 ;
        RECT 371.460 4183.710 371.740 4183.990 ;
        RECT 372.170 4183.710 372.450 4183.990 ;
        RECT 372.880 4183.710 373.160 4183.990 ;
        RECT 373.590 4183.710 373.870 4183.990 ;
        RECT 374.300 4183.710 374.580 4183.990 ;
        RECT 375.010 4183.710 375.290 4183.990 ;
        RECT 375.720 4183.710 376.000 4183.990 ;
        RECT 376.430 4183.710 376.710 4183.990 ;
        RECT 369.330 4183.000 369.610 4183.280 ;
        RECT 370.040 4183.000 370.320 4183.280 ;
        RECT 370.750 4183.000 371.030 4183.280 ;
        RECT 371.460 4183.000 371.740 4183.280 ;
        RECT 372.170 4183.000 372.450 4183.280 ;
        RECT 372.880 4183.000 373.160 4183.280 ;
        RECT 373.590 4183.000 373.870 4183.280 ;
        RECT 374.300 4183.000 374.580 4183.280 ;
        RECT 375.010 4183.000 375.290 4183.280 ;
        RECT 375.720 4183.000 376.000 4183.280 ;
        RECT 376.430 4183.000 376.710 4183.280 ;
        RECT 369.330 4182.290 369.610 4182.570 ;
        RECT 370.040 4182.290 370.320 4182.570 ;
        RECT 370.750 4182.290 371.030 4182.570 ;
        RECT 371.460 4182.290 371.740 4182.570 ;
        RECT 372.170 4182.290 372.450 4182.570 ;
        RECT 372.880 4182.290 373.160 4182.570 ;
        RECT 373.590 4182.290 373.870 4182.570 ;
        RECT 374.300 4182.290 374.580 4182.570 ;
        RECT 375.010 4182.290 375.290 4182.570 ;
        RECT 375.720 4182.290 376.000 4182.570 ;
        RECT 376.430 4182.290 376.710 4182.570 ;
        RECT 369.330 4181.580 369.610 4181.860 ;
        RECT 370.040 4181.580 370.320 4181.860 ;
        RECT 370.750 4181.580 371.030 4181.860 ;
        RECT 371.460 4181.580 371.740 4181.860 ;
        RECT 372.170 4181.580 372.450 4181.860 ;
        RECT 372.880 4181.580 373.160 4181.860 ;
        RECT 373.590 4181.580 373.870 4181.860 ;
        RECT 374.300 4181.580 374.580 4181.860 ;
        RECT 375.010 4181.580 375.290 4181.860 ;
        RECT 375.720 4181.580 376.000 4181.860 ;
        RECT 376.430 4181.580 376.710 4181.860 ;
        RECT 369.330 4180.870 369.610 4181.150 ;
        RECT 370.040 4180.870 370.320 4181.150 ;
        RECT 370.750 4180.870 371.030 4181.150 ;
        RECT 371.460 4180.870 371.740 4181.150 ;
        RECT 372.170 4180.870 372.450 4181.150 ;
        RECT 372.880 4180.870 373.160 4181.150 ;
        RECT 373.590 4180.870 373.870 4181.150 ;
        RECT 374.300 4180.870 374.580 4181.150 ;
        RECT 375.010 4180.870 375.290 4181.150 ;
        RECT 375.720 4180.870 376.000 4181.150 ;
        RECT 376.430 4180.870 376.710 4181.150 ;
        RECT 369.330 4180.160 369.610 4180.440 ;
        RECT 370.040 4180.160 370.320 4180.440 ;
        RECT 370.750 4180.160 371.030 4180.440 ;
        RECT 371.460 4180.160 371.740 4180.440 ;
        RECT 372.170 4180.160 372.450 4180.440 ;
        RECT 372.880 4180.160 373.160 4180.440 ;
        RECT 373.590 4180.160 373.870 4180.440 ;
        RECT 374.300 4180.160 374.580 4180.440 ;
        RECT 375.010 4180.160 375.290 4180.440 ;
        RECT 375.720 4180.160 376.000 4180.440 ;
        RECT 376.430 4180.160 376.710 4180.440 ;
        RECT 369.330 4179.450 369.610 4179.730 ;
        RECT 370.040 4179.450 370.320 4179.730 ;
        RECT 370.750 4179.450 371.030 4179.730 ;
        RECT 371.460 4179.450 371.740 4179.730 ;
        RECT 372.170 4179.450 372.450 4179.730 ;
        RECT 372.880 4179.450 373.160 4179.730 ;
        RECT 373.590 4179.450 373.870 4179.730 ;
        RECT 374.300 4179.450 374.580 4179.730 ;
        RECT 375.010 4179.450 375.290 4179.730 ;
        RECT 375.720 4179.450 376.000 4179.730 ;
        RECT 376.430 4179.450 376.710 4179.730 ;
        RECT 369.275 4175.565 369.555 4175.845 ;
        RECT 369.985 4175.565 370.265 4175.845 ;
        RECT 370.695 4175.565 370.975 4175.845 ;
        RECT 371.405 4175.565 371.685 4175.845 ;
        RECT 372.115 4175.565 372.395 4175.845 ;
        RECT 372.825 4175.565 373.105 4175.845 ;
        RECT 373.535 4175.565 373.815 4175.845 ;
        RECT 374.245 4175.565 374.525 4175.845 ;
        RECT 374.955 4175.565 375.235 4175.845 ;
        RECT 375.665 4175.565 375.945 4175.845 ;
        RECT 376.375 4175.565 376.655 4175.845 ;
        RECT 369.275 4174.855 369.555 4175.135 ;
        RECT 369.985 4174.855 370.265 4175.135 ;
        RECT 370.695 4174.855 370.975 4175.135 ;
        RECT 371.405 4174.855 371.685 4175.135 ;
        RECT 372.115 4174.855 372.395 4175.135 ;
        RECT 372.825 4174.855 373.105 4175.135 ;
        RECT 373.535 4174.855 373.815 4175.135 ;
        RECT 374.245 4174.855 374.525 4175.135 ;
        RECT 374.955 4174.855 375.235 4175.135 ;
        RECT 375.665 4174.855 375.945 4175.135 ;
        RECT 376.375 4174.855 376.655 4175.135 ;
        RECT 369.275 4174.145 369.555 4174.425 ;
        RECT 369.985 4174.145 370.265 4174.425 ;
        RECT 370.695 4174.145 370.975 4174.425 ;
        RECT 371.405 4174.145 371.685 4174.425 ;
        RECT 372.115 4174.145 372.395 4174.425 ;
        RECT 372.825 4174.145 373.105 4174.425 ;
        RECT 373.535 4174.145 373.815 4174.425 ;
        RECT 374.245 4174.145 374.525 4174.425 ;
        RECT 374.955 4174.145 375.235 4174.425 ;
        RECT 375.665 4174.145 375.945 4174.425 ;
        RECT 376.375 4174.145 376.655 4174.425 ;
        RECT 369.275 4173.435 369.555 4173.715 ;
        RECT 369.985 4173.435 370.265 4173.715 ;
        RECT 370.695 4173.435 370.975 4173.715 ;
        RECT 371.405 4173.435 371.685 4173.715 ;
        RECT 372.115 4173.435 372.395 4173.715 ;
        RECT 372.825 4173.435 373.105 4173.715 ;
        RECT 373.535 4173.435 373.815 4173.715 ;
        RECT 374.245 4173.435 374.525 4173.715 ;
        RECT 374.955 4173.435 375.235 4173.715 ;
        RECT 375.665 4173.435 375.945 4173.715 ;
        RECT 376.375 4173.435 376.655 4173.715 ;
        RECT 369.275 4172.725 369.555 4173.005 ;
        RECT 369.985 4172.725 370.265 4173.005 ;
        RECT 370.695 4172.725 370.975 4173.005 ;
        RECT 371.405 4172.725 371.685 4173.005 ;
        RECT 372.115 4172.725 372.395 4173.005 ;
        RECT 372.825 4172.725 373.105 4173.005 ;
        RECT 373.535 4172.725 373.815 4173.005 ;
        RECT 374.245 4172.725 374.525 4173.005 ;
        RECT 374.955 4172.725 375.235 4173.005 ;
        RECT 375.665 4172.725 375.945 4173.005 ;
        RECT 376.375 4172.725 376.655 4173.005 ;
        RECT 369.275 4172.015 369.555 4172.295 ;
        RECT 369.985 4172.015 370.265 4172.295 ;
        RECT 370.695 4172.015 370.975 4172.295 ;
        RECT 371.405 4172.015 371.685 4172.295 ;
        RECT 372.115 4172.015 372.395 4172.295 ;
        RECT 372.825 4172.015 373.105 4172.295 ;
        RECT 373.535 4172.015 373.815 4172.295 ;
        RECT 374.245 4172.015 374.525 4172.295 ;
        RECT 374.955 4172.015 375.235 4172.295 ;
        RECT 375.665 4172.015 375.945 4172.295 ;
        RECT 376.375 4172.015 376.655 4172.295 ;
        RECT 369.275 4171.305 369.555 4171.585 ;
        RECT 369.985 4171.305 370.265 4171.585 ;
        RECT 370.695 4171.305 370.975 4171.585 ;
        RECT 371.405 4171.305 371.685 4171.585 ;
        RECT 372.115 4171.305 372.395 4171.585 ;
        RECT 372.825 4171.305 373.105 4171.585 ;
        RECT 373.535 4171.305 373.815 4171.585 ;
        RECT 374.245 4171.305 374.525 4171.585 ;
        RECT 374.955 4171.305 375.235 4171.585 ;
        RECT 375.665 4171.305 375.945 4171.585 ;
        RECT 376.375 4171.305 376.655 4171.585 ;
        RECT 369.275 4170.595 369.555 4170.875 ;
        RECT 369.985 4170.595 370.265 4170.875 ;
        RECT 370.695 4170.595 370.975 4170.875 ;
        RECT 371.405 4170.595 371.685 4170.875 ;
        RECT 372.115 4170.595 372.395 4170.875 ;
        RECT 372.825 4170.595 373.105 4170.875 ;
        RECT 373.535 4170.595 373.815 4170.875 ;
        RECT 374.245 4170.595 374.525 4170.875 ;
        RECT 374.955 4170.595 375.235 4170.875 ;
        RECT 375.665 4170.595 375.945 4170.875 ;
        RECT 376.375 4170.595 376.655 4170.875 ;
        RECT 369.275 4169.885 369.555 4170.165 ;
        RECT 369.985 4169.885 370.265 4170.165 ;
        RECT 370.695 4169.885 370.975 4170.165 ;
        RECT 371.405 4169.885 371.685 4170.165 ;
        RECT 372.115 4169.885 372.395 4170.165 ;
        RECT 372.825 4169.885 373.105 4170.165 ;
        RECT 373.535 4169.885 373.815 4170.165 ;
        RECT 374.245 4169.885 374.525 4170.165 ;
        RECT 374.955 4169.885 375.235 4170.165 ;
        RECT 375.665 4169.885 375.945 4170.165 ;
        RECT 376.375 4169.885 376.655 4170.165 ;
        RECT 369.275 4169.175 369.555 4169.455 ;
        RECT 369.985 4169.175 370.265 4169.455 ;
        RECT 370.695 4169.175 370.975 4169.455 ;
        RECT 371.405 4169.175 371.685 4169.455 ;
        RECT 372.115 4169.175 372.395 4169.455 ;
        RECT 372.825 4169.175 373.105 4169.455 ;
        RECT 373.535 4169.175 373.815 4169.455 ;
        RECT 374.245 4169.175 374.525 4169.455 ;
        RECT 374.955 4169.175 375.235 4169.455 ;
        RECT 375.665 4169.175 375.945 4169.455 ;
        RECT 376.375 4169.175 376.655 4169.455 ;
        RECT 369.275 4168.465 369.555 4168.745 ;
        RECT 369.985 4168.465 370.265 4168.745 ;
        RECT 370.695 4168.465 370.975 4168.745 ;
        RECT 371.405 4168.465 371.685 4168.745 ;
        RECT 372.115 4168.465 372.395 4168.745 ;
        RECT 372.825 4168.465 373.105 4168.745 ;
        RECT 373.535 4168.465 373.815 4168.745 ;
        RECT 374.245 4168.465 374.525 4168.745 ;
        RECT 374.955 4168.465 375.235 4168.745 ;
        RECT 375.665 4168.465 375.945 4168.745 ;
        RECT 376.375 4168.465 376.655 4168.745 ;
        RECT 369.275 4167.755 369.555 4168.035 ;
        RECT 369.985 4167.755 370.265 4168.035 ;
        RECT 370.695 4167.755 370.975 4168.035 ;
        RECT 371.405 4167.755 371.685 4168.035 ;
        RECT 372.115 4167.755 372.395 4168.035 ;
        RECT 372.825 4167.755 373.105 4168.035 ;
        RECT 373.535 4167.755 373.815 4168.035 ;
        RECT 374.245 4167.755 374.525 4168.035 ;
        RECT 374.955 4167.755 375.235 4168.035 ;
        RECT 375.665 4167.755 375.945 4168.035 ;
        RECT 376.375 4167.755 376.655 4168.035 ;
        RECT 369.275 4167.045 369.555 4167.325 ;
        RECT 369.985 4167.045 370.265 4167.325 ;
        RECT 370.695 4167.045 370.975 4167.325 ;
        RECT 371.405 4167.045 371.685 4167.325 ;
        RECT 372.115 4167.045 372.395 4167.325 ;
        RECT 372.825 4167.045 373.105 4167.325 ;
        RECT 373.535 4167.045 373.815 4167.325 ;
        RECT 374.245 4167.045 374.525 4167.325 ;
        RECT 374.955 4167.045 375.235 4167.325 ;
        RECT 375.665 4167.045 375.945 4167.325 ;
        RECT 376.375 4167.045 376.655 4167.325 ;
        RECT 369.275 4166.335 369.555 4166.615 ;
        RECT 369.985 4166.335 370.265 4166.615 ;
        RECT 370.695 4166.335 370.975 4166.615 ;
        RECT 371.405 4166.335 371.685 4166.615 ;
        RECT 372.115 4166.335 372.395 4166.615 ;
        RECT 372.825 4166.335 373.105 4166.615 ;
        RECT 373.535 4166.335 373.815 4166.615 ;
        RECT 374.245 4166.335 374.525 4166.615 ;
        RECT 374.955 4166.335 375.235 4166.615 ;
        RECT 375.665 4166.335 375.945 4166.615 ;
        RECT 376.375 4166.335 376.655 4166.615 ;
        RECT 369.275 4163.715 369.555 4163.995 ;
        RECT 369.985 4163.715 370.265 4163.995 ;
        RECT 370.695 4163.715 370.975 4163.995 ;
        RECT 371.405 4163.715 371.685 4163.995 ;
        RECT 372.115 4163.715 372.395 4163.995 ;
        RECT 372.825 4163.715 373.105 4163.995 ;
        RECT 373.535 4163.715 373.815 4163.995 ;
        RECT 374.245 4163.715 374.525 4163.995 ;
        RECT 374.955 4163.715 375.235 4163.995 ;
        RECT 375.665 4163.715 375.945 4163.995 ;
        RECT 376.375 4163.715 376.655 4163.995 ;
        RECT 369.275 4163.005 369.555 4163.285 ;
        RECT 369.985 4163.005 370.265 4163.285 ;
        RECT 370.695 4163.005 370.975 4163.285 ;
        RECT 371.405 4163.005 371.685 4163.285 ;
        RECT 372.115 4163.005 372.395 4163.285 ;
        RECT 372.825 4163.005 373.105 4163.285 ;
        RECT 373.535 4163.005 373.815 4163.285 ;
        RECT 374.245 4163.005 374.525 4163.285 ;
        RECT 374.955 4163.005 375.235 4163.285 ;
        RECT 375.665 4163.005 375.945 4163.285 ;
        RECT 376.375 4163.005 376.655 4163.285 ;
        RECT 369.275 4162.295 369.555 4162.575 ;
        RECT 369.985 4162.295 370.265 4162.575 ;
        RECT 370.695 4162.295 370.975 4162.575 ;
        RECT 371.405 4162.295 371.685 4162.575 ;
        RECT 372.115 4162.295 372.395 4162.575 ;
        RECT 372.825 4162.295 373.105 4162.575 ;
        RECT 373.535 4162.295 373.815 4162.575 ;
        RECT 374.245 4162.295 374.525 4162.575 ;
        RECT 374.955 4162.295 375.235 4162.575 ;
        RECT 375.665 4162.295 375.945 4162.575 ;
        RECT 376.375 4162.295 376.655 4162.575 ;
        RECT 369.275 4161.585 369.555 4161.865 ;
        RECT 369.985 4161.585 370.265 4161.865 ;
        RECT 370.695 4161.585 370.975 4161.865 ;
        RECT 371.405 4161.585 371.685 4161.865 ;
        RECT 372.115 4161.585 372.395 4161.865 ;
        RECT 372.825 4161.585 373.105 4161.865 ;
        RECT 373.535 4161.585 373.815 4161.865 ;
        RECT 374.245 4161.585 374.525 4161.865 ;
        RECT 374.955 4161.585 375.235 4161.865 ;
        RECT 375.665 4161.585 375.945 4161.865 ;
        RECT 376.375 4161.585 376.655 4161.865 ;
        RECT 369.275 4160.875 369.555 4161.155 ;
        RECT 369.985 4160.875 370.265 4161.155 ;
        RECT 370.695 4160.875 370.975 4161.155 ;
        RECT 371.405 4160.875 371.685 4161.155 ;
        RECT 372.115 4160.875 372.395 4161.155 ;
        RECT 372.825 4160.875 373.105 4161.155 ;
        RECT 373.535 4160.875 373.815 4161.155 ;
        RECT 374.245 4160.875 374.525 4161.155 ;
        RECT 374.955 4160.875 375.235 4161.155 ;
        RECT 375.665 4160.875 375.945 4161.155 ;
        RECT 376.375 4160.875 376.655 4161.155 ;
        RECT 369.275 4160.165 369.555 4160.445 ;
        RECT 369.985 4160.165 370.265 4160.445 ;
        RECT 370.695 4160.165 370.975 4160.445 ;
        RECT 371.405 4160.165 371.685 4160.445 ;
        RECT 372.115 4160.165 372.395 4160.445 ;
        RECT 372.825 4160.165 373.105 4160.445 ;
        RECT 373.535 4160.165 373.815 4160.445 ;
        RECT 374.245 4160.165 374.525 4160.445 ;
        RECT 374.955 4160.165 375.235 4160.445 ;
        RECT 375.665 4160.165 375.945 4160.445 ;
        RECT 376.375 4160.165 376.655 4160.445 ;
        RECT 369.275 4159.455 369.555 4159.735 ;
        RECT 369.985 4159.455 370.265 4159.735 ;
        RECT 370.695 4159.455 370.975 4159.735 ;
        RECT 371.405 4159.455 371.685 4159.735 ;
        RECT 372.115 4159.455 372.395 4159.735 ;
        RECT 372.825 4159.455 373.105 4159.735 ;
        RECT 373.535 4159.455 373.815 4159.735 ;
        RECT 374.245 4159.455 374.525 4159.735 ;
        RECT 374.955 4159.455 375.235 4159.735 ;
        RECT 375.665 4159.455 375.945 4159.735 ;
        RECT 376.375 4159.455 376.655 4159.735 ;
        RECT 369.275 4158.745 369.555 4159.025 ;
        RECT 369.985 4158.745 370.265 4159.025 ;
        RECT 370.695 4158.745 370.975 4159.025 ;
        RECT 371.405 4158.745 371.685 4159.025 ;
        RECT 372.115 4158.745 372.395 4159.025 ;
        RECT 372.825 4158.745 373.105 4159.025 ;
        RECT 373.535 4158.745 373.815 4159.025 ;
        RECT 374.245 4158.745 374.525 4159.025 ;
        RECT 374.955 4158.745 375.235 4159.025 ;
        RECT 375.665 4158.745 375.945 4159.025 ;
        RECT 376.375 4158.745 376.655 4159.025 ;
        RECT 369.275 4158.035 369.555 4158.315 ;
        RECT 369.985 4158.035 370.265 4158.315 ;
        RECT 370.695 4158.035 370.975 4158.315 ;
        RECT 371.405 4158.035 371.685 4158.315 ;
        RECT 372.115 4158.035 372.395 4158.315 ;
        RECT 372.825 4158.035 373.105 4158.315 ;
        RECT 373.535 4158.035 373.815 4158.315 ;
        RECT 374.245 4158.035 374.525 4158.315 ;
        RECT 374.955 4158.035 375.235 4158.315 ;
        RECT 375.665 4158.035 375.945 4158.315 ;
        RECT 376.375 4158.035 376.655 4158.315 ;
        RECT 369.275 4157.325 369.555 4157.605 ;
        RECT 369.985 4157.325 370.265 4157.605 ;
        RECT 370.695 4157.325 370.975 4157.605 ;
        RECT 371.405 4157.325 371.685 4157.605 ;
        RECT 372.115 4157.325 372.395 4157.605 ;
        RECT 372.825 4157.325 373.105 4157.605 ;
        RECT 373.535 4157.325 373.815 4157.605 ;
        RECT 374.245 4157.325 374.525 4157.605 ;
        RECT 374.955 4157.325 375.235 4157.605 ;
        RECT 375.665 4157.325 375.945 4157.605 ;
        RECT 376.375 4157.325 376.655 4157.605 ;
        RECT 369.275 4156.615 369.555 4156.895 ;
        RECT 369.985 4156.615 370.265 4156.895 ;
        RECT 370.695 4156.615 370.975 4156.895 ;
        RECT 371.405 4156.615 371.685 4156.895 ;
        RECT 372.115 4156.615 372.395 4156.895 ;
        RECT 372.825 4156.615 373.105 4156.895 ;
        RECT 373.535 4156.615 373.815 4156.895 ;
        RECT 374.245 4156.615 374.525 4156.895 ;
        RECT 374.955 4156.615 375.235 4156.895 ;
        RECT 375.665 4156.615 375.945 4156.895 ;
        RECT 376.375 4156.615 376.655 4156.895 ;
        RECT 369.275 4155.905 369.555 4156.185 ;
        RECT 369.985 4155.905 370.265 4156.185 ;
        RECT 370.695 4155.905 370.975 4156.185 ;
        RECT 371.405 4155.905 371.685 4156.185 ;
        RECT 372.115 4155.905 372.395 4156.185 ;
        RECT 372.825 4155.905 373.105 4156.185 ;
        RECT 373.535 4155.905 373.815 4156.185 ;
        RECT 374.245 4155.905 374.525 4156.185 ;
        RECT 374.955 4155.905 375.235 4156.185 ;
        RECT 375.665 4155.905 375.945 4156.185 ;
        RECT 376.375 4155.905 376.655 4156.185 ;
        RECT 369.275 4155.195 369.555 4155.475 ;
        RECT 369.985 4155.195 370.265 4155.475 ;
        RECT 370.695 4155.195 370.975 4155.475 ;
        RECT 371.405 4155.195 371.685 4155.475 ;
        RECT 372.115 4155.195 372.395 4155.475 ;
        RECT 372.825 4155.195 373.105 4155.475 ;
        RECT 373.535 4155.195 373.815 4155.475 ;
        RECT 374.245 4155.195 374.525 4155.475 ;
        RECT 374.955 4155.195 375.235 4155.475 ;
        RECT 375.665 4155.195 375.945 4155.475 ;
        RECT 376.375 4155.195 376.655 4155.475 ;
        RECT 369.275 4154.485 369.555 4154.765 ;
        RECT 369.985 4154.485 370.265 4154.765 ;
        RECT 370.695 4154.485 370.975 4154.765 ;
        RECT 371.405 4154.485 371.685 4154.765 ;
        RECT 372.115 4154.485 372.395 4154.765 ;
        RECT 372.825 4154.485 373.105 4154.765 ;
        RECT 373.535 4154.485 373.815 4154.765 ;
        RECT 374.245 4154.485 374.525 4154.765 ;
        RECT 374.955 4154.485 375.235 4154.765 ;
        RECT 375.665 4154.485 375.945 4154.765 ;
        RECT 376.375 4154.485 376.655 4154.765 ;
        RECT 369.275 4150.185 369.555 4150.465 ;
        RECT 369.985 4150.185 370.265 4150.465 ;
        RECT 370.695 4150.185 370.975 4150.465 ;
        RECT 371.405 4150.185 371.685 4150.465 ;
        RECT 372.115 4150.185 372.395 4150.465 ;
        RECT 372.825 4150.185 373.105 4150.465 ;
        RECT 373.535 4150.185 373.815 4150.465 ;
        RECT 374.245 4150.185 374.525 4150.465 ;
        RECT 374.955 4150.185 375.235 4150.465 ;
        RECT 375.665 4150.185 375.945 4150.465 ;
        RECT 376.375 4150.185 376.655 4150.465 ;
        RECT 369.275 4149.475 369.555 4149.755 ;
        RECT 369.985 4149.475 370.265 4149.755 ;
        RECT 370.695 4149.475 370.975 4149.755 ;
        RECT 371.405 4149.475 371.685 4149.755 ;
        RECT 372.115 4149.475 372.395 4149.755 ;
        RECT 372.825 4149.475 373.105 4149.755 ;
        RECT 373.535 4149.475 373.815 4149.755 ;
        RECT 374.245 4149.475 374.525 4149.755 ;
        RECT 374.955 4149.475 375.235 4149.755 ;
        RECT 375.665 4149.475 375.945 4149.755 ;
        RECT 376.375 4149.475 376.655 4149.755 ;
        RECT 369.275 4148.765 369.555 4149.045 ;
        RECT 369.985 4148.765 370.265 4149.045 ;
        RECT 370.695 4148.765 370.975 4149.045 ;
        RECT 371.405 4148.765 371.685 4149.045 ;
        RECT 372.115 4148.765 372.395 4149.045 ;
        RECT 372.825 4148.765 373.105 4149.045 ;
        RECT 373.535 4148.765 373.815 4149.045 ;
        RECT 374.245 4148.765 374.525 4149.045 ;
        RECT 374.955 4148.765 375.235 4149.045 ;
        RECT 375.665 4148.765 375.945 4149.045 ;
        RECT 376.375 4148.765 376.655 4149.045 ;
        RECT 369.275 4148.055 369.555 4148.335 ;
        RECT 369.985 4148.055 370.265 4148.335 ;
        RECT 370.695 4148.055 370.975 4148.335 ;
        RECT 371.405 4148.055 371.685 4148.335 ;
        RECT 372.115 4148.055 372.395 4148.335 ;
        RECT 372.825 4148.055 373.105 4148.335 ;
        RECT 373.535 4148.055 373.815 4148.335 ;
        RECT 374.245 4148.055 374.525 4148.335 ;
        RECT 374.955 4148.055 375.235 4148.335 ;
        RECT 375.665 4148.055 375.945 4148.335 ;
        RECT 376.375 4148.055 376.655 4148.335 ;
        RECT 369.275 4147.345 369.555 4147.625 ;
        RECT 369.985 4147.345 370.265 4147.625 ;
        RECT 370.695 4147.345 370.975 4147.625 ;
        RECT 371.405 4147.345 371.685 4147.625 ;
        RECT 372.115 4147.345 372.395 4147.625 ;
        RECT 372.825 4147.345 373.105 4147.625 ;
        RECT 373.535 4147.345 373.815 4147.625 ;
        RECT 374.245 4147.345 374.525 4147.625 ;
        RECT 374.955 4147.345 375.235 4147.625 ;
        RECT 375.665 4147.345 375.945 4147.625 ;
        RECT 376.375 4147.345 376.655 4147.625 ;
        RECT 369.275 4146.635 369.555 4146.915 ;
        RECT 369.985 4146.635 370.265 4146.915 ;
        RECT 370.695 4146.635 370.975 4146.915 ;
        RECT 371.405 4146.635 371.685 4146.915 ;
        RECT 372.115 4146.635 372.395 4146.915 ;
        RECT 372.825 4146.635 373.105 4146.915 ;
        RECT 373.535 4146.635 373.815 4146.915 ;
        RECT 374.245 4146.635 374.525 4146.915 ;
        RECT 374.955 4146.635 375.235 4146.915 ;
        RECT 375.665 4146.635 375.945 4146.915 ;
        RECT 376.375 4146.635 376.655 4146.915 ;
        RECT 369.275 4145.925 369.555 4146.205 ;
        RECT 369.985 4145.925 370.265 4146.205 ;
        RECT 370.695 4145.925 370.975 4146.205 ;
        RECT 371.405 4145.925 371.685 4146.205 ;
        RECT 372.115 4145.925 372.395 4146.205 ;
        RECT 372.825 4145.925 373.105 4146.205 ;
        RECT 373.535 4145.925 373.815 4146.205 ;
        RECT 374.245 4145.925 374.525 4146.205 ;
        RECT 374.955 4145.925 375.235 4146.205 ;
        RECT 375.665 4145.925 375.945 4146.205 ;
        RECT 376.375 4145.925 376.655 4146.205 ;
        RECT 369.275 4145.215 369.555 4145.495 ;
        RECT 369.985 4145.215 370.265 4145.495 ;
        RECT 370.695 4145.215 370.975 4145.495 ;
        RECT 371.405 4145.215 371.685 4145.495 ;
        RECT 372.115 4145.215 372.395 4145.495 ;
        RECT 372.825 4145.215 373.105 4145.495 ;
        RECT 373.535 4145.215 373.815 4145.495 ;
        RECT 374.245 4145.215 374.525 4145.495 ;
        RECT 374.955 4145.215 375.235 4145.495 ;
        RECT 375.665 4145.215 375.945 4145.495 ;
        RECT 376.375 4145.215 376.655 4145.495 ;
        RECT 369.275 4144.505 369.555 4144.785 ;
        RECT 369.985 4144.505 370.265 4144.785 ;
        RECT 370.695 4144.505 370.975 4144.785 ;
        RECT 371.405 4144.505 371.685 4144.785 ;
        RECT 372.115 4144.505 372.395 4144.785 ;
        RECT 372.825 4144.505 373.105 4144.785 ;
        RECT 373.535 4144.505 373.815 4144.785 ;
        RECT 374.245 4144.505 374.525 4144.785 ;
        RECT 374.955 4144.505 375.235 4144.785 ;
        RECT 375.665 4144.505 375.945 4144.785 ;
        RECT 376.375 4144.505 376.655 4144.785 ;
        RECT 369.275 4143.795 369.555 4144.075 ;
        RECT 369.985 4143.795 370.265 4144.075 ;
        RECT 370.695 4143.795 370.975 4144.075 ;
        RECT 371.405 4143.795 371.685 4144.075 ;
        RECT 372.115 4143.795 372.395 4144.075 ;
        RECT 372.825 4143.795 373.105 4144.075 ;
        RECT 373.535 4143.795 373.815 4144.075 ;
        RECT 374.245 4143.795 374.525 4144.075 ;
        RECT 374.955 4143.795 375.235 4144.075 ;
        RECT 375.665 4143.795 375.945 4144.075 ;
        RECT 376.375 4143.795 376.655 4144.075 ;
        RECT 369.275 4143.085 369.555 4143.365 ;
        RECT 369.985 4143.085 370.265 4143.365 ;
        RECT 370.695 4143.085 370.975 4143.365 ;
        RECT 371.405 4143.085 371.685 4143.365 ;
        RECT 372.115 4143.085 372.395 4143.365 ;
        RECT 372.825 4143.085 373.105 4143.365 ;
        RECT 373.535 4143.085 373.815 4143.365 ;
        RECT 374.245 4143.085 374.525 4143.365 ;
        RECT 374.955 4143.085 375.235 4143.365 ;
        RECT 375.665 4143.085 375.945 4143.365 ;
        RECT 376.375 4143.085 376.655 4143.365 ;
        RECT 369.275 4142.375 369.555 4142.655 ;
        RECT 369.985 4142.375 370.265 4142.655 ;
        RECT 370.695 4142.375 370.975 4142.655 ;
        RECT 371.405 4142.375 371.685 4142.655 ;
        RECT 372.115 4142.375 372.395 4142.655 ;
        RECT 372.825 4142.375 373.105 4142.655 ;
        RECT 373.535 4142.375 373.815 4142.655 ;
        RECT 374.245 4142.375 374.525 4142.655 ;
        RECT 374.955 4142.375 375.235 4142.655 ;
        RECT 375.665 4142.375 375.945 4142.655 ;
        RECT 376.375 4142.375 376.655 4142.655 ;
        RECT 369.275 4141.665 369.555 4141.945 ;
        RECT 369.985 4141.665 370.265 4141.945 ;
        RECT 370.695 4141.665 370.975 4141.945 ;
        RECT 371.405 4141.665 371.685 4141.945 ;
        RECT 372.115 4141.665 372.395 4141.945 ;
        RECT 372.825 4141.665 373.105 4141.945 ;
        RECT 373.535 4141.665 373.815 4141.945 ;
        RECT 374.245 4141.665 374.525 4141.945 ;
        RECT 374.955 4141.665 375.235 4141.945 ;
        RECT 375.665 4141.665 375.945 4141.945 ;
        RECT 376.375 4141.665 376.655 4141.945 ;
        RECT 369.275 4140.955 369.555 4141.235 ;
        RECT 369.985 4140.955 370.265 4141.235 ;
        RECT 370.695 4140.955 370.975 4141.235 ;
        RECT 371.405 4140.955 371.685 4141.235 ;
        RECT 372.115 4140.955 372.395 4141.235 ;
        RECT 372.825 4140.955 373.105 4141.235 ;
        RECT 373.535 4140.955 373.815 4141.235 ;
        RECT 374.245 4140.955 374.525 4141.235 ;
        RECT 374.955 4140.955 375.235 4141.235 ;
        RECT 375.665 4140.955 375.945 4141.235 ;
        RECT 376.375 4140.955 376.655 4141.235 ;
        RECT 369.275 4138.335 369.555 4138.615 ;
        RECT 369.985 4138.335 370.265 4138.615 ;
        RECT 370.695 4138.335 370.975 4138.615 ;
        RECT 371.405 4138.335 371.685 4138.615 ;
        RECT 372.115 4138.335 372.395 4138.615 ;
        RECT 372.825 4138.335 373.105 4138.615 ;
        RECT 373.535 4138.335 373.815 4138.615 ;
        RECT 374.245 4138.335 374.525 4138.615 ;
        RECT 374.955 4138.335 375.235 4138.615 ;
        RECT 375.665 4138.335 375.945 4138.615 ;
        RECT 376.375 4138.335 376.655 4138.615 ;
        RECT 369.275 4137.625 369.555 4137.905 ;
        RECT 369.985 4137.625 370.265 4137.905 ;
        RECT 370.695 4137.625 370.975 4137.905 ;
        RECT 371.405 4137.625 371.685 4137.905 ;
        RECT 372.115 4137.625 372.395 4137.905 ;
        RECT 372.825 4137.625 373.105 4137.905 ;
        RECT 373.535 4137.625 373.815 4137.905 ;
        RECT 374.245 4137.625 374.525 4137.905 ;
        RECT 374.955 4137.625 375.235 4137.905 ;
        RECT 375.665 4137.625 375.945 4137.905 ;
        RECT 376.375 4137.625 376.655 4137.905 ;
        RECT 369.275 4136.915 369.555 4137.195 ;
        RECT 369.985 4136.915 370.265 4137.195 ;
        RECT 370.695 4136.915 370.975 4137.195 ;
        RECT 371.405 4136.915 371.685 4137.195 ;
        RECT 372.115 4136.915 372.395 4137.195 ;
        RECT 372.825 4136.915 373.105 4137.195 ;
        RECT 373.535 4136.915 373.815 4137.195 ;
        RECT 374.245 4136.915 374.525 4137.195 ;
        RECT 374.955 4136.915 375.235 4137.195 ;
        RECT 375.665 4136.915 375.945 4137.195 ;
        RECT 376.375 4136.915 376.655 4137.195 ;
        RECT 369.275 4136.205 369.555 4136.485 ;
        RECT 369.985 4136.205 370.265 4136.485 ;
        RECT 370.695 4136.205 370.975 4136.485 ;
        RECT 371.405 4136.205 371.685 4136.485 ;
        RECT 372.115 4136.205 372.395 4136.485 ;
        RECT 372.825 4136.205 373.105 4136.485 ;
        RECT 373.535 4136.205 373.815 4136.485 ;
        RECT 374.245 4136.205 374.525 4136.485 ;
        RECT 374.955 4136.205 375.235 4136.485 ;
        RECT 375.665 4136.205 375.945 4136.485 ;
        RECT 376.375 4136.205 376.655 4136.485 ;
        RECT 369.275 4135.495 369.555 4135.775 ;
        RECT 369.985 4135.495 370.265 4135.775 ;
        RECT 370.695 4135.495 370.975 4135.775 ;
        RECT 371.405 4135.495 371.685 4135.775 ;
        RECT 372.115 4135.495 372.395 4135.775 ;
        RECT 372.825 4135.495 373.105 4135.775 ;
        RECT 373.535 4135.495 373.815 4135.775 ;
        RECT 374.245 4135.495 374.525 4135.775 ;
        RECT 374.955 4135.495 375.235 4135.775 ;
        RECT 375.665 4135.495 375.945 4135.775 ;
        RECT 376.375 4135.495 376.655 4135.775 ;
        RECT 369.275 4134.785 369.555 4135.065 ;
        RECT 369.985 4134.785 370.265 4135.065 ;
        RECT 370.695 4134.785 370.975 4135.065 ;
        RECT 371.405 4134.785 371.685 4135.065 ;
        RECT 372.115 4134.785 372.395 4135.065 ;
        RECT 372.825 4134.785 373.105 4135.065 ;
        RECT 373.535 4134.785 373.815 4135.065 ;
        RECT 374.245 4134.785 374.525 4135.065 ;
        RECT 374.955 4134.785 375.235 4135.065 ;
        RECT 375.665 4134.785 375.945 4135.065 ;
        RECT 376.375 4134.785 376.655 4135.065 ;
        RECT 369.275 4134.075 369.555 4134.355 ;
        RECT 369.985 4134.075 370.265 4134.355 ;
        RECT 370.695 4134.075 370.975 4134.355 ;
        RECT 371.405 4134.075 371.685 4134.355 ;
        RECT 372.115 4134.075 372.395 4134.355 ;
        RECT 372.825 4134.075 373.105 4134.355 ;
        RECT 373.535 4134.075 373.815 4134.355 ;
        RECT 374.245 4134.075 374.525 4134.355 ;
        RECT 374.955 4134.075 375.235 4134.355 ;
        RECT 375.665 4134.075 375.945 4134.355 ;
        RECT 376.375 4134.075 376.655 4134.355 ;
        RECT 369.275 4133.365 369.555 4133.645 ;
        RECT 369.985 4133.365 370.265 4133.645 ;
        RECT 370.695 4133.365 370.975 4133.645 ;
        RECT 371.405 4133.365 371.685 4133.645 ;
        RECT 372.115 4133.365 372.395 4133.645 ;
        RECT 372.825 4133.365 373.105 4133.645 ;
        RECT 373.535 4133.365 373.815 4133.645 ;
        RECT 374.245 4133.365 374.525 4133.645 ;
        RECT 374.955 4133.365 375.235 4133.645 ;
        RECT 375.665 4133.365 375.945 4133.645 ;
        RECT 376.375 4133.365 376.655 4133.645 ;
        RECT 369.275 4132.655 369.555 4132.935 ;
        RECT 369.985 4132.655 370.265 4132.935 ;
        RECT 370.695 4132.655 370.975 4132.935 ;
        RECT 371.405 4132.655 371.685 4132.935 ;
        RECT 372.115 4132.655 372.395 4132.935 ;
        RECT 372.825 4132.655 373.105 4132.935 ;
        RECT 373.535 4132.655 373.815 4132.935 ;
        RECT 374.245 4132.655 374.525 4132.935 ;
        RECT 374.955 4132.655 375.235 4132.935 ;
        RECT 375.665 4132.655 375.945 4132.935 ;
        RECT 376.375 4132.655 376.655 4132.935 ;
        RECT 369.275 4131.945 369.555 4132.225 ;
        RECT 369.985 4131.945 370.265 4132.225 ;
        RECT 370.695 4131.945 370.975 4132.225 ;
        RECT 371.405 4131.945 371.685 4132.225 ;
        RECT 372.115 4131.945 372.395 4132.225 ;
        RECT 372.825 4131.945 373.105 4132.225 ;
        RECT 373.535 4131.945 373.815 4132.225 ;
        RECT 374.245 4131.945 374.525 4132.225 ;
        RECT 374.955 4131.945 375.235 4132.225 ;
        RECT 375.665 4131.945 375.945 4132.225 ;
        RECT 376.375 4131.945 376.655 4132.225 ;
        RECT 369.275 4131.235 369.555 4131.515 ;
        RECT 369.985 4131.235 370.265 4131.515 ;
        RECT 370.695 4131.235 370.975 4131.515 ;
        RECT 371.405 4131.235 371.685 4131.515 ;
        RECT 372.115 4131.235 372.395 4131.515 ;
        RECT 372.825 4131.235 373.105 4131.515 ;
        RECT 373.535 4131.235 373.815 4131.515 ;
        RECT 374.245 4131.235 374.525 4131.515 ;
        RECT 374.955 4131.235 375.235 4131.515 ;
        RECT 375.665 4131.235 375.945 4131.515 ;
        RECT 376.375 4131.235 376.655 4131.515 ;
        RECT 369.275 4130.525 369.555 4130.805 ;
        RECT 369.985 4130.525 370.265 4130.805 ;
        RECT 370.695 4130.525 370.975 4130.805 ;
        RECT 371.405 4130.525 371.685 4130.805 ;
        RECT 372.115 4130.525 372.395 4130.805 ;
        RECT 372.825 4130.525 373.105 4130.805 ;
        RECT 373.535 4130.525 373.815 4130.805 ;
        RECT 374.245 4130.525 374.525 4130.805 ;
        RECT 374.955 4130.525 375.235 4130.805 ;
        RECT 375.665 4130.525 375.945 4130.805 ;
        RECT 376.375 4130.525 376.655 4130.805 ;
        RECT 369.275 4129.815 369.555 4130.095 ;
        RECT 369.985 4129.815 370.265 4130.095 ;
        RECT 370.695 4129.815 370.975 4130.095 ;
        RECT 371.405 4129.815 371.685 4130.095 ;
        RECT 372.115 4129.815 372.395 4130.095 ;
        RECT 372.825 4129.815 373.105 4130.095 ;
        RECT 373.535 4129.815 373.815 4130.095 ;
        RECT 374.245 4129.815 374.525 4130.095 ;
        RECT 374.955 4129.815 375.235 4130.095 ;
        RECT 375.665 4129.815 375.945 4130.095 ;
        RECT 376.375 4129.815 376.655 4130.095 ;
        RECT 369.275 4129.105 369.555 4129.385 ;
        RECT 369.985 4129.105 370.265 4129.385 ;
        RECT 370.695 4129.105 370.975 4129.385 ;
        RECT 371.405 4129.105 371.685 4129.385 ;
        RECT 372.115 4129.105 372.395 4129.385 ;
        RECT 372.825 4129.105 373.105 4129.385 ;
        RECT 373.535 4129.105 373.815 4129.385 ;
        RECT 374.245 4129.105 374.525 4129.385 ;
        RECT 374.955 4129.105 375.235 4129.385 ;
        RECT 375.665 4129.105 375.945 4129.385 ;
        RECT 376.375 4129.105 376.655 4129.385 ;
        RECT 369.330 4125.190 369.610 4125.470 ;
        RECT 370.040 4125.190 370.320 4125.470 ;
        RECT 370.750 4125.190 371.030 4125.470 ;
        RECT 371.460 4125.190 371.740 4125.470 ;
        RECT 372.170 4125.190 372.450 4125.470 ;
        RECT 372.880 4125.190 373.160 4125.470 ;
        RECT 373.590 4125.190 373.870 4125.470 ;
        RECT 374.300 4125.190 374.580 4125.470 ;
        RECT 375.010 4125.190 375.290 4125.470 ;
        RECT 375.720 4125.190 376.000 4125.470 ;
        RECT 376.430 4125.190 376.710 4125.470 ;
        RECT 369.330 4124.480 369.610 4124.760 ;
        RECT 370.040 4124.480 370.320 4124.760 ;
        RECT 370.750 4124.480 371.030 4124.760 ;
        RECT 371.460 4124.480 371.740 4124.760 ;
        RECT 372.170 4124.480 372.450 4124.760 ;
        RECT 372.880 4124.480 373.160 4124.760 ;
        RECT 373.590 4124.480 373.870 4124.760 ;
        RECT 374.300 4124.480 374.580 4124.760 ;
        RECT 375.010 4124.480 375.290 4124.760 ;
        RECT 375.720 4124.480 376.000 4124.760 ;
        RECT 376.430 4124.480 376.710 4124.760 ;
        RECT 369.330 4123.770 369.610 4124.050 ;
        RECT 370.040 4123.770 370.320 4124.050 ;
        RECT 370.750 4123.770 371.030 4124.050 ;
        RECT 371.460 4123.770 371.740 4124.050 ;
        RECT 372.170 4123.770 372.450 4124.050 ;
        RECT 372.880 4123.770 373.160 4124.050 ;
        RECT 373.590 4123.770 373.870 4124.050 ;
        RECT 374.300 4123.770 374.580 4124.050 ;
        RECT 375.010 4123.770 375.290 4124.050 ;
        RECT 375.720 4123.770 376.000 4124.050 ;
        RECT 376.430 4123.770 376.710 4124.050 ;
        RECT 369.330 4123.060 369.610 4123.340 ;
        RECT 370.040 4123.060 370.320 4123.340 ;
        RECT 370.750 4123.060 371.030 4123.340 ;
        RECT 371.460 4123.060 371.740 4123.340 ;
        RECT 372.170 4123.060 372.450 4123.340 ;
        RECT 372.880 4123.060 373.160 4123.340 ;
        RECT 373.590 4123.060 373.870 4123.340 ;
        RECT 374.300 4123.060 374.580 4123.340 ;
        RECT 375.010 4123.060 375.290 4123.340 ;
        RECT 375.720 4123.060 376.000 4123.340 ;
        RECT 376.430 4123.060 376.710 4123.340 ;
        RECT 369.330 4122.350 369.610 4122.630 ;
        RECT 370.040 4122.350 370.320 4122.630 ;
        RECT 370.750 4122.350 371.030 4122.630 ;
        RECT 371.460 4122.350 371.740 4122.630 ;
        RECT 372.170 4122.350 372.450 4122.630 ;
        RECT 372.880 4122.350 373.160 4122.630 ;
        RECT 373.590 4122.350 373.870 4122.630 ;
        RECT 374.300 4122.350 374.580 4122.630 ;
        RECT 375.010 4122.350 375.290 4122.630 ;
        RECT 375.720 4122.350 376.000 4122.630 ;
        RECT 376.430 4122.350 376.710 4122.630 ;
        RECT 369.330 4121.640 369.610 4121.920 ;
        RECT 370.040 4121.640 370.320 4121.920 ;
        RECT 370.750 4121.640 371.030 4121.920 ;
        RECT 371.460 4121.640 371.740 4121.920 ;
        RECT 372.170 4121.640 372.450 4121.920 ;
        RECT 372.880 4121.640 373.160 4121.920 ;
        RECT 373.590 4121.640 373.870 4121.920 ;
        RECT 374.300 4121.640 374.580 4121.920 ;
        RECT 375.010 4121.640 375.290 4121.920 ;
        RECT 375.720 4121.640 376.000 4121.920 ;
        RECT 376.430 4121.640 376.710 4121.920 ;
        RECT 369.330 4120.930 369.610 4121.210 ;
        RECT 370.040 4120.930 370.320 4121.210 ;
        RECT 370.750 4120.930 371.030 4121.210 ;
        RECT 371.460 4120.930 371.740 4121.210 ;
        RECT 372.170 4120.930 372.450 4121.210 ;
        RECT 372.880 4120.930 373.160 4121.210 ;
        RECT 373.590 4120.930 373.870 4121.210 ;
        RECT 374.300 4120.930 374.580 4121.210 ;
        RECT 375.010 4120.930 375.290 4121.210 ;
        RECT 375.720 4120.930 376.000 4121.210 ;
        RECT 376.430 4120.930 376.710 4121.210 ;
        RECT 369.330 4120.220 369.610 4120.500 ;
        RECT 370.040 4120.220 370.320 4120.500 ;
        RECT 370.750 4120.220 371.030 4120.500 ;
        RECT 371.460 4120.220 371.740 4120.500 ;
        RECT 372.170 4120.220 372.450 4120.500 ;
        RECT 372.880 4120.220 373.160 4120.500 ;
        RECT 373.590 4120.220 373.870 4120.500 ;
        RECT 374.300 4120.220 374.580 4120.500 ;
        RECT 375.010 4120.220 375.290 4120.500 ;
        RECT 375.720 4120.220 376.000 4120.500 ;
        RECT 376.430 4120.220 376.710 4120.500 ;
        RECT 369.330 4119.510 369.610 4119.790 ;
        RECT 370.040 4119.510 370.320 4119.790 ;
        RECT 370.750 4119.510 371.030 4119.790 ;
        RECT 371.460 4119.510 371.740 4119.790 ;
        RECT 372.170 4119.510 372.450 4119.790 ;
        RECT 372.880 4119.510 373.160 4119.790 ;
        RECT 373.590 4119.510 373.870 4119.790 ;
        RECT 374.300 4119.510 374.580 4119.790 ;
        RECT 375.010 4119.510 375.290 4119.790 ;
        RECT 375.720 4119.510 376.000 4119.790 ;
        RECT 376.430 4119.510 376.710 4119.790 ;
        RECT 369.330 4118.800 369.610 4119.080 ;
        RECT 370.040 4118.800 370.320 4119.080 ;
        RECT 370.750 4118.800 371.030 4119.080 ;
        RECT 371.460 4118.800 371.740 4119.080 ;
        RECT 372.170 4118.800 372.450 4119.080 ;
        RECT 372.880 4118.800 373.160 4119.080 ;
        RECT 373.590 4118.800 373.870 4119.080 ;
        RECT 374.300 4118.800 374.580 4119.080 ;
        RECT 375.010 4118.800 375.290 4119.080 ;
        RECT 375.720 4118.800 376.000 4119.080 ;
        RECT 376.430 4118.800 376.710 4119.080 ;
        RECT 369.330 4118.090 369.610 4118.370 ;
        RECT 370.040 4118.090 370.320 4118.370 ;
        RECT 370.750 4118.090 371.030 4118.370 ;
        RECT 371.460 4118.090 371.740 4118.370 ;
        RECT 372.170 4118.090 372.450 4118.370 ;
        RECT 372.880 4118.090 373.160 4118.370 ;
        RECT 373.590 4118.090 373.870 4118.370 ;
        RECT 374.300 4118.090 374.580 4118.370 ;
        RECT 375.010 4118.090 375.290 4118.370 ;
        RECT 375.720 4118.090 376.000 4118.370 ;
        RECT 376.430 4118.090 376.710 4118.370 ;
        RECT 369.330 4117.380 369.610 4117.660 ;
        RECT 370.040 4117.380 370.320 4117.660 ;
        RECT 370.750 4117.380 371.030 4117.660 ;
        RECT 371.460 4117.380 371.740 4117.660 ;
        RECT 372.170 4117.380 372.450 4117.660 ;
        RECT 372.880 4117.380 373.160 4117.660 ;
        RECT 373.590 4117.380 373.870 4117.660 ;
        RECT 374.300 4117.380 374.580 4117.660 ;
        RECT 375.010 4117.380 375.290 4117.660 ;
        RECT 375.720 4117.380 376.000 4117.660 ;
        RECT 376.430 4117.380 376.710 4117.660 ;
        RECT 369.330 4116.670 369.610 4116.950 ;
        RECT 370.040 4116.670 370.320 4116.950 ;
        RECT 370.750 4116.670 371.030 4116.950 ;
        RECT 371.460 4116.670 371.740 4116.950 ;
        RECT 372.170 4116.670 372.450 4116.950 ;
        RECT 372.880 4116.670 373.160 4116.950 ;
        RECT 373.590 4116.670 373.870 4116.950 ;
        RECT 374.300 4116.670 374.580 4116.950 ;
        RECT 375.010 4116.670 375.290 4116.950 ;
        RECT 375.720 4116.670 376.000 4116.950 ;
        RECT 376.430 4116.670 376.710 4116.950 ;
        RECT 357.330 3982.970 357.610 3983.250 ;
        RECT 358.040 3982.970 358.320 3983.250 ;
        RECT 358.750 3982.970 359.030 3983.250 ;
        RECT 359.460 3982.970 359.740 3983.250 ;
        RECT 360.170 3982.970 360.450 3983.250 ;
        RECT 360.880 3982.970 361.160 3983.250 ;
        RECT 361.590 3982.970 361.870 3983.250 ;
        RECT 362.300 3982.970 362.580 3983.250 ;
        RECT 363.010 3982.970 363.290 3983.250 ;
        RECT 363.720 3982.970 364.000 3983.250 ;
        RECT 364.430 3982.970 364.710 3983.250 ;
        RECT 365.140 3982.970 365.420 3983.250 ;
        RECT 365.850 3982.970 366.130 3983.250 ;
        RECT 366.560 3982.970 366.840 3983.250 ;
        RECT 357.330 3982.260 357.610 3982.540 ;
        RECT 358.040 3982.260 358.320 3982.540 ;
        RECT 358.750 3982.260 359.030 3982.540 ;
        RECT 359.460 3982.260 359.740 3982.540 ;
        RECT 360.170 3982.260 360.450 3982.540 ;
        RECT 360.880 3982.260 361.160 3982.540 ;
        RECT 361.590 3982.260 361.870 3982.540 ;
        RECT 362.300 3982.260 362.580 3982.540 ;
        RECT 363.010 3982.260 363.290 3982.540 ;
        RECT 363.720 3982.260 364.000 3982.540 ;
        RECT 364.430 3982.260 364.710 3982.540 ;
        RECT 365.140 3982.260 365.420 3982.540 ;
        RECT 365.850 3982.260 366.130 3982.540 ;
        RECT 366.560 3982.260 366.840 3982.540 ;
        RECT 357.330 3981.550 357.610 3981.830 ;
        RECT 358.040 3981.550 358.320 3981.830 ;
        RECT 358.750 3981.550 359.030 3981.830 ;
        RECT 359.460 3981.550 359.740 3981.830 ;
        RECT 360.170 3981.550 360.450 3981.830 ;
        RECT 360.880 3981.550 361.160 3981.830 ;
        RECT 361.590 3981.550 361.870 3981.830 ;
        RECT 362.300 3981.550 362.580 3981.830 ;
        RECT 363.010 3981.550 363.290 3981.830 ;
        RECT 363.720 3981.550 364.000 3981.830 ;
        RECT 364.430 3981.550 364.710 3981.830 ;
        RECT 365.140 3981.550 365.420 3981.830 ;
        RECT 365.850 3981.550 366.130 3981.830 ;
        RECT 366.560 3981.550 366.840 3981.830 ;
        RECT 357.330 3980.840 357.610 3981.120 ;
        RECT 358.040 3980.840 358.320 3981.120 ;
        RECT 358.750 3980.840 359.030 3981.120 ;
        RECT 359.460 3980.840 359.740 3981.120 ;
        RECT 360.170 3980.840 360.450 3981.120 ;
        RECT 360.880 3980.840 361.160 3981.120 ;
        RECT 361.590 3980.840 361.870 3981.120 ;
        RECT 362.300 3980.840 362.580 3981.120 ;
        RECT 363.010 3980.840 363.290 3981.120 ;
        RECT 363.720 3980.840 364.000 3981.120 ;
        RECT 364.430 3980.840 364.710 3981.120 ;
        RECT 365.140 3980.840 365.420 3981.120 ;
        RECT 365.850 3980.840 366.130 3981.120 ;
        RECT 366.560 3980.840 366.840 3981.120 ;
        RECT 357.330 3980.130 357.610 3980.410 ;
        RECT 358.040 3980.130 358.320 3980.410 ;
        RECT 358.750 3980.130 359.030 3980.410 ;
        RECT 359.460 3980.130 359.740 3980.410 ;
        RECT 360.170 3980.130 360.450 3980.410 ;
        RECT 360.880 3980.130 361.160 3980.410 ;
        RECT 361.590 3980.130 361.870 3980.410 ;
        RECT 362.300 3980.130 362.580 3980.410 ;
        RECT 363.010 3980.130 363.290 3980.410 ;
        RECT 363.720 3980.130 364.000 3980.410 ;
        RECT 364.430 3980.130 364.710 3980.410 ;
        RECT 365.140 3980.130 365.420 3980.410 ;
        RECT 365.850 3980.130 366.130 3980.410 ;
        RECT 366.560 3980.130 366.840 3980.410 ;
        RECT 357.330 3979.420 357.610 3979.700 ;
        RECT 358.040 3979.420 358.320 3979.700 ;
        RECT 358.750 3979.420 359.030 3979.700 ;
        RECT 359.460 3979.420 359.740 3979.700 ;
        RECT 360.170 3979.420 360.450 3979.700 ;
        RECT 360.880 3979.420 361.160 3979.700 ;
        RECT 361.590 3979.420 361.870 3979.700 ;
        RECT 362.300 3979.420 362.580 3979.700 ;
        RECT 363.010 3979.420 363.290 3979.700 ;
        RECT 363.720 3979.420 364.000 3979.700 ;
        RECT 364.430 3979.420 364.710 3979.700 ;
        RECT 365.140 3979.420 365.420 3979.700 ;
        RECT 365.850 3979.420 366.130 3979.700 ;
        RECT 366.560 3979.420 366.840 3979.700 ;
        RECT 357.330 3978.710 357.610 3978.990 ;
        RECT 358.040 3978.710 358.320 3978.990 ;
        RECT 358.750 3978.710 359.030 3978.990 ;
        RECT 359.460 3978.710 359.740 3978.990 ;
        RECT 360.170 3978.710 360.450 3978.990 ;
        RECT 360.880 3978.710 361.160 3978.990 ;
        RECT 361.590 3978.710 361.870 3978.990 ;
        RECT 362.300 3978.710 362.580 3978.990 ;
        RECT 363.010 3978.710 363.290 3978.990 ;
        RECT 363.720 3978.710 364.000 3978.990 ;
        RECT 364.430 3978.710 364.710 3978.990 ;
        RECT 365.140 3978.710 365.420 3978.990 ;
        RECT 365.850 3978.710 366.130 3978.990 ;
        RECT 366.560 3978.710 366.840 3978.990 ;
        RECT 357.330 3978.000 357.610 3978.280 ;
        RECT 358.040 3978.000 358.320 3978.280 ;
        RECT 358.750 3978.000 359.030 3978.280 ;
        RECT 359.460 3978.000 359.740 3978.280 ;
        RECT 360.170 3978.000 360.450 3978.280 ;
        RECT 360.880 3978.000 361.160 3978.280 ;
        RECT 361.590 3978.000 361.870 3978.280 ;
        RECT 362.300 3978.000 362.580 3978.280 ;
        RECT 363.010 3978.000 363.290 3978.280 ;
        RECT 363.720 3978.000 364.000 3978.280 ;
        RECT 364.430 3978.000 364.710 3978.280 ;
        RECT 365.140 3978.000 365.420 3978.280 ;
        RECT 365.850 3978.000 366.130 3978.280 ;
        RECT 366.560 3978.000 366.840 3978.280 ;
        RECT 357.330 3977.290 357.610 3977.570 ;
        RECT 358.040 3977.290 358.320 3977.570 ;
        RECT 358.750 3977.290 359.030 3977.570 ;
        RECT 359.460 3977.290 359.740 3977.570 ;
        RECT 360.170 3977.290 360.450 3977.570 ;
        RECT 360.880 3977.290 361.160 3977.570 ;
        RECT 361.590 3977.290 361.870 3977.570 ;
        RECT 362.300 3977.290 362.580 3977.570 ;
        RECT 363.010 3977.290 363.290 3977.570 ;
        RECT 363.720 3977.290 364.000 3977.570 ;
        RECT 364.430 3977.290 364.710 3977.570 ;
        RECT 365.140 3977.290 365.420 3977.570 ;
        RECT 365.850 3977.290 366.130 3977.570 ;
        RECT 366.560 3977.290 366.840 3977.570 ;
        RECT 357.330 3976.580 357.610 3976.860 ;
        RECT 358.040 3976.580 358.320 3976.860 ;
        RECT 358.750 3976.580 359.030 3976.860 ;
        RECT 359.460 3976.580 359.740 3976.860 ;
        RECT 360.170 3976.580 360.450 3976.860 ;
        RECT 360.880 3976.580 361.160 3976.860 ;
        RECT 361.590 3976.580 361.870 3976.860 ;
        RECT 362.300 3976.580 362.580 3976.860 ;
        RECT 363.010 3976.580 363.290 3976.860 ;
        RECT 363.720 3976.580 364.000 3976.860 ;
        RECT 364.430 3976.580 364.710 3976.860 ;
        RECT 365.140 3976.580 365.420 3976.860 ;
        RECT 365.850 3976.580 366.130 3976.860 ;
        RECT 366.560 3976.580 366.840 3976.860 ;
        RECT 357.330 3975.870 357.610 3976.150 ;
        RECT 358.040 3975.870 358.320 3976.150 ;
        RECT 358.750 3975.870 359.030 3976.150 ;
        RECT 359.460 3975.870 359.740 3976.150 ;
        RECT 360.170 3975.870 360.450 3976.150 ;
        RECT 360.880 3975.870 361.160 3976.150 ;
        RECT 361.590 3975.870 361.870 3976.150 ;
        RECT 362.300 3975.870 362.580 3976.150 ;
        RECT 363.010 3975.870 363.290 3976.150 ;
        RECT 363.720 3975.870 364.000 3976.150 ;
        RECT 364.430 3975.870 364.710 3976.150 ;
        RECT 365.140 3975.870 365.420 3976.150 ;
        RECT 365.850 3975.870 366.130 3976.150 ;
        RECT 366.560 3975.870 366.840 3976.150 ;
        RECT 357.330 3975.160 357.610 3975.440 ;
        RECT 358.040 3975.160 358.320 3975.440 ;
        RECT 358.750 3975.160 359.030 3975.440 ;
        RECT 359.460 3975.160 359.740 3975.440 ;
        RECT 360.170 3975.160 360.450 3975.440 ;
        RECT 360.880 3975.160 361.160 3975.440 ;
        RECT 361.590 3975.160 361.870 3975.440 ;
        RECT 362.300 3975.160 362.580 3975.440 ;
        RECT 363.010 3975.160 363.290 3975.440 ;
        RECT 363.720 3975.160 364.000 3975.440 ;
        RECT 364.430 3975.160 364.710 3975.440 ;
        RECT 365.140 3975.160 365.420 3975.440 ;
        RECT 365.850 3975.160 366.130 3975.440 ;
        RECT 366.560 3975.160 366.840 3975.440 ;
        RECT 357.330 3974.450 357.610 3974.730 ;
        RECT 358.040 3974.450 358.320 3974.730 ;
        RECT 358.750 3974.450 359.030 3974.730 ;
        RECT 359.460 3974.450 359.740 3974.730 ;
        RECT 360.170 3974.450 360.450 3974.730 ;
        RECT 360.880 3974.450 361.160 3974.730 ;
        RECT 361.590 3974.450 361.870 3974.730 ;
        RECT 362.300 3974.450 362.580 3974.730 ;
        RECT 363.010 3974.450 363.290 3974.730 ;
        RECT 363.720 3974.450 364.000 3974.730 ;
        RECT 364.430 3974.450 364.710 3974.730 ;
        RECT 365.140 3974.450 365.420 3974.730 ;
        RECT 365.850 3974.450 366.130 3974.730 ;
        RECT 366.560 3974.450 366.840 3974.730 ;
        RECT 357.275 3970.565 357.555 3970.845 ;
        RECT 357.985 3970.565 358.265 3970.845 ;
        RECT 358.695 3970.565 358.975 3970.845 ;
        RECT 359.405 3970.565 359.685 3970.845 ;
        RECT 360.115 3970.565 360.395 3970.845 ;
        RECT 360.825 3970.565 361.105 3970.845 ;
        RECT 361.535 3970.565 361.815 3970.845 ;
        RECT 362.245 3970.565 362.525 3970.845 ;
        RECT 362.955 3970.565 363.235 3970.845 ;
        RECT 363.665 3970.565 363.945 3970.845 ;
        RECT 364.375 3970.565 364.655 3970.845 ;
        RECT 365.085 3970.565 365.365 3970.845 ;
        RECT 365.795 3970.565 366.075 3970.845 ;
        RECT 366.505 3970.565 366.785 3970.845 ;
        RECT 357.275 3969.855 357.555 3970.135 ;
        RECT 357.985 3969.855 358.265 3970.135 ;
        RECT 358.695 3969.855 358.975 3970.135 ;
        RECT 359.405 3969.855 359.685 3970.135 ;
        RECT 360.115 3969.855 360.395 3970.135 ;
        RECT 360.825 3969.855 361.105 3970.135 ;
        RECT 361.535 3969.855 361.815 3970.135 ;
        RECT 362.245 3969.855 362.525 3970.135 ;
        RECT 362.955 3969.855 363.235 3970.135 ;
        RECT 363.665 3969.855 363.945 3970.135 ;
        RECT 364.375 3969.855 364.655 3970.135 ;
        RECT 365.085 3969.855 365.365 3970.135 ;
        RECT 365.795 3969.855 366.075 3970.135 ;
        RECT 366.505 3969.855 366.785 3970.135 ;
        RECT 357.275 3969.145 357.555 3969.425 ;
        RECT 357.985 3969.145 358.265 3969.425 ;
        RECT 358.695 3969.145 358.975 3969.425 ;
        RECT 359.405 3969.145 359.685 3969.425 ;
        RECT 360.115 3969.145 360.395 3969.425 ;
        RECT 360.825 3969.145 361.105 3969.425 ;
        RECT 361.535 3969.145 361.815 3969.425 ;
        RECT 362.245 3969.145 362.525 3969.425 ;
        RECT 362.955 3969.145 363.235 3969.425 ;
        RECT 363.665 3969.145 363.945 3969.425 ;
        RECT 364.375 3969.145 364.655 3969.425 ;
        RECT 365.085 3969.145 365.365 3969.425 ;
        RECT 365.795 3969.145 366.075 3969.425 ;
        RECT 366.505 3969.145 366.785 3969.425 ;
        RECT 357.275 3968.435 357.555 3968.715 ;
        RECT 357.985 3968.435 358.265 3968.715 ;
        RECT 358.695 3968.435 358.975 3968.715 ;
        RECT 359.405 3968.435 359.685 3968.715 ;
        RECT 360.115 3968.435 360.395 3968.715 ;
        RECT 360.825 3968.435 361.105 3968.715 ;
        RECT 361.535 3968.435 361.815 3968.715 ;
        RECT 362.245 3968.435 362.525 3968.715 ;
        RECT 362.955 3968.435 363.235 3968.715 ;
        RECT 363.665 3968.435 363.945 3968.715 ;
        RECT 364.375 3968.435 364.655 3968.715 ;
        RECT 365.085 3968.435 365.365 3968.715 ;
        RECT 365.795 3968.435 366.075 3968.715 ;
        RECT 366.505 3968.435 366.785 3968.715 ;
        RECT 357.275 3967.725 357.555 3968.005 ;
        RECT 357.985 3967.725 358.265 3968.005 ;
        RECT 358.695 3967.725 358.975 3968.005 ;
        RECT 359.405 3967.725 359.685 3968.005 ;
        RECT 360.115 3967.725 360.395 3968.005 ;
        RECT 360.825 3967.725 361.105 3968.005 ;
        RECT 361.535 3967.725 361.815 3968.005 ;
        RECT 362.245 3967.725 362.525 3968.005 ;
        RECT 362.955 3967.725 363.235 3968.005 ;
        RECT 363.665 3967.725 363.945 3968.005 ;
        RECT 364.375 3967.725 364.655 3968.005 ;
        RECT 365.085 3967.725 365.365 3968.005 ;
        RECT 365.795 3967.725 366.075 3968.005 ;
        RECT 366.505 3967.725 366.785 3968.005 ;
        RECT 357.275 3967.015 357.555 3967.295 ;
        RECT 357.985 3967.015 358.265 3967.295 ;
        RECT 358.695 3967.015 358.975 3967.295 ;
        RECT 359.405 3967.015 359.685 3967.295 ;
        RECT 360.115 3967.015 360.395 3967.295 ;
        RECT 360.825 3967.015 361.105 3967.295 ;
        RECT 361.535 3967.015 361.815 3967.295 ;
        RECT 362.245 3967.015 362.525 3967.295 ;
        RECT 362.955 3967.015 363.235 3967.295 ;
        RECT 363.665 3967.015 363.945 3967.295 ;
        RECT 364.375 3967.015 364.655 3967.295 ;
        RECT 365.085 3967.015 365.365 3967.295 ;
        RECT 365.795 3967.015 366.075 3967.295 ;
        RECT 366.505 3967.015 366.785 3967.295 ;
        RECT 357.275 3966.305 357.555 3966.585 ;
        RECT 357.985 3966.305 358.265 3966.585 ;
        RECT 358.695 3966.305 358.975 3966.585 ;
        RECT 359.405 3966.305 359.685 3966.585 ;
        RECT 360.115 3966.305 360.395 3966.585 ;
        RECT 360.825 3966.305 361.105 3966.585 ;
        RECT 361.535 3966.305 361.815 3966.585 ;
        RECT 362.245 3966.305 362.525 3966.585 ;
        RECT 362.955 3966.305 363.235 3966.585 ;
        RECT 363.665 3966.305 363.945 3966.585 ;
        RECT 364.375 3966.305 364.655 3966.585 ;
        RECT 365.085 3966.305 365.365 3966.585 ;
        RECT 365.795 3966.305 366.075 3966.585 ;
        RECT 366.505 3966.305 366.785 3966.585 ;
        RECT 357.275 3965.595 357.555 3965.875 ;
        RECT 357.985 3965.595 358.265 3965.875 ;
        RECT 358.695 3965.595 358.975 3965.875 ;
        RECT 359.405 3965.595 359.685 3965.875 ;
        RECT 360.115 3965.595 360.395 3965.875 ;
        RECT 360.825 3965.595 361.105 3965.875 ;
        RECT 361.535 3965.595 361.815 3965.875 ;
        RECT 362.245 3965.595 362.525 3965.875 ;
        RECT 362.955 3965.595 363.235 3965.875 ;
        RECT 363.665 3965.595 363.945 3965.875 ;
        RECT 364.375 3965.595 364.655 3965.875 ;
        RECT 365.085 3965.595 365.365 3965.875 ;
        RECT 365.795 3965.595 366.075 3965.875 ;
        RECT 366.505 3965.595 366.785 3965.875 ;
        RECT 357.275 3964.885 357.555 3965.165 ;
        RECT 357.985 3964.885 358.265 3965.165 ;
        RECT 358.695 3964.885 358.975 3965.165 ;
        RECT 359.405 3964.885 359.685 3965.165 ;
        RECT 360.115 3964.885 360.395 3965.165 ;
        RECT 360.825 3964.885 361.105 3965.165 ;
        RECT 361.535 3964.885 361.815 3965.165 ;
        RECT 362.245 3964.885 362.525 3965.165 ;
        RECT 362.955 3964.885 363.235 3965.165 ;
        RECT 363.665 3964.885 363.945 3965.165 ;
        RECT 364.375 3964.885 364.655 3965.165 ;
        RECT 365.085 3964.885 365.365 3965.165 ;
        RECT 365.795 3964.885 366.075 3965.165 ;
        RECT 366.505 3964.885 366.785 3965.165 ;
        RECT 357.275 3964.175 357.555 3964.455 ;
        RECT 357.985 3964.175 358.265 3964.455 ;
        RECT 358.695 3964.175 358.975 3964.455 ;
        RECT 359.405 3964.175 359.685 3964.455 ;
        RECT 360.115 3964.175 360.395 3964.455 ;
        RECT 360.825 3964.175 361.105 3964.455 ;
        RECT 361.535 3964.175 361.815 3964.455 ;
        RECT 362.245 3964.175 362.525 3964.455 ;
        RECT 362.955 3964.175 363.235 3964.455 ;
        RECT 363.665 3964.175 363.945 3964.455 ;
        RECT 364.375 3964.175 364.655 3964.455 ;
        RECT 365.085 3964.175 365.365 3964.455 ;
        RECT 365.795 3964.175 366.075 3964.455 ;
        RECT 366.505 3964.175 366.785 3964.455 ;
        RECT 357.275 3963.465 357.555 3963.745 ;
        RECT 357.985 3963.465 358.265 3963.745 ;
        RECT 358.695 3963.465 358.975 3963.745 ;
        RECT 359.405 3963.465 359.685 3963.745 ;
        RECT 360.115 3963.465 360.395 3963.745 ;
        RECT 360.825 3963.465 361.105 3963.745 ;
        RECT 361.535 3963.465 361.815 3963.745 ;
        RECT 362.245 3963.465 362.525 3963.745 ;
        RECT 362.955 3963.465 363.235 3963.745 ;
        RECT 363.665 3963.465 363.945 3963.745 ;
        RECT 364.375 3963.465 364.655 3963.745 ;
        RECT 365.085 3963.465 365.365 3963.745 ;
        RECT 365.795 3963.465 366.075 3963.745 ;
        RECT 366.505 3963.465 366.785 3963.745 ;
        RECT 357.275 3962.755 357.555 3963.035 ;
        RECT 357.985 3962.755 358.265 3963.035 ;
        RECT 358.695 3962.755 358.975 3963.035 ;
        RECT 359.405 3962.755 359.685 3963.035 ;
        RECT 360.115 3962.755 360.395 3963.035 ;
        RECT 360.825 3962.755 361.105 3963.035 ;
        RECT 361.535 3962.755 361.815 3963.035 ;
        RECT 362.245 3962.755 362.525 3963.035 ;
        RECT 362.955 3962.755 363.235 3963.035 ;
        RECT 363.665 3962.755 363.945 3963.035 ;
        RECT 364.375 3962.755 364.655 3963.035 ;
        RECT 365.085 3962.755 365.365 3963.035 ;
        RECT 365.795 3962.755 366.075 3963.035 ;
        RECT 366.505 3962.755 366.785 3963.035 ;
        RECT 357.275 3962.045 357.555 3962.325 ;
        RECT 357.985 3962.045 358.265 3962.325 ;
        RECT 358.695 3962.045 358.975 3962.325 ;
        RECT 359.405 3962.045 359.685 3962.325 ;
        RECT 360.115 3962.045 360.395 3962.325 ;
        RECT 360.825 3962.045 361.105 3962.325 ;
        RECT 361.535 3962.045 361.815 3962.325 ;
        RECT 362.245 3962.045 362.525 3962.325 ;
        RECT 362.955 3962.045 363.235 3962.325 ;
        RECT 363.665 3962.045 363.945 3962.325 ;
        RECT 364.375 3962.045 364.655 3962.325 ;
        RECT 365.085 3962.045 365.365 3962.325 ;
        RECT 365.795 3962.045 366.075 3962.325 ;
        RECT 366.505 3962.045 366.785 3962.325 ;
        RECT 357.275 3961.335 357.555 3961.615 ;
        RECT 357.985 3961.335 358.265 3961.615 ;
        RECT 358.695 3961.335 358.975 3961.615 ;
        RECT 359.405 3961.335 359.685 3961.615 ;
        RECT 360.115 3961.335 360.395 3961.615 ;
        RECT 360.825 3961.335 361.105 3961.615 ;
        RECT 361.535 3961.335 361.815 3961.615 ;
        RECT 362.245 3961.335 362.525 3961.615 ;
        RECT 362.955 3961.335 363.235 3961.615 ;
        RECT 363.665 3961.335 363.945 3961.615 ;
        RECT 364.375 3961.335 364.655 3961.615 ;
        RECT 365.085 3961.335 365.365 3961.615 ;
        RECT 365.795 3961.335 366.075 3961.615 ;
        RECT 366.505 3961.335 366.785 3961.615 ;
        RECT 357.275 3958.715 357.555 3958.995 ;
        RECT 357.985 3958.715 358.265 3958.995 ;
        RECT 358.695 3958.715 358.975 3958.995 ;
        RECT 359.405 3958.715 359.685 3958.995 ;
        RECT 360.115 3958.715 360.395 3958.995 ;
        RECT 360.825 3958.715 361.105 3958.995 ;
        RECT 361.535 3958.715 361.815 3958.995 ;
        RECT 362.245 3958.715 362.525 3958.995 ;
        RECT 362.955 3958.715 363.235 3958.995 ;
        RECT 363.665 3958.715 363.945 3958.995 ;
        RECT 364.375 3958.715 364.655 3958.995 ;
        RECT 365.085 3958.715 365.365 3958.995 ;
        RECT 365.795 3958.715 366.075 3958.995 ;
        RECT 366.505 3958.715 366.785 3958.995 ;
        RECT 357.275 3958.005 357.555 3958.285 ;
        RECT 357.985 3958.005 358.265 3958.285 ;
        RECT 358.695 3958.005 358.975 3958.285 ;
        RECT 359.405 3958.005 359.685 3958.285 ;
        RECT 360.115 3958.005 360.395 3958.285 ;
        RECT 360.825 3958.005 361.105 3958.285 ;
        RECT 361.535 3958.005 361.815 3958.285 ;
        RECT 362.245 3958.005 362.525 3958.285 ;
        RECT 362.955 3958.005 363.235 3958.285 ;
        RECT 363.665 3958.005 363.945 3958.285 ;
        RECT 364.375 3958.005 364.655 3958.285 ;
        RECT 365.085 3958.005 365.365 3958.285 ;
        RECT 365.795 3958.005 366.075 3958.285 ;
        RECT 366.505 3958.005 366.785 3958.285 ;
        RECT 357.275 3957.295 357.555 3957.575 ;
        RECT 357.985 3957.295 358.265 3957.575 ;
        RECT 358.695 3957.295 358.975 3957.575 ;
        RECT 359.405 3957.295 359.685 3957.575 ;
        RECT 360.115 3957.295 360.395 3957.575 ;
        RECT 360.825 3957.295 361.105 3957.575 ;
        RECT 361.535 3957.295 361.815 3957.575 ;
        RECT 362.245 3957.295 362.525 3957.575 ;
        RECT 362.955 3957.295 363.235 3957.575 ;
        RECT 363.665 3957.295 363.945 3957.575 ;
        RECT 364.375 3957.295 364.655 3957.575 ;
        RECT 365.085 3957.295 365.365 3957.575 ;
        RECT 365.795 3957.295 366.075 3957.575 ;
        RECT 366.505 3957.295 366.785 3957.575 ;
        RECT 357.275 3956.585 357.555 3956.865 ;
        RECT 357.985 3956.585 358.265 3956.865 ;
        RECT 358.695 3956.585 358.975 3956.865 ;
        RECT 359.405 3956.585 359.685 3956.865 ;
        RECT 360.115 3956.585 360.395 3956.865 ;
        RECT 360.825 3956.585 361.105 3956.865 ;
        RECT 361.535 3956.585 361.815 3956.865 ;
        RECT 362.245 3956.585 362.525 3956.865 ;
        RECT 362.955 3956.585 363.235 3956.865 ;
        RECT 363.665 3956.585 363.945 3956.865 ;
        RECT 364.375 3956.585 364.655 3956.865 ;
        RECT 365.085 3956.585 365.365 3956.865 ;
        RECT 365.795 3956.585 366.075 3956.865 ;
        RECT 366.505 3956.585 366.785 3956.865 ;
        RECT 357.275 3955.875 357.555 3956.155 ;
        RECT 357.985 3955.875 358.265 3956.155 ;
        RECT 358.695 3955.875 358.975 3956.155 ;
        RECT 359.405 3955.875 359.685 3956.155 ;
        RECT 360.115 3955.875 360.395 3956.155 ;
        RECT 360.825 3955.875 361.105 3956.155 ;
        RECT 361.535 3955.875 361.815 3956.155 ;
        RECT 362.245 3955.875 362.525 3956.155 ;
        RECT 362.955 3955.875 363.235 3956.155 ;
        RECT 363.665 3955.875 363.945 3956.155 ;
        RECT 364.375 3955.875 364.655 3956.155 ;
        RECT 365.085 3955.875 365.365 3956.155 ;
        RECT 365.795 3955.875 366.075 3956.155 ;
        RECT 366.505 3955.875 366.785 3956.155 ;
        RECT 357.275 3955.165 357.555 3955.445 ;
        RECT 357.985 3955.165 358.265 3955.445 ;
        RECT 358.695 3955.165 358.975 3955.445 ;
        RECT 359.405 3955.165 359.685 3955.445 ;
        RECT 360.115 3955.165 360.395 3955.445 ;
        RECT 360.825 3955.165 361.105 3955.445 ;
        RECT 361.535 3955.165 361.815 3955.445 ;
        RECT 362.245 3955.165 362.525 3955.445 ;
        RECT 362.955 3955.165 363.235 3955.445 ;
        RECT 363.665 3955.165 363.945 3955.445 ;
        RECT 364.375 3955.165 364.655 3955.445 ;
        RECT 365.085 3955.165 365.365 3955.445 ;
        RECT 365.795 3955.165 366.075 3955.445 ;
        RECT 366.505 3955.165 366.785 3955.445 ;
        RECT 357.275 3954.455 357.555 3954.735 ;
        RECT 357.985 3954.455 358.265 3954.735 ;
        RECT 358.695 3954.455 358.975 3954.735 ;
        RECT 359.405 3954.455 359.685 3954.735 ;
        RECT 360.115 3954.455 360.395 3954.735 ;
        RECT 360.825 3954.455 361.105 3954.735 ;
        RECT 361.535 3954.455 361.815 3954.735 ;
        RECT 362.245 3954.455 362.525 3954.735 ;
        RECT 362.955 3954.455 363.235 3954.735 ;
        RECT 363.665 3954.455 363.945 3954.735 ;
        RECT 364.375 3954.455 364.655 3954.735 ;
        RECT 365.085 3954.455 365.365 3954.735 ;
        RECT 365.795 3954.455 366.075 3954.735 ;
        RECT 366.505 3954.455 366.785 3954.735 ;
        RECT 357.275 3953.745 357.555 3954.025 ;
        RECT 357.985 3953.745 358.265 3954.025 ;
        RECT 358.695 3953.745 358.975 3954.025 ;
        RECT 359.405 3953.745 359.685 3954.025 ;
        RECT 360.115 3953.745 360.395 3954.025 ;
        RECT 360.825 3953.745 361.105 3954.025 ;
        RECT 361.535 3953.745 361.815 3954.025 ;
        RECT 362.245 3953.745 362.525 3954.025 ;
        RECT 362.955 3953.745 363.235 3954.025 ;
        RECT 363.665 3953.745 363.945 3954.025 ;
        RECT 364.375 3953.745 364.655 3954.025 ;
        RECT 365.085 3953.745 365.365 3954.025 ;
        RECT 365.795 3953.745 366.075 3954.025 ;
        RECT 366.505 3953.745 366.785 3954.025 ;
        RECT 357.275 3953.035 357.555 3953.315 ;
        RECT 357.985 3953.035 358.265 3953.315 ;
        RECT 358.695 3953.035 358.975 3953.315 ;
        RECT 359.405 3953.035 359.685 3953.315 ;
        RECT 360.115 3953.035 360.395 3953.315 ;
        RECT 360.825 3953.035 361.105 3953.315 ;
        RECT 361.535 3953.035 361.815 3953.315 ;
        RECT 362.245 3953.035 362.525 3953.315 ;
        RECT 362.955 3953.035 363.235 3953.315 ;
        RECT 363.665 3953.035 363.945 3953.315 ;
        RECT 364.375 3953.035 364.655 3953.315 ;
        RECT 365.085 3953.035 365.365 3953.315 ;
        RECT 365.795 3953.035 366.075 3953.315 ;
        RECT 366.505 3953.035 366.785 3953.315 ;
        RECT 357.275 3952.325 357.555 3952.605 ;
        RECT 357.985 3952.325 358.265 3952.605 ;
        RECT 358.695 3952.325 358.975 3952.605 ;
        RECT 359.405 3952.325 359.685 3952.605 ;
        RECT 360.115 3952.325 360.395 3952.605 ;
        RECT 360.825 3952.325 361.105 3952.605 ;
        RECT 361.535 3952.325 361.815 3952.605 ;
        RECT 362.245 3952.325 362.525 3952.605 ;
        RECT 362.955 3952.325 363.235 3952.605 ;
        RECT 363.665 3952.325 363.945 3952.605 ;
        RECT 364.375 3952.325 364.655 3952.605 ;
        RECT 365.085 3952.325 365.365 3952.605 ;
        RECT 365.795 3952.325 366.075 3952.605 ;
        RECT 366.505 3952.325 366.785 3952.605 ;
        RECT 357.275 3951.615 357.555 3951.895 ;
        RECT 357.985 3951.615 358.265 3951.895 ;
        RECT 358.695 3951.615 358.975 3951.895 ;
        RECT 359.405 3951.615 359.685 3951.895 ;
        RECT 360.115 3951.615 360.395 3951.895 ;
        RECT 360.825 3951.615 361.105 3951.895 ;
        RECT 361.535 3951.615 361.815 3951.895 ;
        RECT 362.245 3951.615 362.525 3951.895 ;
        RECT 362.955 3951.615 363.235 3951.895 ;
        RECT 363.665 3951.615 363.945 3951.895 ;
        RECT 364.375 3951.615 364.655 3951.895 ;
        RECT 365.085 3951.615 365.365 3951.895 ;
        RECT 365.795 3951.615 366.075 3951.895 ;
        RECT 366.505 3951.615 366.785 3951.895 ;
        RECT 357.275 3950.905 357.555 3951.185 ;
        RECT 357.985 3950.905 358.265 3951.185 ;
        RECT 358.695 3950.905 358.975 3951.185 ;
        RECT 359.405 3950.905 359.685 3951.185 ;
        RECT 360.115 3950.905 360.395 3951.185 ;
        RECT 360.825 3950.905 361.105 3951.185 ;
        RECT 361.535 3950.905 361.815 3951.185 ;
        RECT 362.245 3950.905 362.525 3951.185 ;
        RECT 362.955 3950.905 363.235 3951.185 ;
        RECT 363.665 3950.905 363.945 3951.185 ;
        RECT 364.375 3950.905 364.655 3951.185 ;
        RECT 365.085 3950.905 365.365 3951.185 ;
        RECT 365.795 3950.905 366.075 3951.185 ;
        RECT 366.505 3950.905 366.785 3951.185 ;
        RECT 357.275 3950.195 357.555 3950.475 ;
        RECT 357.985 3950.195 358.265 3950.475 ;
        RECT 358.695 3950.195 358.975 3950.475 ;
        RECT 359.405 3950.195 359.685 3950.475 ;
        RECT 360.115 3950.195 360.395 3950.475 ;
        RECT 360.825 3950.195 361.105 3950.475 ;
        RECT 361.535 3950.195 361.815 3950.475 ;
        RECT 362.245 3950.195 362.525 3950.475 ;
        RECT 362.955 3950.195 363.235 3950.475 ;
        RECT 363.665 3950.195 363.945 3950.475 ;
        RECT 364.375 3950.195 364.655 3950.475 ;
        RECT 365.085 3950.195 365.365 3950.475 ;
        RECT 365.795 3950.195 366.075 3950.475 ;
        RECT 366.505 3950.195 366.785 3950.475 ;
        RECT 357.275 3949.485 357.555 3949.765 ;
        RECT 357.985 3949.485 358.265 3949.765 ;
        RECT 358.695 3949.485 358.975 3949.765 ;
        RECT 359.405 3949.485 359.685 3949.765 ;
        RECT 360.115 3949.485 360.395 3949.765 ;
        RECT 360.825 3949.485 361.105 3949.765 ;
        RECT 361.535 3949.485 361.815 3949.765 ;
        RECT 362.245 3949.485 362.525 3949.765 ;
        RECT 362.955 3949.485 363.235 3949.765 ;
        RECT 363.665 3949.485 363.945 3949.765 ;
        RECT 364.375 3949.485 364.655 3949.765 ;
        RECT 365.085 3949.485 365.365 3949.765 ;
        RECT 365.795 3949.485 366.075 3949.765 ;
        RECT 366.505 3949.485 366.785 3949.765 ;
        RECT 3500.200 3958.050 3500.480 3958.330 ;
        RECT 3500.910 3958.050 3501.190 3958.330 ;
        RECT 3501.620 3958.050 3501.900 3958.330 ;
        RECT 3502.330 3958.050 3502.610 3958.330 ;
        RECT 3503.040 3958.050 3503.320 3958.330 ;
        RECT 3503.750 3958.050 3504.030 3958.330 ;
        RECT 3504.460 3958.050 3504.740 3958.330 ;
        RECT 3505.170 3958.050 3505.450 3958.330 ;
        RECT 3505.880 3958.050 3506.160 3958.330 ;
        RECT 3506.590 3958.050 3506.870 3958.330 ;
        RECT 3507.300 3958.050 3507.580 3958.330 ;
        RECT 3508.010 3958.050 3508.290 3958.330 ;
        RECT 3508.720 3958.050 3509.000 3958.330 ;
        RECT 3509.430 3958.050 3509.710 3958.330 ;
        RECT 3500.200 3957.340 3500.480 3957.620 ;
        RECT 3500.910 3957.340 3501.190 3957.620 ;
        RECT 3501.620 3957.340 3501.900 3957.620 ;
        RECT 3502.330 3957.340 3502.610 3957.620 ;
        RECT 3503.040 3957.340 3503.320 3957.620 ;
        RECT 3503.750 3957.340 3504.030 3957.620 ;
        RECT 3504.460 3957.340 3504.740 3957.620 ;
        RECT 3505.170 3957.340 3505.450 3957.620 ;
        RECT 3505.880 3957.340 3506.160 3957.620 ;
        RECT 3506.590 3957.340 3506.870 3957.620 ;
        RECT 3507.300 3957.340 3507.580 3957.620 ;
        RECT 3508.010 3957.340 3508.290 3957.620 ;
        RECT 3508.720 3957.340 3509.000 3957.620 ;
        RECT 3509.430 3957.340 3509.710 3957.620 ;
        RECT 3500.200 3956.630 3500.480 3956.910 ;
        RECT 3500.910 3956.630 3501.190 3956.910 ;
        RECT 3501.620 3956.630 3501.900 3956.910 ;
        RECT 3502.330 3956.630 3502.610 3956.910 ;
        RECT 3503.040 3956.630 3503.320 3956.910 ;
        RECT 3503.750 3956.630 3504.030 3956.910 ;
        RECT 3504.460 3956.630 3504.740 3956.910 ;
        RECT 3505.170 3956.630 3505.450 3956.910 ;
        RECT 3505.880 3956.630 3506.160 3956.910 ;
        RECT 3506.590 3956.630 3506.870 3956.910 ;
        RECT 3507.300 3956.630 3507.580 3956.910 ;
        RECT 3508.010 3956.630 3508.290 3956.910 ;
        RECT 3508.720 3956.630 3509.000 3956.910 ;
        RECT 3509.430 3956.630 3509.710 3956.910 ;
        RECT 3500.200 3955.920 3500.480 3956.200 ;
        RECT 3500.910 3955.920 3501.190 3956.200 ;
        RECT 3501.620 3955.920 3501.900 3956.200 ;
        RECT 3502.330 3955.920 3502.610 3956.200 ;
        RECT 3503.040 3955.920 3503.320 3956.200 ;
        RECT 3503.750 3955.920 3504.030 3956.200 ;
        RECT 3504.460 3955.920 3504.740 3956.200 ;
        RECT 3505.170 3955.920 3505.450 3956.200 ;
        RECT 3505.880 3955.920 3506.160 3956.200 ;
        RECT 3506.590 3955.920 3506.870 3956.200 ;
        RECT 3507.300 3955.920 3507.580 3956.200 ;
        RECT 3508.010 3955.920 3508.290 3956.200 ;
        RECT 3508.720 3955.920 3509.000 3956.200 ;
        RECT 3509.430 3955.920 3509.710 3956.200 ;
        RECT 3500.200 3955.210 3500.480 3955.490 ;
        RECT 3500.910 3955.210 3501.190 3955.490 ;
        RECT 3501.620 3955.210 3501.900 3955.490 ;
        RECT 3502.330 3955.210 3502.610 3955.490 ;
        RECT 3503.040 3955.210 3503.320 3955.490 ;
        RECT 3503.750 3955.210 3504.030 3955.490 ;
        RECT 3504.460 3955.210 3504.740 3955.490 ;
        RECT 3505.170 3955.210 3505.450 3955.490 ;
        RECT 3505.880 3955.210 3506.160 3955.490 ;
        RECT 3506.590 3955.210 3506.870 3955.490 ;
        RECT 3507.300 3955.210 3507.580 3955.490 ;
        RECT 3508.010 3955.210 3508.290 3955.490 ;
        RECT 3508.720 3955.210 3509.000 3955.490 ;
        RECT 3509.430 3955.210 3509.710 3955.490 ;
        RECT 3500.200 3954.500 3500.480 3954.780 ;
        RECT 3500.910 3954.500 3501.190 3954.780 ;
        RECT 3501.620 3954.500 3501.900 3954.780 ;
        RECT 3502.330 3954.500 3502.610 3954.780 ;
        RECT 3503.040 3954.500 3503.320 3954.780 ;
        RECT 3503.750 3954.500 3504.030 3954.780 ;
        RECT 3504.460 3954.500 3504.740 3954.780 ;
        RECT 3505.170 3954.500 3505.450 3954.780 ;
        RECT 3505.880 3954.500 3506.160 3954.780 ;
        RECT 3506.590 3954.500 3506.870 3954.780 ;
        RECT 3507.300 3954.500 3507.580 3954.780 ;
        RECT 3508.010 3954.500 3508.290 3954.780 ;
        RECT 3508.720 3954.500 3509.000 3954.780 ;
        RECT 3509.430 3954.500 3509.710 3954.780 ;
        RECT 3500.200 3953.790 3500.480 3954.070 ;
        RECT 3500.910 3953.790 3501.190 3954.070 ;
        RECT 3501.620 3953.790 3501.900 3954.070 ;
        RECT 3502.330 3953.790 3502.610 3954.070 ;
        RECT 3503.040 3953.790 3503.320 3954.070 ;
        RECT 3503.750 3953.790 3504.030 3954.070 ;
        RECT 3504.460 3953.790 3504.740 3954.070 ;
        RECT 3505.170 3953.790 3505.450 3954.070 ;
        RECT 3505.880 3953.790 3506.160 3954.070 ;
        RECT 3506.590 3953.790 3506.870 3954.070 ;
        RECT 3507.300 3953.790 3507.580 3954.070 ;
        RECT 3508.010 3953.790 3508.290 3954.070 ;
        RECT 3508.720 3953.790 3509.000 3954.070 ;
        RECT 3509.430 3953.790 3509.710 3954.070 ;
        RECT 3500.200 3953.080 3500.480 3953.360 ;
        RECT 3500.910 3953.080 3501.190 3953.360 ;
        RECT 3501.620 3953.080 3501.900 3953.360 ;
        RECT 3502.330 3953.080 3502.610 3953.360 ;
        RECT 3503.040 3953.080 3503.320 3953.360 ;
        RECT 3503.750 3953.080 3504.030 3953.360 ;
        RECT 3504.460 3953.080 3504.740 3953.360 ;
        RECT 3505.170 3953.080 3505.450 3953.360 ;
        RECT 3505.880 3953.080 3506.160 3953.360 ;
        RECT 3506.590 3953.080 3506.870 3953.360 ;
        RECT 3507.300 3953.080 3507.580 3953.360 ;
        RECT 3508.010 3953.080 3508.290 3953.360 ;
        RECT 3508.720 3953.080 3509.000 3953.360 ;
        RECT 3509.430 3953.080 3509.710 3953.360 ;
        RECT 3500.200 3952.370 3500.480 3952.650 ;
        RECT 3500.910 3952.370 3501.190 3952.650 ;
        RECT 3501.620 3952.370 3501.900 3952.650 ;
        RECT 3502.330 3952.370 3502.610 3952.650 ;
        RECT 3503.040 3952.370 3503.320 3952.650 ;
        RECT 3503.750 3952.370 3504.030 3952.650 ;
        RECT 3504.460 3952.370 3504.740 3952.650 ;
        RECT 3505.170 3952.370 3505.450 3952.650 ;
        RECT 3505.880 3952.370 3506.160 3952.650 ;
        RECT 3506.590 3952.370 3506.870 3952.650 ;
        RECT 3507.300 3952.370 3507.580 3952.650 ;
        RECT 3508.010 3952.370 3508.290 3952.650 ;
        RECT 3508.720 3952.370 3509.000 3952.650 ;
        RECT 3509.430 3952.370 3509.710 3952.650 ;
        RECT 3500.200 3951.660 3500.480 3951.940 ;
        RECT 3500.910 3951.660 3501.190 3951.940 ;
        RECT 3501.620 3951.660 3501.900 3951.940 ;
        RECT 3502.330 3951.660 3502.610 3951.940 ;
        RECT 3503.040 3951.660 3503.320 3951.940 ;
        RECT 3503.750 3951.660 3504.030 3951.940 ;
        RECT 3504.460 3951.660 3504.740 3951.940 ;
        RECT 3505.170 3951.660 3505.450 3951.940 ;
        RECT 3505.880 3951.660 3506.160 3951.940 ;
        RECT 3506.590 3951.660 3506.870 3951.940 ;
        RECT 3507.300 3951.660 3507.580 3951.940 ;
        RECT 3508.010 3951.660 3508.290 3951.940 ;
        RECT 3508.720 3951.660 3509.000 3951.940 ;
        RECT 3509.430 3951.660 3509.710 3951.940 ;
        RECT 3500.200 3950.950 3500.480 3951.230 ;
        RECT 3500.910 3950.950 3501.190 3951.230 ;
        RECT 3501.620 3950.950 3501.900 3951.230 ;
        RECT 3502.330 3950.950 3502.610 3951.230 ;
        RECT 3503.040 3950.950 3503.320 3951.230 ;
        RECT 3503.750 3950.950 3504.030 3951.230 ;
        RECT 3504.460 3950.950 3504.740 3951.230 ;
        RECT 3505.170 3950.950 3505.450 3951.230 ;
        RECT 3505.880 3950.950 3506.160 3951.230 ;
        RECT 3506.590 3950.950 3506.870 3951.230 ;
        RECT 3507.300 3950.950 3507.580 3951.230 ;
        RECT 3508.010 3950.950 3508.290 3951.230 ;
        RECT 3508.720 3950.950 3509.000 3951.230 ;
        RECT 3509.430 3950.950 3509.710 3951.230 ;
        RECT 3500.200 3950.240 3500.480 3950.520 ;
        RECT 3500.910 3950.240 3501.190 3950.520 ;
        RECT 3501.620 3950.240 3501.900 3950.520 ;
        RECT 3502.330 3950.240 3502.610 3950.520 ;
        RECT 3503.040 3950.240 3503.320 3950.520 ;
        RECT 3503.750 3950.240 3504.030 3950.520 ;
        RECT 3504.460 3950.240 3504.740 3950.520 ;
        RECT 3505.170 3950.240 3505.450 3950.520 ;
        RECT 3505.880 3950.240 3506.160 3950.520 ;
        RECT 3506.590 3950.240 3506.870 3950.520 ;
        RECT 3507.300 3950.240 3507.580 3950.520 ;
        RECT 3508.010 3950.240 3508.290 3950.520 ;
        RECT 3508.720 3950.240 3509.000 3950.520 ;
        RECT 3509.430 3950.240 3509.710 3950.520 ;
        RECT 3500.200 3949.530 3500.480 3949.810 ;
        RECT 3500.910 3949.530 3501.190 3949.810 ;
        RECT 3501.620 3949.530 3501.900 3949.810 ;
        RECT 3502.330 3949.530 3502.610 3949.810 ;
        RECT 3503.040 3949.530 3503.320 3949.810 ;
        RECT 3503.750 3949.530 3504.030 3949.810 ;
        RECT 3504.460 3949.530 3504.740 3949.810 ;
        RECT 3505.170 3949.530 3505.450 3949.810 ;
        RECT 3505.880 3949.530 3506.160 3949.810 ;
        RECT 3506.590 3949.530 3506.870 3949.810 ;
        RECT 3507.300 3949.530 3507.580 3949.810 ;
        RECT 3508.010 3949.530 3508.290 3949.810 ;
        RECT 3508.720 3949.530 3509.000 3949.810 ;
        RECT 3509.430 3949.530 3509.710 3949.810 ;
        RECT 357.275 3945.185 357.555 3945.465 ;
        RECT 357.985 3945.185 358.265 3945.465 ;
        RECT 358.695 3945.185 358.975 3945.465 ;
        RECT 359.405 3945.185 359.685 3945.465 ;
        RECT 360.115 3945.185 360.395 3945.465 ;
        RECT 360.825 3945.185 361.105 3945.465 ;
        RECT 361.535 3945.185 361.815 3945.465 ;
        RECT 362.245 3945.185 362.525 3945.465 ;
        RECT 362.955 3945.185 363.235 3945.465 ;
        RECT 363.665 3945.185 363.945 3945.465 ;
        RECT 364.375 3945.185 364.655 3945.465 ;
        RECT 365.085 3945.185 365.365 3945.465 ;
        RECT 365.795 3945.185 366.075 3945.465 ;
        RECT 366.505 3945.185 366.785 3945.465 ;
        RECT 357.275 3944.475 357.555 3944.755 ;
        RECT 357.985 3944.475 358.265 3944.755 ;
        RECT 358.695 3944.475 358.975 3944.755 ;
        RECT 359.405 3944.475 359.685 3944.755 ;
        RECT 360.115 3944.475 360.395 3944.755 ;
        RECT 360.825 3944.475 361.105 3944.755 ;
        RECT 361.535 3944.475 361.815 3944.755 ;
        RECT 362.245 3944.475 362.525 3944.755 ;
        RECT 362.955 3944.475 363.235 3944.755 ;
        RECT 363.665 3944.475 363.945 3944.755 ;
        RECT 364.375 3944.475 364.655 3944.755 ;
        RECT 365.085 3944.475 365.365 3944.755 ;
        RECT 365.795 3944.475 366.075 3944.755 ;
        RECT 366.505 3944.475 366.785 3944.755 ;
        RECT 357.275 3943.765 357.555 3944.045 ;
        RECT 357.985 3943.765 358.265 3944.045 ;
        RECT 358.695 3943.765 358.975 3944.045 ;
        RECT 359.405 3943.765 359.685 3944.045 ;
        RECT 360.115 3943.765 360.395 3944.045 ;
        RECT 360.825 3943.765 361.105 3944.045 ;
        RECT 361.535 3943.765 361.815 3944.045 ;
        RECT 362.245 3943.765 362.525 3944.045 ;
        RECT 362.955 3943.765 363.235 3944.045 ;
        RECT 363.665 3943.765 363.945 3944.045 ;
        RECT 364.375 3943.765 364.655 3944.045 ;
        RECT 365.085 3943.765 365.365 3944.045 ;
        RECT 365.795 3943.765 366.075 3944.045 ;
        RECT 366.505 3943.765 366.785 3944.045 ;
        RECT 357.275 3943.055 357.555 3943.335 ;
        RECT 357.985 3943.055 358.265 3943.335 ;
        RECT 358.695 3943.055 358.975 3943.335 ;
        RECT 359.405 3943.055 359.685 3943.335 ;
        RECT 360.115 3943.055 360.395 3943.335 ;
        RECT 360.825 3943.055 361.105 3943.335 ;
        RECT 361.535 3943.055 361.815 3943.335 ;
        RECT 362.245 3943.055 362.525 3943.335 ;
        RECT 362.955 3943.055 363.235 3943.335 ;
        RECT 363.665 3943.055 363.945 3943.335 ;
        RECT 364.375 3943.055 364.655 3943.335 ;
        RECT 365.085 3943.055 365.365 3943.335 ;
        RECT 365.795 3943.055 366.075 3943.335 ;
        RECT 366.505 3943.055 366.785 3943.335 ;
        RECT 357.275 3942.345 357.555 3942.625 ;
        RECT 357.985 3942.345 358.265 3942.625 ;
        RECT 358.695 3942.345 358.975 3942.625 ;
        RECT 359.405 3942.345 359.685 3942.625 ;
        RECT 360.115 3942.345 360.395 3942.625 ;
        RECT 360.825 3942.345 361.105 3942.625 ;
        RECT 361.535 3942.345 361.815 3942.625 ;
        RECT 362.245 3942.345 362.525 3942.625 ;
        RECT 362.955 3942.345 363.235 3942.625 ;
        RECT 363.665 3942.345 363.945 3942.625 ;
        RECT 364.375 3942.345 364.655 3942.625 ;
        RECT 365.085 3942.345 365.365 3942.625 ;
        RECT 365.795 3942.345 366.075 3942.625 ;
        RECT 366.505 3942.345 366.785 3942.625 ;
        RECT 357.275 3941.635 357.555 3941.915 ;
        RECT 357.985 3941.635 358.265 3941.915 ;
        RECT 358.695 3941.635 358.975 3941.915 ;
        RECT 359.405 3941.635 359.685 3941.915 ;
        RECT 360.115 3941.635 360.395 3941.915 ;
        RECT 360.825 3941.635 361.105 3941.915 ;
        RECT 361.535 3941.635 361.815 3941.915 ;
        RECT 362.245 3941.635 362.525 3941.915 ;
        RECT 362.955 3941.635 363.235 3941.915 ;
        RECT 363.665 3941.635 363.945 3941.915 ;
        RECT 364.375 3941.635 364.655 3941.915 ;
        RECT 365.085 3941.635 365.365 3941.915 ;
        RECT 365.795 3941.635 366.075 3941.915 ;
        RECT 366.505 3941.635 366.785 3941.915 ;
        RECT 357.275 3940.925 357.555 3941.205 ;
        RECT 357.985 3940.925 358.265 3941.205 ;
        RECT 358.695 3940.925 358.975 3941.205 ;
        RECT 359.405 3940.925 359.685 3941.205 ;
        RECT 360.115 3940.925 360.395 3941.205 ;
        RECT 360.825 3940.925 361.105 3941.205 ;
        RECT 361.535 3940.925 361.815 3941.205 ;
        RECT 362.245 3940.925 362.525 3941.205 ;
        RECT 362.955 3940.925 363.235 3941.205 ;
        RECT 363.665 3940.925 363.945 3941.205 ;
        RECT 364.375 3940.925 364.655 3941.205 ;
        RECT 365.085 3940.925 365.365 3941.205 ;
        RECT 365.795 3940.925 366.075 3941.205 ;
        RECT 366.505 3940.925 366.785 3941.205 ;
        RECT 357.275 3940.215 357.555 3940.495 ;
        RECT 357.985 3940.215 358.265 3940.495 ;
        RECT 358.695 3940.215 358.975 3940.495 ;
        RECT 359.405 3940.215 359.685 3940.495 ;
        RECT 360.115 3940.215 360.395 3940.495 ;
        RECT 360.825 3940.215 361.105 3940.495 ;
        RECT 361.535 3940.215 361.815 3940.495 ;
        RECT 362.245 3940.215 362.525 3940.495 ;
        RECT 362.955 3940.215 363.235 3940.495 ;
        RECT 363.665 3940.215 363.945 3940.495 ;
        RECT 364.375 3940.215 364.655 3940.495 ;
        RECT 365.085 3940.215 365.365 3940.495 ;
        RECT 365.795 3940.215 366.075 3940.495 ;
        RECT 366.505 3940.215 366.785 3940.495 ;
        RECT 357.275 3939.505 357.555 3939.785 ;
        RECT 357.985 3939.505 358.265 3939.785 ;
        RECT 358.695 3939.505 358.975 3939.785 ;
        RECT 359.405 3939.505 359.685 3939.785 ;
        RECT 360.115 3939.505 360.395 3939.785 ;
        RECT 360.825 3939.505 361.105 3939.785 ;
        RECT 361.535 3939.505 361.815 3939.785 ;
        RECT 362.245 3939.505 362.525 3939.785 ;
        RECT 362.955 3939.505 363.235 3939.785 ;
        RECT 363.665 3939.505 363.945 3939.785 ;
        RECT 364.375 3939.505 364.655 3939.785 ;
        RECT 365.085 3939.505 365.365 3939.785 ;
        RECT 365.795 3939.505 366.075 3939.785 ;
        RECT 366.505 3939.505 366.785 3939.785 ;
        RECT 357.275 3938.795 357.555 3939.075 ;
        RECT 357.985 3938.795 358.265 3939.075 ;
        RECT 358.695 3938.795 358.975 3939.075 ;
        RECT 359.405 3938.795 359.685 3939.075 ;
        RECT 360.115 3938.795 360.395 3939.075 ;
        RECT 360.825 3938.795 361.105 3939.075 ;
        RECT 361.535 3938.795 361.815 3939.075 ;
        RECT 362.245 3938.795 362.525 3939.075 ;
        RECT 362.955 3938.795 363.235 3939.075 ;
        RECT 363.665 3938.795 363.945 3939.075 ;
        RECT 364.375 3938.795 364.655 3939.075 ;
        RECT 365.085 3938.795 365.365 3939.075 ;
        RECT 365.795 3938.795 366.075 3939.075 ;
        RECT 366.505 3938.795 366.785 3939.075 ;
        RECT 357.275 3938.085 357.555 3938.365 ;
        RECT 357.985 3938.085 358.265 3938.365 ;
        RECT 358.695 3938.085 358.975 3938.365 ;
        RECT 359.405 3938.085 359.685 3938.365 ;
        RECT 360.115 3938.085 360.395 3938.365 ;
        RECT 360.825 3938.085 361.105 3938.365 ;
        RECT 361.535 3938.085 361.815 3938.365 ;
        RECT 362.245 3938.085 362.525 3938.365 ;
        RECT 362.955 3938.085 363.235 3938.365 ;
        RECT 363.665 3938.085 363.945 3938.365 ;
        RECT 364.375 3938.085 364.655 3938.365 ;
        RECT 365.085 3938.085 365.365 3938.365 ;
        RECT 365.795 3938.085 366.075 3938.365 ;
        RECT 366.505 3938.085 366.785 3938.365 ;
        RECT 357.275 3937.375 357.555 3937.655 ;
        RECT 357.985 3937.375 358.265 3937.655 ;
        RECT 358.695 3937.375 358.975 3937.655 ;
        RECT 359.405 3937.375 359.685 3937.655 ;
        RECT 360.115 3937.375 360.395 3937.655 ;
        RECT 360.825 3937.375 361.105 3937.655 ;
        RECT 361.535 3937.375 361.815 3937.655 ;
        RECT 362.245 3937.375 362.525 3937.655 ;
        RECT 362.955 3937.375 363.235 3937.655 ;
        RECT 363.665 3937.375 363.945 3937.655 ;
        RECT 364.375 3937.375 364.655 3937.655 ;
        RECT 365.085 3937.375 365.365 3937.655 ;
        RECT 365.795 3937.375 366.075 3937.655 ;
        RECT 366.505 3937.375 366.785 3937.655 ;
        RECT 357.275 3936.665 357.555 3936.945 ;
        RECT 357.985 3936.665 358.265 3936.945 ;
        RECT 358.695 3936.665 358.975 3936.945 ;
        RECT 359.405 3936.665 359.685 3936.945 ;
        RECT 360.115 3936.665 360.395 3936.945 ;
        RECT 360.825 3936.665 361.105 3936.945 ;
        RECT 361.535 3936.665 361.815 3936.945 ;
        RECT 362.245 3936.665 362.525 3936.945 ;
        RECT 362.955 3936.665 363.235 3936.945 ;
        RECT 363.665 3936.665 363.945 3936.945 ;
        RECT 364.375 3936.665 364.655 3936.945 ;
        RECT 365.085 3936.665 365.365 3936.945 ;
        RECT 365.795 3936.665 366.075 3936.945 ;
        RECT 366.505 3936.665 366.785 3936.945 ;
        RECT 357.275 3935.955 357.555 3936.235 ;
        RECT 357.985 3935.955 358.265 3936.235 ;
        RECT 358.695 3935.955 358.975 3936.235 ;
        RECT 359.405 3935.955 359.685 3936.235 ;
        RECT 360.115 3935.955 360.395 3936.235 ;
        RECT 360.825 3935.955 361.105 3936.235 ;
        RECT 361.535 3935.955 361.815 3936.235 ;
        RECT 362.245 3935.955 362.525 3936.235 ;
        RECT 362.955 3935.955 363.235 3936.235 ;
        RECT 363.665 3935.955 363.945 3936.235 ;
        RECT 364.375 3935.955 364.655 3936.235 ;
        RECT 365.085 3935.955 365.365 3936.235 ;
        RECT 365.795 3935.955 366.075 3936.235 ;
        RECT 366.505 3935.955 366.785 3936.235 ;
        RECT 3500.255 3945.615 3500.535 3945.895 ;
        RECT 3500.965 3945.615 3501.245 3945.895 ;
        RECT 3501.675 3945.615 3501.955 3945.895 ;
        RECT 3502.385 3945.615 3502.665 3945.895 ;
        RECT 3503.095 3945.615 3503.375 3945.895 ;
        RECT 3503.805 3945.615 3504.085 3945.895 ;
        RECT 3504.515 3945.615 3504.795 3945.895 ;
        RECT 3505.225 3945.615 3505.505 3945.895 ;
        RECT 3505.935 3945.615 3506.215 3945.895 ;
        RECT 3506.645 3945.615 3506.925 3945.895 ;
        RECT 3507.355 3945.615 3507.635 3945.895 ;
        RECT 3508.065 3945.615 3508.345 3945.895 ;
        RECT 3508.775 3945.615 3509.055 3945.895 ;
        RECT 3509.485 3945.615 3509.765 3945.895 ;
        RECT 3500.255 3944.905 3500.535 3945.185 ;
        RECT 3500.965 3944.905 3501.245 3945.185 ;
        RECT 3501.675 3944.905 3501.955 3945.185 ;
        RECT 3502.385 3944.905 3502.665 3945.185 ;
        RECT 3503.095 3944.905 3503.375 3945.185 ;
        RECT 3503.805 3944.905 3504.085 3945.185 ;
        RECT 3504.515 3944.905 3504.795 3945.185 ;
        RECT 3505.225 3944.905 3505.505 3945.185 ;
        RECT 3505.935 3944.905 3506.215 3945.185 ;
        RECT 3506.645 3944.905 3506.925 3945.185 ;
        RECT 3507.355 3944.905 3507.635 3945.185 ;
        RECT 3508.065 3944.905 3508.345 3945.185 ;
        RECT 3508.775 3944.905 3509.055 3945.185 ;
        RECT 3509.485 3944.905 3509.765 3945.185 ;
        RECT 3500.255 3944.195 3500.535 3944.475 ;
        RECT 3500.965 3944.195 3501.245 3944.475 ;
        RECT 3501.675 3944.195 3501.955 3944.475 ;
        RECT 3502.385 3944.195 3502.665 3944.475 ;
        RECT 3503.095 3944.195 3503.375 3944.475 ;
        RECT 3503.805 3944.195 3504.085 3944.475 ;
        RECT 3504.515 3944.195 3504.795 3944.475 ;
        RECT 3505.225 3944.195 3505.505 3944.475 ;
        RECT 3505.935 3944.195 3506.215 3944.475 ;
        RECT 3506.645 3944.195 3506.925 3944.475 ;
        RECT 3507.355 3944.195 3507.635 3944.475 ;
        RECT 3508.065 3944.195 3508.345 3944.475 ;
        RECT 3508.775 3944.195 3509.055 3944.475 ;
        RECT 3509.485 3944.195 3509.765 3944.475 ;
        RECT 3500.255 3943.485 3500.535 3943.765 ;
        RECT 3500.965 3943.485 3501.245 3943.765 ;
        RECT 3501.675 3943.485 3501.955 3943.765 ;
        RECT 3502.385 3943.485 3502.665 3943.765 ;
        RECT 3503.095 3943.485 3503.375 3943.765 ;
        RECT 3503.805 3943.485 3504.085 3943.765 ;
        RECT 3504.515 3943.485 3504.795 3943.765 ;
        RECT 3505.225 3943.485 3505.505 3943.765 ;
        RECT 3505.935 3943.485 3506.215 3943.765 ;
        RECT 3506.645 3943.485 3506.925 3943.765 ;
        RECT 3507.355 3943.485 3507.635 3943.765 ;
        RECT 3508.065 3943.485 3508.345 3943.765 ;
        RECT 3508.775 3943.485 3509.055 3943.765 ;
        RECT 3509.485 3943.485 3509.765 3943.765 ;
        RECT 3500.255 3942.775 3500.535 3943.055 ;
        RECT 3500.965 3942.775 3501.245 3943.055 ;
        RECT 3501.675 3942.775 3501.955 3943.055 ;
        RECT 3502.385 3942.775 3502.665 3943.055 ;
        RECT 3503.095 3942.775 3503.375 3943.055 ;
        RECT 3503.805 3942.775 3504.085 3943.055 ;
        RECT 3504.515 3942.775 3504.795 3943.055 ;
        RECT 3505.225 3942.775 3505.505 3943.055 ;
        RECT 3505.935 3942.775 3506.215 3943.055 ;
        RECT 3506.645 3942.775 3506.925 3943.055 ;
        RECT 3507.355 3942.775 3507.635 3943.055 ;
        RECT 3508.065 3942.775 3508.345 3943.055 ;
        RECT 3508.775 3942.775 3509.055 3943.055 ;
        RECT 3509.485 3942.775 3509.765 3943.055 ;
        RECT 3500.255 3942.065 3500.535 3942.345 ;
        RECT 3500.965 3942.065 3501.245 3942.345 ;
        RECT 3501.675 3942.065 3501.955 3942.345 ;
        RECT 3502.385 3942.065 3502.665 3942.345 ;
        RECT 3503.095 3942.065 3503.375 3942.345 ;
        RECT 3503.805 3942.065 3504.085 3942.345 ;
        RECT 3504.515 3942.065 3504.795 3942.345 ;
        RECT 3505.225 3942.065 3505.505 3942.345 ;
        RECT 3505.935 3942.065 3506.215 3942.345 ;
        RECT 3506.645 3942.065 3506.925 3942.345 ;
        RECT 3507.355 3942.065 3507.635 3942.345 ;
        RECT 3508.065 3942.065 3508.345 3942.345 ;
        RECT 3508.775 3942.065 3509.055 3942.345 ;
        RECT 3509.485 3942.065 3509.765 3942.345 ;
        RECT 3500.255 3941.355 3500.535 3941.635 ;
        RECT 3500.965 3941.355 3501.245 3941.635 ;
        RECT 3501.675 3941.355 3501.955 3941.635 ;
        RECT 3502.385 3941.355 3502.665 3941.635 ;
        RECT 3503.095 3941.355 3503.375 3941.635 ;
        RECT 3503.805 3941.355 3504.085 3941.635 ;
        RECT 3504.515 3941.355 3504.795 3941.635 ;
        RECT 3505.225 3941.355 3505.505 3941.635 ;
        RECT 3505.935 3941.355 3506.215 3941.635 ;
        RECT 3506.645 3941.355 3506.925 3941.635 ;
        RECT 3507.355 3941.355 3507.635 3941.635 ;
        RECT 3508.065 3941.355 3508.345 3941.635 ;
        RECT 3508.775 3941.355 3509.055 3941.635 ;
        RECT 3509.485 3941.355 3509.765 3941.635 ;
        RECT 3500.255 3940.645 3500.535 3940.925 ;
        RECT 3500.965 3940.645 3501.245 3940.925 ;
        RECT 3501.675 3940.645 3501.955 3940.925 ;
        RECT 3502.385 3940.645 3502.665 3940.925 ;
        RECT 3503.095 3940.645 3503.375 3940.925 ;
        RECT 3503.805 3940.645 3504.085 3940.925 ;
        RECT 3504.515 3940.645 3504.795 3940.925 ;
        RECT 3505.225 3940.645 3505.505 3940.925 ;
        RECT 3505.935 3940.645 3506.215 3940.925 ;
        RECT 3506.645 3940.645 3506.925 3940.925 ;
        RECT 3507.355 3940.645 3507.635 3940.925 ;
        RECT 3508.065 3940.645 3508.345 3940.925 ;
        RECT 3508.775 3940.645 3509.055 3940.925 ;
        RECT 3509.485 3940.645 3509.765 3940.925 ;
        RECT 3500.255 3939.935 3500.535 3940.215 ;
        RECT 3500.965 3939.935 3501.245 3940.215 ;
        RECT 3501.675 3939.935 3501.955 3940.215 ;
        RECT 3502.385 3939.935 3502.665 3940.215 ;
        RECT 3503.095 3939.935 3503.375 3940.215 ;
        RECT 3503.805 3939.935 3504.085 3940.215 ;
        RECT 3504.515 3939.935 3504.795 3940.215 ;
        RECT 3505.225 3939.935 3505.505 3940.215 ;
        RECT 3505.935 3939.935 3506.215 3940.215 ;
        RECT 3506.645 3939.935 3506.925 3940.215 ;
        RECT 3507.355 3939.935 3507.635 3940.215 ;
        RECT 3508.065 3939.935 3508.345 3940.215 ;
        RECT 3508.775 3939.935 3509.055 3940.215 ;
        RECT 3509.485 3939.935 3509.765 3940.215 ;
        RECT 3500.255 3939.225 3500.535 3939.505 ;
        RECT 3500.965 3939.225 3501.245 3939.505 ;
        RECT 3501.675 3939.225 3501.955 3939.505 ;
        RECT 3502.385 3939.225 3502.665 3939.505 ;
        RECT 3503.095 3939.225 3503.375 3939.505 ;
        RECT 3503.805 3939.225 3504.085 3939.505 ;
        RECT 3504.515 3939.225 3504.795 3939.505 ;
        RECT 3505.225 3939.225 3505.505 3939.505 ;
        RECT 3505.935 3939.225 3506.215 3939.505 ;
        RECT 3506.645 3939.225 3506.925 3939.505 ;
        RECT 3507.355 3939.225 3507.635 3939.505 ;
        RECT 3508.065 3939.225 3508.345 3939.505 ;
        RECT 3508.775 3939.225 3509.055 3939.505 ;
        RECT 3509.485 3939.225 3509.765 3939.505 ;
        RECT 3500.255 3938.515 3500.535 3938.795 ;
        RECT 3500.965 3938.515 3501.245 3938.795 ;
        RECT 3501.675 3938.515 3501.955 3938.795 ;
        RECT 3502.385 3938.515 3502.665 3938.795 ;
        RECT 3503.095 3938.515 3503.375 3938.795 ;
        RECT 3503.805 3938.515 3504.085 3938.795 ;
        RECT 3504.515 3938.515 3504.795 3938.795 ;
        RECT 3505.225 3938.515 3505.505 3938.795 ;
        RECT 3505.935 3938.515 3506.215 3938.795 ;
        RECT 3506.645 3938.515 3506.925 3938.795 ;
        RECT 3507.355 3938.515 3507.635 3938.795 ;
        RECT 3508.065 3938.515 3508.345 3938.795 ;
        RECT 3508.775 3938.515 3509.055 3938.795 ;
        RECT 3509.485 3938.515 3509.765 3938.795 ;
        RECT 3500.255 3937.805 3500.535 3938.085 ;
        RECT 3500.965 3937.805 3501.245 3938.085 ;
        RECT 3501.675 3937.805 3501.955 3938.085 ;
        RECT 3502.385 3937.805 3502.665 3938.085 ;
        RECT 3503.095 3937.805 3503.375 3938.085 ;
        RECT 3503.805 3937.805 3504.085 3938.085 ;
        RECT 3504.515 3937.805 3504.795 3938.085 ;
        RECT 3505.225 3937.805 3505.505 3938.085 ;
        RECT 3505.935 3937.805 3506.215 3938.085 ;
        RECT 3506.645 3937.805 3506.925 3938.085 ;
        RECT 3507.355 3937.805 3507.635 3938.085 ;
        RECT 3508.065 3937.805 3508.345 3938.085 ;
        RECT 3508.775 3937.805 3509.055 3938.085 ;
        RECT 3509.485 3937.805 3509.765 3938.085 ;
        RECT 3500.255 3937.095 3500.535 3937.375 ;
        RECT 3500.965 3937.095 3501.245 3937.375 ;
        RECT 3501.675 3937.095 3501.955 3937.375 ;
        RECT 3502.385 3937.095 3502.665 3937.375 ;
        RECT 3503.095 3937.095 3503.375 3937.375 ;
        RECT 3503.805 3937.095 3504.085 3937.375 ;
        RECT 3504.515 3937.095 3504.795 3937.375 ;
        RECT 3505.225 3937.095 3505.505 3937.375 ;
        RECT 3505.935 3937.095 3506.215 3937.375 ;
        RECT 3506.645 3937.095 3506.925 3937.375 ;
        RECT 3507.355 3937.095 3507.635 3937.375 ;
        RECT 3508.065 3937.095 3508.345 3937.375 ;
        RECT 3508.775 3937.095 3509.055 3937.375 ;
        RECT 3509.485 3937.095 3509.765 3937.375 ;
        RECT 3500.255 3936.385 3500.535 3936.665 ;
        RECT 3500.965 3936.385 3501.245 3936.665 ;
        RECT 3501.675 3936.385 3501.955 3936.665 ;
        RECT 3502.385 3936.385 3502.665 3936.665 ;
        RECT 3503.095 3936.385 3503.375 3936.665 ;
        RECT 3503.805 3936.385 3504.085 3936.665 ;
        RECT 3504.515 3936.385 3504.795 3936.665 ;
        RECT 3505.225 3936.385 3505.505 3936.665 ;
        RECT 3505.935 3936.385 3506.215 3936.665 ;
        RECT 3506.645 3936.385 3506.925 3936.665 ;
        RECT 3507.355 3936.385 3507.635 3936.665 ;
        RECT 3508.065 3936.385 3508.345 3936.665 ;
        RECT 3508.775 3936.385 3509.055 3936.665 ;
        RECT 3509.485 3936.385 3509.765 3936.665 ;
        RECT 357.275 3933.335 357.555 3933.615 ;
        RECT 357.985 3933.335 358.265 3933.615 ;
        RECT 358.695 3933.335 358.975 3933.615 ;
        RECT 359.405 3933.335 359.685 3933.615 ;
        RECT 360.115 3933.335 360.395 3933.615 ;
        RECT 360.825 3933.335 361.105 3933.615 ;
        RECT 361.535 3933.335 361.815 3933.615 ;
        RECT 362.245 3933.335 362.525 3933.615 ;
        RECT 362.955 3933.335 363.235 3933.615 ;
        RECT 363.665 3933.335 363.945 3933.615 ;
        RECT 364.375 3933.335 364.655 3933.615 ;
        RECT 365.085 3933.335 365.365 3933.615 ;
        RECT 365.795 3933.335 366.075 3933.615 ;
        RECT 366.505 3933.335 366.785 3933.615 ;
        RECT 357.275 3932.625 357.555 3932.905 ;
        RECT 357.985 3932.625 358.265 3932.905 ;
        RECT 358.695 3932.625 358.975 3932.905 ;
        RECT 359.405 3932.625 359.685 3932.905 ;
        RECT 360.115 3932.625 360.395 3932.905 ;
        RECT 360.825 3932.625 361.105 3932.905 ;
        RECT 361.535 3932.625 361.815 3932.905 ;
        RECT 362.245 3932.625 362.525 3932.905 ;
        RECT 362.955 3932.625 363.235 3932.905 ;
        RECT 363.665 3932.625 363.945 3932.905 ;
        RECT 364.375 3932.625 364.655 3932.905 ;
        RECT 365.085 3932.625 365.365 3932.905 ;
        RECT 365.795 3932.625 366.075 3932.905 ;
        RECT 366.505 3932.625 366.785 3932.905 ;
        RECT 357.275 3931.915 357.555 3932.195 ;
        RECT 357.985 3931.915 358.265 3932.195 ;
        RECT 358.695 3931.915 358.975 3932.195 ;
        RECT 359.405 3931.915 359.685 3932.195 ;
        RECT 360.115 3931.915 360.395 3932.195 ;
        RECT 360.825 3931.915 361.105 3932.195 ;
        RECT 361.535 3931.915 361.815 3932.195 ;
        RECT 362.245 3931.915 362.525 3932.195 ;
        RECT 362.955 3931.915 363.235 3932.195 ;
        RECT 363.665 3931.915 363.945 3932.195 ;
        RECT 364.375 3931.915 364.655 3932.195 ;
        RECT 365.085 3931.915 365.365 3932.195 ;
        RECT 365.795 3931.915 366.075 3932.195 ;
        RECT 366.505 3931.915 366.785 3932.195 ;
        RECT 357.275 3931.205 357.555 3931.485 ;
        RECT 357.985 3931.205 358.265 3931.485 ;
        RECT 358.695 3931.205 358.975 3931.485 ;
        RECT 359.405 3931.205 359.685 3931.485 ;
        RECT 360.115 3931.205 360.395 3931.485 ;
        RECT 360.825 3931.205 361.105 3931.485 ;
        RECT 361.535 3931.205 361.815 3931.485 ;
        RECT 362.245 3931.205 362.525 3931.485 ;
        RECT 362.955 3931.205 363.235 3931.485 ;
        RECT 363.665 3931.205 363.945 3931.485 ;
        RECT 364.375 3931.205 364.655 3931.485 ;
        RECT 365.085 3931.205 365.365 3931.485 ;
        RECT 365.795 3931.205 366.075 3931.485 ;
        RECT 366.505 3931.205 366.785 3931.485 ;
        RECT 357.275 3930.495 357.555 3930.775 ;
        RECT 357.985 3930.495 358.265 3930.775 ;
        RECT 358.695 3930.495 358.975 3930.775 ;
        RECT 359.405 3930.495 359.685 3930.775 ;
        RECT 360.115 3930.495 360.395 3930.775 ;
        RECT 360.825 3930.495 361.105 3930.775 ;
        RECT 361.535 3930.495 361.815 3930.775 ;
        RECT 362.245 3930.495 362.525 3930.775 ;
        RECT 362.955 3930.495 363.235 3930.775 ;
        RECT 363.665 3930.495 363.945 3930.775 ;
        RECT 364.375 3930.495 364.655 3930.775 ;
        RECT 365.085 3930.495 365.365 3930.775 ;
        RECT 365.795 3930.495 366.075 3930.775 ;
        RECT 366.505 3930.495 366.785 3930.775 ;
        RECT 357.275 3929.785 357.555 3930.065 ;
        RECT 357.985 3929.785 358.265 3930.065 ;
        RECT 358.695 3929.785 358.975 3930.065 ;
        RECT 359.405 3929.785 359.685 3930.065 ;
        RECT 360.115 3929.785 360.395 3930.065 ;
        RECT 360.825 3929.785 361.105 3930.065 ;
        RECT 361.535 3929.785 361.815 3930.065 ;
        RECT 362.245 3929.785 362.525 3930.065 ;
        RECT 362.955 3929.785 363.235 3930.065 ;
        RECT 363.665 3929.785 363.945 3930.065 ;
        RECT 364.375 3929.785 364.655 3930.065 ;
        RECT 365.085 3929.785 365.365 3930.065 ;
        RECT 365.795 3929.785 366.075 3930.065 ;
        RECT 366.505 3929.785 366.785 3930.065 ;
        RECT 357.275 3929.075 357.555 3929.355 ;
        RECT 357.985 3929.075 358.265 3929.355 ;
        RECT 358.695 3929.075 358.975 3929.355 ;
        RECT 359.405 3929.075 359.685 3929.355 ;
        RECT 360.115 3929.075 360.395 3929.355 ;
        RECT 360.825 3929.075 361.105 3929.355 ;
        RECT 361.535 3929.075 361.815 3929.355 ;
        RECT 362.245 3929.075 362.525 3929.355 ;
        RECT 362.955 3929.075 363.235 3929.355 ;
        RECT 363.665 3929.075 363.945 3929.355 ;
        RECT 364.375 3929.075 364.655 3929.355 ;
        RECT 365.085 3929.075 365.365 3929.355 ;
        RECT 365.795 3929.075 366.075 3929.355 ;
        RECT 366.505 3929.075 366.785 3929.355 ;
        RECT 357.275 3928.365 357.555 3928.645 ;
        RECT 357.985 3928.365 358.265 3928.645 ;
        RECT 358.695 3928.365 358.975 3928.645 ;
        RECT 359.405 3928.365 359.685 3928.645 ;
        RECT 360.115 3928.365 360.395 3928.645 ;
        RECT 360.825 3928.365 361.105 3928.645 ;
        RECT 361.535 3928.365 361.815 3928.645 ;
        RECT 362.245 3928.365 362.525 3928.645 ;
        RECT 362.955 3928.365 363.235 3928.645 ;
        RECT 363.665 3928.365 363.945 3928.645 ;
        RECT 364.375 3928.365 364.655 3928.645 ;
        RECT 365.085 3928.365 365.365 3928.645 ;
        RECT 365.795 3928.365 366.075 3928.645 ;
        RECT 366.505 3928.365 366.785 3928.645 ;
        RECT 357.275 3927.655 357.555 3927.935 ;
        RECT 357.985 3927.655 358.265 3927.935 ;
        RECT 358.695 3927.655 358.975 3927.935 ;
        RECT 359.405 3927.655 359.685 3927.935 ;
        RECT 360.115 3927.655 360.395 3927.935 ;
        RECT 360.825 3927.655 361.105 3927.935 ;
        RECT 361.535 3927.655 361.815 3927.935 ;
        RECT 362.245 3927.655 362.525 3927.935 ;
        RECT 362.955 3927.655 363.235 3927.935 ;
        RECT 363.665 3927.655 363.945 3927.935 ;
        RECT 364.375 3927.655 364.655 3927.935 ;
        RECT 365.085 3927.655 365.365 3927.935 ;
        RECT 365.795 3927.655 366.075 3927.935 ;
        RECT 366.505 3927.655 366.785 3927.935 ;
        RECT 357.275 3926.945 357.555 3927.225 ;
        RECT 357.985 3926.945 358.265 3927.225 ;
        RECT 358.695 3926.945 358.975 3927.225 ;
        RECT 359.405 3926.945 359.685 3927.225 ;
        RECT 360.115 3926.945 360.395 3927.225 ;
        RECT 360.825 3926.945 361.105 3927.225 ;
        RECT 361.535 3926.945 361.815 3927.225 ;
        RECT 362.245 3926.945 362.525 3927.225 ;
        RECT 362.955 3926.945 363.235 3927.225 ;
        RECT 363.665 3926.945 363.945 3927.225 ;
        RECT 364.375 3926.945 364.655 3927.225 ;
        RECT 365.085 3926.945 365.365 3927.225 ;
        RECT 365.795 3926.945 366.075 3927.225 ;
        RECT 366.505 3926.945 366.785 3927.225 ;
        RECT 357.275 3926.235 357.555 3926.515 ;
        RECT 357.985 3926.235 358.265 3926.515 ;
        RECT 358.695 3926.235 358.975 3926.515 ;
        RECT 359.405 3926.235 359.685 3926.515 ;
        RECT 360.115 3926.235 360.395 3926.515 ;
        RECT 360.825 3926.235 361.105 3926.515 ;
        RECT 361.535 3926.235 361.815 3926.515 ;
        RECT 362.245 3926.235 362.525 3926.515 ;
        RECT 362.955 3926.235 363.235 3926.515 ;
        RECT 363.665 3926.235 363.945 3926.515 ;
        RECT 364.375 3926.235 364.655 3926.515 ;
        RECT 365.085 3926.235 365.365 3926.515 ;
        RECT 365.795 3926.235 366.075 3926.515 ;
        RECT 366.505 3926.235 366.785 3926.515 ;
        RECT 357.275 3925.525 357.555 3925.805 ;
        RECT 357.985 3925.525 358.265 3925.805 ;
        RECT 358.695 3925.525 358.975 3925.805 ;
        RECT 359.405 3925.525 359.685 3925.805 ;
        RECT 360.115 3925.525 360.395 3925.805 ;
        RECT 360.825 3925.525 361.105 3925.805 ;
        RECT 361.535 3925.525 361.815 3925.805 ;
        RECT 362.245 3925.525 362.525 3925.805 ;
        RECT 362.955 3925.525 363.235 3925.805 ;
        RECT 363.665 3925.525 363.945 3925.805 ;
        RECT 364.375 3925.525 364.655 3925.805 ;
        RECT 365.085 3925.525 365.365 3925.805 ;
        RECT 365.795 3925.525 366.075 3925.805 ;
        RECT 366.505 3925.525 366.785 3925.805 ;
        RECT 357.275 3924.815 357.555 3925.095 ;
        RECT 357.985 3924.815 358.265 3925.095 ;
        RECT 358.695 3924.815 358.975 3925.095 ;
        RECT 359.405 3924.815 359.685 3925.095 ;
        RECT 360.115 3924.815 360.395 3925.095 ;
        RECT 360.825 3924.815 361.105 3925.095 ;
        RECT 361.535 3924.815 361.815 3925.095 ;
        RECT 362.245 3924.815 362.525 3925.095 ;
        RECT 362.955 3924.815 363.235 3925.095 ;
        RECT 363.665 3924.815 363.945 3925.095 ;
        RECT 364.375 3924.815 364.655 3925.095 ;
        RECT 365.085 3924.815 365.365 3925.095 ;
        RECT 365.795 3924.815 366.075 3925.095 ;
        RECT 366.505 3924.815 366.785 3925.095 ;
        RECT 357.275 3924.105 357.555 3924.385 ;
        RECT 357.985 3924.105 358.265 3924.385 ;
        RECT 358.695 3924.105 358.975 3924.385 ;
        RECT 359.405 3924.105 359.685 3924.385 ;
        RECT 360.115 3924.105 360.395 3924.385 ;
        RECT 360.825 3924.105 361.105 3924.385 ;
        RECT 361.535 3924.105 361.815 3924.385 ;
        RECT 362.245 3924.105 362.525 3924.385 ;
        RECT 362.955 3924.105 363.235 3924.385 ;
        RECT 363.665 3924.105 363.945 3924.385 ;
        RECT 364.375 3924.105 364.655 3924.385 ;
        RECT 365.085 3924.105 365.365 3924.385 ;
        RECT 365.795 3924.105 366.075 3924.385 ;
        RECT 366.505 3924.105 366.785 3924.385 ;
        RECT 3500.255 3933.765 3500.535 3934.045 ;
        RECT 3500.965 3933.765 3501.245 3934.045 ;
        RECT 3501.675 3933.765 3501.955 3934.045 ;
        RECT 3502.385 3933.765 3502.665 3934.045 ;
        RECT 3503.095 3933.765 3503.375 3934.045 ;
        RECT 3503.805 3933.765 3504.085 3934.045 ;
        RECT 3504.515 3933.765 3504.795 3934.045 ;
        RECT 3505.225 3933.765 3505.505 3934.045 ;
        RECT 3505.935 3933.765 3506.215 3934.045 ;
        RECT 3506.645 3933.765 3506.925 3934.045 ;
        RECT 3507.355 3933.765 3507.635 3934.045 ;
        RECT 3508.065 3933.765 3508.345 3934.045 ;
        RECT 3508.775 3933.765 3509.055 3934.045 ;
        RECT 3509.485 3933.765 3509.765 3934.045 ;
        RECT 3500.255 3933.055 3500.535 3933.335 ;
        RECT 3500.965 3933.055 3501.245 3933.335 ;
        RECT 3501.675 3933.055 3501.955 3933.335 ;
        RECT 3502.385 3933.055 3502.665 3933.335 ;
        RECT 3503.095 3933.055 3503.375 3933.335 ;
        RECT 3503.805 3933.055 3504.085 3933.335 ;
        RECT 3504.515 3933.055 3504.795 3933.335 ;
        RECT 3505.225 3933.055 3505.505 3933.335 ;
        RECT 3505.935 3933.055 3506.215 3933.335 ;
        RECT 3506.645 3933.055 3506.925 3933.335 ;
        RECT 3507.355 3933.055 3507.635 3933.335 ;
        RECT 3508.065 3933.055 3508.345 3933.335 ;
        RECT 3508.775 3933.055 3509.055 3933.335 ;
        RECT 3509.485 3933.055 3509.765 3933.335 ;
        RECT 3500.255 3932.345 3500.535 3932.625 ;
        RECT 3500.965 3932.345 3501.245 3932.625 ;
        RECT 3501.675 3932.345 3501.955 3932.625 ;
        RECT 3502.385 3932.345 3502.665 3932.625 ;
        RECT 3503.095 3932.345 3503.375 3932.625 ;
        RECT 3503.805 3932.345 3504.085 3932.625 ;
        RECT 3504.515 3932.345 3504.795 3932.625 ;
        RECT 3505.225 3932.345 3505.505 3932.625 ;
        RECT 3505.935 3932.345 3506.215 3932.625 ;
        RECT 3506.645 3932.345 3506.925 3932.625 ;
        RECT 3507.355 3932.345 3507.635 3932.625 ;
        RECT 3508.065 3932.345 3508.345 3932.625 ;
        RECT 3508.775 3932.345 3509.055 3932.625 ;
        RECT 3509.485 3932.345 3509.765 3932.625 ;
        RECT 3500.255 3931.635 3500.535 3931.915 ;
        RECT 3500.965 3931.635 3501.245 3931.915 ;
        RECT 3501.675 3931.635 3501.955 3931.915 ;
        RECT 3502.385 3931.635 3502.665 3931.915 ;
        RECT 3503.095 3931.635 3503.375 3931.915 ;
        RECT 3503.805 3931.635 3504.085 3931.915 ;
        RECT 3504.515 3931.635 3504.795 3931.915 ;
        RECT 3505.225 3931.635 3505.505 3931.915 ;
        RECT 3505.935 3931.635 3506.215 3931.915 ;
        RECT 3506.645 3931.635 3506.925 3931.915 ;
        RECT 3507.355 3931.635 3507.635 3931.915 ;
        RECT 3508.065 3931.635 3508.345 3931.915 ;
        RECT 3508.775 3931.635 3509.055 3931.915 ;
        RECT 3509.485 3931.635 3509.765 3931.915 ;
        RECT 3500.255 3930.925 3500.535 3931.205 ;
        RECT 3500.965 3930.925 3501.245 3931.205 ;
        RECT 3501.675 3930.925 3501.955 3931.205 ;
        RECT 3502.385 3930.925 3502.665 3931.205 ;
        RECT 3503.095 3930.925 3503.375 3931.205 ;
        RECT 3503.805 3930.925 3504.085 3931.205 ;
        RECT 3504.515 3930.925 3504.795 3931.205 ;
        RECT 3505.225 3930.925 3505.505 3931.205 ;
        RECT 3505.935 3930.925 3506.215 3931.205 ;
        RECT 3506.645 3930.925 3506.925 3931.205 ;
        RECT 3507.355 3930.925 3507.635 3931.205 ;
        RECT 3508.065 3930.925 3508.345 3931.205 ;
        RECT 3508.775 3930.925 3509.055 3931.205 ;
        RECT 3509.485 3930.925 3509.765 3931.205 ;
        RECT 3500.255 3930.215 3500.535 3930.495 ;
        RECT 3500.965 3930.215 3501.245 3930.495 ;
        RECT 3501.675 3930.215 3501.955 3930.495 ;
        RECT 3502.385 3930.215 3502.665 3930.495 ;
        RECT 3503.095 3930.215 3503.375 3930.495 ;
        RECT 3503.805 3930.215 3504.085 3930.495 ;
        RECT 3504.515 3930.215 3504.795 3930.495 ;
        RECT 3505.225 3930.215 3505.505 3930.495 ;
        RECT 3505.935 3930.215 3506.215 3930.495 ;
        RECT 3506.645 3930.215 3506.925 3930.495 ;
        RECT 3507.355 3930.215 3507.635 3930.495 ;
        RECT 3508.065 3930.215 3508.345 3930.495 ;
        RECT 3508.775 3930.215 3509.055 3930.495 ;
        RECT 3509.485 3930.215 3509.765 3930.495 ;
        RECT 3500.255 3929.505 3500.535 3929.785 ;
        RECT 3500.965 3929.505 3501.245 3929.785 ;
        RECT 3501.675 3929.505 3501.955 3929.785 ;
        RECT 3502.385 3929.505 3502.665 3929.785 ;
        RECT 3503.095 3929.505 3503.375 3929.785 ;
        RECT 3503.805 3929.505 3504.085 3929.785 ;
        RECT 3504.515 3929.505 3504.795 3929.785 ;
        RECT 3505.225 3929.505 3505.505 3929.785 ;
        RECT 3505.935 3929.505 3506.215 3929.785 ;
        RECT 3506.645 3929.505 3506.925 3929.785 ;
        RECT 3507.355 3929.505 3507.635 3929.785 ;
        RECT 3508.065 3929.505 3508.345 3929.785 ;
        RECT 3508.775 3929.505 3509.055 3929.785 ;
        RECT 3509.485 3929.505 3509.765 3929.785 ;
        RECT 3500.255 3928.795 3500.535 3929.075 ;
        RECT 3500.965 3928.795 3501.245 3929.075 ;
        RECT 3501.675 3928.795 3501.955 3929.075 ;
        RECT 3502.385 3928.795 3502.665 3929.075 ;
        RECT 3503.095 3928.795 3503.375 3929.075 ;
        RECT 3503.805 3928.795 3504.085 3929.075 ;
        RECT 3504.515 3928.795 3504.795 3929.075 ;
        RECT 3505.225 3928.795 3505.505 3929.075 ;
        RECT 3505.935 3928.795 3506.215 3929.075 ;
        RECT 3506.645 3928.795 3506.925 3929.075 ;
        RECT 3507.355 3928.795 3507.635 3929.075 ;
        RECT 3508.065 3928.795 3508.345 3929.075 ;
        RECT 3508.775 3928.795 3509.055 3929.075 ;
        RECT 3509.485 3928.795 3509.765 3929.075 ;
        RECT 3500.255 3928.085 3500.535 3928.365 ;
        RECT 3500.965 3928.085 3501.245 3928.365 ;
        RECT 3501.675 3928.085 3501.955 3928.365 ;
        RECT 3502.385 3928.085 3502.665 3928.365 ;
        RECT 3503.095 3928.085 3503.375 3928.365 ;
        RECT 3503.805 3928.085 3504.085 3928.365 ;
        RECT 3504.515 3928.085 3504.795 3928.365 ;
        RECT 3505.225 3928.085 3505.505 3928.365 ;
        RECT 3505.935 3928.085 3506.215 3928.365 ;
        RECT 3506.645 3928.085 3506.925 3928.365 ;
        RECT 3507.355 3928.085 3507.635 3928.365 ;
        RECT 3508.065 3928.085 3508.345 3928.365 ;
        RECT 3508.775 3928.085 3509.055 3928.365 ;
        RECT 3509.485 3928.085 3509.765 3928.365 ;
        RECT 3500.255 3927.375 3500.535 3927.655 ;
        RECT 3500.965 3927.375 3501.245 3927.655 ;
        RECT 3501.675 3927.375 3501.955 3927.655 ;
        RECT 3502.385 3927.375 3502.665 3927.655 ;
        RECT 3503.095 3927.375 3503.375 3927.655 ;
        RECT 3503.805 3927.375 3504.085 3927.655 ;
        RECT 3504.515 3927.375 3504.795 3927.655 ;
        RECT 3505.225 3927.375 3505.505 3927.655 ;
        RECT 3505.935 3927.375 3506.215 3927.655 ;
        RECT 3506.645 3927.375 3506.925 3927.655 ;
        RECT 3507.355 3927.375 3507.635 3927.655 ;
        RECT 3508.065 3927.375 3508.345 3927.655 ;
        RECT 3508.775 3927.375 3509.055 3927.655 ;
        RECT 3509.485 3927.375 3509.765 3927.655 ;
        RECT 3500.255 3926.665 3500.535 3926.945 ;
        RECT 3500.965 3926.665 3501.245 3926.945 ;
        RECT 3501.675 3926.665 3501.955 3926.945 ;
        RECT 3502.385 3926.665 3502.665 3926.945 ;
        RECT 3503.095 3926.665 3503.375 3926.945 ;
        RECT 3503.805 3926.665 3504.085 3926.945 ;
        RECT 3504.515 3926.665 3504.795 3926.945 ;
        RECT 3505.225 3926.665 3505.505 3926.945 ;
        RECT 3505.935 3926.665 3506.215 3926.945 ;
        RECT 3506.645 3926.665 3506.925 3926.945 ;
        RECT 3507.355 3926.665 3507.635 3926.945 ;
        RECT 3508.065 3926.665 3508.345 3926.945 ;
        RECT 3508.775 3926.665 3509.055 3926.945 ;
        RECT 3509.485 3926.665 3509.765 3926.945 ;
        RECT 3500.255 3925.955 3500.535 3926.235 ;
        RECT 3500.965 3925.955 3501.245 3926.235 ;
        RECT 3501.675 3925.955 3501.955 3926.235 ;
        RECT 3502.385 3925.955 3502.665 3926.235 ;
        RECT 3503.095 3925.955 3503.375 3926.235 ;
        RECT 3503.805 3925.955 3504.085 3926.235 ;
        RECT 3504.515 3925.955 3504.795 3926.235 ;
        RECT 3505.225 3925.955 3505.505 3926.235 ;
        RECT 3505.935 3925.955 3506.215 3926.235 ;
        RECT 3506.645 3925.955 3506.925 3926.235 ;
        RECT 3507.355 3925.955 3507.635 3926.235 ;
        RECT 3508.065 3925.955 3508.345 3926.235 ;
        RECT 3508.775 3925.955 3509.055 3926.235 ;
        RECT 3509.485 3925.955 3509.765 3926.235 ;
        RECT 3500.255 3925.245 3500.535 3925.525 ;
        RECT 3500.965 3925.245 3501.245 3925.525 ;
        RECT 3501.675 3925.245 3501.955 3925.525 ;
        RECT 3502.385 3925.245 3502.665 3925.525 ;
        RECT 3503.095 3925.245 3503.375 3925.525 ;
        RECT 3503.805 3925.245 3504.085 3925.525 ;
        RECT 3504.515 3925.245 3504.795 3925.525 ;
        RECT 3505.225 3925.245 3505.505 3925.525 ;
        RECT 3505.935 3925.245 3506.215 3925.525 ;
        RECT 3506.645 3925.245 3506.925 3925.525 ;
        RECT 3507.355 3925.245 3507.635 3925.525 ;
        RECT 3508.065 3925.245 3508.345 3925.525 ;
        RECT 3508.775 3925.245 3509.055 3925.525 ;
        RECT 3509.485 3925.245 3509.765 3925.525 ;
        RECT 3500.255 3924.535 3500.535 3924.815 ;
        RECT 3500.965 3924.535 3501.245 3924.815 ;
        RECT 3501.675 3924.535 3501.955 3924.815 ;
        RECT 3502.385 3924.535 3502.665 3924.815 ;
        RECT 3503.095 3924.535 3503.375 3924.815 ;
        RECT 3503.805 3924.535 3504.085 3924.815 ;
        RECT 3504.515 3924.535 3504.795 3924.815 ;
        RECT 3505.225 3924.535 3505.505 3924.815 ;
        RECT 3505.935 3924.535 3506.215 3924.815 ;
        RECT 3506.645 3924.535 3506.925 3924.815 ;
        RECT 3507.355 3924.535 3507.635 3924.815 ;
        RECT 3508.065 3924.535 3508.345 3924.815 ;
        RECT 3508.775 3924.535 3509.055 3924.815 ;
        RECT 3509.485 3924.535 3509.765 3924.815 ;
        RECT 357.330 3920.190 357.610 3920.470 ;
        RECT 358.040 3920.190 358.320 3920.470 ;
        RECT 358.750 3920.190 359.030 3920.470 ;
        RECT 359.460 3920.190 359.740 3920.470 ;
        RECT 360.170 3920.190 360.450 3920.470 ;
        RECT 360.880 3920.190 361.160 3920.470 ;
        RECT 361.590 3920.190 361.870 3920.470 ;
        RECT 362.300 3920.190 362.580 3920.470 ;
        RECT 363.010 3920.190 363.290 3920.470 ;
        RECT 363.720 3920.190 364.000 3920.470 ;
        RECT 364.430 3920.190 364.710 3920.470 ;
        RECT 365.140 3920.190 365.420 3920.470 ;
        RECT 365.850 3920.190 366.130 3920.470 ;
        RECT 366.560 3920.190 366.840 3920.470 ;
        RECT 357.330 3919.480 357.610 3919.760 ;
        RECT 358.040 3919.480 358.320 3919.760 ;
        RECT 358.750 3919.480 359.030 3919.760 ;
        RECT 359.460 3919.480 359.740 3919.760 ;
        RECT 360.170 3919.480 360.450 3919.760 ;
        RECT 360.880 3919.480 361.160 3919.760 ;
        RECT 361.590 3919.480 361.870 3919.760 ;
        RECT 362.300 3919.480 362.580 3919.760 ;
        RECT 363.010 3919.480 363.290 3919.760 ;
        RECT 363.720 3919.480 364.000 3919.760 ;
        RECT 364.430 3919.480 364.710 3919.760 ;
        RECT 365.140 3919.480 365.420 3919.760 ;
        RECT 365.850 3919.480 366.130 3919.760 ;
        RECT 366.560 3919.480 366.840 3919.760 ;
        RECT 357.330 3918.770 357.610 3919.050 ;
        RECT 358.040 3918.770 358.320 3919.050 ;
        RECT 358.750 3918.770 359.030 3919.050 ;
        RECT 359.460 3918.770 359.740 3919.050 ;
        RECT 360.170 3918.770 360.450 3919.050 ;
        RECT 360.880 3918.770 361.160 3919.050 ;
        RECT 361.590 3918.770 361.870 3919.050 ;
        RECT 362.300 3918.770 362.580 3919.050 ;
        RECT 363.010 3918.770 363.290 3919.050 ;
        RECT 363.720 3918.770 364.000 3919.050 ;
        RECT 364.430 3918.770 364.710 3919.050 ;
        RECT 365.140 3918.770 365.420 3919.050 ;
        RECT 365.850 3918.770 366.130 3919.050 ;
        RECT 366.560 3918.770 366.840 3919.050 ;
        RECT 357.330 3918.060 357.610 3918.340 ;
        RECT 358.040 3918.060 358.320 3918.340 ;
        RECT 358.750 3918.060 359.030 3918.340 ;
        RECT 359.460 3918.060 359.740 3918.340 ;
        RECT 360.170 3918.060 360.450 3918.340 ;
        RECT 360.880 3918.060 361.160 3918.340 ;
        RECT 361.590 3918.060 361.870 3918.340 ;
        RECT 362.300 3918.060 362.580 3918.340 ;
        RECT 363.010 3918.060 363.290 3918.340 ;
        RECT 363.720 3918.060 364.000 3918.340 ;
        RECT 364.430 3918.060 364.710 3918.340 ;
        RECT 365.140 3918.060 365.420 3918.340 ;
        RECT 365.850 3918.060 366.130 3918.340 ;
        RECT 366.560 3918.060 366.840 3918.340 ;
        RECT 357.330 3917.350 357.610 3917.630 ;
        RECT 358.040 3917.350 358.320 3917.630 ;
        RECT 358.750 3917.350 359.030 3917.630 ;
        RECT 359.460 3917.350 359.740 3917.630 ;
        RECT 360.170 3917.350 360.450 3917.630 ;
        RECT 360.880 3917.350 361.160 3917.630 ;
        RECT 361.590 3917.350 361.870 3917.630 ;
        RECT 362.300 3917.350 362.580 3917.630 ;
        RECT 363.010 3917.350 363.290 3917.630 ;
        RECT 363.720 3917.350 364.000 3917.630 ;
        RECT 364.430 3917.350 364.710 3917.630 ;
        RECT 365.140 3917.350 365.420 3917.630 ;
        RECT 365.850 3917.350 366.130 3917.630 ;
        RECT 366.560 3917.350 366.840 3917.630 ;
        RECT 357.330 3916.640 357.610 3916.920 ;
        RECT 358.040 3916.640 358.320 3916.920 ;
        RECT 358.750 3916.640 359.030 3916.920 ;
        RECT 359.460 3916.640 359.740 3916.920 ;
        RECT 360.170 3916.640 360.450 3916.920 ;
        RECT 360.880 3916.640 361.160 3916.920 ;
        RECT 361.590 3916.640 361.870 3916.920 ;
        RECT 362.300 3916.640 362.580 3916.920 ;
        RECT 363.010 3916.640 363.290 3916.920 ;
        RECT 363.720 3916.640 364.000 3916.920 ;
        RECT 364.430 3916.640 364.710 3916.920 ;
        RECT 365.140 3916.640 365.420 3916.920 ;
        RECT 365.850 3916.640 366.130 3916.920 ;
        RECT 366.560 3916.640 366.840 3916.920 ;
        RECT 357.330 3915.930 357.610 3916.210 ;
        RECT 358.040 3915.930 358.320 3916.210 ;
        RECT 358.750 3915.930 359.030 3916.210 ;
        RECT 359.460 3915.930 359.740 3916.210 ;
        RECT 360.170 3915.930 360.450 3916.210 ;
        RECT 360.880 3915.930 361.160 3916.210 ;
        RECT 361.590 3915.930 361.870 3916.210 ;
        RECT 362.300 3915.930 362.580 3916.210 ;
        RECT 363.010 3915.930 363.290 3916.210 ;
        RECT 363.720 3915.930 364.000 3916.210 ;
        RECT 364.430 3915.930 364.710 3916.210 ;
        RECT 365.140 3915.930 365.420 3916.210 ;
        RECT 365.850 3915.930 366.130 3916.210 ;
        RECT 366.560 3915.930 366.840 3916.210 ;
        RECT 357.330 3915.220 357.610 3915.500 ;
        RECT 358.040 3915.220 358.320 3915.500 ;
        RECT 358.750 3915.220 359.030 3915.500 ;
        RECT 359.460 3915.220 359.740 3915.500 ;
        RECT 360.170 3915.220 360.450 3915.500 ;
        RECT 360.880 3915.220 361.160 3915.500 ;
        RECT 361.590 3915.220 361.870 3915.500 ;
        RECT 362.300 3915.220 362.580 3915.500 ;
        RECT 363.010 3915.220 363.290 3915.500 ;
        RECT 363.720 3915.220 364.000 3915.500 ;
        RECT 364.430 3915.220 364.710 3915.500 ;
        RECT 365.140 3915.220 365.420 3915.500 ;
        RECT 365.850 3915.220 366.130 3915.500 ;
        RECT 366.560 3915.220 366.840 3915.500 ;
        RECT 357.330 3914.510 357.610 3914.790 ;
        RECT 358.040 3914.510 358.320 3914.790 ;
        RECT 358.750 3914.510 359.030 3914.790 ;
        RECT 359.460 3914.510 359.740 3914.790 ;
        RECT 360.170 3914.510 360.450 3914.790 ;
        RECT 360.880 3914.510 361.160 3914.790 ;
        RECT 361.590 3914.510 361.870 3914.790 ;
        RECT 362.300 3914.510 362.580 3914.790 ;
        RECT 363.010 3914.510 363.290 3914.790 ;
        RECT 363.720 3914.510 364.000 3914.790 ;
        RECT 364.430 3914.510 364.710 3914.790 ;
        RECT 365.140 3914.510 365.420 3914.790 ;
        RECT 365.850 3914.510 366.130 3914.790 ;
        RECT 366.560 3914.510 366.840 3914.790 ;
        RECT 357.330 3913.800 357.610 3914.080 ;
        RECT 358.040 3913.800 358.320 3914.080 ;
        RECT 358.750 3913.800 359.030 3914.080 ;
        RECT 359.460 3913.800 359.740 3914.080 ;
        RECT 360.170 3913.800 360.450 3914.080 ;
        RECT 360.880 3913.800 361.160 3914.080 ;
        RECT 361.590 3913.800 361.870 3914.080 ;
        RECT 362.300 3913.800 362.580 3914.080 ;
        RECT 363.010 3913.800 363.290 3914.080 ;
        RECT 363.720 3913.800 364.000 3914.080 ;
        RECT 364.430 3913.800 364.710 3914.080 ;
        RECT 365.140 3913.800 365.420 3914.080 ;
        RECT 365.850 3913.800 366.130 3914.080 ;
        RECT 366.560 3913.800 366.840 3914.080 ;
        RECT 357.330 3913.090 357.610 3913.370 ;
        RECT 358.040 3913.090 358.320 3913.370 ;
        RECT 358.750 3913.090 359.030 3913.370 ;
        RECT 359.460 3913.090 359.740 3913.370 ;
        RECT 360.170 3913.090 360.450 3913.370 ;
        RECT 360.880 3913.090 361.160 3913.370 ;
        RECT 361.590 3913.090 361.870 3913.370 ;
        RECT 362.300 3913.090 362.580 3913.370 ;
        RECT 363.010 3913.090 363.290 3913.370 ;
        RECT 363.720 3913.090 364.000 3913.370 ;
        RECT 364.430 3913.090 364.710 3913.370 ;
        RECT 365.140 3913.090 365.420 3913.370 ;
        RECT 365.850 3913.090 366.130 3913.370 ;
        RECT 366.560 3913.090 366.840 3913.370 ;
        RECT 357.330 3912.380 357.610 3912.660 ;
        RECT 358.040 3912.380 358.320 3912.660 ;
        RECT 358.750 3912.380 359.030 3912.660 ;
        RECT 359.460 3912.380 359.740 3912.660 ;
        RECT 360.170 3912.380 360.450 3912.660 ;
        RECT 360.880 3912.380 361.160 3912.660 ;
        RECT 361.590 3912.380 361.870 3912.660 ;
        RECT 362.300 3912.380 362.580 3912.660 ;
        RECT 363.010 3912.380 363.290 3912.660 ;
        RECT 363.720 3912.380 364.000 3912.660 ;
        RECT 364.430 3912.380 364.710 3912.660 ;
        RECT 365.140 3912.380 365.420 3912.660 ;
        RECT 365.850 3912.380 366.130 3912.660 ;
        RECT 366.560 3912.380 366.840 3912.660 ;
        RECT 357.330 3911.670 357.610 3911.950 ;
        RECT 358.040 3911.670 358.320 3911.950 ;
        RECT 358.750 3911.670 359.030 3911.950 ;
        RECT 359.460 3911.670 359.740 3911.950 ;
        RECT 360.170 3911.670 360.450 3911.950 ;
        RECT 360.880 3911.670 361.160 3911.950 ;
        RECT 361.590 3911.670 361.870 3911.950 ;
        RECT 362.300 3911.670 362.580 3911.950 ;
        RECT 363.010 3911.670 363.290 3911.950 ;
        RECT 363.720 3911.670 364.000 3911.950 ;
        RECT 364.430 3911.670 364.710 3911.950 ;
        RECT 365.140 3911.670 365.420 3911.950 ;
        RECT 365.850 3911.670 366.130 3911.950 ;
        RECT 366.560 3911.670 366.840 3911.950 ;
        RECT 3500.255 3920.235 3500.535 3920.515 ;
        RECT 3500.965 3920.235 3501.245 3920.515 ;
        RECT 3501.675 3920.235 3501.955 3920.515 ;
        RECT 3502.385 3920.235 3502.665 3920.515 ;
        RECT 3503.095 3920.235 3503.375 3920.515 ;
        RECT 3503.805 3920.235 3504.085 3920.515 ;
        RECT 3504.515 3920.235 3504.795 3920.515 ;
        RECT 3505.225 3920.235 3505.505 3920.515 ;
        RECT 3505.935 3920.235 3506.215 3920.515 ;
        RECT 3506.645 3920.235 3506.925 3920.515 ;
        RECT 3507.355 3920.235 3507.635 3920.515 ;
        RECT 3508.065 3920.235 3508.345 3920.515 ;
        RECT 3508.775 3920.235 3509.055 3920.515 ;
        RECT 3509.485 3920.235 3509.765 3920.515 ;
        RECT 3500.255 3919.525 3500.535 3919.805 ;
        RECT 3500.965 3919.525 3501.245 3919.805 ;
        RECT 3501.675 3919.525 3501.955 3919.805 ;
        RECT 3502.385 3919.525 3502.665 3919.805 ;
        RECT 3503.095 3919.525 3503.375 3919.805 ;
        RECT 3503.805 3919.525 3504.085 3919.805 ;
        RECT 3504.515 3919.525 3504.795 3919.805 ;
        RECT 3505.225 3919.525 3505.505 3919.805 ;
        RECT 3505.935 3919.525 3506.215 3919.805 ;
        RECT 3506.645 3919.525 3506.925 3919.805 ;
        RECT 3507.355 3919.525 3507.635 3919.805 ;
        RECT 3508.065 3919.525 3508.345 3919.805 ;
        RECT 3508.775 3919.525 3509.055 3919.805 ;
        RECT 3509.485 3919.525 3509.765 3919.805 ;
        RECT 3500.255 3918.815 3500.535 3919.095 ;
        RECT 3500.965 3918.815 3501.245 3919.095 ;
        RECT 3501.675 3918.815 3501.955 3919.095 ;
        RECT 3502.385 3918.815 3502.665 3919.095 ;
        RECT 3503.095 3918.815 3503.375 3919.095 ;
        RECT 3503.805 3918.815 3504.085 3919.095 ;
        RECT 3504.515 3918.815 3504.795 3919.095 ;
        RECT 3505.225 3918.815 3505.505 3919.095 ;
        RECT 3505.935 3918.815 3506.215 3919.095 ;
        RECT 3506.645 3918.815 3506.925 3919.095 ;
        RECT 3507.355 3918.815 3507.635 3919.095 ;
        RECT 3508.065 3918.815 3508.345 3919.095 ;
        RECT 3508.775 3918.815 3509.055 3919.095 ;
        RECT 3509.485 3918.815 3509.765 3919.095 ;
        RECT 3500.255 3918.105 3500.535 3918.385 ;
        RECT 3500.965 3918.105 3501.245 3918.385 ;
        RECT 3501.675 3918.105 3501.955 3918.385 ;
        RECT 3502.385 3918.105 3502.665 3918.385 ;
        RECT 3503.095 3918.105 3503.375 3918.385 ;
        RECT 3503.805 3918.105 3504.085 3918.385 ;
        RECT 3504.515 3918.105 3504.795 3918.385 ;
        RECT 3505.225 3918.105 3505.505 3918.385 ;
        RECT 3505.935 3918.105 3506.215 3918.385 ;
        RECT 3506.645 3918.105 3506.925 3918.385 ;
        RECT 3507.355 3918.105 3507.635 3918.385 ;
        RECT 3508.065 3918.105 3508.345 3918.385 ;
        RECT 3508.775 3918.105 3509.055 3918.385 ;
        RECT 3509.485 3918.105 3509.765 3918.385 ;
        RECT 3500.255 3917.395 3500.535 3917.675 ;
        RECT 3500.965 3917.395 3501.245 3917.675 ;
        RECT 3501.675 3917.395 3501.955 3917.675 ;
        RECT 3502.385 3917.395 3502.665 3917.675 ;
        RECT 3503.095 3917.395 3503.375 3917.675 ;
        RECT 3503.805 3917.395 3504.085 3917.675 ;
        RECT 3504.515 3917.395 3504.795 3917.675 ;
        RECT 3505.225 3917.395 3505.505 3917.675 ;
        RECT 3505.935 3917.395 3506.215 3917.675 ;
        RECT 3506.645 3917.395 3506.925 3917.675 ;
        RECT 3507.355 3917.395 3507.635 3917.675 ;
        RECT 3508.065 3917.395 3508.345 3917.675 ;
        RECT 3508.775 3917.395 3509.055 3917.675 ;
        RECT 3509.485 3917.395 3509.765 3917.675 ;
        RECT 3500.255 3916.685 3500.535 3916.965 ;
        RECT 3500.965 3916.685 3501.245 3916.965 ;
        RECT 3501.675 3916.685 3501.955 3916.965 ;
        RECT 3502.385 3916.685 3502.665 3916.965 ;
        RECT 3503.095 3916.685 3503.375 3916.965 ;
        RECT 3503.805 3916.685 3504.085 3916.965 ;
        RECT 3504.515 3916.685 3504.795 3916.965 ;
        RECT 3505.225 3916.685 3505.505 3916.965 ;
        RECT 3505.935 3916.685 3506.215 3916.965 ;
        RECT 3506.645 3916.685 3506.925 3916.965 ;
        RECT 3507.355 3916.685 3507.635 3916.965 ;
        RECT 3508.065 3916.685 3508.345 3916.965 ;
        RECT 3508.775 3916.685 3509.055 3916.965 ;
        RECT 3509.485 3916.685 3509.765 3916.965 ;
        RECT 3500.255 3915.975 3500.535 3916.255 ;
        RECT 3500.965 3915.975 3501.245 3916.255 ;
        RECT 3501.675 3915.975 3501.955 3916.255 ;
        RECT 3502.385 3915.975 3502.665 3916.255 ;
        RECT 3503.095 3915.975 3503.375 3916.255 ;
        RECT 3503.805 3915.975 3504.085 3916.255 ;
        RECT 3504.515 3915.975 3504.795 3916.255 ;
        RECT 3505.225 3915.975 3505.505 3916.255 ;
        RECT 3505.935 3915.975 3506.215 3916.255 ;
        RECT 3506.645 3915.975 3506.925 3916.255 ;
        RECT 3507.355 3915.975 3507.635 3916.255 ;
        RECT 3508.065 3915.975 3508.345 3916.255 ;
        RECT 3508.775 3915.975 3509.055 3916.255 ;
        RECT 3509.485 3915.975 3509.765 3916.255 ;
        RECT 3500.255 3915.265 3500.535 3915.545 ;
        RECT 3500.965 3915.265 3501.245 3915.545 ;
        RECT 3501.675 3915.265 3501.955 3915.545 ;
        RECT 3502.385 3915.265 3502.665 3915.545 ;
        RECT 3503.095 3915.265 3503.375 3915.545 ;
        RECT 3503.805 3915.265 3504.085 3915.545 ;
        RECT 3504.515 3915.265 3504.795 3915.545 ;
        RECT 3505.225 3915.265 3505.505 3915.545 ;
        RECT 3505.935 3915.265 3506.215 3915.545 ;
        RECT 3506.645 3915.265 3506.925 3915.545 ;
        RECT 3507.355 3915.265 3507.635 3915.545 ;
        RECT 3508.065 3915.265 3508.345 3915.545 ;
        RECT 3508.775 3915.265 3509.055 3915.545 ;
        RECT 3509.485 3915.265 3509.765 3915.545 ;
        RECT 3500.255 3914.555 3500.535 3914.835 ;
        RECT 3500.965 3914.555 3501.245 3914.835 ;
        RECT 3501.675 3914.555 3501.955 3914.835 ;
        RECT 3502.385 3914.555 3502.665 3914.835 ;
        RECT 3503.095 3914.555 3503.375 3914.835 ;
        RECT 3503.805 3914.555 3504.085 3914.835 ;
        RECT 3504.515 3914.555 3504.795 3914.835 ;
        RECT 3505.225 3914.555 3505.505 3914.835 ;
        RECT 3505.935 3914.555 3506.215 3914.835 ;
        RECT 3506.645 3914.555 3506.925 3914.835 ;
        RECT 3507.355 3914.555 3507.635 3914.835 ;
        RECT 3508.065 3914.555 3508.345 3914.835 ;
        RECT 3508.775 3914.555 3509.055 3914.835 ;
        RECT 3509.485 3914.555 3509.765 3914.835 ;
        RECT 3500.255 3913.845 3500.535 3914.125 ;
        RECT 3500.965 3913.845 3501.245 3914.125 ;
        RECT 3501.675 3913.845 3501.955 3914.125 ;
        RECT 3502.385 3913.845 3502.665 3914.125 ;
        RECT 3503.095 3913.845 3503.375 3914.125 ;
        RECT 3503.805 3913.845 3504.085 3914.125 ;
        RECT 3504.515 3913.845 3504.795 3914.125 ;
        RECT 3505.225 3913.845 3505.505 3914.125 ;
        RECT 3505.935 3913.845 3506.215 3914.125 ;
        RECT 3506.645 3913.845 3506.925 3914.125 ;
        RECT 3507.355 3913.845 3507.635 3914.125 ;
        RECT 3508.065 3913.845 3508.345 3914.125 ;
        RECT 3508.775 3913.845 3509.055 3914.125 ;
        RECT 3509.485 3913.845 3509.765 3914.125 ;
        RECT 3500.255 3913.135 3500.535 3913.415 ;
        RECT 3500.965 3913.135 3501.245 3913.415 ;
        RECT 3501.675 3913.135 3501.955 3913.415 ;
        RECT 3502.385 3913.135 3502.665 3913.415 ;
        RECT 3503.095 3913.135 3503.375 3913.415 ;
        RECT 3503.805 3913.135 3504.085 3913.415 ;
        RECT 3504.515 3913.135 3504.795 3913.415 ;
        RECT 3505.225 3913.135 3505.505 3913.415 ;
        RECT 3505.935 3913.135 3506.215 3913.415 ;
        RECT 3506.645 3913.135 3506.925 3913.415 ;
        RECT 3507.355 3913.135 3507.635 3913.415 ;
        RECT 3508.065 3913.135 3508.345 3913.415 ;
        RECT 3508.775 3913.135 3509.055 3913.415 ;
        RECT 3509.485 3913.135 3509.765 3913.415 ;
        RECT 3500.255 3912.425 3500.535 3912.705 ;
        RECT 3500.965 3912.425 3501.245 3912.705 ;
        RECT 3501.675 3912.425 3501.955 3912.705 ;
        RECT 3502.385 3912.425 3502.665 3912.705 ;
        RECT 3503.095 3912.425 3503.375 3912.705 ;
        RECT 3503.805 3912.425 3504.085 3912.705 ;
        RECT 3504.515 3912.425 3504.795 3912.705 ;
        RECT 3505.225 3912.425 3505.505 3912.705 ;
        RECT 3505.935 3912.425 3506.215 3912.705 ;
        RECT 3506.645 3912.425 3506.925 3912.705 ;
        RECT 3507.355 3912.425 3507.635 3912.705 ;
        RECT 3508.065 3912.425 3508.345 3912.705 ;
        RECT 3508.775 3912.425 3509.055 3912.705 ;
        RECT 3509.485 3912.425 3509.765 3912.705 ;
        RECT 3500.255 3911.715 3500.535 3911.995 ;
        RECT 3500.965 3911.715 3501.245 3911.995 ;
        RECT 3501.675 3911.715 3501.955 3911.995 ;
        RECT 3502.385 3911.715 3502.665 3911.995 ;
        RECT 3503.095 3911.715 3503.375 3911.995 ;
        RECT 3503.805 3911.715 3504.085 3911.995 ;
        RECT 3504.515 3911.715 3504.795 3911.995 ;
        RECT 3505.225 3911.715 3505.505 3911.995 ;
        RECT 3505.935 3911.715 3506.215 3911.995 ;
        RECT 3506.645 3911.715 3506.925 3911.995 ;
        RECT 3507.355 3911.715 3507.635 3911.995 ;
        RECT 3508.065 3911.715 3508.345 3911.995 ;
        RECT 3508.775 3911.715 3509.055 3911.995 ;
        RECT 3509.485 3911.715 3509.765 3911.995 ;
        RECT 3500.255 3911.005 3500.535 3911.285 ;
        RECT 3500.965 3911.005 3501.245 3911.285 ;
        RECT 3501.675 3911.005 3501.955 3911.285 ;
        RECT 3502.385 3911.005 3502.665 3911.285 ;
        RECT 3503.095 3911.005 3503.375 3911.285 ;
        RECT 3503.805 3911.005 3504.085 3911.285 ;
        RECT 3504.515 3911.005 3504.795 3911.285 ;
        RECT 3505.225 3911.005 3505.505 3911.285 ;
        RECT 3505.935 3911.005 3506.215 3911.285 ;
        RECT 3506.645 3911.005 3506.925 3911.285 ;
        RECT 3507.355 3911.005 3507.635 3911.285 ;
        RECT 3508.065 3911.005 3508.345 3911.285 ;
        RECT 3508.775 3911.005 3509.055 3911.285 ;
        RECT 3509.485 3911.005 3509.765 3911.285 ;
        RECT 3500.255 3908.385 3500.535 3908.665 ;
        RECT 3500.965 3908.385 3501.245 3908.665 ;
        RECT 3501.675 3908.385 3501.955 3908.665 ;
        RECT 3502.385 3908.385 3502.665 3908.665 ;
        RECT 3503.095 3908.385 3503.375 3908.665 ;
        RECT 3503.805 3908.385 3504.085 3908.665 ;
        RECT 3504.515 3908.385 3504.795 3908.665 ;
        RECT 3505.225 3908.385 3505.505 3908.665 ;
        RECT 3505.935 3908.385 3506.215 3908.665 ;
        RECT 3506.645 3908.385 3506.925 3908.665 ;
        RECT 3507.355 3908.385 3507.635 3908.665 ;
        RECT 3508.065 3908.385 3508.345 3908.665 ;
        RECT 3508.775 3908.385 3509.055 3908.665 ;
        RECT 3509.485 3908.385 3509.765 3908.665 ;
        RECT 3500.255 3907.675 3500.535 3907.955 ;
        RECT 3500.965 3907.675 3501.245 3907.955 ;
        RECT 3501.675 3907.675 3501.955 3907.955 ;
        RECT 3502.385 3907.675 3502.665 3907.955 ;
        RECT 3503.095 3907.675 3503.375 3907.955 ;
        RECT 3503.805 3907.675 3504.085 3907.955 ;
        RECT 3504.515 3907.675 3504.795 3907.955 ;
        RECT 3505.225 3907.675 3505.505 3907.955 ;
        RECT 3505.935 3907.675 3506.215 3907.955 ;
        RECT 3506.645 3907.675 3506.925 3907.955 ;
        RECT 3507.355 3907.675 3507.635 3907.955 ;
        RECT 3508.065 3907.675 3508.345 3907.955 ;
        RECT 3508.775 3907.675 3509.055 3907.955 ;
        RECT 3509.485 3907.675 3509.765 3907.955 ;
        RECT 3500.255 3906.965 3500.535 3907.245 ;
        RECT 3500.965 3906.965 3501.245 3907.245 ;
        RECT 3501.675 3906.965 3501.955 3907.245 ;
        RECT 3502.385 3906.965 3502.665 3907.245 ;
        RECT 3503.095 3906.965 3503.375 3907.245 ;
        RECT 3503.805 3906.965 3504.085 3907.245 ;
        RECT 3504.515 3906.965 3504.795 3907.245 ;
        RECT 3505.225 3906.965 3505.505 3907.245 ;
        RECT 3505.935 3906.965 3506.215 3907.245 ;
        RECT 3506.645 3906.965 3506.925 3907.245 ;
        RECT 3507.355 3906.965 3507.635 3907.245 ;
        RECT 3508.065 3906.965 3508.345 3907.245 ;
        RECT 3508.775 3906.965 3509.055 3907.245 ;
        RECT 3509.485 3906.965 3509.765 3907.245 ;
        RECT 3500.255 3906.255 3500.535 3906.535 ;
        RECT 3500.965 3906.255 3501.245 3906.535 ;
        RECT 3501.675 3906.255 3501.955 3906.535 ;
        RECT 3502.385 3906.255 3502.665 3906.535 ;
        RECT 3503.095 3906.255 3503.375 3906.535 ;
        RECT 3503.805 3906.255 3504.085 3906.535 ;
        RECT 3504.515 3906.255 3504.795 3906.535 ;
        RECT 3505.225 3906.255 3505.505 3906.535 ;
        RECT 3505.935 3906.255 3506.215 3906.535 ;
        RECT 3506.645 3906.255 3506.925 3906.535 ;
        RECT 3507.355 3906.255 3507.635 3906.535 ;
        RECT 3508.065 3906.255 3508.345 3906.535 ;
        RECT 3508.775 3906.255 3509.055 3906.535 ;
        RECT 3509.485 3906.255 3509.765 3906.535 ;
        RECT 3500.255 3905.545 3500.535 3905.825 ;
        RECT 3500.965 3905.545 3501.245 3905.825 ;
        RECT 3501.675 3905.545 3501.955 3905.825 ;
        RECT 3502.385 3905.545 3502.665 3905.825 ;
        RECT 3503.095 3905.545 3503.375 3905.825 ;
        RECT 3503.805 3905.545 3504.085 3905.825 ;
        RECT 3504.515 3905.545 3504.795 3905.825 ;
        RECT 3505.225 3905.545 3505.505 3905.825 ;
        RECT 3505.935 3905.545 3506.215 3905.825 ;
        RECT 3506.645 3905.545 3506.925 3905.825 ;
        RECT 3507.355 3905.545 3507.635 3905.825 ;
        RECT 3508.065 3905.545 3508.345 3905.825 ;
        RECT 3508.775 3905.545 3509.055 3905.825 ;
        RECT 3509.485 3905.545 3509.765 3905.825 ;
        RECT 3500.255 3904.835 3500.535 3905.115 ;
        RECT 3500.965 3904.835 3501.245 3905.115 ;
        RECT 3501.675 3904.835 3501.955 3905.115 ;
        RECT 3502.385 3904.835 3502.665 3905.115 ;
        RECT 3503.095 3904.835 3503.375 3905.115 ;
        RECT 3503.805 3904.835 3504.085 3905.115 ;
        RECT 3504.515 3904.835 3504.795 3905.115 ;
        RECT 3505.225 3904.835 3505.505 3905.115 ;
        RECT 3505.935 3904.835 3506.215 3905.115 ;
        RECT 3506.645 3904.835 3506.925 3905.115 ;
        RECT 3507.355 3904.835 3507.635 3905.115 ;
        RECT 3508.065 3904.835 3508.345 3905.115 ;
        RECT 3508.775 3904.835 3509.055 3905.115 ;
        RECT 3509.485 3904.835 3509.765 3905.115 ;
        RECT 3500.255 3904.125 3500.535 3904.405 ;
        RECT 3500.965 3904.125 3501.245 3904.405 ;
        RECT 3501.675 3904.125 3501.955 3904.405 ;
        RECT 3502.385 3904.125 3502.665 3904.405 ;
        RECT 3503.095 3904.125 3503.375 3904.405 ;
        RECT 3503.805 3904.125 3504.085 3904.405 ;
        RECT 3504.515 3904.125 3504.795 3904.405 ;
        RECT 3505.225 3904.125 3505.505 3904.405 ;
        RECT 3505.935 3904.125 3506.215 3904.405 ;
        RECT 3506.645 3904.125 3506.925 3904.405 ;
        RECT 3507.355 3904.125 3507.635 3904.405 ;
        RECT 3508.065 3904.125 3508.345 3904.405 ;
        RECT 3508.775 3904.125 3509.055 3904.405 ;
        RECT 3509.485 3904.125 3509.765 3904.405 ;
        RECT 3500.255 3903.415 3500.535 3903.695 ;
        RECT 3500.965 3903.415 3501.245 3903.695 ;
        RECT 3501.675 3903.415 3501.955 3903.695 ;
        RECT 3502.385 3903.415 3502.665 3903.695 ;
        RECT 3503.095 3903.415 3503.375 3903.695 ;
        RECT 3503.805 3903.415 3504.085 3903.695 ;
        RECT 3504.515 3903.415 3504.795 3903.695 ;
        RECT 3505.225 3903.415 3505.505 3903.695 ;
        RECT 3505.935 3903.415 3506.215 3903.695 ;
        RECT 3506.645 3903.415 3506.925 3903.695 ;
        RECT 3507.355 3903.415 3507.635 3903.695 ;
        RECT 3508.065 3903.415 3508.345 3903.695 ;
        RECT 3508.775 3903.415 3509.055 3903.695 ;
        RECT 3509.485 3903.415 3509.765 3903.695 ;
        RECT 3500.255 3902.705 3500.535 3902.985 ;
        RECT 3500.965 3902.705 3501.245 3902.985 ;
        RECT 3501.675 3902.705 3501.955 3902.985 ;
        RECT 3502.385 3902.705 3502.665 3902.985 ;
        RECT 3503.095 3902.705 3503.375 3902.985 ;
        RECT 3503.805 3902.705 3504.085 3902.985 ;
        RECT 3504.515 3902.705 3504.795 3902.985 ;
        RECT 3505.225 3902.705 3505.505 3902.985 ;
        RECT 3505.935 3902.705 3506.215 3902.985 ;
        RECT 3506.645 3902.705 3506.925 3902.985 ;
        RECT 3507.355 3902.705 3507.635 3902.985 ;
        RECT 3508.065 3902.705 3508.345 3902.985 ;
        RECT 3508.775 3902.705 3509.055 3902.985 ;
        RECT 3509.485 3902.705 3509.765 3902.985 ;
        RECT 3500.255 3901.995 3500.535 3902.275 ;
        RECT 3500.965 3901.995 3501.245 3902.275 ;
        RECT 3501.675 3901.995 3501.955 3902.275 ;
        RECT 3502.385 3901.995 3502.665 3902.275 ;
        RECT 3503.095 3901.995 3503.375 3902.275 ;
        RECT 3503.805 3901.995 3504.085 3902.275 ;
        RECT 3504.515 3901.995 3504.795 3902.275 ;
        RECT 3505.225 3901.995 3505.505 3902.275 ;
        RECT 3505.935 3901.995 3506.215 3902.275 ;
        RECT 3506.645 3901.995 3506.925 3902.275 ;
        RECT 3507.355 3901.995 3507.635 3902.275 ;
        RECT 3508.065 3901.995 3508.345 3902.275 ;
        RECT 3508.775 3901.995 3509.055 3902.275 ;
        RECT 3509.485 3901.995 3509.765 3902.275 ;
        RECT 3500.255 3901.285 3500.535 3901.565 ;
        RECT 3500.965 3901.285 3501.245 3901.565 ;
        RECT 3501.675 3901.285 3501.955 3901.565 ;
        RECT 3502.385 3901.285 3502.665 3901.565 ;
        RECT 3503.095 3901.285 3503.375 3901.565 ;
        RECT 3503.805 3901.285 3504.085 3901.565 ;
        RECT 3504.515 3901.285 3504.795 3901.565 ;
        RECT 3505.225 3901.285 3505.505 3901.565 ;
        RECT 3505.935 3901.285 3506.215 3901.565 ;
        RECT 3506.645 3901.285 3506.925 3901.565 ;
        RECT 3507.355 3901.285 3507.635 3901.565 ;
        RECT 3508.065 3901.285 3508.345 3901.565 ;
        RECT 3508.775 3901.285 3509.055 3901.565 ;
        RECT 3509.485 3901.285 3509.765 3901.565 ;
        RECT 3500.255 3900.575 3500.535 3900.855 ;
        RECT 3500.965 3900.575 3501.245 3900.855 ;
        RECT 3501.675 3900.575 3501.955 3900.855 ;
        RECT 3502.385 3900.575 3502.665 3900.855 ;
        RECT 3503.095 3900.575 3503.375 3900.855 ;
        RECT 3503.805 3900.575 3504.085 3900.855 ;
        RECT 3504.515 3900.575 3504.795 3900.855 ;
        RECT 3505.225 3900.575 3505.505 3900.855 ;
        RECT 3505.935 3900.575 3506.215 3900.855 ;
        RECT 3506.645 3900.575 3506.925 3900.855 ;
        RECT 3507.355 3900.575 3507.635 3900.855 ;
        RECT 3508.065 3900.575 3508.345 3900.855 ;
        RECT 3508.775 3900.575 3509.055 3900.855 ;
        RECT 3509.485 3900.575 3509.765 3900.855 ;
        RECT 3500.255 3899.865 3500.535 3900.145 ;
        RECT 3500.965 3899.865 3501.245 3900.145 ;
        RECT 3501.675 3899.865 3501.955 3900.145 ;
        RECT 3502.385 3899.865 3502.665 3900.145 ;
        RECT 3503.095 3899.865 3503.375 3900.145 ;
        RECT 3503.805 3899.865 3504.085 3900.145 ;
        RECT 3504.515 3899.865 3504.795 3900.145 ;
        RECT 3505.225 3899.865 3505.505 3900.145 ;
        RECT 3505.935 3899.865 3506.215 3900.145 ;
        RECT 3506.645 3899.865 3506.925 3900.145 ;
        RECT 3507.355 3899.865 3507.635 3900.145 ;
        RECT 3508.065 3899.865 3508.345 3900.145 ;
        RECT 3508.775 3899.865 3509.055 3900.145 ;
        RECT 3509.485 3899.865 3509.765 3900.145 ;
        RECT 3500.255 3899.155 3500.535 3899.435 ;
        RECT 3500.965 3899.155 3501.245 3899.435 ;
        RECT 3501.675 3899.155 3501.955 3899.435 ;
        RECT 3502.385 3899.155 3502.665 3899.435 ;
        RECT 3503.095 3899.155 3503.375 3899.435 ;
        RECT 3503.805 3899.155 3504.085 3899.435 ;
        RECT 3504.515 3899.155 3504.795 3899.435 ;
        RECT 3505.225 3899.155 3505.505 3899.435 ;
        RECT 3505.935 3899.155 3506.215 3899.435 ;
        RECT 3506.645 3899.155 3506.925 3899.435 ;
        RECT 3507.355 3899.155 3507.635 3899.435 ;
        RECT 3508.065 3899.155 3508.345 3899.435 ;
        RECT 3508.775 3899.155 3509.055 3899.435 ;
        RECT 3509.485 3899.155 3509.765 3899.435 ;
        RECT 3500.200 3895.270 3500.480 3895.550 ;
        RECT 3500.910 3895.270 3501.190 3895.550 ;
        RECT 3501.620 3895.270 3501.900 3895.550 ;
        RECT 3502.330 3895.270 3502.610 3895.550 ;
        RECT 3503.040 3895.270 3503.320 3895.550 ;
        RECT 3503.750 3895.270 3504.030 3895.550 ;
        RECT 3504.460 3895.270 3504.740 3895.550 ;
        RECT 3505.170 3895.270 3505.450 3895.550 ;
        RECT 3505.880 3895.270 3506.160 3895.550 ;
        RECT 3506.590 3895.270 3506.870 3895.550 ;
        RECT 3507.300 3895.270 3507.580 3895.550 ;
        RECT 3508.010 3895.270 3508.290 3895.550 ;
        RECT 3508.720 3895.270 3509.000 3895.550 ;
        RECT 3509.430 3895.270 3509.710 3895.550 ;
        RECT 3500.200 3894.560 3500.480 3894.840 ;
        RECT 3500.910 3894.560 3501.190 3894.840 ;
        RECT 3501.620 3894.560 3501.900 3894.840 ;
        RECT 3502.330 3894.560 3502.610 3894.840 ;
        RECT 3503.040 3894.560 3503.320 3894.840 ;
        RECT 3503.750 3894.560 3504.030 3894.840 ;
        RECT 3504.460 3894.560 3504.740 3894.840 ;
        RECT 3505.170 3894.560 3505.450 3894.840 ;
        RECT 3505.880 3894.560 3506.160 3894.840 ;
        RECT 3506.590 3894.560 3506.870 3894.840 ;
        RECT 3507.300 3894.560 3507.580 3894.840 ;
        RECT 3508.010 3894.560 3508.290 3894.840 ;
        RECT 3508.720 3894.560 3509.000 3894.840 ;
        RECT 3509.430 3894.560 3509.710 3894.840 ;
        RECT 3500.200 3893.850 3500.480 3894.130 ;
        RECT 3500.910 3893.850 3501.190 3894.130 ;
        RECT 3501.620 3893.850 3501.900 3894.130 ;
        RECT 3502.330 3893.850 3502.610 3894.130 ;
        RECT 3503.040 3893.850 3503.320 3894.130 ;
        RECT 3503.750 3893.850 3504.030 3894.130 ;
        RECT 3504.460 3893.850 3504.740 3894.130 ;
        RECT 3505.170 3893.850 3505.450 3894.130 ;
        RECT 3505.880 3893.850 3506.160 3894.130 ;
        RECT 3506.590 3893.850 3506.870 3894.130 ;
        RECT 3507.300 3893.850 3507.580 3894.130 ;
        RECT 3508.010 3893.850 3508.290 3894.130 ;
        RECT 3508.720 3893.850 3509.000 3894.130 ;
        RECT 3509.430 3893.850 3509.710 3894.130 ;
        RECT 3500.200 3893.140 3500.480 3893.420 ;
        RECT 3500.910 3893.140 3501.190 3893.420 ;
        RECT 3501.620 3893.140 3501.900 3893.420 ;
        RECT 3502.330 3893.140 3502.610 3893.420 ;
        RECT 3503.040 3893.140 3503.320 3893.420 ;
        RECT 3503.750 3893.140 3504.030 3893.420 ;
        RECT 3504.460 3893.140 3504.740 3893.420 ;
        RECT 3505.170 3893.140 3505.450 3893.420 ;
        RECT 3505.880 3893.140 3506.160 3893.420 ;
        RECT 3506.590 3893.140 3506.870 3893.420 ;
        RECT 3507.300 3893.140 3507.580 3893.420 ;
        RECT 3508.010 3893.140 3508.290 3893.420 ;
        RECT 3508.720 3893.140 3509.000 3893.420 ;
        RECT 3509.430 3893.140 3509.710 3893.420 ;
        RECT 3500.200 3892.430 3500.480 3892.710 ;
        RECT 3500.910 3892.430 3501.190 3892.710 ;
        RECT 3501.620 3892.430 3501.900 3892.710 ;
        RECT 3502.330 3892.430 3502.610 3892.710 ;
        RECT 3503.040 3892.430 3503.320 3892.710 ;
        RECT 3503.750 3892.430 3504.030 3892.710 ;
        RECT 3504.460 3892.430 3504.740 3892.710 ;
        RECT 3505.170 3892.430 3505.450 3892.710 ;
        RECT 3505.880 3892.430 3506.160 3892.710 ;
        RECT 3506.590 3892.430 3506.870 3892.710 ;
        RECT 3507.300 3892.430 3507.580 3892.710 ;
        RECT 3508.010 3892.430 3508.290 3892.710 ;
        RECT 3508.720 3892.430 3509.000 3892.710 ;
        RECT 3509.430 3892.430 3509.710 3892.710 ;
        RECT 3500.200 3891.720 3500.480 3892.000 ;
        RECT 3500.910 3891.720 3501.190 3892.000 ;
        RECT 3501.620 3891.720 3501.900 3892.000 ;
        RECT 3502.330 3891.720 3502.610 3892.000 ;
        RECT 3503.040 3891.720 3503.320 3892.000 ;
        RECT 3503.750 3891.720 3504.030 3892.000 ;
        RECT 3504.460 3891.720 3504.740 3892.000 ;
        RECT 3505.170 3891.720 3505.450 3892.000 ;
        RECT 3505.880 3891.720 3506.160 3892.000 ;
        RECT 3506.590 3891.720 3506.870 3892.000 ;
        RECT 3507.300 3891.720 3507.580 3892.000 ;
        RECT 3508.010 3891.720 3508.290 3892.000 ;
        RECT 3508.720 3891.720 3509.000 3892.000 ;
        RECT 3509.430 3891.720 3509.710 3892.000 ;
        RECT 3500.200 3891.010 3500.480 3891.290 ;
        RECT 3500.910 3891.010 3501.190 3891.290 ;
        RECT 3501.620 3891.010 3501.900 3891.290 ;
        RECT 3502.330 3891.010 3502.610 3891.290 ;
        RECT 3503.040 3891.010 3503.320 3891.290 ;
        RECT 3503.750 3891.010 3504.030 3891.290 ;
        RECT 3504.460 3891.010 3504.740 3891.290 ;
        RECT 3505.170 3891.010 3505.450 3891.290 ;
        RECT 3505.880 3891.010 3506.160 3891.290 ;
        RECT 3506.590 3891.010 3506.870 3891.290 ;
        RECT 3507.300 3891.010 3507.580 3891.290 ;
        RECT 3508.010 3891.010 3508.290 3891.290 ;
        RECT 3508.720 3891.010 3509.000 3891.290 ;
        RECT 3509.430 3891.010 3509.710 3891.290 ;
        RECT 3500.200 3890.300 3500.480 3890.580 ;
        RECT 3500.910 3890.300 3501.190 3890.580 ;
        RECT 3501.620 3890.300 3501.900 3890.580 ;
        RECT 3502.330 3890.300 3502.610 3890.580 ;
        RECT 3503.040 3890.300 3503.320 3890.580 ;
        RECT 3503.750 3890.300 3504.030 3890.580 ;
        RECT 3504.460 3890.300 3504.740 3890.580 ;
        RECT 3505.170 3890.300 3505.450 3890.580 ;
        RECT 3505.880 3890.300 3506.160 3890.580 ;
        RECT 3506.590 3890.300 3506.870 3890.580 ;
        RECT 3507.300 3890.300 3507.580 3890.580 ;
        RECT 3508.010 3890.300 3508.290 3890.580 ;
        RECT 3508.720 3890.300 3509.000 3890.580 ;
        RECT 3509.430 3890.300 3509.710 3890.580 ;
        RECT 3500.200 3889.590 3500.480 3889.870 ;
        RECT 3500.910 3889.590 3501.190 3889.870 ;
        RECT 3501.620 3889.590 3501.900 3889.870 ;
        RECT 3502.330 3889.590 3502.610 3889.870 ;
        RECT 3503.040 3889.590 3503.320 3889.870 ;
        RECT 3503.750 3889.590 3504.030 3889.870 ;
        RECT 3504.460 3889.590 3504.740 3889.870 ;
        RECT 3505.170 3889.590 3505.450 3889.870 ;
        RECT 3505.880 3889.590 3506.160 3889.870 ;
        RECT 3506.590 3889.590 3506.870 3889.870 ;
        RECT 3507.300 3889.590 3507.580 3889.870 ;
        RECT 3508.010 3889.590 3508.290 3889.870 ;
        RECT 3508.720 3889.590 3509.000 3889.870 ;
        RECT 3509.430 3889.590 3509.710 3889.870 ;
        RECT 3500.200 3888.880 3500.480 3889.160 ;
        RECT 3500.910 3888.880 3501.190 3889.160 ;
        RECT 3501.620 3888.880 3501.900 3889.160 ;
        RECT 3502.330 3888.880 3502.610 3889.160 ;
        RECT 3503.040 3888.880 3503.320 3889.160 ;
        RECT 3503.750 3888.880 3504.030 3889.160 ;
        RECT 3504.460 3888.880 3504.740 3889.160 ;
        RECT 3505.170 3888.880 3505.450 3889.160 ;
        RECT 3505.880 3888.880 3506.160 3889.160 ;
        RECT 3506.590 3888.880 3506.870 3889.160 ;
        RECT 3507.300 3888.880 3507.580 3889.160 ;
        RECT 3508.010 3888.880 3508.290 3889.160 ;
        RECT 3508.720 3888.880 3509.000 3889.160 ;
        RECT 3509.430 3888.880 3509.710 3889.160 ;
        RECT 3500.200 3888.170 3500.480 3888.450 ;
        RECT 3500.910 3888.170 3501.190 3888.450 ;
        RECT 3501.620 3888.170 3501.900 3888.450 ;
        RECT 3502.330 3888.170 3502.610 3888.450 ;
        RECT 3503.040 3888.170 3503.320 3888.450 ;
        RECT 3503.750 3888.170 3504.030 3888.450 ;
        RECT 3504.460 3888.170 3504.740 3888.450 ;
        RECT 3505.170 3888.170 3505.450 3888.450 ;
        RECT 3505.880 3888.170 3506.160 3888.450 ;
        RECT 3506.590 3888.170 3506.870 3888.450 ;
        RECT 3507.300 3888.170 3507.580 3888.450 ;
        RECT 3508.010 3888.170 3508.290 3888.450 ;
        RECT 3508.720 3888.170 3509.000 3888.450 ;
        RECT 3509.430 3888.170 3509.710 3888.450 ;
        RECT 3500.200 3887.460 3500.480 3887.740 ;
        RECT 3500.910 3887.460 3501.190 3887.740 ;
        RECT 3501.620 3887.460 3501.900 3887.740 ;
        RECT 3502.330 3887.460 3502.610 3887.740 ;
        RECT 3503.040 3887.460 3503.320 3887.740 ;
        RECT 3503.750 3887.460 3504.030 3887.740 ;
        RECT 3504.460 3887.460 3504.740 3887.740 ;
        RECT 3505.170 3887.460 3505.450 3887.740 ;
        RECT 3505.880 3887.460 3506.160 3887.740 ;
        RECT 3506.590 3887.460 3506.870 3887.740 ;
        RECT 3507.300 3887.460 3507.580 3887.740 ;
        RECT 3508.010 3887.460 3508.290 3887.740 ;
        RECT 3508.720 3887.460 3509.000 3887.740 ;
        RECT 3509.430 3887.460 3509.710 3887.740 ;
        RECT 3500.200 3886.750 3500.480 3887.030 ;
        RECT 3500.910 3886.750 3501.190 3887.030 ;
        RECT 3501.620 3886.750 3501.900 3887.030 ;
        RECT 3502.330 3886.750 3502.610 3887.030 ;
        RECT 3503.040 3886.750 3503.320 3887.030 ;
        RECT 3503.750 3886.750 3504.030 3887.030 ;
        RECT 3504.460 3886.750 3504.740 3887.030 ;
        RECT 3505.170 3886.750 3505.450 3887.030 ;
        RECT 3505.880 3886.750 3506.160 3887.030 ;
        RECT 3506.590 3886.750 3506.870 3887.030 ;
        RECT 3507.300 3886.750 3507.580 3887.030 ;
        RECT 3508.010 3886.750 3508.290 3887.030 ;
        RECT 3508.720 3886.750 3509.000 3887.030 ;
        RECT 3509.430 3886.750 3509.710 3887.030 ;
        RECT 3500.200 2453.050 3500.480 2453.330 ;
        RECT 3500.910 2453.050 3501.190 2453.330 ;
        RECT 3501.620 2453.050 3501.900 2453.330 ;
        RECT 3502.330 2453.050 3502.610 2453.330 ;
        RECT 3503.040 2453.050 3503.320 2453.330 ;
        RECT 3503.750 2453.050 3504.030 2453.330 ;
        RECT 3504.460 2453.050 3504.740 2453.330 ;
        RECT 3505.170 2453.050 3505.450 2453.330 ;
        RECT 3505.880 2453.050 3506.160 2453.330 ;
        RECT 3506.590 2453.050 3506.870 2453.330 ;
        RECT 3507.300 2453.050 3507.580 2453.330 ;
        RECT 3508.010 2453.050 3508.290 2453.330 ;
        RECT 3508.720 2453.050 3509.000 2453.330 ;
        RECT 3509.430 2453.050 3509.710 2453.330 ;
        RECT 3500.200 2452.340 3500.480 2452.620 ;
        RECT 3500.910 2452.340 3501.190 2452.620 ;
        RECT 3501.620 2452.340 3501.900 2452.620 ;
        RECT 3502.330 2452.340 3502.610 2452.620 ;
        RECT 3503.040 2452.340 3503.320 2452.620 ;
        RECT 3503.750 2452.340 3504.030 2452.620 ;
        RECT 3504.460 2452.340 3504.740 2452.620 ;
        RECT 3505.170 2452.340 3505.450 2452.620 ;
        RECT 3505.880 2452.340 3506.160 2452.620 ;
        RECT 3506.590 2452.340 3506.870 2452.620 ;
        RECT 3507.300 2452.340 3507.580 2452.620 ;
        RECT 3508.010 2452.340 3508.290 2452.620 ;
        RECT 3508.720 2452.340 3509.000 2452.620 ;
        RECT 3509.430 2452.340 3509.710 2452.620 ;
        RECT 3500.200 2451.630 3500.480 2451.910 ;
        RECT 3500.910 2451.630 3501.190 2451.910 ;
        RECT 3501.620 2451.630 3501.900 2451.910 ;
        RECT 3502.330 2451.630 3502.610 2451.910 ;
        RECT 3503.040 2451.630 3503.320 2451.910 ;
        RECT 3503.750 2451.630 3504.030 2451.910 ;
        RECT 3504.460 2451.630 3504.740 2451.910 ;
        RECT 3505.170 2451.630 3505.450 2451.910 ;
        RECT 3505.880 2451.630 3506.160 2451.910 ;
        RECT 3506.590 2451.630 3506.870 2451.910 ;
        RECT 3507.300 2451.630 3507.580 2451.910 ;
        RECT 3508.010 2451.630 3508.290 2451.910 ;
        RECT 3508.720 2451.630 3509.000 2451.910 ;
        RECT 3509.430 2451.630 3509.710 2451.910 ;
        RECT 3500.200 2450.920 3500.480 2451.200 ;
        RECT 3500.910 2450.920 3501.190 2451.200 ;
        RECT 3501.620 2450.920 3501.900 2451.200 ;
        RECT 3502.330 2450.920 3502.610 2451.200 ;
        RECT 3503.040 2450.920 3503.320 2451.200 ;
        RECT 3503.750 2450.920 3504.030 2451.200 ;
        RECT 3504.460 2450.920 3504.740 2451.200 ;
        RECT 3505.170 2450.920 3505.450 2451.200 ;
        RECT 3505.880 2450.920 3506.160 2451.200 ;
        RECT 3506.590 2450.920 3506.870 2451.200 ;
        RECT 3507.300 2450.920 3507.580 2451.200 ;
        RECT 3508.010 2450.920 3508.290 2451.200 ;
        RECT 3508.720 2450.920 3509.000 2451.200 ;
        RECT 3509.430 2450.920 3509.710 2451.200 ;
        RECT 3500.200 2450.210 3500.480 2450.490 ;
        RECT 3500.910 2450.210 3501.190 2450.490 ;
        RECT 3501.620 2450.210 3501.900 2450.490 ;
        RECT 3502.330 2450.210 3502.610 2450.490 ;
        RECT 3503.040 2450.210 3503.320 2450.490 ;
        RECT 3503.750 2450.210 3504.030 2450.490 ;
        RECT 3504.460 2450.210 3504.740 2450.490 ;
        RECT 3505.170 2450.210 3505.450 2450.490 ;
        RECT 3505.880 2450.210 3506.160 2450.490 ;
        RECT 3506.590 2450.210 3506.870 2450.490 ;
        RECT 3507.300 2450.210 3507.580 2450.490 ;
        RECT 3508.010 2450.210 3508.290 2450.490 ;
        RECT 3508.720 2450.210 3509.000 2450.490 ;
        RECT 3509.430 2450.210 3509.710 2450.490 ;
        RECT 3500.200 2449.500 3500.480 2449.780 ;
        RECT 3500.910 2449.500 3501.190 2449.780 ;
        RECT 3501.620 2449.500 3501.900 2449.780 ;
        RECT 3502.330 2449.500 3502.610 2449.780 ;
        RECT 3503.040 2449.500 3503.320 2449.780 ;
        RECT 3503.750 2449.500 3504.030 2449.780 ;
        RECT 3504.460 2449.500 3504.740 2449.780 ;
        RECT 3505.170 2449.500 3505.450 2449.780 ;
        RECT 3505.880 2449.500 3506.160 2449.780 ;
        RECT 3506.590 2449.500 3506.870 2449.780 ;
        RECT 3507.300 2449.500 3507.580 2449.780 ;
        RECT 3508.010 2449.500 3508.290 2449.780 ;
        RECT 3508.720 2449.500 3509.000 2449.780 ;
        RECT 3509.430 2449.500 3509.710 2449.780 ;
        RECT 3500.200 2448.790 3500.480 2449.070 ;
        RECT 3500.910 2448.790 3501.190 2449.070 ;
        RECT 3501.620 2448.790 3501.900 2449.070 ;
        RECT 3502.330 2448.790 3502.610 2449.070 ;
        RECT 3503.040 2448.790 3503.320 2449.070 ;
        RECT 3503.750 2448.790 3504.030 2449.070 ;
        RECT 3504.460 2448.790 3504.740 2449.070 ;
        RECT 3505.170 2448.790 3505.450 2449.070 ;
        RECT 3505.880 2448.790 3506.160 2449.070 ;
        RECT 3506.590 2448.790 3506.870 2449.070 ;
        RECT 3507.300 2448.790 3507.580 2449.070 ;
        RECT 3508.010 2448.790 3508.290 2449.070 ;
        RECT 3508.720 2448.790 3509.000 2449.070 ;
        RECT 3509.430 2448.790 3509.710 2449.070 ;
        RECT 3500.200 2448.080 3500.480 2448.360 ;
        RECT 3500.910 2448.080 3501.190 2448.360 ;
        RECT 3501.620 2448.080 3501.900 2448.360 ;
        RECT 3502.330 2448.080 3502.610 2448.360 ;
        RECT 3503.040 2448.080 3503.320 2448.360 ;
        RECT 3503.750 2448.080 3504.030 2448.360 ;
        RECT 3504.460 2448.080 3504.740 2448.360 ;
        RECT 3505.170 2448.080 3505.450 2448.360 ;
        RECT 3505.880 2448.080 3506.160 2448.360 ;
        RECT 3506.590 2448.080 3506.870 2448.360 ;
        RECT 3507.300 2448.080 3507.580 2448.360 ;
        RECT 3508.010 2448.080 3508.290 2448.360 ;
        RECT 3508.720 2448.080 3509.000 2448.360 ;
        RECT 3509.430 2448.080 3509.710 2448.360 ;
        RECT 3500.200 2447.370 3500.480 2447.650 ;
        RECT 3500.910 2447.370 3501.190 2447.650 ;
        RECT 3501.620 2447.370 3501.900 2447.650 ;
        RECT 3502.330 2447.370 3502.610 2447.650 ;
        RECT 3503.040 2447.370 3503.320 2447.650 ;
        RECT 3503.750 2447.370 3504.030 2447.650 ;
        RECT 3504.460 2447.370 3504.740 2447.650 ;
        RECT 3505.170 2447.370 3505.450 2447.650 ;
        RECT 3505.880 2447.370 3506.160 2447.650 ;
        RECT 3506.590 2447.370 3506.870 2447.650 ;
        RECT 3507.300 2447.370 3507.580 2447.650 ;
        RECT 3508.010 2447.370 3508.290 2447.650 ;
        RECT 3508.720 2447.370 3509.000 2447.650 ;
        RECT 3509.430 2447.370 3509.710 2447.650 ;
        RECT 3500.200 2446.660 3500.480 2446.940 ;
        RECT 3500.910 2446.660 3501.190 2446.940 ;
        RECT 3501.620 2446.660 3501.900 2446.940 ;
        RECT 3502.330 2446.660 3502.610 2446.940 ;
        RECT 3503.040 2446.660 3503.320 2446.940 ;
        RECT 3503.750 2446.660 3504.030 2446.940 ;
        RECT 3504.460 2446.660 3504.740 2446.940 ;
        RECT 3505.170 2446.660 3505.450 2446.940 ;
        RECT 3505.880 2446.660 3506.160 2446.940 ;
        RECT 3506.590 2446.660 3506.870 2446.940 ;
        RECT 3507.300 2446.660 3507.580 2446.940 ;
        RECT 3508.010 2446.660 3508.290 2446.940 ;
        RECT 3508.720 2446.660 3509.000 2446.940 ;
        RECT 3509.430 2446.660 3509.710 2446.940 ;
        RECT 3500.200 2445.950 3500.480 2446.230 ;
        RECT 3500.910 2445.950 3501.190 2446.230 ;
        RECT 3501.620 2445.950 3501.900 2446.230 ;
        RECT 3502.330 2445.950 3502.610 2446.230 ;
        RECT 3503.040 2445.950 3503.320 2446.230 ;
        RECT 3503.750 2445.950 3504.030 2446.230 ;
        RECT 3504.460 2445.950 3504.740 2446.230 ;
        RECT 3505.170 2445.950 3505.450 2446.230 ;
        RECT 3505.880 2445.950 3506.160 2446.230 ;
        RECT 3506.590 2445.950 3506.870 2446.230 ;
        RECT 3507.300 2445.950 3507.580 2446.230 ;
        RECT 3508.010 2445.950 3508.290 2446.230 ;
        RECT 3508.720 2445.950 3509.000 2446.230 ;
        RECT 3509.430 2445.950 3509.710 2446.230 ;
        RECT 3500.200 2445.240 3500.480 2445.520 ;
        RECT 3500.910 2445.240 3501.190 2445.520 ;
        RECT 3501.620 2445.240 3501.900 2445.520 ;
        RECT 3502.330 2445.240 3502.610 2445.520 ;
        RECT 3503.040 2445.240 3503.320 2445.520 ;
        RECT 3503.750 2445.240 3504.030 2445.520 ;
        RECT 3504.460 2445.240 3504.740 2445.520 ;
        RECT 3505.170 2445.240 3505.450 2445.520 ;
        RECT 3505.880 2445.240 3506.160 2445.520 ;
        RECT 3506.590 2445.240 3506.870 2445.520 ;
        RECT 3507.300 2445.240 3507.580 2445.520 ;
        RECT 3508.010 2445.240 3508.290 2445.520 ;
        RECT 3508.720 2445.240 3509.000 2445.520 ;
        RECT 3509.430 2445.240 3509.710 2445.520 ;
        RECT 3500.200 2444.530 3500.480 2444.810 ;
        RECT 3500.910 2444.530 3501.190 2444.810 ;
        RECT 3501.620 2444.530 3501.900 2444.810 ;
        RECT 3502.330 2444.530 3502.610 2444.810 ;
        RECT 3503.040 2444.530 3503.320 2444.810 ;
        RECT 3503.750 2444.530 3504.030 2444.810 ;
        RECT 3504.460 2444.530 3504.740 2444.810 ;
        RECT 3505.170 2444.530 3505.450 2444.810 ;
        RECT 3505.880 2444.530 3506.160 2444.810 ;
        RECT 3506.590 2444.530 3506.870 2444.810 ;
        RECT 3507.300 2444.530 3507.580 2444.810 ;
        RECT 3508.010 2444.530 3508.290 2444.810 ;
        RECT 3508.720 2444.530 3509.000 2444.810 ;
        RECT 3509.430 2444.530 3509.710 2444.810 ;
        RECT 3500.255 2440.615 3500.535 2440.895 ;
        RECT 3500.965 2440.615 3501.245 2440.895 ;
        RECT 3501.675 2440.615 3501.955 2440.895 ;
        RECT 3502.385 2440.615 3502.665 2440.895 ;
        RECT 3503.095 2440.615 3503.375 2440.895 ;
        RECT 3503.805 2440.615 3504.085 2440.895 ;
        RECT 3504.515 2440.615 3504.795 2440.895 ;
        RECT 3505.225 2440.615 3505.505 2440.895 ;
        RECT 3505.935 2440.615 3506.215 2440.895 ;
        RECT 3506.645 2440.615 3506.925 2440.895 ;
        RECT 3507.355 2440.615 3507.635 2440.895 ;
        RECT 3508.065 2440.615 3508.345 2440.895 ;
        RECT 3508.775 2440.615 3509.055 2440.895 ;
        RECT 3509.485 2440.615 3509.765 2440.895 ;
        RECT 3500.255 2439.905 3500.535 2440.185 ;
        RECT 3500.965 2439.905 3501.245 2440.185 ;
        RECT 3501.675 2439.905 3501.955 2440.185 ;
        RECT 3502.385 2439.905 3502.665 2440.185 ;
        RECT 3503.095 2439.905 3503.375 2440.185 ;
        RECT 3503.805 2439.905 3504.085 2440.185 ;
        RECT 3504.515 2439.905 3504.795 2440.185 ;
        RECT 3505.225 2439.905 3505.505 2440.185 ;
        RECT 3505.935 2439.905 3506.215 2440.185 ;
        RECT 3506.645 2439.905 3506.925 2440.185 ;
        RECT 3507.355 2439.905 3507.635 2440.185 ;
        RECT 3508.065 2439.905 3508.345 2440.185 ;
        RECT 3508.775 2439.905 3509.055 2440.185 ;
        RECT 3509.485 2439.905 3509.765 2440.185 ;
        RECT 3500.255 2439.195 3500.535 2439.475 ;
        RECT 3500.965 2439.195 3501.245 2439.475 ;
        RECT 3501.675 2439.195 3501.955 2439.475 ;
        RECT 3502.385 2439.195 3502.665 2439.475 ;
        RECT 3503.095 2439.195 3503.375 2439.475 ;
        RECT 3503.805 2439.195 3504.085 2439.475 ;
        RECT 3504.515 2439.195 3504.795 2439.475 ;
        RECT 3505.225 2439.195 3505.505 2439.475 ;
        RECT 3505.935 2439.195 3506.215 2439.475 ;
        RECT 3506.645 2439.195 3506.925 2439.475 ;
        RECT 3507.355 2439.195 3507.635 2439.475 ;
        RECT 3508.065 2439.195 3508.345 2439.475 ;
        RECT 3508.775 2439.195 3509.055 2439.475 ;
        RECT 3509.485 2439.195 3509.765 2439.475 ;
        RECT 3500.255 2438.485 3500.535 2438.765 ;
        RECT 3500.965 2438.485 3501.245 2438.765 ;
        RECT 3501.675 2438.485 3501.955 2438.765 ;
        RECT 3502.385 2438.485 3502.665 2438.765 ;
        RECT 3503.095 2438.485 3503.375 2438.765 ;
        RECT 3503.805 2438.485 3504.085 2438.765 ;
        RECT 3504.515 2438.485 3504.795 2438.765 ;
        RECT 3505.225 2438.485 3505.505 2438.765 ;
        RECT 3505.935 2438.485 3506.215 2438.765 ;
        RECT 3506.645 2438.485 3506.925 2438.765 ;
        RECT 3507.355 2438.485 3507.635 2438.765 ;
        RECT 3508.065 2438.485 3508.345 2438.765 ;
        RECT 3508.775 2438.485 3509.055 2438.765 ;
        RECT 3509.485 2438.485 3509.765 2438.765 ;
        RECT 3500.255 2437.775 3500.535 2438.055 ;
        RECT 3500.965 2437.775 3501.245 2438.055 ;
        RECT 3501.675 2437.775 3501.955 2438.055 ;
        RECT 3502.385 2437.775 3502.665 2438.055 ;
        RECT 3503.095 2437.775 3503.375 2438.055 ;
        RECT 3503.805 2437.775 3504.085 2438.055 ;
        RECT 3504.515 2437.775 3504.795 2438.055 ;
        RECT 3505.225 2437.775 3505.505 2438.055 ;
        RECT 3505.935 2437.775 3506.215 2438.055 ;
        RECT 3506.645 2437.775 3506.925 2438.055 ;
        RECT 3507.355 2437.775 3507.635 2438.055 ;
        RECT 3508.065 2437.775 3508.345 2438.055 ;
        RECT 3508.775 2437.775 3509.055 2438.055 ;
        RECT 3509.485 2437.775 3509.765 2438.055 ;
        RECT 3500.255 2437.065 3500.535 2437.345 ;
        RECT 3500.965 2437.065 3501.245 2437.345 ;
        RECT 3501.675 2437.065 3501.955 2437.345 ;
        RECT 3502.385 2437.065 3502.665 2437.345 ;
        RECT 3503.095 2437.065 3503.375 2437.345 ;
        RECT 3503.805 2437.065 3504.085 2437.345 ;
        RECT 3504.515 2437.065 3504.795 2437.345 ;
        RECT 3505.225 2437.065 3505.505 2437.345 ;
        RECT 3505.935 2437.065 3506.215 2437.345 ;
        RECT 3506.645 2437.065 3506.925 2437.345 ;
        RECT 3507.355 2437.065 3507.635 2437.345 ;
        RECT 3508.065 2437.065 3508.345 2437.345 ;
        RECT 3508.775 2437.065 3509.055 2437.345 ;
        RECT 3509.485 2437.065 3509.765 2437.345 ;
        RECT 3500.255 2436.355 3500.535 2436.635 ;
        RECT 3500.965 2436.355 3501.245 2436.635 ;
        RECT 3501.675 2436.355 3501.955 2436.635 ;
        RECT 3502.385 2436.355 3502.665 2436.635 ;
        RECT 3503.095 2436.355 3503.375 2436.635 ;
        RECT 3503.805 2436.355 3504.085 2436.635 ;
        RECT 3504.515 2436.355 3504.795 2436.635 ;
        RECT 3505.225 2436.355 3505.505 2436.635 ;
        RECT 3505.935 2436.355 3506.215 2436.635 ;
        RECT 3506.645 2436.355 3506.925 2436.635 ;
        RECT 3507.355 2436.355 3507.635 2436.635 ;
        RECT 3508.065 2436.355 3508.345 2436.635 ;
        RECT 3508.775 2436.355 3509.055 2436.635 ;
        RECT 3509.485 2436.355 3509.765 2436.635 ;
        RECT 3500.255 2435.645 3500.535 2435.925 ;
        RECT 3500.965 2435.645 3501.245 2435.925 ;
        RECT 3501.675 2435.645 3501.955 2435.925 ;
        RECT 3502.385 2435.645 3502.665 2435.925 ;
        RECT 3503.095 2435.645 3503.375 2435.925 ;
        RECT 3503.805 2435.645 3504.085 2435.925 ;
        RECT 3504.515 2435.645 3504.795 2435.925 ;
        RECT 3505.225 2435.645 3505.505 2435.925 ;
        RECT 3505.935 2435.645 3506.215 2435.925 ;
        RECT 3506.645 2435.645 3506.925 2435.925 ;
        RECT 3507.355 2435.645 3507.635 2435.925 ;
        RECT 3508.065 2435.645 3508.345 2435.925 ;
        RECT 3508.775 2435.645 3509.055 2435.925 ;
        RECT 3509.485 2435.645 3509.765 2435.925 ;
        RECT 3500.255 2434.935 3500.535 2435.215 ;
        RECT 3500.965 2434.935 3501.245 2435.215 ;
        RECT 3501.675 2434.935 3501.955 2435.215 ;
        RECT 3502.385 2434.935 3502.665 2435.215 ;
        RECT 3503.095 2434.935 3503.375 2435.215 ;
        RECT 3503.805 2434.935 3504.085 2435.215 ;
        RECT 3504.515 2434.935 3504.795 2435.215 ;
        RECT 3505.225 2434.935 3505.505 2435.215 ;
        RECT 3505.935 2434.935 3506.215 2435.215 ;
        RECT 3506.645 2434.935 3506.925 2435.215 ;
        RECT 3507.355 2434.935 3507.635 2435.215 ;
        RECT 3508.065 2434.935 3508.345 2435.215 ;
        RECT 3508.775 2434.935 3509.055 2435.215 ;
        RECT 3509.485 2434.935 3509.765 2435.215 ;
        RECT 3500.255 2434.225 3500.535 2434.505 ;
        RECT 3500.965 2434.225 3501.245 2434.505 ;
        RECT 3501.675 2434.225 3501.955 2434.505 ;
        RECT 3502.385 2434.225 3502.665 2434.505 ;
        RECT 3503.095 2434.225 3503.375 2434.505 ;
        RECT 3503.805 2434.225 3504.085 2434.505 ;
        RECT 3504.515 2434.225 3504.795 2434.505 ;
        RECT 3505.225 2434.225 3505.505 2434.505 ;
        RECT 3505.935 2434.225 3506.215 2434.505 ;
        RECT 3506.645 2434.225 3506.925 2434.505 ;
        RECT 3507.355 2434.225 3507.635 2434.505 ;
        RECT 3508.065 2434.225 3508.345 2434.505 ;
        RECT 3508.775 2434.225 3509.055 2434.505 ;
        RECT 3509.485 2434.225 3509.765 2434.505 ;
        RECT 3500.255 2433.515 3500.535 2433.795 ;
        RECT 3500.965 2433.515 3501.245 2433.795 ;
        RECT 3501.675 2433.515 3501.955 2433.795 ;
        RECT 3502.385 2433.515 3502.665 2433.795 ;
        RECT 3503.095 2433.515 3503.375 2433.795 ;
        RECT 3503.805 2433.515 3504.085 2433.795 ;
        RECT 3504.515 2433.515 3504.795 2433.795 ;
        RECT 3505.225 2433.515 3505.505 2433.795 ;
        RECT 3505.935 2433.515 3506.215 2433.795 ;
        RECT 3506.645 2433.515 3506.925 2433.795 ;
        RECT 3507.355 2433.515 3507.635 2433.795 ;
        RECT 3508.065 2433.515 3508.345 2433.795 ;
        RECT 3508.775 2433.515 3509.055 2433.795 ;
        RECT 3509.485 2433.515 3509.765 2433.795 ;
        RECT 3500.255 2432.805 3500.535 2433.085 ;
        RECT 3500.965 2432.805 3501.245 2433.085 ;
        RECT 3501.675 2432.805 3501.955 2433.085 ;
        RECT 3502.385 2432.805 3502.665 2433.085 ;
        RECT 3503.095 2432.805 3503.375 2433.085 ;
        RECT 3503.805 2432.805 3504.085 2433.085 ;
        RECT 3504.515 2432.805 3504.795 2433.085 ;
        RECT 3505.225 2432.805 3505.505 2433.085 ;
        RECT 3505.935 2432.805 3506.215 2433.085 ;
        RECT 3506.645 2432.805 3506.925 2433.085 ;
        RECT 3507.355 2432.805 3507.635 2433.085 ;
        RECT 3508.065 2432.805 3508.345 2433.085 ;
        RECT 3508.775 2432.805 3509.055 2433.085 ;
        RECT 3509.485 2432.805 3509.765 2433.085 ;
        RECT 3500.255 2432.095 3500.535 2432.375 ;
        RECT 3500.965 2432.095 3501.245 2432.375 ;
        RECT 3501.675 2432.095 3501.955 2432.375 ;
        RECT 3502.385 2432.095 3502.665 2432.375 ;
        RECT 3503.095 2432.095 3503.375 2432.375 ;
        RECT 3503.805 2432.095 3504.085 2432.375 ;
        RECT 3504.515 2432.095 3504.795 2432.375 ;
        RECT 3505.225 2432.095 3505.505 2432.375 ;
        RECT 3505.935 2432.095 3506.215 2432.375 ;
        RECT 3506.645 2432.095 3506.925 2432.375 ;
        RECT 3507.355 2432.095 3507.635 2432.375 ;
        RECT 3508.065 2432.095 3508.345 2432.375 ;
        RECT 3508.775 2432.095 3509.055 2432.375 ;
        RECT 3509.485 2432.095 3509.765 2432.375 ;
        RECT 3500.255 2431.385 3500.535 2431.665 ;
        RECT 3500.965 2431.385 3501.245 2431.665 ;
        RECT 3501.675 2431.385 3501.955 2431.665 ;
        RECT 3502.385 2431.385 3502.665 2431.665 ;
        RECT 3503.095 2431.385 3503.375 2431.665 ;
        RECT 3503.805 2431.385 3504.085 2431.665 ;
        RECT 3504.515 2431.385 3504.795 2431.665 ;
        RECT 3505.225 2431.385 3505.505 2431.665 ;
        RECT 3505.935 2431.385 3506.215 2431.665 ;
        RECT 3506.645 2431.385 3506.925 2431.665 ;
        RECT 3507.355 2431.385 3507.635 2431.665 ;
        RECT 3508.065 2431.385 3508.345 2431.665 ;
        RECT 3508.775 2431.385 3509.055 2431.665 ;
        RECT 3509.485 2431.385 3509.765 2431.665 ;
        RECT 3500.255 2428.765 3500.535 2429.045 ;
        RECT 3500.965 2428.765 3501.245 2429.045 ;
        RECT 3501.675 2428.765 3501.955 2429.045 ;
        RECT 3502.385 2428.765 3502.665 2429.045 ;
        RECT 3503.095 2428.765 3503.375 2429.045 ;
        RECT 3503.805 2428.765 3504.085 2429.045 ;
        RECT 3504.515 2428.765 3504.795 2429.045 ;
        RECT 3505.225 2428.765 3505.505 2429.045 ;
        RECT 3505.935 2428.765 3506.215 2429.045 ;
        RECT 3506.645 2428.765 3506.925 2429.045 ;
        RECT 3507.355 2428.765 3507.635 2429.045 ;
        RECT 3508.065 2428.765 3508.345 2429.045 ;
        RECT 3508.775 2428.765 3509.055 2429.045 ;
        RECT 3509.485 2428.765 3509.765 2429.045 ;
        RECT 3500.255 2428.055 3500.535 2428.335 ;
        RECT 3500.965 2428.055 3501.245 2428.335 ;
        RECT 3501.675 2428.055 3501.955 2428.335 ;
        RECT 3502.385 2428.055 3502.665 2428.335 ;
        RECT 3503.095 2428.055 3503.375 2428.335 ;
        RECT 3503.805 2428.055 3504.085 2428.335 ;
        RECT 3504.515 2428.055 3504.795 2428.335 ;
        RECT 3505.225 2428.055 3505.505 2428.335 ;
        RECT 3505.935 2428.055 3506.215 2428.335 ;
        RECT 3506.645 2428.055 3506.925 2428.335 ;
        RECT 3507.355 2428.055 3507.635 2428.335 ;
        RECT 3508.065 2428.055 3508.345 2428.335 ;
        RECT 3508.775 2428.055 3509.055 2428.335 ;
        RECT 3509.485 2428.055 3509.765 2428.335 ;
        RECT 3500.255 2427.345 3500.535 2427.625 ;
        RECT 3500.965 2427.345 3501.245 2427.625 ;
        RECT 3501.675 2427.345 3501.955 2427.625 ;
        RECT 3502.385 2427.345 3502.665 2427.625 ;
        RECT 3503.095 2427.345 3503.375 2427.625 ;
        RECT 3503.805 2427.345 3504.085 2427.625 ;
        RECT 3504.515 2427.345 3504.795 2427.625 ;
        RECT 3505.225 2427.345 3505.505 2427.625 ;
        RECT 3505.935 2427.345 3506.215 2427.625 ;
        RECT 3506.645 2427.345 3506.925 2427.625 ;
        RECT 3507.355 2427.345 3507.635 2427.625 ;
        RECT 3508.065 2427.345 3508.345 2427.625 ;
        RECT 3508.775 2427.345 3509.055 2427.625 ;
        RECT 3509.485 2427.345 3509.765 2427.625 ;
        RECT 3500.255 2426.635 3500.535 2426.915 ;
        RECT 3500.965 2426.635 3501.245 2426.915 ;
        RECT 3501.675 2426.635 3501.955 2426.915 ;
        RECT 3502.385 2426.635 3502.665 2426.915 ;
        RECT 3503.095 2426.635 3503.375 2426.915 ;
        RECT 3503.805 2426.635 3504.085 2426.915 ;
        RECT 3504.515 2426.635 3504.795 2426.915 ;
        RECT 3505.225 2426.635 3505.505 2426.915 ;
        RECT 3505.935 2426.635 3506.215 2426.915 ;
        RECT 3506.645 2426.635 3506.925 2426.915 ;
        RECT 3507.355 2426.635 3507.635 2426.915 ;
        RECT 3508.065 2426.635 3508.345 2426.915 ;
        RECT 3508.775 2426.635 3509.055 2426.915 ;
        RECT 3509.485 2426.635 3509.765 2426.915 ;
        RECT 3500.255 2425.925 3500.535 2426.205 ;
        RECT 3500.965 2425.925 3501.245 2426.205 ;
        RECT 3501.675 2425.925 3501.955 2426.205 ;
        RECT 3502.385 2425.925 3502.665 2426.205 ;
        RECT 3503.095 2425.925 3503.375 2426.205 ;
        RECT 3503.805 2425.925 3504.085 2426.205 ;
        RECT 3504.515 2425.925 3504.795 2426.205 ;
        RECT 3505.225 2425.925 3505.505 2426.205 ;
        RECT 3505.935 2425.925 3506.215 2426.205 ;
        RECT 3506.645 2425.925 3506.925 2426.205 ;
        RECT 3507.355 2425.925 3507.635 2426.205 ;
        RECT 3508.065 2425.925 3508.345 2426.205 ;
        RECT 3508.775 2425.925 3509.055 2426.205 ;
        RECT 3509.485 2425.925 3509.765 2426.205 ;
        RECT 3500.255 2425.215 3500.535 2425.495 ;
        RECT 3500.965 2425.215 3501.245 2425.495 ;
        RECT 3501.675 2425.215 3501.955 2425.495 ;
        RECT 3502.385 2425.215 3502.665 2425.495 ;
        RECT 3503.095 2425.215 3503.375 2425.495 ;
        RECT 3503.805 2425.215 3504.085 2425.495 ;
        RECT 3504.515 2425.215 3504.795 2425.495 ;
        RECT 3505.225 2425.215 3505.505 2425.495 ;
        RECT 3505.935 2425.215 3506.215 2425.495 ;
        RECT 3506.645 2425.215 3506.925 2425.495 ;
        RECT 3507.355 2425.215 3507.635 2425.495 ;
        RECT 3508.065 2425.215 3508.345 2425.495 ;
        RECT 3508.775 2425.215 3509.055 2425.495 ;
        RECT 3509.485 2425.215 3509.765 2425.495 ;
        RECT 3500.255 2424.505 3500.535 2424.785 ;
        RECT 3500.965 2424.505 3501.245 2424.785 ;
        RECT 3501.675 2424.505 3501.955 2424.785 ;
        RECT 3502.385 2424.505 3502.665 2424.785 ;
        RECT 3503.095 2424.505 3503.375 2424.785 ;
        RECT 3503.805 2424.505 3504.085 2424.785 ;
        RECT 3504.515 2424.505 3504.795 2424.785 ;
        RECT 3505.225 2424.505 3505.505 2424.785 ;
        RECT 3505.935 2424.505 3506.215 2424.785 ;
        RECT 3506.645 2424.505 3506.925 2424.785 ;
        RECT 3507.355 2424.505 3507.635 2424.785 ;
        RECT 3508.065 2424.505 3508.345 2424.785 ;
        RECT 3508.775 2424.505 3509.055 2424.785 ;
        RECT 3509.485 2424.505 3509.765 2424.785 ;
        RECT 3500.255 2423.795 3500.535 2424.075 ;
        RECT 3500.965 2423.795 3501.245 2424.075 ;
        RECT 3501.675 2423.795 3501.955 2424.075 ;
        RECT 3502.385 2423.795 3502.665 2424.075 ;
        RECT 3503.095 2423.795 3503.375 2424.075 ;
        RECT 3503.805 2423.795 3504.085 2424.075 ;
        RECT 3504.515 2423.795 3504.795 2424.075 ;
        RECT 3505.225 2423.795 3505.505 2424.075 ;
        RECT 3505.935 2423.795 3506.215 2424.075 ;
        RECT 3506.645 2423.795 3506.925 2424.075 ;
        RECT 3507.355 2423.795 3507.635 2424.075 ;
        RECT 3508.065 2423.795 3508.345 2424.075 ;
        RECT 3508.775 2423.795 3509.055 2424.075 ;
        RECT 3509.485 2423.795 3509.765 2424.075 ;
        RECT 3500.255 2423.085 3500.535 2423.365 ;
        RECT 3500.965 2423.085 3501.245 2423.365 ;
        RECT 3501.675 2423.085 3501.955 2423.365 ;
        RECT 3502.385 2423.085 3502.665 2423.365 ;
        RECT 3503.095 2423.085 3503.375 2423.365 ;
        RECT 3503.805 2423.085 3504.085 2423.365 ;
        RECT 3504.515 2423.085 3504.795 2423.365 ;
        RECT 3505.225 2423.085 3505.505 2423.365 ;
        RECT 3505.935 2423.085 3506.215 2423.365 ;
        RECT 3506.645 2423.085 3506.925 2423.365 ;
        RECT 3507.355 2423.085 3507.635 2423.365 ;
        RECT 3508.065 2423.085 3508.345 2423.365 ;
        RECT 3508.775 2423.085 3509.055 2423.365 ;
        RECT 3509.485 2423.085 3509.765 2423.365 ;
        RECT 3500.255 2422.375 3500.535 2422.655 ;
        RECT 3500.965 2422.375 3501.245 2422.655 ;
        RECT 3501.675 2422.375 3501.955 2422.655 ;
        RECT 3502.385 2422.375 3502.665 2422.655 ;
        RECT 3503.095 2422.375 3503.375 2422.655 ;
        RECT 3503.805 2422.375 3504.085 2422.655 ;
        RECT 3504.515 2422.375 3504.795 2422.655 ;
        RECT 3505.225 2422.375 3505.505 2422.655 ;
        RECT 3505.935 2422.375 3506.215 2422.655 ;
        RECT 3506.645 2422.375 3506.925 2422.655 ;
        RECT 3507.355 2422.375 3507.635 2422.655 ;
        RECT 3508.065 2422.375 3508.345 2422.655 ;
        RECT 3508.775 2422.375 3509.055 2422.655 ;
        RECT 3509.485 2422.375 3509.765 2422.655 ;
        RECT 3500.255 2421.665 3500.535 2421.945 ;
        RECT 3500.965 2421.665 3501.245 2421.945 ;
        RECT 3501.675 2421.665 3501.955 2421.945 ;
        RECT 3502.385 2421.665 3502.665 2421.945 ;
        RECT 3503.095 2421.665 3503.375 2421.945 ;
        RECT 3503.805 2421.665 3504.085 2421.945 ;
        RECT 3504.515 2421.665 3504.795 2421.945 ;
        RECT 3505.225 2421.665 3505.505 2421.945 ;
        RECT 3505.935 2421.665 3506.215 2421.945 ;
        RECT 3506.645 2421.665 3506.925 2421.945 ;
        RECT 3507.355 2421.665 3507.635 2421.945 ;
        RECT 3508.065 2421.665 3508.345 2421.945 ;
        RECT 3508.775 2421.665 3509.055 2421.945 ;
        RECT 3509.485 2421.665 3509.765 2421.945 ;
        RECT 3500.255 2420.955 3500.535 2421.235 ;
        RECT 3500.965 2420.955 3501.245 2421.235 ;
        RECT 3501.675 2420.955 3501.955 2421.235 ;
        RECT 3502.385 2420.955 3502.665 2421.235 ;
        RECT 3503.095 2420.955 3503.375 2421.235 ;
        RECT 3503.805 2420.955 3504.085 2421.235 ;
        RECT 3504.515 2420.955 3504.795 2421.235 ;
        RECT 3505.225 2420.955 3505.505 2421.235 ;
        RECT 3505.935 2420.955 3506.215 2421.235 ;
        RECT 3506.645 2420.955 3506.925 2421.235 ;
        RECT 3507.355 2420.955 3507.635 2421.235 ;
        RECT 3508.065 2420.955 3508.345 2421.235 ;
        RECT 3508.775 2420.955 3509.055 2421.235 ;
        RECT 3509.485 2420.955 3509.765 2421.235 ;
        RECT 3500.255 2420.245 3500.535 2420.525 ;
        RECT 3500.965 2420.245 3501.245 2420.525 ;
        RECT 3501.675 2420.245 3501.955 2420.525 ;
        RECT 3502.385 2420.245 3502.665 2420.525 ;
        RECT 3503.095 2420.245 3503.375 2420.525 ;
        RECT 3503.805 2420.245 3504.085 2420.525 ;
        RECT 3504.515 2420.245 3504.795 2420.525 ;
        RECT 3505.225 2420.245 3505.505 2420.525 ;
        RECT 3505.935 2420.245 3506.215 2420.525 ;
        RECT 3506.645 2420.245 3506.925 2420.525 ;
        RECT 3507.355 2420.245 3507.635 2420.525 ;
        RECT 3508.065 2420.245 3508.345 2420.525 ;
        RECT 3508.775 2420.245 3509.055 2420.525 ;
        RECT 3509.485 2420.245 3509.765 2420.525 ;
        RECT 3500.255 2419.535 3500.535 2419.815 ;
        RECT 3500.965 2419.535 3501.245 2419.815 ;
        RECT 3501.675 2419.535 3501.955 2419.815 ;
        RECT 3502.385 2419.535 3502.665 2419.815 ;
        RECT 3503.095 2419.535 3503.375 2419.815 ;
        RECT 3503.805 2419.535 3504.085 2419.815 ;
        RECT 3504.515 2419.535 3504.795 2419.815 ;
        RECT 3505.225 2419.535 3505.505 2419.815 ;
        RECT 3505.935 2419.535 3506.215 2419.815 ;
        RECT 3506.645 2419.535 3506.925 2419.815 ;
        RECT 3507.355 2419.535 3507.635 2419.815 ;
        RECT 3508.065 2419.535 3508.345 2419.815 ;
        RECT 3508.775 2419.535 3509.055 2419.815 ;
        RECT 3509.485 2419.535 3509.765 2419.815 ;
        RECT 3500.255 2415.235 3500.535 2415.515 ;
        RECT 3500.965 2415.235 3501.245 2415.515 ;
        RECT 3501.675 2415.235 3501.955 2415.515 ;
        RECT 3502.385 2415.235 3502.665 2415.515 ;
        RECT 3503.095 2415.235 3503.375 2415.515 ;
        RECT 3503.805 2415.235 3504.085 2415.515 ;
        RECT 3504.515 2415.235 3504.795 2415.515 ;
        RECT 3505.225 2415.235 3505.505 2415.515 ;
        RECT 3505.935 2415.235 3506.215 2415.515 ;
        RECT 3506.645 2415.235 3506.925 2415.515 ;
        RECT 3507.355 2415.235 3507.635 2415.515 ;
        RECT 3508.065 2415.235 3508.345 2415.515 ;
        RECT 3508.775 2415.235 3509.055 2415.515 ;
        RECT 3509.485 2415.235 3509.765 2415.515 ;
        RECT 3500.255 2414.525 3500.535 2414.805 ;
        RECT 3500.965 2414.525 3501.245 2414.805 ;
        RECT 3501.675 2414.525 3501.955 2414.805 ;
        RECT 3502.385 2414.525 3502.665 2414.805 ;
        RECT 3503.095 2414.525 3503.375 2414.805 ;
        RECT 3503.805 2414.525 3504.085 2414.805 ;
        RECT 3504.515 2414.525 3504.795 2414.805 ;
        RECT 3505.225 2414.525 3505.505 2414.805 ;
        RECT 3505.935 2414.525 3506.215 2414.805 ;
        RECT 3506.645 2414.525 3506.925 2414.805 ;
        RECT 3507.355 2414.525 3507.635 2414.805 ;
        RECT 3508.065 2414.525 3508.345 2414.805 ;
        RECT 3508.775 2414.525 3509.055 2414.805 ;
        RECT 3509.485 2414.525 3509.765 2414.805 ;
        RECT 3500.255 2413.815 3500.535 2414.095 ;
        RECT 3500.965 2413.815 3501.245 2414.095 ;
        RECT 3501.675 2413.815 3501.955 2414.095 ;
        RECT 3502.385 2413.815 3502.665 2414.095 ;
        RECT 3503.095 2413.815 3503.375 2414.095 ;
        RECT 3503.805 2413.815 3504.085 2414.095 ;
        RECT 3504.515 2413.815 3504.795 2414.095 ;
        RECT 3505.225 2413.815 3505.505 2414.095 ;
        RECT 3505.935 2413.815 3506.215 2414.095 ;
        RECT 3506.645 2413.815 3506.925 2414.095 ;
        RECT 3507.355 2413.815 3507.635 2414.095 ;
        RECT 3508.065 2413.815 3508.345 2414.095 ;
        RECT 3508.775 2413.815 3509.055 2414.095 ;
        RECT 3509.485 2413.815 3509.765 2414.095 ;
        RECT 3500.255 2413.105 3500.535 2413.385 ;
        RECT 3500.965 2413.105 3501.245 2413.385 ;
        RECT 3501.675 2413.105 3501.955 2413.385 ;
        RECT 3502.385 2413.105 3502.665 2413.385 ;
        RECT 3503.095 2413.105 3503.375 2413.385 ;
        RECT 3503.805 2413.105 3504.085 2413.385 ;
        RECT 3504.515 2413.105 3504.795 2413.385 ;
        RECT 3505.225 2413.105 3505.505 2413.385 ;
        RECT 3505.935 2413.105 3506.215 2413.385 ;
        RECT 3506.645 2413.105 3506.925 2413.385 ;
        RECT 3507.355 2413.105 3507.635 2413.385 ;
        RECT 3508.065 2413.105 3508.345 2413.385 ;
        RECT 3508.775 2413.105 3509.055 2413.385 ;
        RECT 3509.485 2413.105 3509.765 2413.385 ;
        RECT 3500.255 2412.395 3500.535 2412.675 ;
        RECT 3500.965 2412.395 3501.245 2412.675 ;
        RECT 3501.675 2412.395 3501.955 2412.675 ;
        RECT 3502.385 2412.395 3502.665 2412.675 ;
        RECT 3503.095 2412.395 3503.375 2412.675 ;
        RECT 3503.805 2412.395 3504.085 2412.675 ;
        RECT 3504.515 2412.395 3504.795 2412.675 ;
        RECT 3505.225 2412.395 3505.505 2412.675 ;
        RECT 3505.935 2412.395 3506.215 2412.675 ;
        RECT 3506.645 2412.395 3506.925 2412.675 ;
        RECT 3507.355 2412.395 3507.635 2412.675 ;
        RECT 3508.065 2412.395 3508.345 2412.675 ;
        RECT 3508.775 2412.395 3509.055 2412.675 ;
        RECT 3509.485 2412.395 3509.765 2412.675 ;
        RECT 3500.255 2411.685 3500.535 2411.965 ;
        RECT 3500.965 2411.685 3501.245 2411.965 ;
        RECT 3501.675 2411.685 3501.955 2411.965 ;
        RECT 3502.385 2411.685 3502.665 2411.965 ;
        RECT 3503.095 2411.685 3503.375 2411.965 ;
        RECT 3503.805 2411.685 3504.085 2411.965 ;
        RECT 3504.515 2411.685 3504.795 2411.965 ;
        RECT 3505.225 2411.685 3505.505 2411.965 ;
        RECT 3505.935 2411.685 3506.215 2411.965 ;
        RECT 3506.645 2411.685 3506.925 2411.965 ;
        RECT 3507.355 2411.685 3507.635 2411.965 ;
        RECT 3508.065 2411.685 3508.345 2411.965 ;
        RECT 3508.775 2411.685 3509.055 2411.965 ;
        RECT 3509.485 2411.685 3509.765 2411.965 ;
        RECT 3500.255 2410.975 3500.535 2411.255 ;
        RECT 3500.965 2410.975 3501.245 2411.255 ;
        RECT 3501.675 2410.975 3501.955 2411.255 ;
        RECT 3502.385 2410.975 3502.665 2411.255 ;
        RECT 3503.095 2410.975 3503.375 2411.255 ;
        RECT 3503.805 2410.975 3504.085 2411.255 ;
        RECT 3504.515 2410.975 3504.795 2411.255 ;
        RECT 3505.225 2410.975 3505.505 2411.255 ;
        RECT 3505.935 2410.975 3506.215 2411.255 ;
        RECT 3506.645 2410.975 3506.925 2411.255 ;
        RECT 3507.355 2410.975 3507.635 2411.255 ;
        RECT 3508.065 2410.975 3508.345 2411.255 ;
        RECT 3508.775 2410.975 3509.055 2411.255 ;
        RECT 3509.485 2410.975 3509.765 2411.255 ;
        RECT 3500.255 2410.265 3500.535 2410.545 ;
        RECT 3500.965 2410.265 3501.245 2410.545 ;
        RECT 3501.675 2410.265 3501.955 2410.545 ;
        RECT 3502.385 2410.265 3502.665 2410.545 ;
        RECT 3503.095 2410.265 3503.375 2410.545 ;
        RECT 3503.805 2410.265 3504.085 2410.545 ;
        RECT 3504.515 2410.265 3504.795 2410.545 ;
        RECT 3505.225 2410.265 3505.505 2410.545 ;
        RECT 3505.935 2410.265 3506.215 2410.545 ;
        RECT 3506.645 2410.265 3506.925 2410.545 ;
        RECT 3507.355 2410.265 3507.635 2410.545 ;
        RECT 3508.065 2410.265 3508.345 2410.545 ;
        RECT 3508.775 2410.265 3509.055 2410.545 ;
        RECT 3509.485 2410.265 3509.765 2410.545 ;
        RECT 3500.255 2409.555 3500.535 2409.835 ;
        RECT 3500.965 2409.555 3501.245 2409.835 ;
        RECT 3501.675 2409.555 3501.955 2409.835 ;
        RECT 3502.385 2409.555 3502.665 2409.835 ;
        RECT 3503.095 2409.555 3503.375 2409.835 ;
        RECT 3503.805 2409.555 3504.085 2409.835 ;
        RECT 3504.515 2409.555 3504.795 2409.835 ;
        RECT 3505.225 2409.555 3505.505 2409.835 ;
        RECT 3505.935 2409.555 3506.215 2409.835 ;
        RECT 3506.645 2409.555 3506.925 2409.835 ;
        RECT 3507.355 2409.555 3507.635 2409.835 ;
        RECT 3508.065 2409.555 3508.345 2409.835 ;
        RECT 3508.775 2409.555 3509.055 2409.835 ;
        RECT 3509.485 2409.555 3509.765 2409.835 ;
        RECT 3500.255 2408.845 3500.535 2409.125 ;
        RECT 3500.965 2408.845 3501.245 2409.125 ;
        RECT 3501.675 2408.845 3501.955 2409.125 ;
        RECT 3502.385 2408.845 3502.665 2409.125 ;
        RECT 3503.095 2408.845 3503.375 2409.125 ;
        RECT 3503.805 2408.845 3504.085 2409.125 ;
        RECT 3504.515 2408.845 3504.795 2409.125 ;
        RECT 3505.225 2408.845 3505.505 2409.125 ;
        RECT 3505.935 2408.845 3506.215 2409.125 ;
        RECT 3506.645 2408.845 3506.925 2409.125 ;
        RECT 3507.355 2408.845 3507.635 2409.125 ;
        RECT 3508.065 2408.845 3508.345 2409.125 ;
        RECT 3508.775 2408.845 3509.055 2409.125 ;
        RECT 3509.485 2408.845 3509.765 2409.125 ;
        RECT 3500.255 2408.135 3500.535 2408.415 ;
        RECT 3500.965 2408.135 3501.245 2408.415 ;
        RECT 3501.675 2408.135 3501.955 2408.415 ;
        RECT 3502.385 2408.135 3502.665 2408.415 ;
        RECT 3503.095 2408.135 3503.375 2408.415 ;
        RECT 3503.805 2408.135 3504.085 2408.415 ;
        RECT 3504.515 2408.135 3504.795 2408.415 ;
        RECT 3505.225 2408.135 3505.505 2408.415 ;
        RECT 3505.935 2408.135 3506.215 2408.415 ;
        RECT 3506.645 2408.135 3506.925 2408.415 ;
        RECT 3507.355 2408.135 3507.635 2408.415 ;
        RECT 3508.065 2408.135 3508.345 2408.415 ;
        RECT 3508.775 2408.135 3509.055 2408.415 ;
        RECT 3509.485 2408.135 3509.765 2408.415 ;
        RECT 3500.255 2407.425 3500.535 2407.705 ;
        RECT 3500.965 2407.425 3501.245 2407.705 ;
        RECT 3501.675 2407.425 3501.955 2407.705 ;
        RECT 3502.385 2407.425 3502.665 2407.705 ;
        RECT 3503.095 2407.425 3503.375 2407.705 ;
        RECT 3503.805 2407.425 3504.085 2407.705 ;
        RECT 3504.515 2407.425 3504.795 2407.705 ;
        RECT 3505.225 2407.425 3505.505 2407.705 ;
        RECT 3505.935 2407.425 3506.215 2407.705 ;
        RECT 3506.645 2407.425 3506.925 2407.705 ;
        RECT 3507.355 2407.425 3507.635 2407.705 ;
        RECT 3508.065 2407.425 3508.345 2407.705 ;
        RECT 3508.775 2407.425 3509.055 2407.705 ;
        RECT 3509.485 2407.425 3509.765 2407.705 ;
        RECT 3500.255 2406.715 3500.535 2406.995 ;
        RECT 3500.965 2406.715 3501.245 2406.995 ;
        RECT 3501.675 2406.715 3501.955 2406.995 ;
        RECT 3502.385 2406.715 3502.665 2406.995 ;
        RECT 3503.095 2406.715 3503.375 2406.995 ;
        RECT 3503.805 2406.715 3504.085 2406.995 ;
        RECT 3504.515 2406.715 3504.795 2406.995 ;
        RECT 3505.225 2406.715 3505.505 2406.995 ;
        RECT 3505.935 2406.715 3506.215 2406.995 ;
        RECT 3506.645 2406.715 3506.925 2406.995 ;
        RECT 3507.355 2406.715 3507.635 2406.995 ;
        RECT 3508.065 2406.715 3508.345 2406.995 ;
        RECT 3508.775 2406.715 3509.055 2406.995 ;
        RECT 3509.485 2406.715 3509.765 2406.995 ;
        RECT 3500.255 2406.005 3500.535 2406.285 ;
        RECT 3500.965 2406.005 3501.245 2406.285 ;
        RECT 3501.675 2406.005 3501.955 2406.285 ;
        RECT 3502.385 2406.005 3502.665 2406.285 ;
        RECT 3503.095 2406.005 3503.375 2406.285 ;
        RECT 3503.805 2406.005 3504.085 2406.285 ;
        RECT 3504.515 2406.005 3504.795 2406.285 ;
        RECT 3505.225 2406.005 3505.505 2406.285 ;
        RECT 3505.935 2406.005 3506.215 2406.285 ;
        RECT 3506.645 2406.005 3506.925 2406.285 ;
        RECT 3507.355 2406.005 3507.635 2406.285 ;
        RECT 3508.065 2406.005 3508.345 2406.285 ;
        RECT 3508.775 2406.005 3509.055 2406.285 ;
        RECT 3509.485 2406.005 3509.765 2406.285 ;
        RECT 3500.255 2403.385 3500.535 2403.665 ;
        RECT 3500.965 2403.385 3501.245 2403.665 ;
        RECT 3501.675 2403.385 3501.955 2403.665 ;
        RECT 3502.385 2403.385 3502.665 2403.665 ;
        RECT 3503.095 2403.385 3503.375 2403.665 ;
        RECT 3503.805 2403.385 3504.085 2403.665 ;
        RECT 3504.515 2403.385 3504.795 2403.665 ;
        RECT 3505.225 2403.385 3505.505 2403.665 ;
        RECT 3505.935 2403.385 3506.215 2403.665 ;
        RECT 3506.645 2403.385 3506.925 2403.665 ;
        RECT 3507.355 2403.385 3507.635 2403.665 ;
        RECT 3508.065 2403.385 3508.345 2403.665 ;
        RECT 3508.775 2403.385 3509.055 2403.665 ;
        RECT 3509.485 2403.385 3509.765 2403.665 ;
        RECT 3500.255 2402.675 3500.535 2402.955 ;
        RECT 3500.965 2402.675 3501.245 2402.955 ;
        RECT 3501.675 2402.675 3501.955 2402.955 ;
        RECT 3502.385 2402.675 3502.665 2402.955 ;
        RECT 3503.095 2402.675 3503.375 2402.955 ;
        RECT 3503.805 2402.675 3504.085 2402.955 ;
        RECT 3504.515 2402.675 3504.795 2402.955 ;
        RECT 3505.225 2402.675 3505.505 2402.955 ;
        RECT 3505.935 2402.675 3506.215 2402.955 ;
        RECT 3506.645 2402.675 3506.925 2402.955 ;
        RECT 3507.355 2402.675 3507.635 2402.955 ;
        RECT 3508.065 2402.675 3508.345 2402.955 ;
        RECT 3508.775 2402.675 3509.055 2402.955 ;
        RECT 3509.485 2402.675 3509.765 2402.955 ;
        RECT 3500.255 2401.965 3500.535 2402.245 ;
        RECT 3500.965 2401.965 3501.245 2402.245 ;
        RECT 3501.675 2401.965 3501.955 2402.245 ;
        RECT 3502.385 2401.965 3502.665 2402.245 ;
        RECT 3503.095 2401.965 3503.375 2402.245 ;
        RECT 3503.805 2401.965 3504.085 2402.245 ;
        RECT 3504.515 2401.965 3504.795 2402.245 ;
        RECT 3505.225 2401.965 3505.505 2402.245 ;
        RECT 3505.935 2401.965 3506.215 2402.245 ;
        RECT 3506.645 2401.965 3506.925 2402.245 ;
        RECT 3507.355 2401.965 3507.635 2402.245 ;
        RECT 3508.065 2401.965 3508.345 2402.245 ;
        RECT 3508.775 2401.965 3509.055 2402.245 ;
        RECT 3509.485 2401.965 3509.765 2402.245 ;
        RECT 3500.255 2401.255 3500.535 2401.535 ;
        RECT 3500.965 2401.255 3501.245 2401.535 ;
        RECT 3501.675 2401.255 3501.955 2401.535 ;
        RECT 3502.385 2401.255 3502.665 2401.535 ;
        RECT 3503.095 2401.255 3503.375 2401.535 ;
        RECT 3503.805 2401.255 3504.085 2401.535 ;
        RECT 3504.515 2401.255 3504.795 2401.535 ;
        RECT 3505.225 2401.255 3505.505 2401.535 ;
        RECT 3505.935 2401.255 3506.215 2401.535 ;
        RECT 3506.645 2401.255 3506.925 2401.535 ;
        RECT 3507.355 2401.255 3507.635 2401.535 ;
        RECT 3508.065 2401.255 3508.345 2401.535 ;
        RECT 3508.775 2401.255 3509.055 2401.535 ;
        RECT 3509.485 2401.255 3509.765 2401.535 ;
        RECT 3500.255 2400.545 3500.535 2400.825 ;
        RECT 3500.965 2400.545 3501.245 2400.825 ;
        RECT 3501.675 2400.545 3501.955 2400.825 ;
        RECT 3502.385 2400.545 3502.665 2400.825 ;
        RECT 3503.095 2400.545 3503.375 2400.825 ;
        RECT 3503.805 2400.545 3504.085 2400.825 ;
        RECT 3504.515 2400.545 3504.795 2400.825 ;
        RECT 3505.225 2400.545 3505.505 2400.825 ;
        RECT 3505.935 2400.545 3506.215 2400.825 ;
        RECT 3506.645 2400.545 3506.925 2400.825 ;
        RECT 3507.355 2400.545 3507.635 2400.825 ;
        RECT 3508.065 2400.545 3508.345 2400.825 ;
        RECT 3508.775 2400.545 3509.055 2400.825 ;
        RECT 3509.485 2400.545 3509.765 2400.825 ;
        RECT 3500.255 2399.835 3500.535 2400.115 ;
        RECT 3500.965 2399.835 3501.245 2400.115 ;
        RECT 3501.675 2399.835 3501.955 2400.115 ;
        RECT 3502.385 2399.835 3502.665 2400.115 ;
        RECT 3503.095 2399.835 3503.375 2400.115 ;
        RECT 3503.805 2399.835 3504.085 2400.115 ;
        RECT 3504.515 2399.835 3504.795 2400.115 ;
        RECT 3505.225 2399.835 3505.505 2400.115 ;
        RECT 3505.935 2399.835 3506.215 2400.115 ;
        RECT 3506.645 2399.835 3506.925 2400.115 ;
        RECT 3507.355 2399.835 3507.635 2400.115 ;
        RECT 3508.065 2399.835 3508.345 2400.115 ;
        RECT 3508.775 2399.835 3509.055 2400.115 ;
        RECT 3509.485 2399.835 3509.765 2400.115 ;
        RECT 3500.255 2399.125 3500.535 2399.405 ;
        RECT 3500.965 2399.125 3501.245 2399.405 ;
        RECT 3501.675 2399.125 3501.955 2399.405 ;
        RECT 3502.385 2399.125 3502.665 2399.405 ;
        RECT 3503.095 2399.125 3503.375 2399.405 ;
        RECT 3503.805 2399.125 3504.085 2399.405 ;
        RECT 3504.515 2399.125 3504.795 2399.405 ;
        RECT 3505.225 2399.125 3505.505 2399.405 ;
        RECT 3505.935 2399.125 3506.215 2399.405 ;
        RECT 3506.645 2399.125 3506.925 2399.405 ;
        RECT 3507.355 2399.125 3507.635 2399.405 ;
        RECT 3508.065 2399.125 3508.345 2399.405 ;
        RECT 3508.775 2399.125 3509.055 2399.405 ;
        RECT 3509.485 2399.125 3509.765 2399.405 ;
        RECT 3500.255 2398.415 3500.535 2398.695 ;
        RECT 3500.965 2398.415 3501.245 2398.695 ;
        RECT 3501.675 2398.415 3501.955 2398.695 ;
        RECT 3502.385 2398.415 3502.665 2398.695 ;
        RECT 3503.095 2398.415 3503.375 2398.695 ;
        RECT 3503.805 2398.415 3504.085 2398.695 ;
        RECT 3504.515 2398.415 3504.795 2398.695 ;
        RECT 3505.225 2398.415 3505.505 2398.695 ;
        RECT 3505.935 2398.415 3506.215 2398.695 ;
        RECT 3506.645 2398.415 3506.925 2398.695 ;
        RECT 3507.355 2398.415 3507.635 2398.695 ;
        RECT 3508.065 2398.415 3508.345 2398.695 ;
        RECT 3508.775 2398.415 3509.055 2398.695 ;
        RECT 3509.485 2398.415 3509.765 2398.695 ;
        RECT 3500.255 2397.705 3500.535 2397.985 ;
        RECT 3500.965 2397.705 3501.245 2397.985 ;
        RECT 3501.675 2397.705 3501.955 2397.985 ;
        RECT 3502.385 2397.705 3502.665 2397.985 ;
        RECT 3503.095 2397.705 3503.375 2397.985 ;
        RECT 3503.805 2397.705 3504.085 2397.985 ;
        RECT 3504.515 2397.705 3504.795 2397.985 ;
        RECT 3505.225 2397.705 3505.505 2397.985 ;
        RECT 3505.935 2397.705 3506.215 2397.985 ;
        RECT 3506.645 2397.705 3506.925 2397.985 ;
        RECT 3507.355 2397.705 3507.635 2397.985 ;
        RECT 3508.065 2397.705 3508.345 2397.985 ;
        RECT 3508.775 2397.705 3509.055 2397.985 ;
        RECT 3509.485 2397.705 3509.765 2397.985 ;
        RECT 3500.255 2396.995 3500.535 2397.275 ;
        RECT 3500.965 2396.995 3501.245 2397.275 ;
        RECT 3501.675 2396.995 3501.955 2397.275 ;
        RECT 3502.385 2396.995 3502.665 2397.275 ;
        RECT 3503.095 2396.995 3503.375 2397.275 ;
        RECT 3503.805 2396.995 3504.085 2397.275 ;
        RECT 3504.515 2396.995 3504.795 2397.275 ;
        RECT 3505.225 2396.995 3505.505 2397.275 ;
        RECT 3505.935 2396.995 3506.215 2397.275 ;
        RECT 3506.645 2396.995 3506.925 2397.275 ;
        RECT 3507.355 2396.995 3507.635 2397.275 ;
        RECT 3508.065 2396.995 3508.345 2397.275 ;
        RECT 3508.775 2396.995 3509.055 2397.275 ;
        RECT 3509.485 2396.995 3509.765 2397.275 ;
        RECT 3500.255 2396.285 3500.535 2396.565 ;
        RECT 3500.965 2396.285 3501.245 2396.565 ;
        RECT 3501.675 2396.285 3501.955 2396.565 ;
        RECT 3502.385 2396.285 3502.665 2396.565 ;
        RECT 3503.095 2396.285 3503.375 2396.565 ;
        RECT 3503.805 2396.285 3504.085 2396.565 ;
        RECT 3504.515 2396.285 3504.795 2396.565 ;
        RECT 3505.225 2396.285 3505.505 2396.565 ;
        RECT 3505.935 2396.285 3506.215 2396.565 ;
        RECT 3506.645 2396.285 3506.925 2396.565 ;
        RECT 3507.355 2396.285 3507.635 2396.565 ;
        RECT 3508.065 2396.285 3508.345 2396.565 ;
        RECT 3508.775 2396.285 3509.055 2396.565 ;
        RECT 3509.485 2396.285 3509.765 2396.565 ;
        RECT 3500.255 2395.575 3500.535 2395.855 ;
        RECT 3500.965 2395.575 3501.245 2395.855 ;
        RECT 3501.675 2395.575 3501.955 2395.855 ;
        RECT 3502.385 2395.575 3502.665 2395.855 ;
        RECT 3503.095 2395.575 3503.375 2395.855 ;
        RECT 3503.805 2395.575 3504.085 2395.855 ;
        RECT 3504.515 2395.575 3504.795 2395.855 ;
        RECT 3505.225 2395.575 3505.505 2395.855 ;
        RECT 3505.935 2395.575 3506.215 2395.855 ;
        RECT 3506.645 2395.575 3506.925 2395.855 ;
        RECT 3507.355 2395.575 3507.635 2395.855 ;
        RECT 3508.065 2395.575 3508.345 2395.855 ;
        RECT 3508.775 2395.575 3509.055 2395.855 ;
        RECT 3509.485 2395.575 3509.765 2395.855 ;
        RECT 3500.255 2394.865 3500.535 2395.145 ;
        RECT 3500.965 2394.865 3501.245 2395.145 ;
        RECT 3501.675 2394.865 3501.955 2395.145 ;
        RECT 3502.385 2394.865 3502.665 2395.145 ;
        RECT 3503.095 2394.865 3503.375 2395.145 ;
        RECT 3503.805 2394.865 3504.085 2395.145 ;
        RECT 3504.515 2394.865 3504.795 2395.145 ;
        RECT 3505.225 2394.865 3505.505 2395.145 ;
        RECT 3505.935 2394.865 3506.215 2395.145 ;
        RECT 3506.645 2394.865 3506.925 2395.145 ;
        RECT 3507.355 2394.865 3507.635 2395.145 ;
        RECT 3508.065 2394.865 3508.345 2395.145 ;
        RECT 3508.775 2394.865 3509.055 2395.145 ;
        RECT 3509.485 2394.865 3509.765 2395.145 ;
        RECT 3500.255 2394.155 3500.535 2394.435 ;
        RECT 3500.965 2394.155 3501.245 2394.435 ;
        RECT 3501.675 2394.155 3501.955 2394.435 ;
        RECT 3502.385 2394.155 3502.665 2394.435 ;
        RECT 3503.095 2394.155 3503.375 2394.435 ;
        RECT 3503.805 2394.155 3504.085 2394.435 ;
        RECT 3504.515 2394.155 3504.795 2394.435 ;
        RECT 3505.225 2394.155 3505.505 2394.435 ;
        RECT 3505.935 2394.155 3506.215 2394.435 ;
        RECT 3506.645 2394.155 3506.925 2394.435 ;
        RECT 3507.355 2394.155 3507.635 2394.435 ;
        RECT 3508.065 2394.155 3508.345 2394.435 ;
        RECT 3508.775 2394.155 3509.055 2394.435 ;
        RECT 3509.485 2394.155 3509.765 2394.435 ;
        RECT 3500.200 2390.270 3500.480 2390.550 ;
        RECT 3500.910 2390.270 3501.190 2390.550 ;
        RECT 3501.620 2390.270 3501.900 2390.550 ;
        RECT 3502.330 2390.270 3502.610 2390.550 ;
        RECT 3503.040 2390.270 3503.320 2390.550 ;
        RECT 3503.750 2390.270 3504.030 2390.550 ;
        RECT 3504.460 2390.270 3504.740 2390.550 ;
        RECT 3505.170 2390.270 3505.450 2390.550 ;
        RECT 3505.880 2390.270 3506.160 2390.550 ;
        RECT 3506.590 2390.270 3506.870 2390.550 ;
        RECT 3507.300 2390.270 3507.580 2390.550 ;
        RECT 3508.010 2390.270 3508.290 2390.550 ;
        RECT 3508.720 2390.270 3509.000 2390.550 ;
        RECT 3509.430 2390.270 3509.710 2390.550 ;
        RECT 3500.200 2389.560 3500.480 2389.840 ;
        RECT 3500.910 2389.560 3501.190 2389.840 ;
        RECT 3501.620 2389.560 3501.900 2389.840 ;
        RECT 3502.330 2389.560 3502.610 2389.840 ;
        RECT 3503.040 2389.560 3503.320 2389.840 ;
        RECT 3503.750 2389.560 3504.030 2389.840 ;
        RECT 3504.460 2389.560 3504.740 2389.840 ;
        RECT 3505.170 2389.560 3505.450 2389.840 ;
        RECT 3505.880 2389.560 3506.160 2389.840 ;
        RECT 3506.590 2389.560 3506.870 2389.840 ;
        RECT 3507.300 2389.560 3507.580 2389.840 ;
        RECT 3508.010 2389.560 3508.290 2389.840 ;
        RECT 3508.720 2389.560 3509.000 2389.840 ;
        RECT 3509.430 2389.560 3509.710 2389.840 ;
        RECT 3500.200 2388.850 3500.480 2389.130 ;
        RECT 3500.910 2388.850 3501.190 2389.130 ;
        RECT 3501.620 2388.850 3501.900 2389.130 ;
        RECT 3502.330 2388.850 3502.610 2389.130 ;
        RECT 3503.040 2388.850 3503.320 2389.130 ;
        RECT 3503.750 2388.850 3504.030 2389.130 ;
        RECT 3504.460 2388.850 3504.740 2389.130 ;
        RECT 3505.170 2388.850 3505.450 2389.130 ;
        RECT 3505.880 2388.850 3506.160 2389.130 ;
        RECT 3506.590 2388.850 3506.870 2389.130 ;
        RECT 3507.300 2388.850 3507.580 2389.130 ;
        RECT 3508.010 2388.850 3508.290 2389.130 ;
        RECT 3508.720 2388.850 3509.000 2389.130 ;
        RECT 3509.430 2388.850 3509.710 2389.130 ;
        RECT 3500.200 2388.140 3500.480 2388.420 ;
        RECT 3500.910 2388.140 3501.190 2388.420 ;
        RECT 3501.620 2388.140 3501.900 2388.420 ;
        RECT 3502.330 2388.140 3502.610 2388.420 ;
        RECT 3503.040 2388.140 3503.320 2388.420 ;
        RECT 3503.750 2388.140 3504.030 2388.420 ;
        RECT 3504.460 2388.140 3504.740 2388.420 ;
        RECT 3505.170 2388.140 3505.450 2388.420 ;
        RECT 3505.880 2388.140 3506.160 2388.420 ;
        RECT 3506.590 2388.140 3506.870 2388.420 ;
        RECT 3507.300 2388.140 3507.580 2388.420 ;
        RECT 3508.010 2388.140 3508.290 2388.420 ;
        RECT 3508.720 2388.140 3509.000 2388.420 ;
        RECT 3509.430 2388.140 3509.710 2388.420 ;
        RECT 3500.200 2387.430 3500.480 2387.710 ;
        RECT 3500.910 2387.430 3501.190 2387.710 ;
        RECT 3501.620 2387.430 3501.900 2387.710 ;
        RECT 3502.330 2387.430 3502.610 2387.710 ;
        RECT 3503.040 2387.430 3503.320 2387.710 ;
        RECT 3503.750 2387.430 3504.030 2387.710 ;
        RECT 3504.460 2387.430 3504.740 2387.710 ;
        RECT 3505.170 2387.430 3505.450 2387.710 ;
        RECT 3505.880 2387.430 3506.160 2387.710 ;
        RECT 3506.590 2387.430 3506.870 2387.710 ;
        RECT 3507.300 2387.430 3507.580 2387.710 ;
        RECT 3508.010 2387.430 3508.290 2387.710 ;
        RECT 3508.720 2387.430 3509.000 2387.710 ;
        RECT 3509.430 2387.430 3509.710 2387.710 ;
        RECT 3500.200 2386.720 3500.480 2387.000 ;
        RECT 3500.910 2386.720 3501.190 2387.000 ;
        RECT 3501.620 2386.720 3501.900 2387.000 ;
        RECT 3502.330 2386.720 3502.610 2387.000 ;
        RECT 3503.040 2386.720 3503.320 2387.000 ;
        RECT 3503.750 2386.720 3504.030 2387.000 ;
        RECT 3504.460 2386.720 3504.740 2387.000 ;
        RECT 3505.170 2386.720 3505.450 2387.000 ;
        RECT 3505.880 2386.720 3506.160 2387.000 ;
        RECT 3506.590 2386.720 3506.870 2387.000 ;
        RECT 3507.300 2386.720 3507.580 2387.000 ;
        RECT 3508.010 2386.720 3508.290 2387.000 ;
        RECT 3508.720 2386.720 3509.000 2387.000 ;
        RECT 3509.430 2386.720 3509.710 2387.000 ;
        RECT 3500.200 2386.010 3500.480 2386.290 ;
        RECT 3500.910 2386.010 3501.190 2386.290 ;
        RECT 3501.620 2386.010 3501.900 2386.290 ;
        RECT 3502.330 2386.010 3502.610 2386.290 ;
        RECT 3503.040 2386.010 3503.320 2386.290 ;
        RECT 3503.750 2386.010 3504.030 2386.290 ;
        RECT 3504.460 2386.010 3504.740 2386.290 ;
        RECT 3505.170 2386.010 3505.450 2386.290 ;
        RECT 3505.880 2386.010 3506.160 2386.290 ;
        RECT 3506.590 2386.010 3506.870 2386.290 ;
        RECT 3507.300 2386.010 3507.580 2386.290 ;
        RECT 3508.010 2386.010 3508.290 2386.290 ;
        RECT 3508.720 2386.010 3509.000 2386.290 ;
        RECT 3509.430 2386.010 3509.710 2386.290 ;
        RECT 3500.200 2385.300 3500.480 2385.580 ;
        RECT 3500.910 2385.300 3501.190 2385.580 ;
        RECT 3501.620 2385.300 3501.900 2385.580 ;
        RECT 3502.330 2385.300 3502.610 2385.580 ;
        RECT 3503.040 2385.300 3503.320 2385.580 ;
        RECT 3503.750 2385.300 3504.030 2385.580 ;
        RECT 3504.460 2385.300 3504.740 2385.580 ;
        RECT 3505.170 2385.300 3505.450 2385.580 ;
        RECT 3505.880 2385.300 3506.160 2385.580 ;
        RECT 3506.590 2385.300 3506.870 2385.580 ;
        RECT 3507.300 2385.300 3507.580 2385.580 ;
        RECT 3508.010 2385.300 3508.290 2385.580 ;
        RECT 3508.720 2385.300 3509.000 2385.580 ;
        RECT 3509.430 2385.300 3509.710 2385.580 ;
        RECT 3500.200 2384.590 3500.480 2384.870 ;
        RECT 3500.910 2384.590 3501.190 2384.870 ;
        RECT 3501.620 2384.590 3501.900 2384.870 ;
        RECT 3502.330 2384.590 3502.610 2384.870 ;
        RECT 3503.040 2384.590 3503.320 2384.870 ;
        RECT 3503.750 2384.590 3504.030 2384.870 ;
        RECT 3504.460 2384.590 3504.740 2384.870 ;
        RECT 3505.170 2384.590 3505.450 2384.870 ;
        RECT 3505.880 2384.590 3506.160 2384.870 ;
        RECT 3506.590 2384.590 3506.870 2384.870 ;
        RECT 3507.300 2384.590 3507.580 2384.870 ;
        RECT 3508.010 2384.590 3508.290 2384.870 ;
        RECT 3508.720 2384.590 3509.000 2384.870 ;
        RECT 3509.430 2384.590 3509.710 2384.870 ;
        RECT 3500.200 2383.880 3500.480 2384.160 ;
        RECT 3500.910 2383.880 3501.190 2384.160 ;
        RECT 3501.620 2383.880 3501.900 2384.160 ;
        RECT 3502.330 2383.880 3502.610 2384.160 ;
        RECT 3503.040 2383.880 3503.320 2384.160 ;
        RECT 3503.750 2383.880 3504.030 2384.160 ;
        RECT 3504.460 2383.880 3504.740 2384.160 ;
        RECT 3505.170 2383.880 3505.450 2384.160 ;
        RECT 3505.880 2383.880 3506.160 2384.160 ;
        RECT 3506.590 2383.880 3506.870 2384.160 ;
        RECT 3507.300 2383.880 3507.580 2384.160 ;
        RECT 3508.010 2383.880 3508.290 2384.160 ;
        RECT 3508.720 2383.880 3509.000 2384.160 ;
        RECT 3509.430 2383.880 3509.710 2384.160 ;
        RECT 3500.200 2383.170 3500.480 2383.450 ;
        RECT 3500.910 2383.170 3501.190 2383.450 ;
        RECT 3501.620 2383.170 3501.900 2383.450 ;
        RECT 3502.330 2383.170 3502.610 2383.450 ;
        RECT 3503.040 2383.170 3503.320 2383.450 ;
        RECT 3503.750 2383.170 3504.030 2383.450 ;
        RECT 3504.460 2383.170 3504.740 2383.450 ;
        RECT 3505.170 2383.170 3505.450 2383.450 ;
        RECT 3505.880 2383.170 3506.160 2383.450 ;
        RECT 3506.590 2383.170 3506.870 2383.450 ;
        RECT 3507.300 2383.170 3507.580 2383.450 ;
        RECT 3508.010 2383.170 3508.290 2383.450 ;
        RECT 3508.720 2383.170 3509.000 2383.450 ;
        RECT 3509.430 2383.170 3509.710 2383.450 ;
        RECT 3500.200 2382.460 3500.480 2382.740 ;
        RECT 3500.910 2382.460 3501.190 2382.740 ;
        RECT 3501.620 2382.460 3501.900 2382.740 ;
        RECT 3502.330 2382.460 3502.610 2382.740 ;
        RECT 3503.040 2382.460 3503.320 2382.740 ;
        RECT 3503.750 2382.460 3504.030 2382.740 ;
        RECT 3504.460 2382.460 3504.740 2382.740 ;
        RECT 3505.170 2382.460 3505.450 2382.740 ;
        RECT 3505.880 2382.460 3506.160 2382.740 ;
        RECT 3506.590 2382.460 3506.870 2382.740 ;
        RECT 3507.300 2382.460 3507.580 2382.740 ;
        RECT 3508.010 2382.460 3508.290 2382.740 ;
        RECT 3508.720 2382.460 3509.000 2382.740 ;
        RECT 3509.430 2382.460 3509.710 2382.740 ;
        RECT 3500.200 2381.750 3500.480 2382.030 ;
        RECT 3500.910 2381.750 3501.190 2382.030 ;
        RECT 3501.620 2381.750 3501.900 2382.030 ;
        RECT 3502.330 2381.750 3502.610 2382.030 ;
        RECT 3503.040 2381.750 3503.320 2382.030 ;
        RECT 3503.750 2381.750 3504.030 2382.030 ;
        RECT 3504.460 2381.750 3504.740 2382.030 ;
        RECT 3505.170 2381.750 3505.450 2382.030 ;
        RECT 3505.880 2381.750 3506.160 2382.030 ;
        RECT 3506.590 2381.750 3506.870 2382.030 ;
        RECT 3507.300 2381.750 3507.580 2382.030 ;
        RECT 3508.010 2381.750 3508.290 2382.030 ;
        RECT 3508.720 2381.750 3509.000 2382.030 ;
        RECT 3509.430 2381.750 3509.710 2382.030 ;
        RECT 369.330 2342.970 369.610 2343.250 ;
        RECT 370.040 2342.970 370.320 2343.250 ;
        RECT 370.750 2342.970 371.030 2343.250 ;
        RECT 371.460 2342.970 371.740 2343.250 ;
        RECT 372.170 2342.970 372.450 2343.250 ;
        RECT 372.880 2342.970 373.160 2343.250 ;
        RECT 373.590 2342.970 373.870 2343.250 ;
        RECT 374.300 2342.970 374.580 2343.250 ;
        RECT 375.010 2342.970 375.290 2343.250 ;
        RECT 375.720 2342.970 376.000 2343.250 ;
        RECT 376.430 2342.970 376.710 2343.250 ;
        RECT 369.330 2342.260 369.610 2342.540 ;
        RECT 370.040 2342.260 370.320 2342.540 ;
        RECT 370.750 2342.260 371.030 2342.540 ;
        RECT 371.460 2342.260 371.740 2342.540 ;
        RECT 372.170 2342.260 372.450 2342.540 ;
        RECT 372.880 2342.260 373.160 2342.540 ;
        RECT 373.590 2342.260 373.870 2342.540 ;
        RECT 374.300 2342.260 374.580 2342.540 ;
        RECT 375.010 2342.260 375.290 2342.540 ;
        RECT 375.720 2342.260 376.000 2342.540 ;
        RECT 376.430 2342.260 376.710 2342.540 ;
        RECT 369.330 2341.550 369.610 2341.830 ;
        RECT 370.040 2341.550 370.320 2341.830 ;
        RECT 370.750 2341.550 371.030 2341.830 ;
        RECT 371.460 2341.550 371.740 2341.830 ;
        RECT 372.170 2341.550 372.450 2341.830 ;
        RECT 372.880 2341.550 373.160 2341.830 ;
        RECT 373.590 2341.550 373.870 2341.830 ;
        RECT 374.300 2341.550 374.580 2341.830 ;
        RECT 375.010 2341.550 375.290 2341.830 ;
        RECT 375.720 2341.550 376.000 2341.830 ;
        RECT 376.430 2341.550 376.710 2341.830 ;
        RECT 369.330 2340.840 369.610 2341.120 ;
        RECT 370.040 2340.840 370.320 2341.120 ;
        RECT 370.750 2340.840 371.030 2341.120 ;
        RECT 371.460 2340.840 371.740 2341.120 ;
        RECT 372.170 2340.840 372.450 2341.120 ;
        RECT 372.880 2340.840 373.160 2341.120 ;
        RECT 373.590 2340.840 373.870 2341.120 ;
        RECT 374.300 2340.840 374.580 2341.120 ;
        RECT 375.010 2340.840 375.290 2341.120 ;
        RECT 375.720 2340.840 376.000 2341.120 ;
        RECT 376.430 2340.840 376.710 2341.120 ;
        RECT 369.330 2340.130 369.610 2340.410 ;
        RECT 370.040 2340.130 370.320 2340.410 ;
        RECT 370.750 2340.130 371.030 2340.410 ;
        RECT 371.460 2340.130 371.740 2340.410 ;
        RECT 372.170 2340.130 372.450 2340.410 ;
        RECT 372.880 2340.130 373.160 2340.410 ;
        RECT 373.590 2340.130 373.870 2340.410 ;
        RECT 374.300 2340.130 374.580 2340.410 ;
        RECT 375.010 2340.130 375.290 2340.410 ;
        RECT 375.720 2340.130 376.000 2340.410 ;
        RECT 376.430 2340.130 376.710 2340.410 ;
        RECT 369.330 2339.420 369.610 2339.700 ;
        RECT 370.040 2339.420 370.320 2339.700 ;
        RECT 370.750 2339.420 371.030 2339.700 ;
        RECT 371.460 2339.420 371.740 2339.700 ;
        RECT 372.170 2339.420 372.450 2339.700 ;
        RECT 372.880 2339.420 373.160 2339.700 ;
        RECT 373.590 2339.420 373.870 2339.700 ;
        RECT 374.300 2339.420 374.580 2339.700 ;
        RECT 375.010 2339.420 375.290 2339.700 ;
        RECT 375.720 2339.420 376.000 2339.700 ;
        RECT 376.430 2339.420 376.710 2339.700 ;
        RECT 369.330 2338.710 369.610 2338.990 ;
        RECT 370.040 2338.710 370.320 2338.990 ;
        RECT 370.750 2338.710 371.030 2338.990 ;
        RECT 371.460 2338.710 371.740 2338.990 ;
        RECT 372.170 2338.710 372.450 2338.990 ;
        RECT 372.880 2338.710 373.160 2338.990 ;
        RECT 373.590 2338.710 373.870 2338.990 ;
        RECT 374.300 2338.710 374.580 2338.990 ;
        RECT 375.010 2338.710 375.290 2338.990 ;
        RECT 375.720 2338.710 376.000 2338.990 ;
        RECT 376.430 2338.710 376.710 2338.990 ;
        RECT 369.330 2338.000 369.610 2338.280 ;
        RECT 370.040 2338.000 370.320 2338.280 ;
        RECT 370.750 2338.000 371.030 2338.280 ;
        RECT 371.460 2338.000 371.740 2338.280 ;
        RECT 372.170 2338.000 372.450 2338.280 ;
        RECT 372.880 2338.000 373.160 2338.280 ;
        RECT 373.590 2338.000 373.870 2338.280 ;
        RECT 374.300 2338.000 374.580 2338.280 ;
        RECT 375.010 2338.000 375.290 2338.280 ;
        RECT 375.720 2338.000 376.000 2338.280 ;
        RECT 376.430 2338.000 376.710 2338.280 ;
        RECT 369.330 2337.290 369.610 2337.570 ;
        RECT 370.040 2337.290 370.320 2337.570 ;
        RECT 370.750 2337.290 371.030 2337.570 ;
        RECT 371.460 2337.290 371.740 2337.570 ;
        RECT 372.170 2337.290 372.450 2337.570 ;
        RECT 372.880 2337.290 373.160 2337.570 ;
        RECT 373.590 2337.290 373.870 2337.570 ;
        RECT 374.300 2337.290 374.580 2337.570 ;
        RECT 375.010 2337.290 375.290 2337.570 ;
        RECT 375.720 2337.290 376.000 2337.570 ;
        RECT 376.430 2337.290 376.710 2337.570 ;
        RECT 369.330 2336.580 369.610 2336.860 ;
        RECT 370.040 2336.580 370.320 2336.860 ;
        RECT 370.750 2336.580 371.030 2336.860 ;
        RECT 371.460 2336.580 371.740 2336.860 ;
        RECT 372.170 2336.580 372.450 2336.860 ;
        RECT 372.880 2336.580 373.160 2336.860 ;
        RECT 373.590 2336.580 373.870 2336.860 ;
        RECT 374.300 2336.580 374.580 2336.860 ;
        RECT 375.010 2336.580 375.290 2336.860 ;
        RECT 375.720 2336.580 376.000 2336.860 ;
        RECT 376.430 2336.580 376.710 2336.860 ;
        RECT 369.330 2335.870 369.610 2336.150 ;
        RECT 370.040 2335.870 370.320 2336.150 ;
        RECT 370.750 2335.870 371.030 2336.150 ;
        RECT 371.460 2335.870 371.740 2336.150 ;
        RECT 372.170 2335.870 372.450 2336.150 ;
        RECT 372.880 2335.870 373.160 2336.150 ;
        RECT 373.590 2335.870 373.870 2336.150 ;
        RECT 374.300 2335.870 374.580 2336.150 ;
        RECT 375.010 2335.870 375.290 2336.150 ;
        RECT 375.720 2335.870 376.000 2336.150 ;
        RECT 376.430 2335.870 376.710 2336.150 ;
        RECT 369.330 2335.160 369.610 2335.440 ;
        RECT 370.040 2335.160 370.320 2335.440 ;
        RECT 370.750 2335.160 371.030 2335.440 ;
        RECT 371.460 2335.160 371.740 2335.440 ;
        RECT 372.170 2335.160 372.450 2335.440 ;
        RECT 372.880 2335.160 373.160 2335.440 ;
        RECT 373.590 2335.160 373.870 2335.440 ;
        RECT 374.300 2335.160 374.580 2335.440 ;
        RECT 375.010 2335.160 375.290 2335.440 ;
        RECT 375.720 2335.160 376.000 2335.440 ;
        RECT 376.430 2335.160 376.710 2335.440 ;
        RECT 369.330 2334.450 369.610 2334.730 ;
        RECT 370.040 2334.450 370.320 2334.730 ;
        RECT 370.750 2334.450 371.030 2334.730 ;
        RECT 371.460 2334.450 371.740 2334.730 ;
        RECT 372.170 2334.450 372.450 2334.730 ;
        RECT 372.880 2334.450 373.160 2334.730 ;
        RECT 373.590 2334.450 373.870 2334.730 ;
        RECT 374.300 2334.450 374.580 2334.730 ;
        RECT 375.010 2334.450 375.290 2334.730 ;
        RECT 375.720 2334.450 376.000 2334.730 ;
        RECT 376.430 2334.450 376.710 2334.730 ;
        RECT 369.275 2330.565 369.555 2330.845 ;
        RECT 369.985 2330.565 370.265 2330.845 ;
        RECT 370.695 2330.565 370.975 2330.845 ;
        RECT 371.405 2330.565 371.685 2330.845 ;
        RECT 372.115 2330.565 372.395 2330.845 ;
        RECT 372.825 2330.565 373.105 2330.845 ;
        RECT 373.535 2330.565 373.815 2330.845 ;
        RECT 374.245 2330.565 374.525 2330.845 ;
        RECT 374.955 2330.565 375.235 2330.845 ;
        RECT 375.665 2330.565 375.945 2330.845 ;
        RECT 376.375 2330.565 376.655 2330.845 ;
        RECT 369.275 2329.855 369.555 2330.135 ;
        RECT 369.985 2329.855 370.265 2330.135 ;
        RECT 370.695 2329.855 370.975 2330.135 ;
        RECT 371.405 2329.855 371.685 2330.135 ;
        RECT 372.115 2329.855 372.395 2330.135 ;
        RECT 372.825 2329.855 373.105 2330.135 ;
        RECT 373.535 2329.855 373.815 2330.135 ;
        RECT 374.245 2329.855 374.525 2330.135 ;
        RECT 374.955 2329.855 375.235 2330.135 ;
        RECT 375.665 2329.855 375.945 2330.135 ;
        RECT 376.375 2329.855 376.655 2330.135 ;
        RECT 369.275 2329.145 369.555 2329.425 ;
        RECT 369.985 2329.145 370.265 2329.425 ;
        RECT 370.695 2329.145 370.975 2329.425 ;
        RECT 371.405 2329.145 371.685 2329.425 ;
        RECT 372.115 2329.145 372.395 2329.425 ;
        RECT 372.825 2329.145 373.105 2329.425 ;
        RECT 373.535 2329.145 373.815 2329.425 ;
        RECT 374.245 2329.145 374.525 2329.425 ;
        RECT 374.955 2329.145 375.235 2329.425 ;
        RECT 375.665 2329.145 375.945 2329.425 ;
        RECT 376.375 2329.145 376.655 2329.425 ;
        RECT 369.275 2328.435 369.555 2328.715 ;
        RECT 369.985 2328.435 370.265 2328.715 ;
        RECT 370.695 2328.435 370.975 2328.715 ;
        RECT 371.405 2328.435 371.685 2328.715 ;
        RECT 372.115 2328.435 372.395 2328.715 ;
        RECT 372.825 2328.435 373.105 2328.715 ;
        RECT 373.535 2328.435 373.815 2328.715 ;
        RECT 374.245 2328.435 374.525 2328.715 ;
        RECT 374.955 2328.435 375.235 2328.715 ;
        RECT 375.665 2328.435 375.945 2328.715 ;
        RECT 376.375 2328.435 376.655 2328.715 ;
        RECT 369.275 2327.725 369.555 2328.005 ;
        RECT 369.985 2327.725 370.265 2328.005 ;
        RECT 370.695 2327.725 370.975 2328.005 ;
        RECT 371.405 2327.725 371.685 2328.005 ;
        RECT 372.115 2327.725 372.395 2328.005 ;
        RECT 372.825 2327.725 373.105 2328.005 ;
        RECT 373.535 2327.725 373.815 2328.005 ;
        RECT 374.245 2327.725 374.525 2328.005 ;
        RECT 374.955 2327.725 375.235 2328.005 ;
        RECT 375.665 2327.725 375.945 2328.005 ;
        RECT 376.375 2327.725 376.655 2328.005 ;
        RECT 369.275 2327.015 369.555 2327.295 ;
        RECT 369.985 2327.015 370.265 2327.295 ;
        RECT 370.695 2327.015 370.975 2327.295 ;
        RECT 371.405 2327.015 371.685 2327.295 ;
        RECT 372.115 2327.015 372.395 2327.295 ;
        RECT 372.825 2327.015 373.105 2327.295 ;
        RECT 373.535 2327.015 373.815 2327.295 ;
        RECT 374.245 2327.015 374.525 2327.295 ;
        RECT 374.955 2327.015 375.235 2327.295 ;
        RECT 375.665 2327.015 375.945 2327.295 ;
        RECT 376.375 2327.015 376.655 2327.295 ;
        RECT 369.275 2326.305 369.555 2326.585 ;
        RECT 369.985 2326.305 370.265 2326.585 ;
        RECT 370.695 2326.305 370.975 2326.585 ;
        RECT 371.405 2326.305 371.685 2326.585 ;
        RECT 372.115 2326.305 372.395 2326.585 ;
        RECT 372.825 2326.305 373.105 2326.585 ;
        RECT 373.535 2326.305 373.815 2326.585 ;
        RECT 374.245 2326.305 374.525 2326.585 ;
        RECT 374.955 2326.305 375.235 2326.585 ;
        RECT 375.665 2326.305 375.945 2326.585 ;
        RECT 376.375 2326.305 376.655 2326.585 ;
        RECT 369.275 2325.595 369.555 2325.875 ;
        RECT 369.985 2325.595 370.265 2325.875 ;
        RECT 370.695 2325.595 370.975 2325.875 ;
        RECT 371.405 2325.595 371.685 2325.875 ;
        RECT 372.115 2325.595 372.395 2325.875 ;
        RECT 372.825 2325.595 373.105 2325.875 ;
        RECT 373.535 2325.595 373.815 2325.875 ;
        RECT 374.245 2325.595 374.525 2325.875 ;
        RECT 374.955 2325.595 375.235 2325.875 ;
        RECT 375.665 2325.595 375.945 2325.875 ;
        RECT 376.375 2325.595 376.655 2325.875 ;
        RECT 369.275 2324.885 369.555 2325.165 ;
        RECT 369.985 2324.885 370.265 2325.165 ;
        RECT 370.695 2324.885 370.975 2325.165 ;
        RECT 371.405 2324.885 371.685 2325.165 ;
        RECT 372.115 2324.885 372.395 2325.165 ;
        RECT 372.825 2324.885 373.105 2325.165 ;
        RECT 373.535 2324.885 373.815 2325.165 ;
        RECT 374.245 2324.885 374.525 2325.165 ;
        RECT 374.955 2324.885 375.235 2325.165 ;
        RECT 375.665 2324.885 375.945 2325.165 ;
        RECT 376.375 2324.885 376.655 2325.165 ;
        RECT 369.275 2324.175 369.555 2324.455 ;
        RECT 369.985 2324.175 370.265 2324.455 ;
        RECT 370.695 2324.175 370.975 2324.455 ;
        RECT 371.405 2324.175 371.685 2324.455 ;
        RECT 372.115 2324.175 372.395 2324.455 ;
        RECT 372.825 2324.175 373.105 2324.455 ;
        RECT 373.535 2324.175 373.815 2324.455 ;
        RECT 374.245 2324.175 374.525 2324.455 ;
        RECT 374.955 2324.175 375.235 2324.455 ;
        RECT 375.665 2324.175 375.945 2324.455 ;
        RECT 376.375 2324.175 376.655 2324.455 ;
        RECT 369.275 2323.465 369.555 2323.745 ;
        RECT 369.985 2323.465 370.265 2323.745 ;
        RECT 370.695 2323.465 370.975 2323.745 ;
        RECT 371.405 2323.465 371.685 2323.745 ;
        RECT 372.115 2323.465 372.395 2323.745 ;
        RECT 372.825 2323.465 373.105 2323.745 ;
        RECT 373.535 2323.465 373.815 2323.745 ;
        RECT 374.245 2323.465 374.525 2323.745 ;
        RECT 374.955 2323.465 375.235 2323.745 ;
        RECT 375.665 2323.465 375.945 2323.745 ;
        RECT 376.375 2323.465 376.655 2323.745 ;
        RECT 369.275 2322.755 369.555 2323.035 ;
        RECT 369.985 2322.755 370.265 2323.035 ;
        RECT 370.695 2322.755 370.975 2323.035 ;
        RECT 371.405 2322.755 371.685 2323.035 ;
        RECT 372.115 2322.755 372.395 2323.035 ;
        RECT 372.825 2322.755 373.105 2323.035 ;
        RECT 373.535 2322.755 373.815 2323.035 ;
        RECT 374.245 2322.755 374.525 2323.035 ;
        RECT 374.955 2322.755 375.235 2323.035 ;
        RECT 375.665 2322.755 375.945 2323.035 ;
        RECT 376.375 2322.755 376.655 2323.035 ;
        RECT 369.275 2322.045 369.555 2322.325 ;
        RECT 369.985 2322.045 370.265 2322.325 ;
        RECT 370.695 2322.045 370.975 2322.325 ;
        RECT 371.405 2322.045 371.685 2322.325 ;
        RECT 372.115 2322.045 372.395 2322.325 ;
        RECT 372.825 2322.045 373.105 2322.325 ;
        RECT 373.535 2322.045 373.815 2322.325 ;
        RECT 374.245 2322.045 374.525 2322.325 ;
        RECT 374.955 2322.045 375.235 2322.325 ;
        RECT 375.665 2322.045 375.945 2322.325 ;
        RECT 376.375 2322.045 376.655 2322.325 ;
        RECT 369.275 2321.335 369.555 2321.615 ;
        RECT 369.985 2321.335 370.265 2321.615 ;
        RECT 370.695 2321.335 370.975 2321.615 ;
        RECT 371.405 2321.335 371.685 2321.615 ;
        RECT 372.115 2321.335 372.395 2321.615 ;
        RECT 372.825 2321.335 373.105 2321.615 ;
        RECT 373.535 2321.335 373.815 2321.615 ;
        RECT 374.245 2321.335 374.525 2321.615 ;
        RECT 374.955 2321.335 375.235 2321.615 ;
        RECT 375.665 2321.335 375.945 2321.615 ;
        RECT 376.375 2321.335 376.655 2321.615 ;
        RECT 369.275 2318.715 369.555 2318.995 ;
        RECT 369.985 2318.715 370.265 2318.995 ;
        RECT 370.695 2318.715 370.975 2318.995 ;
        RECT 371.405 2318.715 371.685 2318.995 ;
        RECT 372.115 2318.715 372.395 2318.995 ;
        RECT 372.825 2318.715 373.105 2318.995 ;
        RECT 373.535 2318.715 373.815 2318.995 ;
        RECT 374.245 2318.715 374.525 2318.995 ;
        RECT 374.955 2318.715 375.235 2318.995 ;
        RECT 375.665 2318.715 375.945 2318.995 ;
        RECT 376.375 2318.715 376.655 2318.995 ;
        RECT 369.275 2318.005 369.555 2318.285 ;
        RECT 369.985 2318.005 370.265 2318.285 ;
        RECT 370.695 2318.005 370.975 2318.285 ;
        RECT 371.405 2318.005 371.685 2318.285 ;
        RECT 372.115 2318.005 372.395 2318.285 ;
        RECT 372.825 2318.005 373.105 2318.285 ;
        RECT 373.535 2318.005 373.815 2318.285 ;
        RECT 374.245 2318.005 374.525 2318.285 ;
        RECT 374.955 2318.005 375.235 2318.285 ;
        RECT 375.665 2318.005 375.945 2318.285 ;
        RECT 376.375 2318.005 376.655 2318.285 ;
        RECT 369.275 2317.295 369.555 2317.575 ;
        RECT 369.985 2317.295 370.265 2317.575 ;
        RECT 370.695 2317.295 370.975 2317.575 ;
        RECT 371.405 2317.295 371.685 2317.575 ;
        RECT 372.115 2317.295 372.395 2317.575 ;
        RECT 372.825 2317.295 373.105 2317.575 ;
        RECT 373.535 2317.295 373.815 2317.575 ;
        RECT 374.245 2317.295 374.525 2317.575 ;
        RECT 374.955 2317.295 375.235 2317.575 ;
        RECT 375.665 2317.295 375.945 2317.575 ;
        RECT 376.375 2317.295 376.655 2317.575 ;
        RECT 369.275 2316.585 369.555 2316.865 ;
        RECT 369.985 2316.585 370.265 2316.865 ;
        RECT 370.695 2316.585 370.975 2316.865 ;
        RECT 371.405 2316.585 371.685 2316.865 ;
        RECT 372.115 2316.585 372.395 2316.865 ;
        RECT 372.825 2316.585 373.105 2316.865 ;
        RECT 373.535 2316.585 373.815 2316.865 ;
        RECT 374.245 2316.585 374.525 2316.865 ;
        RECT 374.955 2316.585 375.235 2316.865 ;
        RECT 375.665 2316.585 375.945 2316.865 ;
        RECT 376.375 2316.585 376.655 2316.865 ;
        RECT 369.275 2315.875 369.555 2316.155 ;
        RECT 369.985 2315.875 370.265 2316.155 ;
        RECT 370.695 2315.875 370.975 2316.155 ;
        RECT 371.405 2315.875 371.685 2316.155 ;
        RECT 372.115 2315.875 372.395 2316.155 ;
        RECT 372.825 2315.875 373.105 2316.155 ;
        RECT 373.535 2315.875 373.815 2316.155 ;
        RECT 374.245 2315.875 374.525 2316.155 ;
        RECT 374.955 2315.875 375.235 2316.155 ;
        RECT 375.665 2315.875 375.945 2316.155 ;
        RECT 376.375 2315.875 376.655 2316.155 ;
        RECT 369.275 2315.165 369.555 2315.445 ;
        RECT 369.985 2315.165 370.265 2315.445 ;
        RECT 370.695 2315.165 370.975 2315.445 ;
        RECT 371.405 2315.165 371.685 2315.445 ;
        RECT 372.115 2315.165 372.395 2315.445 ;
        RECT 372.825 2315.165 373.105 2315.445 ;
        RECT 373.535 2315.165 373.815 2315.445 ;
        RECT 374.245 2315.165 374.525 2315.445 ;
        RECT 374.955 2315.165 375.235 2315.445 ;
        RECT 375.665 2315.165 375.945 2315.445 ;
        RECT 376.375 2315.165 376.655 2315.445 ;
        RECT 369.275 2314.455 369.555 2314.735 ;
        RECT 369.985 2314.455 370.265 2314.735 ;
        RECT 370.695 2314.455 370.975 2314.735 ;
        RECT 371.405 2314.455 371.685 2314.735 ;
        RECT 372.115 2314.455 372.395 2314.735 ;
        RECT 372.825 2314.455 373.105 2314.735 ;
        RECT 373.535 2314.455 373.815 2314.735 ;
        RECT 374.245 2314.455 374.525 2314.735 ;
        RECT 374.955 2314.455 375.235 2314.735 ;
        RECT 375.665 2314.455 375.945 2314.735 ;
        RECT 376.375 2314.455 376.655 2314.735 ;
        RECT 369.275 2313.745 369.555 2314.025 ;
        RECT 369.985 2313.745 370.265 2314.025 ;
        RECT 370.695 2313.745 370.975 2314.025 ;
        RECT 371.405 2313.745 371.685 2314.025 ;
        RECT 372.115 2313.745 372.395 2314.025 ;
        RECT 372.825 2313.745 373.105 2314.025 ;
        RECT 373.535 2313.745 373.815 2314.025 ;
        RECT 374.245 2313.745 374.525 2314.025 ;
        RECT 374.955 2313.745 375.235 2314.025 ;
        RECT 375.665 2313.745 375.945 2314.025 ;
        RECT 376.375 2313.745 376.655 2314.025 ;
        RECT 369.275 2313.035 369.555 2313.315 ;
        RECT 369.985 2313.035 370.265 2313.315 ;
        RECT 370.695 2313.035 370.975 2313.315 ;
        RECT 371.405 2313.035 371.685 2313.315 ;
        RECT 372.115 2313.035 372.395 2313.315 ;
        RECT 372.825 2313.035 373.105 2313.315 ;
        RECT 373.535 2313.035 373.815 2313.315 ;
        RECT 374.245 2313.035 374.525 2313.315 ;
        RECT 374.955 2313.035 375.235 2313.315 ;
        RECT 375.665 2313.035 375.945 2313.315 ;
        RECT 376.375 2313.035 376.655 2313.315 ;
        RECT 369.275 2312.325 369.555 2312.605 ;
        RECT 369.985 2312.325 370.265 2312.605 ;
        RECT 370.695 2312.325 370.975 2312.605 ;
        RECT 371.405 2312.325 371.685 2312.605 ;
        RECT 372.115 2312.325 372.395 2312.605 ;
        RECT 372.825 2312.325 373.105 2312.605 ;
        RECT 373.535 2312.325 373.815 2312.605 ;
        RECT 374.245 2312.325 374.525 2312.605 ;
        RECT 374.955 2312.325 375.235 2312.605 ;
        RECT 375.665 2312.325 375.945 2312.605 ;
        RECT 376.375 2312.325 376.655 2312.605 ;
        RECT 369.275 2311.615 369.555 2311.895 ;
        RECT 369.985 2311.615 370.265 2311.895 ;
        RECT 370.695 2311.615 370.975 2311.895 ;
        RECT 371.405 2311.615 371.685 2311.895 ;
        RECT 372.115 2311.615 372.395 2311.895 ;
        RECT 372.825 2311.615 373.105 2311.895 ;
        RECT 373.535 2311.615 373.815 2311.895 ;
        RECT 374.245 2311.615 374.525 2311.895 ;
        RECT 374.955 2311.615 375.235 2311.895 ;
        RECT 375.665 2311.615 375.945 2311.895 ;
        RECT 376.375 2311.615 376.655 2311.895 ;
        RECT 369.275 2310.905 369.555 2311.185 ;
        RECT 369.985 2310.905 370.265 2311.185 ;
        RECT 370.695 2310.905 370.975 2311.185 ;
        RECT 371.405 2310.905 371.685 2311.185 ;
        RECT 372.115 2310.905 372.395 2311.185 ;
        RECT 372.825 2310.905 373.105 2311.185 ;
        RECT 373.535 2310.905 373.815 2311.185 ;
        RECT 374.245 2310.905 374.525 2311.185 ;
        RECT 374.955 2310.905 375.235 2311.185 ;
        RECT 375.665 2310.905 375.945 2311.185 ;
        RECT 376.375 2310.905 376.655 2311.185 ;
        RECT 369.275 2310.195 369.555 2310.475 ;
        RECT 369.985 2310.195 370.265 2310.475 ;
        RECT 370.695 2310.195 370.975 2310.475 ;
        RECT 371.405 2310.195 371.685 2310.475 ;
        RECT 372.115 2310.195 372.395 2310.475 ;
        RECT 372.825 2310.195 373.105 2310.475 ;
        RECT 373.535 2310.195 373.815 2310.475 ;
        RECT 374.245 2310.195 374.525 2310.475 ;
        RECT 374.955 2310.195 375.235 2310.475 ;
        RECT 375.665 2310.195 375.945 2310.475 ;
        RECT 376.375 2310.195 376.655 2310.475 ;
        RECT 369.275 2309.485 369.555 2309.765 ;
        RECT 369.985 2309.485 370.265 2309.765 ;
        RECT 370.695 2309.485 370.975 2309.765 ;
        RECT 371.405 2309.485 371.685 2309.765 ;
        RECT 372.115 2309.485 372.395 2309.765 ;
        RECT 372.825 2309.485 373.105 2309.765 ;
        RECT 373.535 2309.485 373.815 2309.765 ;
        RECT 374.245 2309.485 374.525 2309.765 ;
        RECT 374.955 2309.485 375.235 2309.765 ;
        RECT 375.665 2309.485 375.945 2309.765 ;
        RECT 376.375 2309.485 376.655 2309.765 ;
        RECT 369.275 2305.185 369.555 2305.465 ;
        RECT 369.985 2305.185 370.265 2305.465 ;
        RECT 370.695 2305.185 370.975 2305.465 ;
        RECT 371.405 2305.185 371.685 2305.465 ;
        RECT 372.115 2305.185 372.395 2305.465 ;
        RECT 372.825 2305.185 373.105 2305.465 ;
        RECT 373.535 2305.185 373.815 2305.465 ;
        RECT 374.245 2305.185 374.525 2305.465 ;
        RECT 374.955 2305.185 375.235 2305.465 ;
        RECT 375.665 2305.185 375.945 2305.465 ;
        RECT 376.375 2305.185 376.655 2305.465 ;
        RECT 369.275 2304.475 369.555 2304.755 ;
        RECT 369.985 2304.475 370.265 2304.755 ;
        RECT 370.695 2304.475 370.975 2304.755 ;
        RECT 371.405 2304.475 371.685 2304.755 ;
        RECT 372.115 2304.475 372.395 2304.755 ;
        RECT 372.825 2304.475 373.105 2304.755 ;
        RECT 373.535 2304.475 373.815 2304.755 ;
        RECT 374.245 2304.475 374.525 2304.755 ;
        RECT 374.955 2304.475 375.235 2304.755 ;
        RECT 375.665 2304.475 375.945 2304.755 ;
        RECT 376.375 2304.475 376.655 2304.755 ;
        RECT 369.275 2303.765 369.555 2304.045 ;
        RECT 369.985 2303.765 370.265 2304.045 ;
        RECT 370.695 2303.765 370.975 2304.045 ;
        RECT 371.405 2303.765 371.685 2304.045 ;
        RECT 372.115 2303.765 372.395 2304.045 ;
        RECT 372.825 2303.765 373.105 2304.045 ;
        RECT 373.535 2303.765 373.815 2304.045 ;
        RECT 374.245 2303.765 374.525 2304.045 ;
        RECT 374.955 2303.765 375.235 2304.045 ;
        RECT 375.665 2303.765 375.945 2304.045 ;
        RECT 376.375 2303.765 376.655 2304.045 ;
        RECT 369.275 2303.055 369.555 2303.335 ;
        RECT 369.985 2303.055 370.265 2303.335 ;
        RECT 370.695 2303.055 370.975 2303.335 ;
        RECT 371.405 2303.055 371.685 2303.335 ;
        RECT 372.115 2303.055 372.395 2303.335 ;
        RECT 372.825 2303.055 373.105 2303.335 ;
        RECT 373.535 2303.055 373.815 2303.335 ;
        RECT 374.245 2303.055 374.525 2303.335 ;
        RECT 374.955 2303.055 375.235 2303.335 ;
        RECT 375.665 2303.055 375.945 2303.335 ;
        RECT 376.375 2303.055 376.655 2303.335 ;
        RECT 369.275 2302.345 369.555 2302.625 ;
        RECT 369.985 2302.345 370.265 2302.625 ;
        RECT 370.695 2302.345 370.975 2302.625 ;
        RECT 371.405 2302.345 371.685 2302.625 ;
        RECT 372.115 2302.345 372.395 2302.625 ;
        RECT 372.825 2302.345 373.105 2302.625 ;
        RECT 373.535 2302.345 373.815 2302.625 ;
        RECT 374.245 2302.345 374.525 2302.625 ;
        RECT 374.955 2302.345 375.235 2302.625 ;
        RECT 375.665 2302.345 375.945 2302.625 ;
        RECT 376.375 2302.345 376.655 2302.625 ;
        RECT 369.275 2301.635 369.555 2301.915 ;
        RECT 369.985 2301.635 370.265 2301.915 ;
        RECT 370.695 2301.635 370.975 2301.915 ;
        RECT 371.405 2301.635 371.685 2301.915 ;
        RECT 372.115 2301.635 372.395 2301.915 ;
        RECT 372.825 2301.635 373.105 2301.915 ;
        RECT 373.535 2301.635 373.815 2301.915 ;
        RECT 374.245 2301.635 374.525 2301.915 ;
        RECT 374.955 2301.635 375.235 2301.915 ;
        RECT 375.665 2301.635 375.945 2301.915 ;
        RECT 376.375 2301.635 376.655 2301.915 ;
        RECT 369.275 2300.925 369.555 2301.205 ;
        RECT 369.985 2300.925 370.265 2301.205 ;
        RECT 370.695 2300.925 370.975 2301.205 ;
        RECT 371.405 2300.925 371.685 2301.205 ;
        RECT 372.115 2300.925 372.395 2301.205 ;
        RECT 372.825 2300.925 373.105 2301.205 ;
        RECT 373.535 2300.925 373.815 2301.205 ;
        RECT 374.245 2300.925 374.525 2301.205 ;
        RECT 374.955 2300.925 375.235 2301.205 ;
        RECT 375.665 2300.925 375.945 2301.205 ;
        RECT 376.375 2300.925 376.655 2301.205 ;
        RECT 369.275 2300.215 369.555 2300.495 ;
        RECT 369.985 2300.215 370.265 2300.495 ;
        RECT 370.695 2300.215 370.975 2300.495 ;
        RECT 371.405 2300.215 371.685 2300.495 ;
        RECT 372.115 2300.215 372.395 2300.495 ;
        RECT 372.825 2300.215 373.105 2300.495 ;
        RECT 373.535 2300.215 373.815 2300.495 ;
        RECT 374.245 2300.215 374.525 2300.495 ;
        RECT 374.955 2300.215 375.235 2300.495 ;
        RECT 375.665 2300.215 375.945 2300.495 ;
        RECT 376.375 2300.215 376.655 2300.495 ;
        RECT 369.275 2299.505 369.555 2299.785 ;
        RECT 369.985 2299.505 370.265 2299.785 ;
        RECT 370.695 2299.505 370.975 2299.785 ;
        RECT 371.405 2299.505 371.685 2299.785 ;
        RECT 372.115 2299.505 372.395 2299.785 ;
        RECT 372.825 2299.505 373.105 2299.785 ;
        RECT 373.535 2299.505 373.815 2299.785 ;
        RECT 374.245 2299.505 374.525 2299.785 ;
        RECT 374.955 2299.505 375.235 2299.785 ;
        RECT 375.665 2299.505 375.945 2299.785 ;
        RECT 376.375 2299.505 376.655 2299.785 ;
        RECT 369.275 2298.795 369.555 2299.075 ;
        RECT 369.985 2298.795 370.265 2299.075 ;
        RECT 370.695 2298.795 370.975 2299.075 ;
        RECT 371.405 2298.795 371.685 2299.075 ;
        RECT 372.115 2298.795 372.395 2299.075 ;
        RECT 372.825 2298.795 373.105 2299.075 ;
        RECT 373.535 2298.795 373.815 2299.075 ;
        RECT 374.245 2298.795 374.525 2299.075 ;
        RECT 374.955 2298.795 375.235 2299.075 ;
        RECT 375.665 2298.795 375.945 2299.075 ;
        RECT 376.375 2298.795 376.655 2299.075 ;
        RECT 369.275 2298.085 369.555 2298.365 ;
        RECT 369.985 2298.085 370.265 2298.365 ;
        RECT 370.695 2298.085 370.975 2298.365 ;
        RECT 371.405 2298.085 371.685 2298.365 ;
        RECT 372.115 2298.085 372.395 2298.365 ;
        RECT 372.825 2298.085 373.105 2298.365 ;
        RECT 373.535 2298.085 373.815 2298.365 ;
        RECT 374.245 2298.085 374.525 2298.365 ;
        RECT 374.955 2298.085 375.235 2298.365 ;
        RECT 375.665 2298.085 375.945 2298.365 ;
        RECT 376.375 2298.085 376.655 2298.365 ;
        RECT 369.275 2297.375 369.555 2297.655 ;
        RECT 369.985 2297.375 370.265 2297.655 ;
        RECT 370.695 2297.375 370.975 2297.655 ;
        RECT 371.405 2297.375 371.685 2297.655 ;
        RECT 372.115 2297.375 372.395 2297.655 ;
        RECT 372.825 2297.375 373.105 2297.655 ;
        RECT 373.535 2297.375 373.815 2297.655 ;
        RECT 374.245 2297.375 374.525 2297.655 ;
        RECT 374.955 2297.375 375.235 2297.655 ;
        RECT 375.665 2297.375 375.945 2297.655 ;
        RECT 376.375 2297.375 376.655 2297.655 ;
        RECT 369.275 2296.665 369.555 2296.945 ;
        RECT 369.985 2296.665 370.265 2296.945 ;
        RECT 370.695 2296.665 370.975 2296.945 ;
        RECT 371.405 2296.665 371.685 2296.945 ;
        RECT 372.115 2296.665 372.395 2296.945 ;
        RECT 372.825 2296.665 373.105 2296.945 ;
        RECT 373.535 2296.665 373.815 2296.945 ;
        RECT 374.245 2296.665 374.525 2296.945 ;
        RECT 374.955 2296.665 375.235 2296.945 ;
        RECT 375.665 2296.665 375.945 2296.945 ;
        RECT 376.375 2296.665 376.655 2296.945 ;
        RECT 369.275 2295.955 369.555 2296.235 ;
        RECT 369.985 2295.955 370.265 2296.235 ;
        RECT 370.695 2295.955 370.975 2296.235 ;
        RECT 371.405 2295.955 371.685 2296.235 ;
        RECT 372.115 2295.955 372.395 2296.235 ;
        RECT 372.825 2295.955 373.105 2296.235 ;
        RECT 373.535 2295.955 373.815 2296.235 ;
        RECT 374.245 2295.955 374.525 2296.235 ;
        RECT 374.955 2295.955 375.235 2296.235 ;
        RECT 375.665 2295.955 375.945 2296.235 ;
        RECT 376.375 2295.955 376.655 2296.235 ;
        RECT 369.275 2293.335 369.555 2293.615 ;
        RECT 369.985 2293.335 370.265 2293.615 ;
        RECT 370.695 2293.335 370.975 2293.615 ;
        RECT 371.405 2293.335 371.685 2293.615 ;
        RECT 372.115 2293.335 372.395 2293.615 ;
        RECT 372.825 2293.335 373.105 2293.615 ;
        RECT 373.535 2293.335 373.815 2293.615 ;
        RECT 374.245 2293.335 374.525 2293.615 ;
        RECT 374.955 2293.335 375.235 2293.615 ;
        RECT 375.665 2293.335 375.945 2293.615 ;
        RECT 376.375 2293.335 376.655 2293.615 ;
        RECT 369.275 2292.625 369.555 2292.905 ;
        RECT 369.985 2292.625 370.265 2292.905 ;
        RECT 370.695 2292.625 370.975 2292.905 ;
        RECT 371.405 2292.625 371.685 2292.905 ;
        RECT 372.115 2292.625 372.395 2292.905 ;
        RECT 372.825 2292.625 373.105 2292.905 ;
        RECT 373.535 2292.625 373.815 2292.905 ;
        RECT 374.245 2292.625 374.525 2292.905 ;
        RECT 374.955 2292.625 375.235 2292.905 ;
        RECT 375.665 2292.625 375.945 2292.905 ;
        RECT 376.375 2292.625 376.655 2292.905 ;
        RECT 369.275 2291.915 369.555 2292.195 ;
        RECT 369.985 2291.915 370.265 2292.195 ;
        RECT 370.695 2291.915 370.975 2292.195 ;
        RECT 371.405 2291.915 371.685 2292.195 ;
        RECT 372.115 2291.915 372.395 2292.195 ;
        RECT 372.825 2291.915 373.105 2292.195 ;
        RECT 373.535 2291.915 373.815 2292.195 ;
        RECT 374.245 2291.915 374.525 2292.195 ;
        RECT 374.955 2291.915 375.235 2292.195 ;
        RECT 375.665 2291.915 375.945 2292.195 ;
        RECT 376.375 2291.915 376.655 2292.195 ;
        RECT 369.275 2291.205 369.555 2291.485 ;
        RECT 369.985 2291.205 370.265 2291.485 ;
        RECT 370.695 2291.205 370.975 2291.485 ;
        RECT 371.405 2291.205 371.685 2291.485 ;
        RECT 372.115 2291.205 372.395 2291.485 ;
        RECT 372.825 2291.205 373.105 2291.485 ;
        RECT 373.535 2291.205 373.815 2291.485 ;
        RECT 374.245 2291.205 374.525 2291.485 ;
        RECT 374.955 2291.205 375.235 2291.485 ;
        RECT 375.665 2291.205 375.945 2291.485 ;
        RECT 376.375 2291.205 376.655 2291.485 ;
        RECT 369.275 2290.495 369.555 2290.775 ;
        RECT 369.985 2290.495 370.265 2290.775 ;
        RECT 370.695 2290.495 370.975 2290.775 ;
        RECT 371.405 2290.495 371.685 2290.775 ;
        RECT 372.115 2290.495 372.395 2290.775 ;
        RECT 372.825 2290.495 373.105 2290.775 ;
        RECT 373.535 2290.495 373.815 2290.775 ;
        RECT 374.245 2290.495 374.525 2290.775 ;
        RECT 374.955 2290.495 375.235 2290.775 ;
        RECT 375.665 2290.495 375.945 2290.775 ;
        RECT 376.375 2290.495 376.655 2290.775 ;
        RECT 369.275 2289.785 369.555 2290.065 ;
        RECT 369.985 2289.785 370.265 2290.065 ;
        RECT 370.695 2289.785 370.975 2290.065 ;
        RECT 371.405 2289.785 371.685 2290.065 ;
        RECT 372.115 2289.785 372.395 2290.065 ;
        RECT 372.825 2289.785 373.105 2290.065 ;
        RECT 373.535 2289.785 373.815 2290.065 ;
        RECT 374.245 2289.785 374.525 2290.065 ;
        RECT 374.955 2289.785 375.235 2290.065 ;
        RECT 375.665 2289.785 375.945 2290.065 ;
        RECT 376.375 2289.785 376.655 2290.065 ;
        RECT 369.275 2289.075 369.555 2289.355 ;
        RECT 369.985 2289.075 370.265 2289.355 ;
        RECT 370.695 2289.075 370.975 2289.355 ;
        RECT 371.405 2289.075 371.685 2289.355 ;
        RECT 372.115 2289.075 372.395 2289.355 ;
        RECT 372.825 2289.075 373.105 2289.355 ;
        RECT 373.535 2289.075 373.815 2289.355 ;
        RECT 374.245 2289.075 374.525 2289.355 ;
        RECT 374.955 2289.075 375.235 2289.355 ;
        RECT 375.665 2289.075 375.945 2289.355 ;
        RECT 376.375 2289.075 376.655 2289.355 ;
        RECT 369.275 2288.365 369.555 2288.645 ;
        RECT 369.985 2288.365 370.265 2288.645 ;
        RECT 370.695 2288.365 370.975 2288.645 ;
        RECT 371.405 2288.365 371.685 2288.645 ;
        RECT 372.115 2288.365 372.395 2288.645 ;
        RECT 372.825 2288.365 373.105 2288.645 ;
        RECT 373.535 2288.365 373.815 2288.645 ;
        RECT 374.245 2288.365 374.525 2288.645 ;
        RECT 374.955 2288.365 375.235 2288.645 ;
        RECT 375.665 2288.365 375.945 2288.645 ;
        RECT 376.375 2288.365 376.655 2288.645 ;
        RECT 369.275 2287.655 369.555 2287.935 ;
        RECT 369.985 2287.655 370.265 2287.935 ;
        RECT 370.695 2287.655 370.975 2287.935 ;
        RECT 371.405 2287.655 371.685 2287.935 ;
        RECT 372.115 2287.655 372.395 2287.935 ;
        RECT 372.825 2287.655 373.105 2287.935 ;
        RECT 373.535 2287.655 373.815 2287.935 ;
        RECT 374.245 2287.655 374.525 2287.935 ;
        RECT 374.955 2287.655 375.235 2287.935 ;
        RECT 375.665 2287.655 375.945 2287.935 ;
        RECT 376.375 2287.655 376.655 2287.935 ;
        RECT 369.275 2286.945 369.555 2287.225 ;
        RECT 369.985 2286.945 370.265 2287.225 ;
        RECT 370.695 2286.945 370.975 2287.225 ;
        RECT 371.405 2286.945 371.685 2287.225 ;
        RECT 372.115 2286.945 372.395 2287.225 ;
        RECT 372.825 2286.945 373.105 2287.225 ;
        RECT 373.535 2286.945 373.815 2287.225 ;
        RECT 374.245 2286.945 374.525 2287.225 ;
        RECT 374.955 2286.945 375.235 2287.225 ;
        RECT 375.665 2286.945 375.945 2287.225 ;
        RECT 376.375 2286.945 376.655 2287.225 ;
        RECT 369.275 2286.235 369.555 2286.515 ;
        RECT 369.985 2286.235 370.265 2286.515 ;
        RECT 370.695 2286.235 370.975 2286.515 ;
        RECT 371.405 2286.235 371.685 2286.515 ;
        RECT 372.115 2286.235 372.395 2286.515 ;
        RECT 372.825 2286.235 373.105 2286.515 ;
        RECT 373.535 2286.235 373.815 2286.515 ;
        RECT 374.245 2286.235 374.525 2286.515 ;
        RECT 374.955 2286.235 375.235 2286.515 ;
        RECT 375.665 2286.235 375.945 2286.515 ;
        RECT 376.375 2286.235 376.655 2286.515 ;
        RECT 369.275 2285.525 369.555 2285.805 ;
        RECT 369.985 2285.525 370.265 2285.805 ;
        RECT 370.695 2285.525 370.975 2285.805 ;
        RECT 371.405 2285.525 371.685 2285.805 ;
        RECT 372.115 2285.525 372.395 2285.805 ;
        RECT 372.825 2285.525 373.105 2285.805 ;
        RECT 373.535 2285.525 373.815 2285.805 ;
        RECT 374.245 2285.525 374.525 2285.805 ;
        RECT 374.955 2285.525 375.235 2285.805 ;
        RECT 375.665 2285.525 375.945 2285.805 ;
        RECT 376.375 2285.525 376.655 2285.805 ;
        RECT 369.275 2284.815 369.555 2285.095 ;
        RECT 369.985 2284.815 370.265 2285.095 ;
        RECT 370.695 2284.815 370.975 2285.095 ;
        RECT 371.405 2284.815 371.685 2285.095 ;
        RECT 372.115 2284.815 372.395 2285.095 ;
        RECT 372.825 2284.815 373.105 2285.095 ;
        RECT 373.535 2284.815 373.815 2285.095 ;
        RECT 374.245 2284.815 374.525 2285.095 ;
        RECT 374.955 2284.815 375.235 2285.095 ;
        RECT 375.665 2284.815 375.945 2285.095 ;
        RECT 376.375 2284.815 376.655 2285.095 ;
        RECT 369.275 2284.105 369.555 2284.385 ;
        RECT 369.985 2284.105 370.265 2284.385 ;
        RECT 370.695 2284.105 370.975 2284.385 ;
        RECT 371.405 2284.105 371.685 2284.385 ;
        RECT 372.115 2284.105 372.395 2284.385 ;
        RECT 372.825 2284.105 373.105 2284.385 ;
        RECT 373.535 2284.105 373.815 2284.385 ;
        RECT 374.245 2284.105 374.525 2284.385 ;
        RECT 374.955 2284.105 375.235 2284.385 ;
        RECT 375.665 2284.105 375.945 2284.385 ;
        RECT 376.375 2284.105 376.655 2284.385 ;
        RECT 369.330 2280.190 369.610 2280.470 ;
        RECT 370.040 2280.190 370.320 2280.470 ;
        RECT 370.750 2280.190 371.030 2280.470 ;
        RECT 371.460 2280.190 371.740 2280.470 ;
        RECT 372.170 2280.190 372.450 2280.470 ;
        RECT 372.880 2280.190 373.160 2280.470 ;
        RECT 373.590 2280.190 373.870 2280.470 ;
        RECT 374.300 2280.190 374.580 2280.470 ;
        RECT 375.010 2280.190 375.290 2280.470 ;
        RECT 375.720 2280.190 376.000 2280.470 ;
        RECT 376.430 2280.190 376.710 2280.470 ;
        RECT 369.330 2279.480 369.610 2279.760 ;
        RECT 370.040 2279.480 370.320 2279.760 ;
        RECT 370.750 2279.480 371.030 2279.760 ;
        RECT 371.460 2279.480 371.740 2279.760 ;
        RECT 372.170 2279.480 372.450 2279.760 ;
        RECT 372.880 2279.480 373.160 2279.760 ;
        RECT 373.590 2279.480 373.870 2279.760 ;
        RECT 374.300 2279.480 374.580 2279.760 ;
        RECT 375.010 2279.480 375.290 2279.760 ;
        RECT 375.720 2279.480 376.000 2279.760 ;
        RECT 376.430 2279.480 376.710 2279.760 ;
        RECT 369.330 2278.770 369.610 2279.050 ;
        RECT 370.040 2278.770 370.320 2279.050 ;
        RECT 370.750 2278.770 371.030 2279.050 ;
        RECT 371.460 2278.770 371.740 2279.050 ;
        RECT 372.170 2278.770 372.450 2279.050 ;
        RECT 372.880 2278.770 373.160 2279.050 ;
        RECT 373.590 2278.770 373.870 2279.050 ;
        RECT 374.300 2278.770 374.580 2279.050 ;
        RECT 375.010 2278.770 375.290 2279.050 ;
        RECT 375.720 2278.770 376.000 2279.050 ;
        RECT 376.430 2278.770 376.710 2279.050 ;
        RECT 369.330 2278.060 369.610 2278.340 ;
        RECT 370.040 2278.060 370.320 2278.340 ;
        RECT 370.750 2278.060 371.030 2278.340 ;
        RECT 371.460 2278.060 371.740 2278.340 ;
        RECT 372.170 2278.060 372.450 2278.340 ;
        RECT 372.880 2278.060 373.160 2278.340 ;
        RECT 373.590 2278.060 373.870 2278.340 ;
        RECT 374.300 2278.060 374.580 2278.340 ;
        RECT 375.010 2278.060 375.290 2278.340 ;
        RECT 375.720 2278.060 376.000 2278.340 ;
        RECT 376.430 2278.060 376.710 2278.340 ;
        RECT 369.330 2277.350 369.610 2277.630 ;
        RECT 370.040 2277.350 370.320 2277.630 ;
        RECT 370.750 2277.350 371.030 2277.630 ;
        RECT 371.460 2277.350 371.740 2277.630 ;
        RECT 372.170 2277.350 372.450 2277.630 ;
        RECT 372.880 2277.350 373.160 2277.630 ;
        RECT 373.590 2277.350 373.870 2277.630 ;
        RECT 374.300 2277.350 374.580 2277.630 ;
        RECT 375.010 2277.350 375.290 2277.630 ;
        RECT 375.720 2277.350 376.000 2277.630 ;
        RECT 376.430 2277.350 376.710 2277.630 ;
        RECT 369.330 2276.640 369.610 2276.920 ;
        RECT 370.040 2276.640 370.320 2276.920 ;
        RECT 370.750 2276.640 371.030 2276.920 ;
        RECT 371.460 2276.640 371.740 2276.920 ;
        RECT 372.170 2276.640 372.450 2276.920 ;
        RECT 372.880 2276.640 373.160 2276.920 ;
        RECT 373.590 2276.640 373.870 2276.920 ;
        RECT 374.300 2276.640 374.580 2276.920 ;
        RECT 375.010 2276.640 375.290 2276.920 ;
        RECT 375.720 2276.640 376.000 2276.920 ;
        RECT 376.430 2276.640 376.710 2276.920 ;
        RECT 369.330 2275.930 369.610 2276.210 ;
        RECT 370.040 2275.930 370.320 2276.210 ;
        RECT 370.750 2275.930 371.030 2276.210 ;
        RECT 371.460 2275.930 371.740 2276.210 ;
        RECT 372.170 2275.930 372.450 2276.210 ;
        RECT 372.880 2275.930 373.160 2276.210 ;
        RECT 373.590 2275.930 373.870 2276.210 ;
        RECT 374.300 2275.930 374.580 2276.210 ;
        RECT 375.010 2275.930 375.290 2276.210 ;
        RECT 375.720 2275.930 376.000 2276.210 ;
        RECT 376.430 2275.930 376.710 2276.210 ;
        RECT 369.330 2275.220 369.610 2275.500 ;
        RECT 370.040 2275.220 370.320 2275.500 ;
        RECT 370.750 2275.220 371.030 2275.500 ;
        RECT 371.460 2275.220 371.740 2275.500 ;
        RECT 372.170 2275.220 372.450 2275.500 ;
        RECT 372.880 2275.220 373.160 2275.500 ;
        RECT 373.590 2275.220 373.870 2275.500 ;
        RECT 374.300 2275.220 374.580 2275.500 ;
        RECT 375.010 2275.220 375.290 2275.500 ;
        RECT 375.720 2275.220 376.000 2275.500 ;
        RECT 376.430 2275.220 376.710 2275.500 ;
        RECT 369.330 2274.510 369.610 2274.790 ;
        RECT 370.040 2274.510 370.320 2274.790 ;
        RECT 370.750 2274.510 371.030 2274.790 ;
        RECT 371.460 2274.510 371.740 2274.790 ;
        RECT 372.170 2274.510 372.450 2274.790 ;
        RECT 372.880 2274.510 373.160 2274.790 ;
        RECT 373.590 2274.510 373.870 2274.790 ;
        RECT 374.300 2274.510 374.580 2274.790 ;
        RECT 375.010 2274.510 375.290 2274.790 ;
        RECT 375.720 2274.510 376.000 2274.790 ;
        RECT 376.430 2274.510 376.710 2274.790 ;
        RECT 369.330 2273.800 369.610 2274.080 ;
        RECT 370.040 2273.800 370.320 2274.080 ;
        RECT 370.750 2273.800 371.030 2274.080 ;
        RECT 371.460 2273.800 371.740 2274.080 ;
        RECT 372.170 2273.800 372.450 2274.080 ;
        RECT 372.880 2273.800 373.160 2274.080 ;
        RECT 373.590 2273.800 373.870 2274.080 ;
        RECT 374.300 2273.800 374.580 2274.080 ;
        RECT 375.010 2273.800 375.290 2274.080 ;
        RECT 375.720 2273.800 376.000 2274.080 ;
        RECT 376.430 2273.800 376.710 2274.080 ;
        RECT 369.330 2273.090 369.610 2273.370 ;
        RECT 370.040 2273.090 370.320 2273.370 ;
        RECT 370.750 2273.090 371.030 2273.370 ;
        RECT 371.460 2273.090 371.740 2273.370 ;
        RECT 372.170 2273.090 372.450 2273.370 ;
        RECT 372.880 2273.090 373.160 2273.370 ;
        RECT 373.590 2273.090 373.870 2273.370 ;
        RECT 374.300 2273.090 374.580 2273.370 ;
        RECT 375.010 2273.090 375.290 2273.370 ;
        RECT 375.720 2273.090 376.000 2273.370 ;
        RECT 376.430 2273.090 376.710 2273.370 ;
        RECT 369.330 2272.380 369.610 2272.660 ;
        RECT 370.040 2272.380 370.320 2272.660 ;
        RECT 370.750 2272.380 371.030 2272.660 ;
        RECT 371.460 2272.380 371.740 2272.660 ;
        RECT 372.170 2272.380 372.450 2272.660 ;
        RECT 372.880 2272.380 373.160 2272.660 ;
        RECT 373.590 2272.380 373.870 2272.660 ;
        RECT 374.300 2272.380 374.580 2272.660 ;
        RECT 375.010 2272.380 375.290 2272.660 ;
        RECT 375.720 2272.380 376.000 2272.660 ;
        RECT 376.430 2272.380 376.710 2272.660 ;
        RECT 369.330 2271.670 369.610 2271.950 ;
        RECT 370.040 2271.670 370.320 2271.950 ;
        RECT 370.750 2271.670 371.030 2271.950 ;
        RECT 371.460 2271.670 371.740 2271.950 ;
        RECT 372.170 2271.670 372.450 2271.950 ;
        RECT 372.880 2271.670 373.160 2271.950 ;
        RECT 373.590 2271.670 373.870 2271.950 ;
        RECT 374.300 2271.670 374.580 2271.950 ;
        RECT 375.010 2271.670 375.290 2271.950 ;
        RECT 375.720 2271.670 376.000 2271.950 ;
        RECT 376.430 2271.670 376.710 2271.950 ;
        RECT 3512.200 2238.050 3512.480 2238.330 ;
        RECT 3512.910 2238.050 3513.190 2238.330 ;
        RECT 3513.620 2238.050 3513.900 2238.330 ;
        RECT 3514.330 2238.050 3514.610 2238.330 ;
        RECT 3515.040 2238.050 3515.320 2238.330 ;
        RECT 3515.750 2238.050 3516.030 2238.330 ;
        RECT 3516.460 2238.050 3516.740 2238.330 ;
        RECT 3517.170 2238.050 3517.450 2238.330 ;
        RECT 3517.880 2238.050 3518.160 2238.330 ;
        RECT 3518.590 2238.050 3518.870 2238.330 ;
        RECT 3519.300 2238.050 3519.580 2238.330 ;
        RECT 3520.010 2238.050 3520.290 2238.330 ;
        RECT 3520.720 2238.050 3521.000 2238.330 ;
        RECT 3521.430 2238.050 3521.710 2238.330 ;
        RECT 3512.200 2237.340 3512.480 2237.620 ;
        RECT 3512.910 2237.340 3513.190 2237.620 ;
        RECT 3513.620 2237.340 3513.900 2237.620 ;
        RECT 3514.330 2237.340 3514.610 2237.620 ;
        RECT 3515.040 2237.340 3515.320 2237.620 ;
        RECT 3515.750 2237.340 3516.030 2237.620 ;
        RECT 3516.460 2237.340 3516.740 2237.620 ;
        RECT 3517.170 2237.340 3517.450 2237.620 ;
        RECT 3517.880 2237.340 3518.160 2237.620 ;
        RECT 3518.590 2237.340 3518.870 2237.620 ;
        RECT 3519.300 2237.340 3519.580 2237.620 ;
        RECT 3520.010 2237.340 3520.290 2237.620 ;
        RECT 3520.720 2237.340 3521.000 2237.620 ;
        RECT 3521.430 2237.340 3521.710 2237.620 ;
        RECT 3512.200 2236.630 3512.480 2236.910 ;
        RECT 3512.910 2236.630 3513.190 2236.910 ;
        RECT 3513.620 2236.630 3513.900 2236.910 ;
        RECT 3514.330 2236.630 3514.610 2236.910 ;
        RECT 3515.040 2236.630 3515.320 2236.910 ;
        RECT 3515.750 2236.630 3516.030 2236.910 ;
        RECT 3516.460 2236.630 3516.740 2236.910 ;
        RECT 3517.170 2236.630 3517.450 2236.910 ;
        RECT 3517.880 2236.630 3518.160 2236.910 ;
        RECT 3518.590 2236.630 3518.870 2236.910 ;
        RECT 3519.300 2236.630 3519.580 2236.910 ;
        RECT 3520.010 2236.630 3520.290 2236.910 ;
        RECT 3520.720 2236.630 3521.000 2236.910 ;
        RECT 3521.430 2236.630 3521.710 2236.910 ;
        RECT 3512.200 2235.920 3512.480 2236.200 ;
        RECT 3512.910 2235.920 3513.190 2236.200 ;
        RECT 3513.620 2235.920 3513.900 2236.200 ;
        RECT 3514.330 2235.920 3514.610 2236.200 ;
        RECT 3515.040 2235.920 3515.320 2236.200 ;
        RECT 3515.750 2235.920 3516.030 2236.200 ;
        RECT 3516.460 2235.920 3516.740 2236.200 ;
        RECT 3517.170 2235.920 3517.450 2236.200 ;
        RECT 3517.880 2235.920 3518.160 2236.200 ;
        RECT 3518.590 2235.920 3518.870 2236.200 ;
        RECT 3519.300 2235.920 3519.580 2236.200 ;
        RECT 3520.010 2235.920 3520.290 2236.200 ;
        RECT 3520.720 2235.920 3521.000 2236.200 ;
        RECT 3521.430 2235.920 3521.710 2236.200 ;
        RECT 3512.200 2235.210 3512.480 2235.490 ;
        RECT 3512.910 2235.210 3513.190 2235.490 ;
        RECT 3513.620 2235.210 3513.900 2235.490 ;
        RECT 3514.330 2235.210 3514.610 2235.490 ;
        RECT 3515.040 2235.210 3515.320 2235.490 ;
        RECT 3515.750 2235.210 3516.030 2235.490 ;
        RECT 3516.460 2235.210 3516.740 2235.490 ;
        RECT 3517.170 2235.210 3517.450 2235.490 ;
        RECT 3517.880 2235.210 3518.160 2235.490 ;
        RECT 3518.590 2235.210 3518.870 2235.490 ;
        RECT 3519.300 2235.210 3519.580 2235.490 ;
        RECT 3520.010 2235.210 3520.290 2235.490 ;
        RECT 3520.720 2235.210 3521.000 2235.490 ;
        RECT 3521.430 2235.210 3521.710 2235.490 ;
        RECT 3512.200 2234.500 3512.480 2234.780 ;
        RECT 3512.910 2234.500 3513.190 2234.780 ;
        RECT 3513.620 2234.500 3513.900 2234.780 ;
        RECT 3514.330 2234.500 3514.610 2234.780 ;
        RECT 3515.040 2234.500 3515.320 2234.780 ;
        RECT 3515.750 2234.500 3516.030 2234.780 ;
        RECT 3516.460 2234.500 3516.740 2234.780 ;
        RECT 3517.170 2234.500 3517.450 2234.780 ;
        RECT 3517.880 2234.500 3518.160 2234.780 ;
        RECT 3518.590 2234.500 3518.870 2234.780 ;
        RECT 3519.300 2234.500 3519.580 2234.780 ;
        RECT 3520.010 2234.500 3520.290 2234.780 ;
        RECT 3520.720 2234.500 3521.000 2234.780 ;
        RECT 3521.430 2234.500 3521.710 2234.780 ;
        RECT 3512.200 2233.790 3512.480 2234.070 ;
        RECT 3512.910 2233.790 3513.190 2234.070 ;
        RECT 3513.620 2233.790 3513.900 2234.070 ;
        RECT 3514.330 2233.790 3514.610 2234.070 ;
        RECT 3515.040 2233.790 3515.320 2234.070 ;
        RECT 3515.750 2233.790 3516.030 2234.070 ;
        RECT 3516.460 2233.790 3516.740 2234.070 ;
        RECT 3517.170 2233.790 3517.450 2234.070 ;
        RECT 3517.880 2233.790 3518.160 2234.070 ;
        RECT 3518.590 2233.790 3518.870 2234.070 ;
        RECT 3519.300 2233.790 3519.580 2234.070 ;
        RECT 3520.010 2233.790 3520.290 2234.070 ;
        RECT 3520.720 2233.790 3521.000 2234.070 ;
        RECT 3521.430 2233.790 3521.710 2234.070 ;
        RECT 3512.200 2233.080 3512.480 2233.360 ;
        RECT 3512.910 2233.080 3513.190 2233.360 ;
        RECT 3513.620 2233.080 3513.900 2233.360 ;
        RECT 3514.330 2233.080 3514.610 2233.360 ;
        RECT 3515.040 2233.080 3515.320 2233.360 ;
        RECT 3515.750 2233.080 3516.030 2233.360 ;
        RECT 3516.460 2233.080 3516.740 2233.360 ;
        RECT 3517.170 2233.080 3517.450 2233.360 ;
        RECT 3517.880 2233.080 3518.160 2233.360 ;
        RECT 3518.590 2233.080 3518.870 2233.360 ;
        RECT 3519.300 2233.080 3519.580 2233.360 ;
        RECT 3520.010 2233.080 3520.290 2233.360 ;
        RECT 3520.720 2233.080 3521.000 2233.360 ;
        RECT 3521.430 2233.080 3521.710 2233.360 ;
        RECT 3512.200 2232.370 3512.480 2232.650 ;
        RECT 3512.910 2232.370 3513.190 2232.650 ;
        RECT 3513.620 2232.370 3513.900 2232.650 ;
        RECT 3514.330 2232.370 3514.610 2232.650 ;
        RECT 3515.040 2232.370 3515.320 2232.650 ;
        RECT 3515.750 2232.370 3516.030 2232.650 ;
        RECT 3516.460 2232.370 3516.740 2232.650 ;
        RECT 3517.170 2232.370 3517.450 2232.650 ;
        RECT 3517.880 2232.370 3518.160 2232.650 ;
        RECT 3518.590 2232.370 3518.870 2232.650 ;
        RECT 3519.300 2232.370 3519.580 2232.650 ;
        RECT 3520.010 2232.370 3520.290 2232.650 ;
        RECT 3520.720 2232.370 3521.000 2232.650 ;
        RECT 3521.430 2232.370 3521.710 2232.650 ;
        RECT 3512.200 2231.660 3512.480 2231.940 ;
        RECT 3512.910 2231.660 3513.190 2231.940 ;
        RECT 3513.620 2231.660 3513.900 2231.940 ;
        RECT 3514.330 2231.660 3514.610 2231.940 ;
        RECT 3515.040 2231.660 3515.320 2231.940 ;
        RECT 3515.750 2231.660 3516.030 2231.940 ;
        RECT 3516.460 2231.660 3516.740 2231.940 ;
        RECT 3517.170 2231.660 3517.450 2231.940 ;
        RECT 3517.880 2231.660 3518.160 2231.940 ;
        RECT 3518.590 2231.660 3518.870 2231.940 ;
        RECT 3519.300 2231.660 3519.580 2231.940 ;
        RECT 3520.010 2231.660 3520.290 2231.940 ;
        RECT 3520.720 2231.660 3521.000 2231.940 ;
        RECT 3521.430 2231.660 3521.710 2231.940 ;
        RECT 3512.200 2230.950 3512.480 2231.230 ;
        RECT 3512.910 2230.950 3513.190 2231.230 ;
        RECT 3513.620 2230.950 3513.900 2231.230 ;
        RECT 3514.330 2230.950 3514.610 2231.230 ;
        RECT 3515.040 2230.950 3515.320 2231.230 ;
        RECT 3515.750 2230.950 3516.030 2231.230 ;
        RECT 3516.460 2230.950 3516.740 2231.230 ;
        RECT 3517.170 2230.950 3517.450 2231.230 ;
        RECT 3517.880 2230.950 3518.160 2231.230 ;
        RECT 3518.590 2230.950 3518.870 2231.230 ;
        RECT 3519.300 2230.950 3519.580 2231.230 ;
        RECT 3520.010 2230.950 3520.290 2231.230 ;
        RECT 3520.720 2230.950 3521.000 2231.230 ;
        RECT 3521.430 2230.950 3521.710 2231.230 ;
        RECT 3512.200 2230.240 3512.480 2230.520 ;
        RECT 3512.910 2230.240 3513.190 2230.520 ;
        RECT 3513.620 2230.240 3513.900 2230.520 ;
        RECT 3514.330 2230.240 3514.610 2230.520 ;
        RECT 3515.040 2230.240 3515.320 2230.520 ;
        RECT 3515.750 2230.240 3516.030 2230.520 ;
        RECT 3516.460 2230.240 3516.740 2230.520 ;
        RECT 3517.170 2230.240 3517.450 2230.520 ;
        RECT 3517.880 2230.240 3518.160 2230.520 ;
        RECT 3518.590 2230.240 3518.870 2230.520 ;
        RECT 3519.300 2230.240 3519.580 2230.520 ;
        RECT 3520.010 2230.240 3520.290 2230.520 ;
        RECT 3520.720 2230.240 3521.000 2230.520 ;
        RECT 3521.430 2230.240 3521.710 2230.520 ;
        RECT 3512.200 2229.530 3512.480 2229.810 ;
        RECT 3512.910 2229.530 3513.190 2229.810 ;
        RECT 3513.620 2229.530 3513.900 2229.810 ;
        RECT 3514.330 2229.530 3514.610 2229.810 ;
        RECT 3515.040 2229.530 3515.320 2229.810 ;
        RECT 3515.750 2229.530 3516.030 2229.810 ;
        RECT 3516.460 2229.530 3516.740 2229.810 ;
        RECT 3517.170 2229.530 3517.450 2229.810 ;
        RECT 3517.880 2229.530 3518.160 2229.810 ;
        RECT 3518.590 2229.530 3518.870 2229.810 ;
        RECT 3519.300 2229.530 3519.580 2229.810 ;
        RECT 3520.010 2229.530 3520.290 2229.810 ;
        RECT 3520.720 2229.530 3521.000 2229.810 ;
        RECT 3521.430 2229.530 3521.710 2229.810 ;
        RECT 3512.255 2225.615 3512.535 2225.895 ;
        RECT 3512.965 2225.615 3513.245 2225.895 ;
        RECT 3513.675 2225.615 3513.955 2225.895 ;
        RECT 3514.385 2225.615 3514.665 2225.895 ;
        RECT 3515.095 2225.615 3515.375 2225.895 ;
        RECT 3515.805 2225.615 3516.085 2225.895 ;
        RECT 3516.515 2225.615 3516.795 2225.895 ;
        RECT 3517.225 2225.615 3517.505 2225.895 ;
        RECT 3517.935 2225.615 3518.215 2225.895 ;
        RECT 3518.645 2225.615 3518.925 2225.895 ;
        RECT 3519.355 2225.615 3519.635 2225.895 ;
        RECT 3520.065 2225.615 3520.345 2225.895 ;
        RECT 3520.775 2225.615 3521.055 2225.895 ;
        RECT 3521.485 2225.615 3521.765 2225.895 ;
        RECT 3512.255 2224.905 3512.535 2225.185 ;
        RECT 3512.965 2224.905 3513.245 2225.185 ;
        RECT 3513.675 2224.905 3513.955 2225.185 ;
        RECT 3514.385 2224.905 3514.665 2225.185 ;
        RECT 3515.095 2224.905 3515.375 2225.185 ;
        RECT 3515.805 2224.905 3516.085 2225.185 ;
        RECT 3516.515 2224.905 3516.795 2225.185 ;
        RECT 3517.225 2224.905 3517.505 2225.185 ;
        RECT 3517.935 2224.905 3518.215 2225.185 ;
        RECT 3518.645 2224.905 3518.925 2225.185 ;
        RECT 3519.355 2224.905 3519.635 2225.185 ;
        RECT 3520.065 2224.905 3520.345 2225.185 ;
        RECT 3520.775 2224.905 3521.055 2225.185 ;
        RECT 3521.485 2224.905 3521.765 2225.185 ;
        RECT 3512.255 2224.195 3512.535 2224.475 ;
        RECT 3512.965 2224.195 3513.245 2224.475 ;
        RECT 3513.675 2224.195 3513.955 2224.475 ;
        RECT 3514.385 2224.195 3514.665 2224.475 ;
        RECT 3515.095 2224.195 3515.375 2224.475 ;
        RECT 3515.805 2224.195 3516.085 2224.475 ;
        RECT 3516.515 2224.195 3516.795 2224.475 ;
        RECT 3517.225 2224.195 3517.505 2224.475 ;
        RECT 3517.935 2224.195 3518.215 2224.475 ;
        RECT 3518.645 2224.195 3518.925 2224.475 ;
        RECT 3519.355 2224.195 3519.635 2224.475 ;
        RECT 3520.065 2224.195 3520.345 2224.475 ;
        RECT 3520.775 2224.195 3521.055 2224.475 ;
        RECT 3521.485 2224.195 3521.765 2224.475 ;
        RECT 3512.255 2223.485 3512.535 2223.765 ;
        RECT 3512.965 2223.485 3513.245 2223.765 ;
        RECT 3513.675 2223.485 3513.955 2223.765 ;
        RECT 3514.385 2223.485 3514.665 2223.765 ;
        RECT 3515.095 2223.485 3515.375 2223.765 ;
        RECT 3515.805 2223.485 3516.085 2223.765 ;
        RECT 3516.515 2223.485 3516.795 2223.765 ;
        RECT 3517.225 2223.485 3517.505 2223.765 ;
        RECT 3517.935 2223.485 3518.215 2223.765 ;
        RECT 3518.645 2223.485 3518.925 2223.765 ;
        RECT 3519.355 2223.485 3519.635 2223.765 ;
        RECT 3520.065 2223.485 3520.345 2223.765 ;
        RECT 3520.775 2223.485 3521.055 2223.765 ;
        RECT 3521.485 2223.485 3521.765 2223.765 ;
        RECT 3512.255 2222.775 3512.535 2223.055 ;
        RECT 3512.965 2222.775 3513.245 2223.055 ;
        RECT 3513.675 2222.775 3513.955 2223.055 ;
        RECT 3514.385 2222.775 3514.665 2223.055 ;
        RECT 3515.095 2222.775 3515.375 2223.055 ;
        RECT 3515.805 2222.775 3516.085 2223.055 ;
        RECT 3516.515 2222.775 3516.795 2223.055 ;
        RECT 3517.225 2222.775 3517.505 2223.055 ;
        RECT 3517.935 2222.775 3518.215 2223.055 ;
        RECT 3518.645 2222.775 3518.925 2223.055 ;
        RECT 3519.355 2222.775 3519.635 2223.055 ;
        RECT 3520.065 2222.775 3520.345 2223.055 ;
        RECT 3520.775 2222.775 3521.055 2223.055 ;
        RECT 3521.485 2222.775 3521.765 2223.055 ;
        RECT 3512.255 2222.065 3512.535 2222.345 ;
        RECT 3512.965 2222.065 3513.245 2222.345 ;
        RECT 3513.675 2222.065 3513.955 2222.345 ;
        RECT 3514.385 2222.065 3514.665 2222.345 ;
        RECT 3515.095 2222.065 3515.375 2222.345 ;
        RECT 3515.805 2222.065 3516.085 2222.345 ;
        RECT 3516.515 2222.065 3516.795 2222.345 ;
        RECT 3517.225 2222.065 3517.505 2222.345 ;
        RECT 3517.935 2222.065 3518.215 2222.345 ;
        RECT 3518.645 2222.065 3518.925 2222.345 ;
        RECT 3519.355 2222.065 3519.635 2222.345 ;
        RECT 3520.065 2222.065 3520.345 2222.345 ;
        RECT 3520.775 2222.065 3521.055 2222.345 ;
        RECT 3521.485 2222.065 3521.765 2222.345 ;
        RECT 3512.255 2221.355 3512.535 2221.635 ;
        RECT 3512.965 2221.355 3513.245 2221.635 ;
        RECT 3513.675 2221.355 3513.955 2221.635 ;
        RECT 3514.385 2221.355 3514.665 2221.635 ;
        RECT 3515.095 2221.355 3515.375 2221.635 ;
        RECT 3515.805 2221.355 3516.085 2221.635 ;
        RECT 3516.515 2221.355 3516.795 2221.635 ;
        RECT 3517.225 2221.355 3517.505 2221.635 ;
        RECT 3517.935 2221.355 3518.215 2221.635 ;
        RECT 3518.645 2221.355 3518.925 2221.635 ;
        RECT 3519.355 2221.355 3519.635 2221.635 ;
        RECT 3520.065 2221.355 3520.345 2221.635 ;
        RECT 3520.775 2221.355 3521.055 2221.635 ;
        RECT 3521.485 2221.355 3521.765 2221.635 ;
        RECT 3512.255 2220.645 3512.535 2220.925 ;
        RECT 3512.965 2220.645 3513.245 2220.925 ;
        RECT 3513.675 2220.645 3513.955 2220.925 ;
        RECT 3514.385 2220.645 3514.665 2220.925 ;
        RECT 3515.095 2220.645 3515.375 2220.925 ;
        RECT 3515.805 2220.645 3516.085 2220.925 ;
        RECT 3516.515 2220.645 3516.795 2220.925 ;
        RECT 3517.225 2220.645 3517.505 2220.925 ;
        RECT 3517.935 2220.645 3518.215 2220.925 ;
        RECT 3518.645 2220.645 3518.925 2220.925 ;
        RECT 3519.355 2220.645 3519.635 2220.925 ;
        RECT 3520.065 2220.645 3520.345 2220.925 ;
        RECT 3520.775 2220.645 3521.055 2220.925 ;
        RECT 3521.485 2220.645 3521.765 2220.925 ;
        RECT 3512.255 2219.935 3512.535 2220.215 ;
        RECT 3512.965 2219.935 3513.245 2220.215 ;
        RECT 3513.675 2219.935 3513.955 2220.215 ;
        RECT 3514.385 2219.935 3514.665 2220.215 ;
        RECT 3515.095 2219.935 3515.375 2220.215 ;
        RECT 3515.805 2219.935 3516.085 2220.215 ;
        RECT 3516.515 2219.935 3516.795 2220.215 ;
        RECT 3517.225 2219.935 3517.505 2220.215 ;
        RECT 3517.935 2219.935 3518.215 2220.215 ;
        RECT 3518.645 2219.935 3518.925 2220.215 ;
        RECT 3519.355 2219.935 3519.635 2220.215 ;
        RECT 3520.065 2219.935 3520.345 2220.215 ;
        RECT 3520.775 2219.935 3521.055 2220.215 ;
        RECT 3521.485 2219.935 3521.765 2220.215 ;
        RECT 3512.255 2219.225 3512.535 2219.505 ;
        RECT 3512.965 2219.225 3513.245 2219.505 ;
        RECT 3513.675 2219.225 3513.955 2219.505 ;
        RECT 3514.385 2219.225 3514.665 2219.505 ;
        RECT 3515.095 2219.225 3515.375 2219.505 ;
        RECT 3515.805 2219.225 3516.085 2219.505 ;
        RECT 3516.515 2219.225 3516.795 2219.505 ;
        RECT 3517.225 2219.225 3517.505 2219.505 ;
        RECT 3517.935 2219.225 3518.215 2219.505 ;
        RECT 3518.645 2219.225 3518.925 2219.505 ;
        RECT 3519.355 2219.225 3519.635 2219.505 ;
        RECT 3520.065 2219.225 3520.345 2219.505 ;
        RECT 3520.775 2219.225 3521.055 2219.505 ;
        RECT 3521.485 2219.225 3521.765 2219.505 ;
        RECT 3512.255 2218.515 3512.535 2218.795 ;
        RECT 3512.965 2218.515 3513.245 2218.795 ;
        RECT 3513.675 2218.515 3513.955 2218.795 ;
        RECT 3514.385 2218.515 3514.665 2218.795 ;
        RECT 3515.095 2218.515 3515.375 2218.795 ;
        RECT 3515.805 2218.515 3516.085 2218.795 ;
        RECT 3516.515 2218.515 3516.795 2218.795 ;
        RECT 3517.225 2218.515 3517.505 2218.795 ;
        RECT 3517.935 2218.515 3518.215 2218.795 ;
        RECT 3518.645 2218.515 3518.925 2218.795 ;
        RECT 3519.355 2218.515 3519.635 2218.795 ;
        RECT 3520.065 2218.515 3520.345 2218.795 ;
        RECT 3520.775 2218.515 3521.055 2218.795 ;
        RECT 3521.485 2218.515 3521.765 2218.795 ;
        RECT 3512.255 2217.805 3512.535 2218.085 ;
        RECT 3512.965 2217.805 3513.245 2218.085 ;
        RECT 3513.675 2217.805 3513.955 2218.085 ;
        RECT 3514.385 2217.805 3514.665 2218.085 ;
        RECT 3515.095 2217.805 3515.375 2218.085 ;
        RECT 3515.805 2217.805 3516.085 2218.085 ;
        RECT 3516.515 2217.805 3516.795 2218.085 ;
        RECT 3517.225 2217.805 3517.505 2218.085 ;
        RECT 3517.935 2217.805 3518.215 2218.085 ;
        RECT 3518.645 2217.805 3518.925 2218.085 ;
        RECT 3519.355 2217.805 3519.635 2218.085 ;
        RECT 3520.065 2217.805 3520.345 2218.085 ;
        RECT 3520.775 2217.805 3521.055 2218.085 ;
        RECT 3521.485 2217.805 3521.765 2218.085 ;
        RECT 3512.255 2217.095 3512.535 2217.375 ;
        RECT 3512.965 2217.095 3513.245 2217.375 ;
        RECT 3513.675 2217.095 3513.955 2217.375 ;
        RECT 3514.385 2217.095 3514.665 2217.375 ;
        RECT 3515.095 2217.095 3515.375 2217.375 ;
        RECT 3515.805 2217.095 3516.085 2217.375 ;
        RECT 3516.515 2217.095 3516.795 2217.375 ;
        RECT 3517.225 2217.095 3517.505 2217.375 ;
        RECT 3517.935 2217.095 3518.215 2217.375 ;
        RECT 3518.645 2217.095 3518.925 2217.375 ;
        RECT 3519.355 2217.095 3519.635 2217.375 ;
        RECT 3520.065 2217.095 3520.345 2217.375 ;
        RECT 3520.775 2217.095 3521.055 2217.375 ;
        RECT 3521.485 2217.095 3521.765 2217.375 ;
        RECT 3512.255 2216.385 3512.535 2216.665 ;
        RECT 3512.965 2216.385 3513.245 2216.665 ;
        RECT 3513.675 2216.385 3513.955 2216.665 ;
        RECT 3514.385 2216.385 3514.665 2216.665 ;
        RECT 3515.095 2216.385 3515.375 2216.665 ;
        RECT 3515.805 2216.385 3516.085 2216.665 ;
        RECT 3516.515 2216.385 3516.795 2216.665 ;
        RECT 3517.225 2216.385 3517.505 2216.665 ;
        RECT 3517.935 2216.385 3518.215 2216.665 ;
        RECT 3518.645 2216.385 3518.925 2216.665 ;
        RECT 3519.355 2216.385 3519.635 2216.665 ;
        RECT 3520.065 2216.385 3520.345 2216.665 ;
        RECT 3520.775 2216.385 3521.055 2216.665 ;
        RECT 3521.485 2216.385 3521.765 2216.665 ;
        RECT 3512.255 2213.765 3512.535 2214.045 ;
        RECT 3512.965 2213.765 3513.245 2214.045 ;
        RECT 3513.675 2213.765 3513.955 2214.045 ;
        RECT 3514.385 2213.765 3514.665 2214.045 ;
        RECT 3515.095 2213.765 3515.375 2214.045 ;
        RECT 3515.805 2213.765 3516.085 2214.045 ;
        RECT 3516.515 2213.765 3516.795 2214.045 ;
        RECT 3517.225 2213.765 3517.505 2214.045 ;
        RECT 3517.935 2213.765 3518.215 2214.045 ;
        RECT 3518.645 2213.765 3518.925 2214.045 ;
        RECT 3519.355 2213.765 3519.635 2214.045 ;
        RECT 3520.065 2213.765 3520.345 2214.045 ;
        RECT 3520.775 2213.765 3521.055 2214.045 ;
        RECT 3521.485 2213.765 3521.765 2214.045 ;
        RECT 3512.255 2213.055 3512.535 2213.335 ;
        RECT 3512.965 2213.055 3513.245 2213.335 ;
        RECT 3513.675 2213.055 3513.955 2213.335 ;
        RECT 3514.385 2213.055 3514.665 2213.335 ;
        RECT 3515.095 2213.055 3515.375 2213.335 ;
        RECT 3515.805 2213.055 3516.085 2213.335 ;
        RECT 3516.515 2213.055 3516.795 2213.335 ;
        RECT 3517.225 2213.055 3517.505 2213.335 ;
        RECT 3517.935 2213.055 3518.215 2213.335 ;
        RECT 3518.645 2213.055 3518.925 2213.335 ;
        RECT 3519.355 2213.055 3519.635 2213.335 ;
        RECT 3520.065 2213.055 3520.345 2213.335 ;
        RECT 3520.775 2213.055 3521.055 2213.335 ;
        RECT 3521.485 2213.055 3521.765 2213.335 ;
        RECT 3512.255 2212.345 3512.535 2212.625 ;
        RECT 3512.965 2212.345 3513.245 2212.625 ;
        RECT 3513.675 2212.345 3513.955 2212.625 ;
        RECT 3514.385 2212.345 3514.665 2212.625 ;
        RECT 3515.095 2212.345 3515.375 2212.625 ;
        RECT 3515.805 2212.345 3516.085 2212.625 ;
        RECT 3516.515 2212.345 3516.795 2212.625 ;
        RECT 3517.225 2212.345 3517.505 2212.625 ;
        RECT 3517.935 2212.345 3518.215 2212.625 ;
        RECT 3518.645 2212.345 3518.925 2212.625 ;
        RECT 3519.355 2212.345 3519.635 2212.625 ;
        RECT 3520.065 2212.345 3520.345 2212.625 ;
        RECT 3520.775 2212.345 3521.055 2212.625 ;
        RECT 3521.485 2212.345 3521.765 2212.625 ;
        RECT 3512.255 2211.635 3512.535 2211.915 ;
        RECT 3512.965 2211.635 3513.245 2211.915 ;
        RECT 3513.675 2211.635 3513.955 2211.915 ;
        RECT 3514.385 2211.635 3514.665 2211.915 ;
        RECT 3515.095 2211.635 3515.375 2211.915 ;
        RECT 3515.805 2211.635 3516.085 2211.915 ;
        RECT 3516.515 2211.635 3516.795 2211.915 ;
        RECT 3517.225 2211.635 3517.505 2211.915 ;
        RECT 3517.935 2211.635 3518.215 2211.915 ;
        RECT 3518.645 2211.635 3518.925 2211.915 ;
        RECT 3519.355 2211.635 3519.635 2211.915 ;
        RECT 3520.065 2211.635 3520.345 2211.915 ;
        RECT 3520.775 2211.635 3521.055 2211.915 ;
        RECT 3521.485 2211.635 3521.765 2211.915 ;
        RECT 3512.255 2210.925 3512.535 2211.205 ;
        RECT 3512.965 2210.925 3513.245 2211.205 ;
        RECT 3513.675 2210.925 3513.955 2211.205 ;
        RECT 3514.385 2210.925 3514.665 2211.205 ;
        RECT 3515.095 2210.925 3515.375 2211.205 ;
        RECT 3515.805 2210.925 3516.085 2211.205 ;
        RECT 3516.515 2210.925 3516.795 2211.205 ;
        RECT 3517.225 2210.925 3517.505 2211.205 ;
        RECT 3517.935 2210.925 3518.215 2211.205 ;
        RECT 3518.645 2210.925 3518.925 2211.205 ;
        RECT 3519.355 2210.925 3519.635 2211.205 ;
        RECT 3520.065 2210.925 3520.345 2211.205 ;
        RECT 3520.775 2210.925 3521.055 2211.205 ;
        RECT 3521.485 2210.925 3521.765 2211.205 ;
        RECT 3512.255 2210.215 3512.535 2210.495 ;
        RECT 3512.965 2210.215 3513.245 2210.495 ;
        RECT 3513.675 2210.215 3513.955 2210.495 ;
        RECT 3514.385 2210.215 3514.665 2210.495 ;
        RECT 3515.095 2210.215 3515.375 2210.495 ;
        RECT 3515.805 2210.215 3516.085 2210.495 ;
        RECT 3516.515 2210.215 3516.795 2210.495 ;
        RECT 3517.225 2210.215 3517.505 2210.495 ;
        RECT 3517.935 2210.215 3518.215 2210.495 ;
        RECT 3518.645 2210.215 3518.925 2210.495 ;
        RECT 3519.355 2210.215 3519.635 2210.495 ;
        RECT 3520.065 2210.215 3520.345 2210.495 ;
        RECT 3520.775 2210.215 3521.055 2210.495 ;
        RECT 3521.485 2210.215 3521.765 2210.495 ;
        RECT 3512.255 2209.505 3512.535 2209.785 ;
        RECT 3512.965 2209.505 3513.245 2209.785 ;
        RECT 3513.675 2209.505 3513.955 2209.785 ;
        RECT 3514.385 2209.505 3514.665 2209.785 ;
        RECT 3515.095 2209.505 3515.375 2209.785 ;
        RECT 3515.805 2209.505 3516.085 2209.785 ;
        RECT 3516.515 2209.505 3516.795 2209.785 ;
        RECT 3517.225 2209.505 3517.505 2209.785 ;
        RECT 3517.935 2209.505 3518.215 2209.785 ;
        RECT 3518.645 2209.505 3518.925 2209.785 ;
        RECT 3519.355 2209.505 3519.635 2209.785 ;
        RECT 3520.065 2209.505 3520.345 2209.785 ;
        RECT 3520.775 2209.505 3521.055 2209.785 ;
        RECT 3521.485 2209.505 3521.765 2209.785 ;
        RECT 3512.255 2208.795 3512.535 2209.075 ;
        RECT 3512.965 2208.795 3513.245 2209.075 ;
        RECT 3513.675 2208.795 3513.955 2209.075 ;
        RECT 3514.385 2208.795 3514.665 2209.075 ;
        RECT 3515.095 2208.795 3515.375 2209.075 ;
        RECT 3515.805 2208.795 3516.085 2209.075 ;
        RECT 3516.515 2208.795 3516.795 2209.075 ;
        RECT 3517.225 2208.795 3517.505 2209.075 ;
        RECT 3517.935 2208.795 3518.215 2209.075 ;
        RECT 3518.645 2208.795 3518.925 2209.075 ;
        RECT 3519.355 2208.795 3519.635 2209.075 ;
        RECT 3520.065 2208.795 3520.345 2209.075 ;
        RECT 3520.775 2208.795 3521.055 2209.075 ;
        RECT 3521.485 2208.795 3521.765 2209.075 ;
        RECT 3512.255 2208.085 3512.535 2208.365 ;
        RECT 3512.965 2208.085 3513.245 2208.365 ;
        RECT 3513.675 2208.085 3513.955 2208.365 ;
        RECT 3514.385 2208.085 3514.665 2208.365 ;
        RECT 3515.095 2208.085 3515.375 2208.365 ;
        RECT 3515.805 2208.085 3516.085 2208.365 ;
        RECT 3516.515 2208.085 3516.795 2208.365 ;
        RECT 3517.225 2208.085 3517.505 2208.365 ;
        RECT 3517.935 2208.085 3518.215 2208.365 ;
        RECT 3518.645 2208.085 3518.925 2208.365 ;
        RECT 3519.355 2208.085 3519.635 2208.365 ;
        RECT 3520.065 2208.085 3520.345 2208.365 ;
        RECT 3520.775 2208.085 3521.055 2208.365 ;
        RECT 3521.485 2208.085 3521.765 2208.365 ;
        RECT 3512.255 2207.375 3512.535 2207.655 ;
        RECT 3512.965 2207.375 3513.245 2207.655 ;
        RECT 3513.675 2207.375 3513.955 2207.655 ;
        RECT 3514.385 2207.375 3514.665 2207.655 ;
        RECT 3515.095 2207.375 3515.375 2207.655 ;
        RECT 3515.805 2207.375 3516.085 2207.655 ;
        RECT 3516.515 2207.375 3516.795 2207.655 ;
        RECT 3517.225 2207.375 3517.505 2207.655 ;
        RECT 3517.935 2207.375 3518.215 2207.655 ;
        RECT 3518.645 2207.375 3518.925 2207.655 ;
        RECT 3519.355 2207.375 3519.635 2207.655 ;
        RECT 3520.065 2207.375 3520.345 2207.655 ;
        RECT 3520.775 2207.375 3521.055 2207.655 ;
        RECT 3521.485 2207.375 3521.765 2207.655 ;
        RECT 3512.255 2206.665 3512.535 2206.945 ;
        RECT 3512.965 2206.665 3513.245 2206.945 ;
        RECT 3513.675 2206.665 3513.955 2206.945 ;
        RECT 3514.385 2206.665 3514.665 2206.945 ;
        RECT 3515.095 2206.665 3515.375 2206.945 ;
        RECT 3515.805 2206.665 3516.085 2206.945 ;
        RECT 3516.515 2206.665 3516.795 2206.945 ;
        RECT 3517.225 2206.665 3517.505 2206.945 ;
        RECT 3517.935 2206.665 3518.215 2206.945 ;
        RECT 3518.645 2206.665 3518.925 2206.945 ;
        RECT 3519.355 2206.665 3519.635 2206.945 ;
        RECT 3520.065 2206.665 3520.345 2206.945 ;
        RECT 3520.775 2206.665 3521.055 2206.945 ;
        RECT 3521.485 2206.665 3521.765 2206.945 ;
        RECT 3512.255 2205.955 3512.535 2206.235 ;
        RECT 3512.965 2205.955 3513.245 2206.235 ;
        RECT 3513.675 2205.955 3513.955 2206.235 ;
        RECT 3514.385 2205.955 3514.665 2206.235 ;
        RECT 3515.095 2205.955 3515.375 2206.235 ;
        RECT 3515.805 2205.955 3516.085 2206.235 ;
        RECT 3516.515 2205.955 3516.795 2206.235 ;
        RECT 3517.225 2205.955 3517.505 2206.235 ;
        RECT 3517.935 2205.955 3518.215 2206.235 ;
        RECT 3518.645 2205.955 3518.925 2206.235 ;
        RECT 3519.355 2205.955 3519.635 2206.235 ;
        RECT 3520.065 2205.955 3520.345 2206.235 ;
        RECT 3520.775 2205.955 3521.055 2206.235 ;
        RECT 3521.485 2205.955 3521.765 2206.235 ;
        RECT 3512.255 2205.245 3512.535 2205.525 ;
        RECT 3512.965 2205.245 3513.245 2205.525 ;
        RECT 3513.675 2205.245 3513.955 2205.525 ;
        RECT 3514.385 2205.245 3514.665 2205.525 ;
        RECT 3515.095 2205.245 3515.375 2205.525 ;
        RECT 3515.805 2205.245 3516.085 2205.525 ;
        RECT 3516.515 2205.245 3516.795 2205.525 ;
        RECT 3517.225 2205.245 3517.505 2205.525 ;
        RECT 3517.935 2205.245 3518.215 2205.525 ;
        RECT 3518.645 2205.245 3518.925 2205.525 ;
        RECT 3519.355 2205.245 3519.635 2205.525 ;
        RECT 3520.065 2205.245 3520.345 2205.525 ;
        RECT 3520.775 2205.245 3521.055 2205.525 ;
        RECT 3521.485 2205.245 3521.765 2205.525 ;
        RECT 3512.255 2204.535 3512.535 2204.815 ;
        RECT 3512.965 2204.535 3513.245 2204.815 ;
        RECT 3513.675 2204.535 3513.955 2204.815 ;
        RECT 3514.385 2204.535 3514.665 2204.815 ;
        RECT 3515.095 2204.535 3515.375 2204.815 ;
        RECT 3515.805 2204.535 3516.085 2204.815 ;
        RECT 3516.515 2204.535 3516.795 2204.815 ;
        RECT 3517.225 2204.535 3517.505 2204.815 ;
        RECT 3517.935 2204.535 3518.215 2204.815 ;
        RECT 3518.645 2204.535 3518.925 2204.815 ;
        RECT 3519.355 2204.535 3519.635 2204.815 ;
        RECT 3520.065 2204.535 3520.345 2204.815 ;
        RECT 3520.775 2204.535 3521.055 2204.815 ;
        RECT 3521.485 2204.535 3521.765 2204.815 ;
        RECT 3512.255 2200.235 3512.535 2200.515 ;
        RECT 3512.965 2200.235 3513.245 2200.515 ;
        RECT 3513.675 2200.235 3513.955 2200.515 ;
        RECT 3514.385 2200.235 3514.665 2200.515 ;
        RECT 3515.095 2200.235 3515.375 2200.515 ;
        RECT 3515.805 2200.235 3516.085 2200.515 ;
        RECT 3516.515 2200.235 3516.795 2200.515 ;
        RECT 3517.225 2200.235 3517.505 2200.515 ;
        RECT 3517.935 2200.235 3518.215 2200.515 ;
        RECT 3518.645 2200.235 3518.925 2200.515 ;
        RECT 3519.355 2200.235 3519.635 2200.515 ;
        RECT 3520.065 2200.235 3520.345 2200.515 ;
        RECT 3520.775 2200.235 3521.055 2200.515 ;
        RECT 3521.485 2200.235 3521.765 2200.515 ;
        RECT 3512.255 2199.525 3512.535 2199.805 ;
        RECT 3512.965 2199.525 3513.245 2199.805 ;
        RECT 3513.675 2199.525 3513.955 2199.805 ;
        RECT 3514.385 2199.525 3514.665 2199.805 ;
        RECT 3515.095 2199.525 3515.375 2199.805 ;
        RECT 3515.805 2199.525 3516.085 2199.805 ;
        RECT 3516.515 2199.525 3516.795 2199.805 ;
        RECT 3517.225 2199.525 3517.505 2199.805 ;
        RECT 3517.935 2199.525 3518.215 2199.805 ;
        RECT 3518.645 2199.525 3518.925 2199.805 ;
        RECT 3519.355 2199.525 3519.635 2199.805 ;
        RECT 3520.065 2199.525 3520.345 2199.805 ;
        RECT 3520.775 2199.525 3521.055 2199.805 ;
        RECT 3521.485 2199.525 3521.765 2199.805 ;
        RECT 3512.255 2198.815 3512.535 2199.095 ;
        RECT 3512.965 2198.815 3513.245 2199.095 ;
        RECT 3513.675 2198.815 3513.955 2199.095 ;
        RECT 3514.385 2198.815 3514.665 2199.095 ;
        RECT 3515.095 2198.815 3515.375 2199.095 ;
        RECT 3515.805 2198.815 3516.085 2199.095 ;
        RECT 3516.515 2198.815 3516.795 2199.095 ;
        RECT 3517.225 2198.815 3517.505 2199.095 ;
        RECT 3517.935 2198.815 3518.215 2199.095 ;
        RECT 3518.645 2198.815 3518.925 2199.095 ;
        RECT 3519.355 2198.815 3519.635 2199.095 ;
        RECT 3520.065 2198.815 3520.345 2199.095 ;
        RECT 3520.775 2198.815 3521.055 2199.095 ;
        RECT 3521.485 2198.815 3521.765 2199.095 ;
        RECT 3512.255 2198.105 3512.535 2198.385 ;
        RECT 3512.965 2198.105 3513.245 2198.385 ;
        RECT 3513.675 2198.105 3513.955 2198.385 ;
        RECT 3514.385 2198.105 3514.665 2198.385 ;
        RECT 3515.095 2198.105 3515.375 2198.385 ;
        RECT 3515.805 2198.105 3516.085 2198.385 ;
        RECT 3516.515 2198.105 3516.795 2198.385 ;
        RECT 3517.225 2198.105 3517.505 2198.385 ;
        RECT 3517.935 2198.105 3518.215 2198.385 ;
        RECT 3518.645 2198.105 3518.925 2198.385 ;
        RECT 3519.355 2198.105 3519.635 2198.385 ;
        RECT 3520.065 2198.105 3520.345 2198.385 ;
        RECT 3520.775 2198.105 3521.055 2198.385 ;
        RECT 3521.485 2198.105 3521.765 2198.385 ;
        RECT 3512.255 2197.395 3512.535 2197.675 ;
        RECT 3512.965 2197.395 3513.245 2197.675 ;
        RECT 3513.675 2197.395 3513.955 2197.675 ;
        RECT 3514.385 2197.395 3514.665 2197.675 ;
        RECT 3515.095 2197.395 3515.375 2197.675 ;
        RECT 3515.805 2197.395 3516.085 2197.675 ;
        RECT 3516.515 2197.395 3516.795 2197.675 ;
        RECT 3517.225 2197.395 3517.505 2197.675 ;
        RECT 3517.935 2197.395 3518.215 2197.675 ;
        RECT 3518.645 2197.395 3518.925 2197.675 ;
        RECT 3519.355 2197.395 3519.635 2197.675 ;
        RECT 3520.065 2197.395 3520.345 2197.675 ;
        RECT 3520.775 2197.395 3521.055 2197.675 ;
        RECT 3521.485 2197.395 3521.765 2197.675 ;
        RECT 3512.255 2196.685 3512.535 2196.965 ;
        RECT 3512.965 2196.685 3513.245 2196.965 ;
        RECT 3513.675 2196.685 3513.955 2196.965 ;
        RECT 3514.385 2196.685 3514.665 2196.965 ;
        RECT 3515.095 2196.685 3515.375 2196.965 ;
        RECT 3515.805 2196.685 3516.085 2196.965 ;
        RECT 3516.515 2196.685 3516.795 2196.965 ;
        RECT 3517.225 2196.685 3517.505 2196.965 ;
        RECT 3517.935 2196.685 3518.215 2196.965 ;
        RECT 3518.645 2196.685 3518.925 2196.965 ;
        RECT 3519.355 2196.685 3519.635 2196.965 ;
        RECT 3520.065 2196.685 3520.345 2196.965 ;
        RECT 3520.775 2196.685 3521.055 2196.965 ;
        RECT 3521.485 2196.685 3521.765 2196.965 ;
        RECT 3512.255 2195.975 3512.535 2196.255 ;
        RECT 3512.965 2195.975 3513.245 2196.255 ;
        RECT 3513.675 2195.975 3513.955 2196.255 ;
        RECT 3514.385 2195.975 3514.665 2196.255 ;
        RECT 3515.095 2195.975 3515.375 2196.255 ;
        RECT 3515.805 2195.975 3516.085 2196.255 ;
        RECT 3516.515 2195.975 3516.795 2196.255 ;
        RECT 3517.225 2195.975 3517.505 2196.255 ;
        RECT 3517.935 2195.975 3518.215 2196.255 ;
        RECT 3518.645 2195.975 3518.925 2196.255 ;
        RECT 3519.355 2195.975 3519.635 2196.255 ;
        RECT 3520.065 2195.975 3520.345 2196.255 ;
        RECT 3520.775 2195.975 3521.055 2196.255 ;
        RECT 3521.485 2195.975 3521.765 2196.255 ;
        RECT 3512.255 2195.265 3512.535 2195.545 ;
        RECT 3512.965 2195.265 3513.245 2195.545 ;
        RECT 3513.675 2195.265 3513.955 2195.545 ;
        RECT 3514.385 2195.265 3514.665 2195.545 ;
        RECT 3515.095 2195.265 3515.375 2195.545 ;
        RECT 3515.805 2195.265 3516.085 2195.545 ;
        RECT 3516.515 2195.265 3516.795 2195.545 ;
        RECT 3517.225 2195.265 3517.505 2195.545 ;
        RECT 3517.935 2195.265 3518.215 2195.545 ;
        RECT 3518.645 2195.265 3518.925 2195.545 ;
        RECT 3519.355 2195.265 3519.635 2195.545 ;
        RECT 3520.065 2195.265 3520.345 2195.545 ;
        RECT 3520.775 2195.265 3521.055 2195.545 ;
        RECT 3521.485 2195.265 3521.765 2195.545 ;
        RECT 3512.255 2194.555 3512.535 2194.835 ;
        RECT 3512.965 2194.555 3513.245 2194.835 ;
        RECT 3513.675 2194.555 3513.955 2194.835 ;
        RECT 3514.385 2194.555 3514.665 2194.835 ;
        RECT 3515.095 2194.555 3515.375 2194.835 ;
        RECT 3515.805 2194.555 3516.085 2194.835 ;
        RECT 3516.515 2194.555 3516.795 2194.835 ;
        RECT 3517.225 2194.555 3517.505 2194.835 ;
        RECT 3517.935 2194.555 3518.215 2194.835 ;
        RECT 3518.645 2194.555 3518.925 2194.835 ;
        RECT 3519.355 2194.555 3519.635 2194.835 ;
        RECT 3520.065 2194.555 3520.345 2194.835 ;
        RECT 3520.775 2194.555 3521.055 2194.835 ;
        RECT 3521.485 2194.555 3521.765 2194.835 ;
        RECT 3512.255 2193.845 3512.535 2194.125 ;
        RECT 3512.965 2193.845 3513.245 2194.125 ;
        RECT 3513.675 2193.845 3513.955 2194.125 ;
        RECT 3514.385 2193.845 3514.665 2194.125 ;
        RECT 3515.095 2193.845 3515.375 2194.125 ;
        RECT 3515.805 2193.845 3516.085 2194.125 ;
        RECT 3516.515 2193.845 3516.795 2194.125 ;
        RECT 3517.225 2193.845 3517.505 2194.125 ;
        RECT 3517.935 2193.845 3518.215 2194.125 ;
        RECT 3518.645 2193.845 3518.925 2194.125 ;
        RECT 3519.355 2193.845 3519.635 2194.125 ;
        RECT 3520.065 2193.845 3520.345 2194.125 ;
        RECT 3520.775 2193.845 3521.055 2194.125 ;
        RECT 3521.485 2193.845 3521.765 2194.125 ;
        RECT 3512.255 2193.135 3512.535 2193.415 ;
        RECT 3512.965 2193.135 3513.245 2193.415 ;
        RECT 3513.675 2193.135 3513.955 2193.415 ;
        RECT 3514.385 2193.135 3514.665 2193.415 ;
        RECT 3515.095 2193.135 3515.375 2193.415 ;
        RECT 3515.805 2193.135 3516.085 2193.415 ;
        RECT 3516.515 2193.135 3516.795 2193.415 ;
        RECT 3517.225 2193.135 3517.505 2193.415 ;
        RECT 3517.935 2193.135 3518.215 2193.415 ;
        RECT 3518.645 2193.135 3518.925 2193.415 ;
        RECT 3519.355 2193.135 3519.635 2193.415 ;
        RECT 3520.065 2193.135 3520.345 2193.415 ;
        RECT 3520.775 2193.135 3521.055 2193.415 ;
        RECT 3521.485 2193.135 3521.765 2193.415 ;
        RECT 3512.255 2192.425 3512.535 2192.705 ;
        RECT 3512.965 2192.425 3513.245 2192.705 ;
        RECT 3513.675 2192.425 3513.955 2192.705 ;
        RECT 3514.385 2192.425 3514.665 2192.705 ;
        RECT 3515.095 2192.425 3515.375 2192.705 ;
        RECT 3515.805 2192.425 3516.085 2192.705 ;
        RECT 3516.515 2192.425 3516.795 2192.705 ;
        RECT 3517.225 2192.425 3517.505 2192.705 ;
        RECT 3517.935 2192.425 3518.215 2192.705 ;
        RECT 3518.645 2192.425 3518.925 2192.705 ;
        RECT 3519.355 2192.425 3519.635 2192.705 ;
        RECT 3520.065 2192.425 3520.345 2192.705 ;
        RECT 3520.775 2192.425 3521.055 2192.705 ;
        RECT 3521.485 2192.425 3521.765 2192.705 ;
        RECT 3512.255 2191.715 3512.535 2191.995 ;
        RECT 3512.965 2191.715 3513.245 2191.995 ;
        RECT 3513.675 2191.715 3513.955 2191.995 ;
        RECT 3514.385 2191.715 3514.665 2191.995 ;
        RECT 3515.095 2191.715 3515.375 2191.995 ;
        RECT 3515.805 2191.715 3516.085 2191.995 ;
        RECT 3516.515 2191.715 3516.795 2191.995 ;
        RECT 3517.225 2191.715 3517.505 2191.995 ;
        RECT 3517.935 2191.715 3518.215 2191.995 ;
        RECT 3518.645 2191.715 3518.925 2191.995 ;
        RECT 3519.355 2191.715 3519.635 2191.995 ;
        RECT 3520.065 2191.715 3520.345 2191.995 ;
        RECT 3520.775 2191.715 3521.055 2191.995 ;
        RECT 3521.485 2191.715 3521.765 2191.995 ;
        RECT 3512.255 2191.005 3512.535 2191.285 ;
        RECT 3512.965 2191.005 3513.245 2191.285 ;
        RECT 3513.675 2191.005 3513.955 2191.285 ;
        RECT 3514.385 2191.005 3514.665 2191.285 ;
        RECT 3515.095 2191.005 3515.375 2191.285 ;
        RECT 3515.805 2191.005 3516.085 2191.285 ;
        RECT 3516.515 2191.005 3516.795 2191.285 ;
        RECT 3517.225 2191.005 3517.505 2191.285 ;
        RECT 3517.935 2191.005 3518.215 2191.285 ;
        RECT 3518.645 2191.005 3518.925 2191.285 ;
        RECT 3519.355 2191.005 3519.635 2191.285 ;
        RECT 3520.065 2191.005 3520.345 2191.285 ;
        RECT 3520.775 2191.005 3521.055 2191.285 ;
        RECT 3521.485 2191.005 3521.765 2191.285 ;
        RECT 3512.255 2188.385 3512.535 2188.665 ;
        RECT 3512.965 2188.385 3513.245 2188.665 ;
        RECT 3513.675 2188.385 3513.955 2188.665 ;
        RECT 3514.385 2188.385 3514.665 2188.665 ;
        RECT 3515.095 2188.385 3515.375 2188.665 ;
        RECT 3515.805 2188.385 3516.085 2188.665 ;
        RECT 3516.515 2188.385 3516.795 2188.665 ;
        RECT 3517.225 2188.385 3517.505 2188.665 ;
        RECT 3517.935 2188.385 3518.215 2188.665 ;
        RECT 3518.645 2188.385 3518.925 2188.665 ;
        RECT 3519.355 2188.385 3519.635 2188.665 ;
        RECT 3520.065 2188.385 3520.345 2188.665 ;
        RECT 3520.775 2188.385 3521.055 2188.665 ;
        RECT 3521.485 2188.385 3521.765 2188.665 ;
        RECT 3512.255 2187.675 3512.535 2187.955 ;
        RECT 3512.965 2187.675 3513.245 2187.955 ;
        RECT 3513.675 2187.675 3513.955 2187.955 ;
        RECT 3514.385 2187.675 3514.665 2187.955 ;
        RECT 3515.095 2187.675 3515.375 2187.955 ;
        RECT 3515.805 2187.675 3516.085 2187.955 ;
        RECT 3516.515 2187.675 3516.795 2187.955 ;
        RECT 3517.225 2187.675 3517.505 2187.955 ;
        RECT 3517.935 2187.675 3518.215 2187.955 ;
        RECT 3518.645 2187.675 3518.925 2187.955 ;
        RECT 3519.355 2187.675 3519.635 2187.955 ;
        RECT 3520.065 2187.675 3520.345 2187.955 ;
        RECT 3520.775 2187.675 3521.055 2187.955 ;
        RECT 3521.485 2187.675 3521.765 2187.955 ;
        RECT 3512.255 2186.965 3512.535 2187.245 ;
        RECT 3512.965 2186.965 3513.245 2187.245 ;
        RECT 3513.675 2186.965 3513.955 2187.245 ;
        RECT 3514.385 2186.965 3514.665 2187.245 ;
        RECT 3515.095 2186.965 3515.375 2187.245 ;
        RECT 3515.805 2186.965 3516.085 2187.245 ;
        RECT 3516.515 2186.965 3516.795 2187.245 ;
        RECT 3517.225 2186.965 3517.505 2187.245 ;
        RECT 3517.935 2186.965 3518.215 2187.245 ;
        RECT 3518.645 2186.965 3518.925 2187.245 ;
        RECT 3519.355 2186.965 3519.635 2187.245 ;
        RECT 3520.065 2186.965 3520.345 2187.245 ;
        RECT 3520.775 2186.965 3521.055 2187.245 ;
        RECT 3521.485 2186.965 3521.765 2187.245 ;
        RECT 3512.255 2186.255 3512.535 2186.535 ;
        RECT 3512.965 2186.255 3513.245 2186.535 ;
        RECT 3513.675 2186.255 3513.955 2186.535 ;
        RECT 3514.385 2186.255 3514.665 2186.535 ;
        RECT 3515.095 2186.255 3515.375 2186.535 ;
        RECT 3515.805 2186.255 3516.085 2186.535 ;
        RECT 3516.515 2186.255 3516.795 2186.535 ;
        RECT 3517.225 2186.255 3517.505 2186.535 ;
        RECT 3517.935 2186.255 3518.215 2186.535 ;
        RECT 3518.645 2186.255 3518.925 2186.535 ;
        RECT 3519.355 2186.255 3519.635 2186.535 ;
        RECT 3520.065 2186.255 3520.345 2186.535 ;
        RECT 3520.775 2186.255 3521.055 2186.535 ;
        RECT 3521.485 2186.255 3521.765 2186.535 ;
        RECT 3512.255 2185.545 3512.535 2185.825 ;
        RECT 3512.965 2185.545 3513.245 2185.825 ;
        RECT 3513.675 2185.545 3513.955 2185.825 ;
        RECT 3514.385 2185.545 3514.665 2185.825 ;
        RECT 3515.095 2185.545 3515.375 2185.825 ;
        RECT 3515.805 2185.545 3516.085 2185.825 ;
        RECT 3516.515 2185.545 3516.795 2185.825 ;
        RECT 3517.225 2185.545 3517.505 2185.825 ;
        RECT 3517.935 2185.545 3518.215 2185.825 ;
        RECT 3518.645 2185.545 3518.925 2185.825 ;
        RECT 3519.355 2185.545 3519.635 2185.825 ;
        RECT 3520.065 2185.545 3520.345 2185.825 ;
        RECT 3520.775 2185.545 3521.055 2185.825 ;
        RECT 3521.485 2185.545 3521.765 2185.825 ;
        RECT 3512.255 2184.835 3512.535 2185.115 ;
        RECT 3512.965 2184.835 3513.245 2185.115 ;
        RECT 3513.675 2184.835 3513.955 2185.115 ;
        RECT 3514.385 2184.835 3514.665 2185.115 ;
        RECT 3515.095 2184.835 3515.375 2185.115 ;
        RECT 3515.805 2184.835 3516.085 2185.115 ;
        RECT 3516.515 2184.835 3516.795 2185.115 ;
        RECT 3517.225 2184.835 3517.505 2185.115 ;
        RECT 3517.935 2184.835 3518.215 2185.115 ;
        RECT 3518.645 2184.835 3518.925 2185.115 ;
        RECT 3519.355 2184.835 3519.635 2185.115 ;
        RECT 3520.065 2184.835 3520.345 2185.115 ;
        RECT 3520.775 2184.835 3521.055 2185.115 ;
        RECT 3521.485 2184.835 3521.765 2185.115 ;
        RECT 3512.255 2184.125 3512.535 2184.405 ;
        RECT 3512.965 2184.125 3513.245 2184.405 ;
        RECT 3513.675 2184.125 3513.955 2184.405 ;
        RECT 3514.385 2184.125 3514.665 2184.405 ;
        RECT 3515.095 2184.125 3515.375 2184.405 ;
        RECT 3515.805 2184.125 3516.085 2184.405 ;
        RECT 3516.515 2184.125 3516.795 2184.405 ;
        RECT 3517.225 2184.125 3517.505 2184.405 ;
        RECT 3517.935 2184.125 3518.215 2184.405 ;
        RECT 3518.645 2184.125 3518.925 2184.405 ;
        RECT 3519.355 2184.125 3519.635 2184.405 ;
        RECT 3520.065 2184.125 3520.345 2184.405 ;
        RECT 3520.775 2184.125 3521.055 2184.405 ;
        RECT 3521.485 2184.125 3521.765 2184.405 ;
        RECT 3512.255 2183.415 3512.535 2183.695 ;
        RECT 3512.965 2183.415 3513.245 2183.695 ;
        RECT 3513.675 2183.415 3513.955 2183.695 ;
        RECT 3514.385 2183.415 3514.665 2183.695 ;
        RECT 3515.095 2183.415 3515.375 2183.695 ;
        RECT 3515.805 2183.415 3516.085 2183.695 ;
        RECT 3516.515 2183.415 3516.795 2183.695 ;
        RECT 3517.225 2183.415 3517.505 2183.695 ;
        RECT 3517.935 2183.415 3518.215 2183.695 ;
        RECT 3518.645 2183.415 3518.925 2183.695 ;
        RECT 3519.355 2183.415 3519.635 2183.695 ;
        RECT 3520.065 2183.415 3520.345 2183.695 ;
        RECT 3520.775 2183.415 3521.055 2183.695 ;
        RECT 3521.485 2183.415 3521.765 2183.695 ;
        RECT 3512.255 2182.705 3512.535 2182.985 ;
        RECT 3512.965 2182.705 3513.245 2182.985 ;
        RECT 3513.675 2182.705 3513.955 2182.985 ;
        RECT 3514.385 2182.705 3514.665 2182.985 ;
        RECT 3515.095 2182.705 3515.375 2182.985 ;
        RECT 3515.805 2182.705 3516.085 2182.985 ;
        RECT 3516.515 2182.705 3516.795 2182.985 ;
        RECT 3517.225 2182.705 3517.505 2182.985 ;
        RECT 3517.935 2182.705 3518.215 2182.985 ;
        RECT 3518.645 2182.705 3518.925 2182.985 ;
        RECT 3519.355 2182.705 3519.635 2182.985 ;
        RECT 3520.065 2182.705 3520.345 2182.985 ;
        RECT 3520.775 2182.705 3521.055 2182.985 ;
        RECT 3521.485 2182.705 3521.765 2182.985 ;
        RECT 3512.255 2181.995 3512.535 2182.275 ;
        RECT 3512.965 2181.995 3513.245 2182.275 ;
        RECT 3513.675 2181.995 3513.955 2182.275 ;
        RECT 3514.385 2181.995 3514.665 2182.275 ;
        RECT 3515.095 2181.995 3515.375 2182.275 ;
        RECT 3515.805 2181.995 3516.085 2182.275 ;
        RECT 3516.515 2181.995 3516.795 2182.275 ;
        RECT 3517.225 2181.995 3517.505 2182.275 ;
        RECT 3517.935 2181.995 3518.215 2182.275 ;
        RECT 3518.645 2181.995 3518.925 2182.275 ;
        RECT 3519.355 2181.995 3519.635 2182.275 ;
        RECT 3520.065 2181.995 3520.345 2182.275 ;
        RECT 3520.775 2181.995 3521.055 2182.275 ;
        RECT 3521.485 2181.995 3521.765 2182.275 ;
        RECT 3512.255 2181.285 3512.535 2181.565 ;
        RECT 3512.965 2181.285 3513.245 2181.565 ;
        RECT 3513.675 2181.285 3513.955 2181.565 ;
        RECT 3514.385 2181.285 3514.665 2181.565 ;
        RECT 3515.095 2181.285 3515.375 2181.565 ;
        RECT 3515.805 2181.285 3516.085 2181.565 ;
        RECT 3516.515 2181.285 3516.795 2181.565 ;
        RECT 3517.225 2181.285 3517.505 2181.565 ;
        RECT 3517.935 2181.285 3518.215 2181.565 ;
        RECT 3518.645 2181.285 3518.925 2181.565 ;
        RECT 3519.355 2181.285 3519.635 2181.565 ;
        RECT 3520.065 2181.285 3520.345 2181.565 ;
        RECT 3520.775 2181.285 3521.055 2181.565 ;
        RECT 3521.485 2181.285 3521.765 2181.565 ;
        RECT 3512.255 2180.575 3512.535 2180.855 ;
        RECT 3512.965 2180.575 3513.245 2180.855 ;
        RECT 3513.675 2180.575 3513.955 2180.855 ;
        RECT 3514.385 2180.575 3514.665 2180.855 ;
        RECT 3515.095 2180.575 3515.375 2180.855 ;
        RECT 3515.805 2180.575 3516.085 2180.855 ;
        RECT 3516.515 2180.575 3516.795 2180.855 ;
        RECT 3517.225 2180.575 3517.505 2180.855 ;
        RECT 3517.935 2180.575 3518.215 2180.855 ;
        RECT 3518.645 2180.575 3518.925 2180.855 ;
        RECT 3519.355 2180.575 3519.635 2180.855 ;
        RECT 3520.065 2180.575 3520.345 2180.855 ;
        RECT 3520.775 2180.575 3521.055 2180.855 ;
        RECT 3521.485 2180.575 3521.765 2180.855 ;
        RECT 3512.200 2175.270 3512.480 2175.550 ;
        RECT 3512.910 2175.270 3513.190 2175.550 ;
        RECT 3513.620 2175.270 3513.900 2175.550 ;
        RECT 3514.330 2175.270 3514.610 2175.550 ;
        RECT 3515.040 2175.270 3515.320 2175.550 ;
        RECT 3515.750 2175.270 3516.030 2175.550 ;
        RECT 3516.460 2175.270 3516.740 2175.550 ;
        RECT 3517.170 2175.270 3517.450 2175.550 ;
        RECT 3517.880 2175.270 3518.160 2175.550 ;
        RECT 3518.590 2175.270 3518.870 2175.550 ;
        RECT 3519.300 2175.270 3519.580 2175.550 ;
        RECT 3520.010 2175.270 3520.290 2175.550 ;
        RECT 3520.720 2175.270 3521.000 2175.550 ;
        RECT 3521.430 2175.270 3521.710 2175.550 ;
        RECT 3512.200 2174.560 3512.480 2174.840 ;
        RECT 3512.910 2174.560 3513.190 2174.840 ;
        RECT 3513.620 2174.560 3513.900 2174.840 ;
        RECT 3514.330 2174.560 3514.610 2174.840 ;
        RECT 3515.040 2174.560 3515.320 2174.840 ;
        RECT 3515.750 2174.560 3516.030 2174.840 ;
        RECT 3516.460 2174.560 3516.740 2174.840 ;
        RECT 3517.170 2174.560 3517.450 2174.840 ;
        RECT 3517.880 2174.560 3518.160 2174.840 ;
        RECT 3518.590 2174.560 3518.870 2174.840 ;
        RECT 3519.300 2174.560 3519.580 2174.840 ;
        RECT 3520.010 2174.560 3520.290 2174.840 ;
        RECT 3520.720 2174.560 3521.000 2174.840 ;
        RECT 3521.430 2174.560 3521.710 2174.840 ;
        RECT 3512.200 2173.850 3512.480 2174.130 ;
        RECT 3512.910 2173.850 3513.190 2174.130 ;
        RECT 3513.620 2173.850 3513.900 2174.130 ;
        RECT 3514.330 2173.850 3514.610 2174.130 ;
        RECT 3515.040 2173.850 3515.320 2174.130 ;
        RECT 3515.750 2173.850 3516.030 2174.130 ;
        RECT 3516.460 2173.850 3516.740 2174.130 ;
        RECT 3517.170 2173.850 3517.450 2174.130 ;
        RECT 3517.880 2173.850 3518.160 2174.130 ;
        RECT 3518.590 2173.850 3518.870 2174.130 ;
        RECT 3519.300 2173.850 3519.580 2174.130 ;
        RECT 3520.010 2173.850 3520.290 2174.130 ;
        RECT 3520.720 2173.850 3521.000 2174.130 ;
        RECT 3521.430 2173.850 3521.710 2174.130 ;
        RECT 3512.200 2173.140 3512.480 2173.420 ;
        RECT 3512.910 2173.140 3513.190 2173.420 ;
        RECT 3513.620 2173.140 3513.900 2173.420 ;
        RECT 3514.330 2173.140 3514.610 2173.420 ;
        RECT 3515.040 2173.140 3515.320 2173.420 ;
        RECT 3515.750 2173.140 3516.030 2173.420 ;
        RECT 3516.460 2173.140 3516.740 2173.420 ;
        RECT 3517.170 2173.140 3517.450 2173.420 ;
        RECT 3517.880 2173.140 3518.160 2173.420 ;
        RECT 3518.590 2173.140 3518.870 2173.420 ;
        RECT 3519.300 2173.140 3519.580 2173.420 ;
        RECT 3520.010 2173.140 3520.290 2173.420 ;
        RECT 3520.720 2173.140 3521.000 2173.420 ;
        RECT 3521.430 2173.140 3521.710 2173.420 ;
        RECT 3512.200 2172.430 3512.480 2172.710 ;
        RECT 3512.910 2172.430 3513.190 2172.710 ;
        RECT 3513.620 2172.430 3513.900 2172.710 ;
        RECT 3514.330 2172.430 3514.610 2172.710 ;
        RECT 3515.040 2172.430 3515.320 2172.710 ;
        RECT 3515.750 2172.430 3516.030 2172.710 ;
        RECT 3516.460 2172.430 3516.740 2172.710 ;
        RECT 3517.170 2172.430 3517.450 2172.710 ;
        RECT 3517.880 2172.430 3518.160 2172.710 ;
        RECT 3518.590 2172.430 3518.870 2172.710 ;
        RECT 3519.300 2172.430 3519.580 2172.710 ;
        RECT 3520.010 2172.430 3520.290 2172.710 ;
        RECT 3520.720 2172.430 3521.000 2172.710 ;
        RECT 3521.430 2172.430 3521.710 2172.710 ;
        RECT 3512.200 2171.720 3512.480 2172.000 ;
        RECT 3512.910 2171.720 3513.190 2172.000 ;
        RECT 3513.620 2171.720 3513.900 2172.000 ;
        RECT 3514.330 2171.720 3514.610 2172.000 ;
        RECT 3515.040 2171.720 3515.320 2172.000 ;
        RECT 3515.750 2171.720 3516.030 2172.000 ;
        RECT 3516.460 2171.720 3516.740 2172.000 ;
        RECT 3517.170 2171.720 3517.450 2172.000 ;
        RECT 3517.880 2171.720 3518.160 2172.000 ;
        RECT 3518.590 2171.720 3518.870 2172.000 ;
        RECT 3519.300 2171.720 3519.580 2172.000 ;
        RECT 3520.010 2171.720 3520.290 2172.000 ;
        RECT 3520.720 2171.720 3521.000 2172.000 ;
        RECT 3521.430 2171.720 3521.710 2172.000 ;
        RECT 3512.200 2171.010 3512.480 2171.290 ;
        RECT 3512.910 2171.010 3513.190 2171.290 ;
        RECT 3513.620 2171.010 3513.900 2171.290 ;
        RECT 3514.330 2171.010 3514.610 2171.290 ;
        RECT 3515.040 2171.010 3515.320 2171.290 ;
        RECT 3515.750 2171.010 3516.030 2171.290 ;
        RECT 3516.460 2171.010 3516.740 2171.290 ;
        RECT 3517.170 2171.010 3517.450 2171.290 ;
        RECT 3517.880 2171.010 3518.160 2171.290 ;
        RECT 3518.590 2171.010 3518.870 2171.290 ;
        RECT 3519.300 2171.010 3519.580 2171.290 ;
        RECT 3520.010 2171.010 3520.290 2171.290 ;
        RECT 3520.720 2171.010 3521.000 2171.290 ;
        RECT 3521.430 2171.010 3521.710 2171.290 ;
        RECT 3512.200 2170.300 3512.480 2170.580 ;
        RECT 3512.910 2170.300 3513.190 2170.580 ;
        RECT 3513.620 2170.300 3513.900 2170.580 ;
        RECT 3514.330 2170.300 3514.610 2170.580 ;
        RECT 3515.040 2170.300 3515.320 2170.580 ;
        RECT 3515.750 2170.300 3516.030 2170.580 ;
        RECT 3516.460 2170.300 3516.740 2170.580 ;
        RECT 3517.170 2170.300 3517.450 2170.580 ;
        RECT 3517.880 2170.300 3518.160 2170.580 ;
        RECT 3518.590 2170.300 3518.870 2170.580 ;
        RECT 3519.300 2170.300 3519.580 2170.580 ;
        RECT 3520.010 2170.300 3520.290 2170.580 ;
        RECT 3520.720 2170.300 3521.000 2170.580 ;
        RECT 3521.430 2170.300 3521.710 2170.580 ;
        RECT 3512.200 2169.590 3512.480 2169.870 ;
        RECT 3512.910 2169.590 3513.190 2169.870 ;
        RECT 3513.620 2169.590 3513.900 2169.870 ;
        RECT 3514.330 2169.590 3514.610 2169.870 ;
        RECT 3515.040 2169.590 3515.320 2169.870 ;
        RECT 3515.750 2169.590 3516.030 2169.870 ;
        RECT 3516.460 2169.590 3516.740 2169.870 ;
        RECT 3517.170 2169.590 3517.450 2169.870 ;
        RECT 3517.880 2169.590 3518.160 2169.870 ;
        RECT 3518.590 2169.590 3518.870 2169.870 ;
        RECT 3519.300 2169.590 3519.580 2169.870 ;
        RECT 3520.010 2169.590 3520.290 2169.870 ;
        RECT 3520.720 2169.590 3521.000 2169.870 ;
        RECT 3521.430 2169.590 3521.710 2169.870 ;
        RECT 3512.200 2168.880 3512.480 2169.160 ;
        RECT 3512.910 2168.880 3513.190 2169.160 ;
        RECT 3513.620 2168.880 3513.900 2169.160 ;
        RECT 3514.330 2168.880 3514.610 2169.160 ;
        RECT 3515.040 2168.880 3515.320 2169.160 ;
        RECT 3515.750 2168.880 3516.030 2169.160 ;
        RECT 3516.460 2168.880 3516.740 2169.160 ;
        RECT 3517.170 2168.880 3517.450 2169.160 ;
        RECT 3517.880 2168.880 3518.160 2169.160 ;
        RECT 3518.590 2168.880 3518.870 2169.160 ;
        RECT 3519.300 2168.880 3519.580 2169.160 ;
        RECT 3520.010 2168.880 3520.290 2169.160 ;
        RECT 3520.720 2168.880 3521.000 2169.160 ;
        RECT 3521.430 2168.880 3521.710 2169.160 ;
        RECT 3512.200 2168.170 3512.480 2168.450 ;
        RECT 3512.910 2168.170 3513.190 2168.450 ;
        RECT 3513.620 2168.170 3513.900 2168.450 ;
        RECT 3514.330 2168.170 3514.610 2168.450 ;
        RECT 3515.040 2168.170 3515.320 2168.450 ;
        RECT 3515.750 2168.170 3516.030 2168.450 ;
        RECT 3516.460 2168.170 3516.740 2168.450 ;
        RECT 3517.170 2168.170 3517.450 2168.450 ;
        RECT 3517.880 2168.170 3518.160 2168.450 ;
        RECT 3518.590 2168.170 3518.870 2168.450 ;
        RECT 3519.300 2168.170 3519.580 2168.450 ;
        RECT 3520.010 2168.170 3520.290 2168.450 ;
        RECT 3520.720 2168.170 3521.000 2168.450 ;
        RECT 3521.430 2168.170 3521.710 2168.450 ;
        RECT 3512.200 2167.460 3512.480 2167.740 ;
        RECT 3512.910 2167.460 3513.190 2167.740 ;
        RECT 3513.620 2167.460 3513.900 2167.740 ;
        RECT 3514.330 2167.460 3514.610 2167.740 ;
        RECT 3515.040 2167.460 3515.320 2167.740 ;
        RECT 3515.750 2167.460 3516.030 2167.740 ;
        RECT 3516.460 2167.460 3516.740 2167.740 ;
        RECT 3517.170 2167.460 3517.450 2167.740 ;
        RECT 3517.880 2167.460 3518.160 2167.740 ;
        RECT 3518.590 2167.460 3518.870 2167.740 ;
        RECT 3519.300 2167.460 3519.580 2167.740 ;
        RECT 3520.010 2167.460 3520.290 2167.740 ;
        RECT 3520.720 2167.460 3521.000 2167.740 ;
        RECT 3521.430 2167.460 3521.710 2167.740 ;
        RECT 3512.200 2166.750 3512.480 2167.030 ;
        RECT 3512.910 2166.750 3513.190 2167.030 ;
        RECT 3513.620 2166.750 3513.900 2167.030 ;
        RECT 3514.330 2166.750 3514.610 2167.030 ;
        RECT 3515.040 2166.750 3515.320 2167.030 ;
        RECT 3515.750 2166.750 3516.030 2167.030 ;
        RECT 3516.460 2166.750 3516.740 2167.030 ;
        RECT 3517.170 2166.750 3517.450 2167.030 ;
        RECT 3517.880 2166.750 3518.160 2167.030 ;
        RECT 3518.590 2166.750 3518.870 2167.030 ;
        RECT 3519.300 2166.750 3519.580 2167.030 ;
        RECT 3520.010 2166.750 3520.290 2167.030 ;
        RECT 3520.720 2166.750 3521.000 2167.030 ;
        RECT 3521.430 2166.750 3521.710 2167.030 ;
        RECT 357.330 2137.970 357.610 2138.250 ;
        RECT 358.040 2137.970 358.320 2138.250 ;
        RECT 358.750 2137.970 359.030 2138.250 ;
        RECT 359.460 2137.970 359.740 2138.250 ;
        RECT 360.170 2137.970 360.450 2138.250 ;
        RECT 360.880 2137.970 361.160 2138.250 ;
        RECT 361.590 2137.970 361.870 2138.250 ;
        RECT 362.300 2137.970 362.580 2138.250 ;
        RECT 363.010 2137.970 363.290 2138.250 ;
        RECT 363.720 2137.970 364.000 2138.250 ;
        RECT 364.430 2137.970 364.710 2138.250 ;
        RECT 365.140 2137.970 365.420 2138.250 ;
        RECT 365.850 2137.970 366.130 2138.250 ;
        RECT 366.560 2137.970 366.840 2138.250 ;
        RECT 357.330 2137.260 357.610 2137.540 ;
        RECT 358.040 2137.260 358.320 2137.540 ;
        RECT 358.750 2137.260 359.030 2137.540 ;
        RECT 359.460 2137.260 359.740 2137.540 ;
        RECT 360.170 2137.260 360.450 2137.540 ;
        RECT 360.880 2137.260 361.160 2137.540 ;
        RECT 361.590 2137.260 361.870 2137.540 ;
        RECT 362.300 2137.260 362.580 2137.540 ;
        RECT 363.010 2137.260 363.290 2137.540 ;
        RECT 363.720 2137.260 364.000 2137.540 ;
        RECT 364.430 2137.260 364.710 2137.540 ;
        RECT 365.140 2137.260 365.420 2137.540 ;
        RECT 365.850 2137.260 366.130 2137.540 ;
        RECT 366.560 2137.260 366.840 2137.540 ;
        RECT 357.330 2136.550 357.610 2136.830 ;
        RECT 358.040 2136.550 358.320 2136.830 ;
        RECT 358.750 2136.550 359.030 2136.830 ;
        RECT 359.460 2136.550 359.740 2136.830 ;
        RECT 360.170 2136.550 360.450 2136.830 ;
        RECT 360.880 2136.550 361.160 2136.830 ;
        RECT 361.590 2136.550 361.870 2136.830 ;
        RECT 362.300 2136.550 362.580 2136.830 ;
        RECT 363.010 2136.550 363.290 2136.830 ;
        RECT 363.720 2136.550 364.000 2136.830 ;
        RECT 364.430 2136.550 364.710 2136.830 ;
        RECT 365.140 2136.550 365.420 2136.830 ;
        RECT 365.850 2136.550 366.130 2136.830 ;
        RECT 366.560 2136.550 366.840 2136.830 ;
        RECT 357.330 2135.840 357.610 2136.120 ;
        RECT 358.040 2135.840 358.320 2136.120 ;
        RECT 358.750 2135.840 359.030 2136.120 ;
        RECT 359.460 2135.840 359.740 2136.120 ;
        RECT 360.170 2135.840 360.450 2136.120 ;
        RECT 360.880 2135.840 361.160 2136.120 ;
        RECT 361.590 2135.840 361.870 2136.120 ;
        RECT 362.300 2135.840 362.580 2136.120 ;
        RECT 363.010 2135.840 363.290 2136.120 ;
        RECT 363.720 2135.840 364.000 2136.120 ;
        RECT 364.430 2135.840 364.710 2136.120 ;
        RECT 365.140 2135.840 365.420 2136.120 ;
        RECT 365.850 2135.840 366.130 2136.120 ;
        RECT 366.560 2135.840 366.840 2136.120 ;
        RECT 357.330 2135.130 357.610 2135.410 ;
        RECT 358.040 2135.130 358.320 2135.410 ;
        RECT 358.750 2135.130 359.030 2135.410 ;
        RECT 359.460 2135.130 359.740 2135.410 ;
        RECT 360.170 2135.130 360.450 2135.410 ;
        RECT 360.880 2135.130 361.160 2135.410 ;
        RECT 361.590 2135.130 361.870 2135.410 ;
        RECT 362.300 2135.130 362.580 2135.410 ;
        RECT 363.010 2135.130 363.290 2135.410 ;
        RECT 363.720 2135.130 364.000 2135.410 ;
        RECT 364.430 2135.130 364.710 2135.410 ;
        RECT 365.140 2135.130 365.420 2135.410 ;
        RECT 365.850 2135.130 366.130 2135.410 ;
        RECT 366.560 2135.130 366.840 2135.410 ;
        RECT 357.330 2134.420 357.610 2134.700 ;
        RECT 358.040 2134.420 358.320 2134.700 ;
        RECT 358.750 2134.420 359.030 2134.700 ;
        RECT 359.460 2134.420 359.740 2134.700 ;
        RECT 360.170 2134.420 360.450 2134.700 ;
        RECT 360.880 2134.420 361.160 2134.700 ;
        RECT 361.590 2134.420 361.870 2134.700 ;
        RECT 362.300 2134.420 362.580 2134.700 ;
        RECT 363.010 2134.420 363.290 2134.700 ;
        RECT 363.720 2134.420 364.000 2134.700 ;
        RECT 364.430 2134.420 364.710 2134.700 ;
        RECT 365.140 2134.420 365.420 2134.700 ;
        RECT 365.850 2134.420 366.130 2134.700 ;
        RECT 366.560 2134.420 366.840 2134.700 ;
        RECT 357.330 2133.710 357.610 2133.990 ;
        RECT 358.040 2133.710 358.320 2133.990 ;
        RECT 358.750 2133.710 359.030 2133.990 ;
        RECT 359.460 2133.710 359.740 2133.990 ;
        RECT 360.170 2133.710 360.450 2133.990 ;
        RECT 360.880 2133.710 361.160 2133.990 ;
        RECT 361.590 2133.710 361.870 2133.990 ;
        RECT 362.300 2133.710 362.580 2133.990 ;
        RECT 363.010 2133.710 363.290 2133.990 ;
        RECT 363.720 2133.710 364.000 2133.990 ;
        RECT 364.430 2133.710 364.710 2133.990 ;
        RECT 365.140 2133.710 365.420 2133.990 ;
        RECT 365.850 2133.710 366.130 2133.990 ;
        RECT 366.560 2133.710 366.840 2133.990 ;
        RECT 357.330 2133.000 357.610 2133.280 ;
        RECT 358.040 2133.000 358.320 2133.280 ;
        RECT 358.750 2133.000 359.030 2133.280 ;
        RECT 359.460 2133.000 359.740 2133.280 ;
        RECT 360.170 2133.000 360.450 2133.280 ;
        RECT 360.880 2133.000 361.160 2133.280 ;
        RECT 361.590 2133.000 361.870 2133.280 ;
        RECT 362.300 2133.000 362.580 2133.280 ;
        RECT 363.010 2133.000 363.290 2133.280 ;
        RECT 363.720 2133.000 364.000 2133.280 ;
        RECT 364.430 2133.000 364.710 2133.280 ;
        RECT 365.140 2133.000 365.420 2133.280 ;
        RECT 365.850 2133.000 366.130 2133.280 ;
        RECT 366.560 2133.000 366.840 2133.280 ;
        RECT 357.330 2132.290 357.610 2132.570 ;
        RECT 358.040 2132.290 358.320 2132.570 ;
        RECT 358.750 2132.290 359.030 2132.570 ;
        RECT 359.460 2132.290 359.740 2132.570 ;
        RECT 360.170 2132.290 360.450 2132.570 ;
        RECT 360.880 2132.290 361.160 2132.570 ;
        RECT 361.590 2132.290 361.870 2132.570 ;
        RECT 362.300 2132.290 362.580 2132.570 ;
        RECT 363.010 2132.290 363.290 2132.570 ;
        RECT 363.720 2132.290 364.000 2132.570 ;
        RECT 364.430 2132.290 364.710 2132.570 ;
        RECT 365.140 2132.290 365.420 2132.570 ;
        RECT 365.850 2132.290 366.130 2132.570 ;
        RECT 366.560 2132.290 366.840 2132.570 ;
        RECT 357.330 2131.580 357.610 2131.860 ;
        RECT 358.040 2131.580 358.320 2131.860 ;
        RECT 358.750 2131.580 359.030 2131.860 ;
        RECT 359.460 2131.580 359.740 2131.860 ;
        RECT 360.170 2131.580 360.450 2131.860 ;
        RECT 360.880 2131.580 361.160 2131.860 ;
        RECT 361.590 2131.580 361.870 2131.860 ;
        RECT 362.300 2131.580 362.580 2131.860 ;
        RECT 363.010 2131.580 363.290 2131.860 ;
        RECT 363.720 2131.580 364.000 2131.860 ;
        RECT 364.430 2131.580 364.710 2131.860 ;
        RECT 365.140 2131.580 365.420 2131.860 ;
        RECT 365.850 2131.580 366.130 2131.860 ;
        RECT 366.560 2131.580 366.840 2131.860 ;
        RECT 357.330 2130.870 357.610 2131.150 ;
        RECT 358.040 2130.870 358.320 2131.150 ;
        RECT 358.750 2130.870 359.030 2131.150 ;
        RECT 359.460 2130.870 359.740 2131.150 ;
        RECT 360.170 2130.870 360.450 2131.150 ;
        RECT 360.880 2130.870 361.160 2131.150 ;
        RECT 361.590 2130.870 361.870 2131.150 ;
        RECT 362.300 2130.870 362.580 2131.150 ;
        RECT 363.010 2130.870 363.290 2131.150 ;
        RECT 363.720 2130.870 364.000 2131.150 ;
        RECT 364.430 2130.870 364.710 2131.150 ;
        RECT 365.140 2130.870 365.420 2131.150 ;
        RECT 365.850 2130.870 366.130 2131.150 ;
        RECT 366.560 2130.870 366.840 2131.150 ;
        RECT 357.330 2130.160 357.610 2130.440 ;
        RECT 358.040 2130.160 358.320 2130.440 ;
        RECT 358.750 2130.160 359.030 2130.440 ;
        RECT 359.460 2130.160 359.740 2130.440 ;
        RECT 360.170 2130.160 360.450 2130.440 ;
        RECT 360.880 2130.160 361.160 2130.440 ;
        RECT 361.590 2130.160 361.870 2130.440 ;
        RECT 362.300 2130.160 362.580 2130.440 ;
        RECT 363.010 2130.160 363.290 2130.440 ;
        RECT 363.720 2130.160 364.000 2130.440 ;
        RECT 364.430 2130.160 364.710 2130.440 ;
        RECT 365.140 2130.160 365.420 2130.440 ;
        RECT 365.850 2130.160 366.130 2130.440 ;
        RECT 366.560 2130.160 366.840 2130.440 ;
        RECT 357.330 2129.450 357.610 2129.730 ;
        RECT 358.040 2129.450 358.320 2129.730 ;
        RECT 358.750 2129.450 359.030 2129.730 ;
        RECT 359.460 2129.450 359.740 2129.730 ;
        RECT 360.170 2129.450 360.450 2129.730 ;
        RECT 360.880 2129.450 361.160 2129.730 ;
        RECT 361.590 2129.450 361.870 2129.730 ;
        RECT 362.300 2129.450 362.580 2129.730 ;
        RECT 363.010 2129.450 363.290 2129.730 ;
        RECT 363.720 2129.450 364.000 2129.730 ;
        RECT 364.430 2129.450 364.710 2129.730 ;
        RECT 365.140 2129.450 365.420 2129.730 ;
        RECT 365.850 2129.450 366.130 2129.730 ;
        RECT 366.560 2129.450 366.840 2129.730 ;
        RECT 357.275 2125.565 357.555 2125.845 ;
        RECT 357.985 2125.565 358.265 2125.845 ;
        RECT 358.695 2125.565 358.975 2125.845 ;
        RECT 359.405 2125.565 359.685 2125.845 ;
        RECT 360.115 2125.565 360.395 2125.845 ;
        RECT 360.825 2125.565 361.105 2125.845 ;
        RECT 361.535 2125.565 361.815 2125.845 ;
        RECT 362.245 2125.565 362.525 2125.845 ;
        RECT 362.955 2125.565 363.235 2125.845 ;
        RECT 363.665 2125.565 363.945 2125.845 ;
        RECT 364.375 2125.565 364.655 2125.845 ;
        RECT 365.085 2125.565 365.365 2125.845 ;
        RECT 365.795 2125.565 366.075 2125.845 ;
        RECT 366.505 2125.565 366.785 2125.845 ;
        RECT 357.275 2124.855 357.555 2125.135 ;
        RECT 357.985 2124.855 358.265 2125.135 ;
        RECT 358.695 2124.855 358.975 2125.135 ;
        RECT 359.405 2124.855 359.685 2125.135 ;
        RECT 360.115 2124.855 360.395 2125.135 ;
        RECT 360.825 2124.855 361.105 2125.135 ;
        RECT 361.535 2124.855 361.815 2125.135 ;
        RECT 362.245 2124.855 362.525 2125.135 ;
        RECT 362.955 2124.855 363.235 2125.135 ;
        RECT 363.665 2124.855 363.945 2125.135 ;
        RECT 364.375 2124.855 364.655 2125.135 ;
        RECT 365.085 2124.855 365.365 2125.135 ;
        RECT 365.795 2124.855 366.075 2125.135 ;
        RECT 366.505 2124.855 366.785 2125.135 ;
        RECT 357.275 2124.145 357.555 2124.425 ;
        RECT 357.985 2124.145 358.265 2124.425 ;
        RECT 358.695 2124.145 358.975 2124.425 ;
        RECT 359.405 2124.145 359.685 2124.425 ;
        RECT 360.115 2124.145 360.395 2124.425 ;
        RECT 360.825 2124.145 361.105 2124.425 ;
        RECT 361.535 2124.145 361.815 2124.425 ;
        RECT 362.245 2124.145 362.525 2124.425 ;
        RECT 362.955 2124.145 363.235 2124.425 ;
        RECT 363.665 2124.145 363.945 2124.425 ;
        RECT 364.375 2124.145 364.655 2124.425 ;
        RECT 365.085 2124.145 365.365 2124.425 ;
        RECT 365.795 2124.145 366.075 2124.425 ;
        RECT 366.505 2124.145 366.785 2124.425 ;
        RECT 357.275 2123.435 357.555 2123.715 ;
        RECT 357.985 2123.435 358.265 2123.715 ;
        RECT 358.695 2123.435 358.975 2123.715 ;
        RECT 359.405 2123.435 359.685 2123.715 ;
        RECT 360.115 2123.435 360.395 2123.715 ;
        RECT 360.825 2123.435 361.105 2123.715 ;
        RECT 361.535 2123.435 361.815 2123.715 ;
        RECT 362.245 2123.435 362.525 2123.715 ;
        RECT 362.955 2123.435 363.235 2123.715 ;
        RECT 363.665 2123.435 363.945 2123.715 ;
        RECT 364.375 2123.435 364.655 2123.715 ;
        RECT 365.085 2123.435 365.365 2123.715 ;
        RECT 365.795 2123.435 366.075 2123.715 ;
        RECT 366.505 2123.435 366.785 2123.715 ;
        RECT 357.275 2122.725 357.555 2123.005 ;
        RECT 357.985 2122.725 358.265 2123.005 ;
        RECT 358.695 2122.725 358.975 2123.005 ;
        RECT 359.405 2122.725 359.685 2123.005 ;
        RECT 360.115 2122.725 360.395 2123.005 ;
        RECT 360.825 2122.725 361.105 2123.005 ;
        RECT 361.535 2122.725 361.815 2123.005 ;
        RECT 362.245 2122.725 362.525 2123.005 ;
        RECT 362.955 2122.725 363.235 2123.005 ;
        RECT 363.665 2122.725 363.945 2123.005 ;
        RECT 364.375 2122.725 364.655 2123.005 ;
        RECT 365.085 2122.725 365.365 2123.005 ;
        RECT 365.795 2122.725 366.075 2123.005 ;
        RECT 366.505 2122.725 366.785 2123.005 ;
        RECT 357.275 2122.015 357.555 2122.295 ;
        RECT 357.985 2122.015 358.265 2122.295 ;
        RECT 358.695 2122.015 358.975 2122.295 ;
        RECT 359.405 2122.015 359.685 2122.295 ;
        RECT 360.115 2122.015 360.395 2122.295 ;
        RECT 360.825 2122.015 361.105 2122.295 ;
        RECT 361.535 2122.015 361.815 2122.295 ;
        RECT 362.245 2122.015 362.525 2122.295 ;
        RECT 362.955 2122.015 363.235 2122.295 ;
        RECT 363.665 2122.015 363.945 2122.295 ;
        RECT 364.375 2122.015 364.655 2122.295 ;
        RECT 365.085 2122.015 365.365 2122.295 ;
        RECT 365.795 2122.015 366.075 2122.295 ;
        RECT 366.505 2122.015 366.785 2122.295 ;
        RECT 357.275 2121.305 357.555 2121.585 ;
        RECT 357.985 2121.305 358.265 2121.585 ;
        RECT 358.695 2121.305 358.975 2121.585 ;
        RECT 359.405 2121.305 359.685 2121.585 ;
        RECT 360.115 2121.305 360.395 2121.585 ;
        RECT 360.825 2121.305 361.105 2121.585 ;
        RECT 361.535 2121.305 361.815 2121.585 ;
        RECT 362.245 2121.305 362.525 2121.585 ;
        RECT 362.955 2121.305 363.235 2121.585 ;
        RECT 363.665 2121.305 363.945 2121.585 ;
        RECT 364.375 2121.305 364.655 2121.585 ;
        RECT 365.085 2121.305 365.365 2121.585 ;
        RECT 365.795 2121.305 366.075 2121.585 ;
        RECT 366.505 2121.305 366.785 2121.585 ;
        RECT 357.275 2120.595 357.555 2120.875 ;
        RECT 357.985 2120.595 358.265 2120.875 ;
        RECT 358.695 2120.595 358.975 2120.875 ;
        RECT 359.405 2120.595 359.685 2120.875 ;
        RECT 360.115 2120.595 360.395 2120.875 ;
        RECT 360.825 2120.595 361.105 2120.875 ;
        RECT 361.535 2120.595 361.815 2120.875 ;
        RECT 362.245 2120.595 362.525 2120.875 ;
        RECT 362.955 2120.595 363.235 2120.875 ;
        RECT 363.665 2120.595 363.945 2120.875 ;
        RECT 364.375 2120.595 364.655 2120.875 ;
        RECT 365.085 2120.595 365.365 2120.875 ;
        RECT 365.795 2120.595 366.075 2120.875 ;
        RECT 366.505 2120.595 366.785 2120.875 ;
        RECT 357.275 2119.885 357.555 2120.165 ;
        RECT 357.985 2119.885 358.265 2120.165 ;
        RECT 358.695 2119.885 358.975 2120.165 ;
        RECT 359.405 2119.885 359.685 2120.165 ;
        RECT 360.115 2119.885 360.395 2120.165 ;
        RECT 360.825 2119.885 361.105 2120.165 ;
        RECT 361.535 2119.885 361.815 2120.165 ;
        RECT 362.245 2119.885 362.525 2120.165 ;
        RECT 362.955 2119.885 363.235 2120.165 ;
        RECT 363.665 2119.885 363.945 2120.165 ;
        RECT 364.375 2119.885 364.655 2120.165 ;
        RECT 365.085 2119.885 365.365 2120.165 ;
        RECT 365.795 2119.885 366.075 2120.165 ;
        RECT 366.505 2119.885 366.785 2120.165 ;
        RECT 357.275 2119.175 357.555 2119.455 ;
        RECT 357.985 2119.175 358.265 2119.455 ;
        RECT 358.695 2119.175 358.975 2119.455 ;
        RECT 359.405 2119.175 359.685 2119.455 ;
        RECT 360.115 2119.175 360.395 2119.455 ;
        RECT 360.825 2119.175 361.105 2119.455 ;
        RECT 361.535 2119.175 361.815 2119.455 ;
        RECT 362.245 2119.175 362.525 2119.455 ;
        RECT 362.955 2119.175 363.235 2119.455 ;
        RECT 363.665 2119.175 363.945 2119.455 ;
        RECT 364.375 2119.175 364.655 2119.455 ;
        RECT 365.085 2119.175 365.365 2119.455 ;
        RECT 365.795 2119.175 366.075 2119.455 ;
        RECT 366.505 2119.175 366.785 2119.455 ;
        RECT 357.275 2118.465 357.555 2118.745 ;
        RECT 357.985 2118.465 358.265 2118.745 ;
        RECT 358.695 2118.465 358.975 2118.745 ;
        RECT 359.405 2118.465 359.685 2118.745 ;
        RECT 360.115 2118.465 360.395 2118.745 ;
        RECT 360.825 2118.465 361.105 2118.745 ;
        RECT 361.535 2118.465 361.815 2118.745 ;
        RECT 362.245 2118.465 362.525 2118.745 ;
        RECT 362.955 2118.465 363.235 2118.745 ;
        RECT 363.665 2118.465 363.945 2118.745 ;
        RECT 364.375 2118.465 364.655 2118.745 ;
        RECT 365.085 2118.465 365.365 2118.745 ;
        RECT 365.795 2118.465 366.075 2118.745 ;
        RECT 366.505 2118.465 366.785 2118.745 ;
        RECT 357.275 2117.755 357.555 2118.035 ;
        RECT 357.985 2117.755 358.265 2118.035 ;
        RECT 358.695 2117.755 358.975 2118.035 ;
        RECT 359.405 2117.755 359.685 2118.035 ;
        RECT 360.115 2117.755 360.395 2118.035 ;
        RECT 360.825 2117.755 361.105 2118.035 ;
        RECT 361.535 2117.755 361.815 2118.035 ;
        RECT 362.245 2117.755 362.525 2118.035 ;
        RECT 362.955 2117.755 363.235 2118.035 ;
        RECT 363.665 2117.755 363.945 2118.035 ;
        RECT 364.375 2117.755 364.655 2118.035 ;
        RECT 365.085 2117.755 365.365 2118.035 ;
        RECT 365.795 2117.755 366.075 2118.035 ;
        RECT 366.505 2117.755 366.785 2118.035 ;
        RECT 357.275 2117.045 357.555 2117.325 ;
        RECT 357.985 2117.045 358.265 2117.325 ;
        RECT 358.695 2117.045 358.975 2117.325 ;
        RECT 359.405 2117.045 359.685 2117.325 ;
        RECT 360.115 2117.045 360.395 2117.325 ;
        RECT 360.825 2117.045 361.105 2117.325 ;
        RECT 361.535 2117.045 361.815 2117.325 ;
        RECT 362.245 2117.045 362.525 2117.325 ;
        RECT 362.955 2117.045 363.235 2117.325 ;
        RECT 363.665 2117.045 363.945 2117.325 ;
        RECT 364.375 2117.045 364.655 2117.325 ;
        RECT 365.085 2117.045 365.365 2117.325 ;
        RECT 365.795 2117.045 366.075 2117.325 ;
        RECT 366.505 2117.045 366.785 2117.325 ;
        RECT 357.275 2116.335 357.555 2116.615 ;
        RECT 357.985 2116.335 358.265 2116.615 ;
        RECT 358.695 2116.335 358.975 2116.615 ;
        RECT 359.405 2116.335 359.685 2116.615 ;
        RECT 360.115 2116.335 360.395 2116.615 ;
        RECT 360.825 2116.335 361.105 2116.615 ;
        RECT 361.535 2116.335 361.815 2116.615 ;
        RECT 362.245 2116.335 362.525 2116.615 ;
        RECT 362.955 2116.335 363.235 2116.615 ;
        RECT 363.665 2116.335 363.945 2116.615 ;
        RECT 364.375 2116.335 364.655 2116.615 ;
        RECT 365.085 2116.335 365.365 2116.615 ;
        RECT 365.795 2116.335 366.075 2116.615 ;
        RECT 366.505 2116.335 366.785 2116.615 ;
        RECT 357.275 2113.715 357.555 2113.995 ;
        RECT 357.985 2113.715 358.265 2113.995 ;
        RECT 358.695 2113.715 358.975 2113.995 ;
        RECT 359.405 2113.715 359.685 2113.995 ;
        RECT 360.115 2113.715 360.395 2113.995 ;
        RECT 360.825 2113.715 361.105 2113.995 ;
        RECT 361.535 2113.715 361.815 2113.995 ;
        RECT 362.245 2113.715 362.525 2113.995 ;
        RECT 362.955 2113.715 363.235 2113.995 ;
        RECT 363.665 2113.715 363.945 2113.995 ;
        RECT 364.375 2113.715 364.655 2113.995 ;
        RECT 365.085 2113.715 365.365 2113.995 ;
        RECT 365.795 2113.715 366.075 2113.995 ;
        RECT 366.505 2113.715 366.785 2113.995 ;
        RECT 357.275 2113.005 357.555 2113.285 ;
        RECT 357.985 2113.005 358.265 2113.285 ;
        RECT 358.695 2113.005 358.975 2113.285 ;
        RECT 359.405 2113.005 359.685 2113.285 ;
        RECT 360.115 2113.005 360.395 2113.285 ;
        RECT 360.825 2113.005 361.105 2113.285 ;
        RECT 361.535 2113.005 361.815 2113.285 ;
        RECT 362.245 2113.005 362.525 2113.285 ;
        RECT 362.955 2113.005 363.235 2113.285 ;
        RECT 363.665 2113.005 363.945 2113.285 ;
        RECT 364.375 2113.005 364.655 2113.285 ;
        RECT 365.085 2113.005 365.365 2113.285 ;
        RECT 365.795 2113.005 366.075 2113.285 ;
        RECT 366.505 2113.005 366.785 2113.285 ;
        RECT 357.275 2112.295 357.555 2112.575 ;
        RECT 357.985 2112.295 358.265 2112.575 ;
        RECT 358.695 2112.295 358.975 2112.575 ;
        RECT 359.405 2112.295 359.685 2112.575 ;
        RECT 360.115 2112.295 360.395 2112.575 ;
        RECT 360.825 2112.295 361.105 2112.575 ;
        RECT 361.535 2112.295 361.815 2112.575 ;
        RECT 362.245 2112.295 362.525 2112.575 ;
        RECT 362.955 2112.295 363.235 2112.575 ;
        RECT 363.665 2112.295 363.945 2112.575 ;
        RECT 364.375 2112.295 364.655 2112.575 ;
        RECT 365.085 2112.295 365.365 2112.575 ;
        RECT 365.795 2112.295 366.075 2112.575 ;
        RECT 366.505 2112.295 366.785 2112.575 ;
        RECT 357.275 2111.585 357.555 2111.865 ;
        RECT 357.985 2111.585 358.265 2111.865 ;
        RECT 358.695 2111.585 358.975 2111.865 ;
        RECT 359.405 2111.585 359.685 2111.865 ;
        RECT 360.115 2111.585 360.395 2111.865 ;
        RECT 360.825 2111.585 361.105 2111.865 ;
        RECT 361.535 2111.585 361.815 2111.865 ;
        RECT 362.245 2111.585 362.525 2111.865 ;
        RECT 362.955 2111.585 363.235 2111.865 ;
        RECT 363.665 2111.585 363.945 2111.865 ;
        RECT 364.375 2111.585 364.655 2111.865 ;
        RECT 365.085 2111.585 365.365 2111.865 ;
        RECT 365.795 2111.585 366.075 2111.865 ;
        RECT 366.505 2111.585 366.785 2111.865 ;
        RECT 357.275 2110.875 357.555 2111.155 ;
        RECT 357.985 2110.875 358.265 2111.155 ;
        RECT 358.695 2110.875 358.975 2111.155 ;
        RECT 359.405 2110.875 359.685 2111.155 ;
        RECT 360.115 2110.875 360.395 2111.155 ;
        RECT 360.825 2110.875 361.105 2111.155 ;
        RECT 361.535 2110.875 361.815 2111.155 ;
        RECT 362.245 2110.875 362.525 2111.155 ;
        RECT 362.955 2110.875 363.235 2111.155 ;
        RECT 363.665 2110.875 363.945 2111.155 ;
        RECT 364.375 2110.875 364.655 2111.155 ;
        RECT 365.085 2110.875 365.365 2111.155 ;
        RECT 365.795 2110.875 366.075 2111.155 ;
        RECT 366.505 2110.875 366.785 2111.155 ;
        RECT 357.275 2110.165 357.555 2110.445 ;
        RECT 357.985 2110.165 358.265 2110.445 ;
        RECT 358.695 2110.165 358.975 2110.445 ;
        RECT 359.405 2110.165 359.685 2110.445 ;
        RECT 360.115 2110.165 360.395 2110.445 ;
        RECT 360.825 2110.165 361.105 2110.445 ;
        RECT 361.535 2110.165 361.815 2110.445 ;
        RECT 362.245 2110.165 362.525 2110.445 ;
        RECT 362.955 2110.165 363.235 2110.445 ;
        RECT 363.665 2110.165 363.945 2110.445 ;
        RECT 364.375 2110.165 364.655 2110.445 ;
        RECT 365.085 2110.165 365.365 2110.445 ;
        RECT 365.795 2110.165 366.075 2110.445 ;
        RECT 366.505 2110.165 366.785 2110.445 ;
        RECT 357.275 2109.455 357.555 2109.735 ;
        RECT 357.985 2109.455 358.265 2109.735 ;
        RECT 358.695 2109.455 358.975 2109.735 ;
        RECT 359.405 2109.455 359.685 2109.735 ;
        RECT 360.115 2109.455 360.395 2109.735 ;
        RECT 360.825 2109.455 361.105 2109.735 ;
        RECT 361.535 2109.455 361.815 2109.735 ;
        RECT 362.245 2109.455 362.525 2109.735 ;
        RECT 362.955 2109.455 363.235 2109.735 ;
        RECT 363.665 2109.455 363.945 2109.735 ;
        RECT 364.375 2109.455 364.655 2109.735 ;
        RECT 365.085 2109.455 365.365 2109.735 ;
        RECT 365.795 2109.455 366.075 2109.735 ;
        RECT 366.505 2109.455 366.785 2109.735 ;
        RECT 357.275 2108.745 357.555 2109.025 ;
        RECT 357.985 2108.745 358.265 2109.025 ;
        RECT 358.695 2108.745 358.975 2109.025 ;
        RECT 359.405 2108.745 359.685 2109.025 ;
        RECT 360.115 2108.745 360.395 2109.025 ;
        RECT 360.825 2108.745 361.105 2109.025 ;
        RECT 361.535 2108.745 361.815 2109.025 ;
        RECT 362.245 2108.745 362.525 2109.025 ;
        RECT 362.955 2108.745 363.235 2109.025 ;
        RECT 363.665 2108.745 363.945 2109.025 ;
        RECT 364.375 2108.745 364.655 2109.025 ;
        RECT 365.085 2108.745 365.365 2109.025 ;
        RECT 365.795 2108.745 366.075 2109.025 ;
        RECT 366.505 2108.745 366.785 2109.025 ;
        RECT 357.275 2108.035 357.555 2108.315 ;
        RECT 357.985 2108.035 358.265 2108.315 ;
        RECT 358.695 2108.035 358.975 2108.315 ;
        RECT 359.405 2108.035 359.685 2108.315 ;
        RECT 360.115 2108.035 360.395 2108.315 ;
        RECT 360.825 2108.035 361.105 2108.315 ;
        RECT 361.535 2108.035 361.815 2108.315 ;
        RECT 362.245 2108.035 362.525 2108.315 ;
        RECT 362.955 2108.035 363.235 2108.315 ;
        RECT 363.665 2108.035 363.945 2108.315 ;
        RECT 364.375 2108.035 364.655 2108.315 ;
        RECT 365.085 2108.035 365.365 2108.315 ;
        RECT 365.795 2108.035 366.075 2108.315 ;
        RECT 366.505 2108.035 366.785 2108.315 ;
        RECT 357.275 2107.325 357.555 2107.605 ;
        RECT 357.985 2107.325 358.265 2107.605 ;
        RECT 358.695 2107.325 358.975 2107.605 ;
        RECT 359.405 2107.325 359.685 2107.605 ;
        RECT 360.115 2107.325 360.395 2107.605 ;
        RECT 360.825 2107.325 361.105 2107.605 ;
        RECT 361.535 2107.325 361.815 2107.605 ;
        RECT 362.245 2107.325 362.525 2107.605 ;
        RECT 362.955 2107.325 363.235 2107.605 ;
        RECT 363.665 2107.325 363.945 2107.605 ;
        RECT 364.375 2107.325 364.655 2107.605 ;
        RECT 365.085 2107.325 365.365 2107.605 ;
        RECT 365.795 2107.325 366.075 2107.605 ;
        RECT 366.505 2107.325 366.785 2107.605 ;
        RECT 357.275 2106.615 357.555 2106.895 ;
        RECT 357.985 2106.615 358.265 2106.895 ;
        RECT 358.695 2106.615 358.975 2106.895 ;
        RECT 359.405 2106.615 359.685 2106.895 ;
        RECT 360.115 2106.615 360.395 2106.895 ;
        RECT 360.825 2106.615 361.105 2106.895 ;
        RECT 361.535 2106.615 361.815 2106.895 ;
        RECT 362.245 2106.615 362.525 2106.895 ;
        RECT 362.955 2106.615 363.235 2106.895 ;
        RECT 363.665 2106.615 363.945 2106.895 ;
        RECT 364.375 2106.615 364.655 2106.895 ;
        RECT 365.085 2106.615 365.365 2106.895 ;
        RECT 365.795 2106.615 366.075 2106.895 ;
        RECT 366.505 2106.615 366.785 2106.895 ;
        RECT 357.275 2105.905 357.555 2106.185 ;
        RECT 357.985 2105.905 358.265 2106.185 ;
        RECT 358.695 2105.905 358.975 2106.185 ;
        RECT 359.405 2105.905 359.685 2106.185 ;
        RECT 360.115 2105.905 360.395 2106.185 ;
        RECT 360.825 2105.905 361.105 2106.185 ;
        RECT 361.535 2105.905 361.815 2106.185 ;
        RECT 362.245 2105.905 362.525 2106.185 ;
        RECT 362.955 2105.905 363.235 2106.185 ;
        RECT 363.665 2105.905 363.945 2106.185 ;
        RECT 364.375 2105.905 364.655 2106.185 ;
        RECT 365.085 2105.905 365.365 2106.185 ;
        RECT 365.795 2105.905 366.075 2106.185 ;
        RECT 366.505 2105.905 366.785 2106.185 ;
        RECT 357.275 2105.195 357.555 2105.475 ;
        RECT 357.985 2105.195 358.265 2105.475 ;
        RECT 358.695 2105.195 358.975 2105.475 ;
        RECT 359.405 2105.195 359.685 2105.475 ;
        RECT 360.115 2105.195 360.395 2105.475 ;
        RECT 360.825 2105.195 361.105 2105.475 ;
        RECT 361.535 2105.195 361.815 2105.475 ;
        RECT 362.245 2105.195 362.525 2105.475 ;
        RECT 362.955 2105.195 363.235 2105.475 ;
        RECT 363.665 2105.195 363.945 2105.475 ;
        RECT 364.375 2105.195 364.655 2105.475 ;
        RECT 365.085 2105.195 365.365 2105.475 ;
        RECT 365.795 2105.195 366.075 2105.475 ;
        RECT 366.505 2105.195 366.785 2105.475 ;
        RECT 357.275 2104.485 357.555 2104.765 ;
        RECT 357.985 2104.485 358.265 2104.765 ;
        RECT 358.695 2104.485 358.975 2104.765 ;
        RECT 359.405 2104.485 359.685 2104.765 ;
        RECT 360.115 2104.485 360.395 2104.765 ;
        RECT 360.825 2104.485 361.105 2104.765 ;
        RECT 361.535 2104.485 361.815 2104.765 ;
        RECT 362.245 2104.485 362.525 2104.765 ;
        RECT 362.955 2104.485 363.235 2104.765 ;
        RECT 363.665 2104.485 363.945 2104.765 ;
        RECT 364.375 2104.485 364.655 2104.765 ;
        RECT 365.085 2104.485 365.365 2104.765 ;
        RECT 365.795 2104.485 366.075 2104.765 ;
        RECT 366.505 2104.485 366.785 2104.765 ;
        RECT 357.275 2100.185 357.555 2100.465 ;
        RECT 357.985 2100.185 358.265 2100.465 ;
        RECT 358.695 2100.185 358.975 2100.465 ;
        RECT 359.405 2100.185 359.685 2100.465 ;
        RECT 360.115 2100.185 360.395 2100.465 ;
        RECT 360.825 2100.185 361.105 2100.465 ;
        RECT 361.535 2100.185 361.815 2100.465 ;
        RECT 362.245 2100.185 362.525 2100.465 ;
        RECT 362.955 2100.185 363.235 2100.465 ;
        RECT 363.665 2100.185 363.945 2100.465 ;
        RECT 364.375 2100.185 364.655 2100.465 ;
        RECT 365.085 2100.185 365.365 2100.465 ;
        RECT 365.795 2100.185 366.075 2100.465 ;
        RECT 366.505 2100.185 366.785 2100.465 ;
        RECT 357.275 2099.475 357.555 2099.755 ;
        RECT 357.985 2099.475 358.265 2099.755 ;
        RECT 358.695 2099.475 358.975 2099.755 ;
        RECT 359.405 2099.475 359.685 2099.755 ;
        RECT 360.115 2099.475 360.395 2099.755 ;
        RECT 360.825 2099.475 361.105 2099.755 ;
        RECT 361.535 2099.475 361.815 2099.755 ;
        RECT 362.245 2099.475 362.525 2099.755 ;
        RECT 362.955 2099.475 363.235 2099.755 ;
        RECT 363.665 2099.475 363.945 2099.755 ;
        RECT 364.375 2099.475 364.655 2099.755 ;
        RECT 365.085 2099.475 365.365 2099.755 ;
        RECT 365.795 2099.475 366.075 2099.755 ;
        RECT 366.505 2099.475 366.785 2099.755 ;
        RECT 357.275 2098.765 357.555 2099.045 ;
        RECT 357.985 2098.765 358.265 2099.045 ;
        RECT 358.695 2098.765 358.975 2099.045 ;
        RECT 359.405 2098.765 359.685 2099.045 ;
        RECT 360.115 2098.765 360.395 2099.045 ;
        RECT 360.825 2098.765 361.105 2099.045 ;
        RECT 361.535 2098.765 361.815 2099.045 ;
        RECT 362.245 2098.765 362.525 2099.045 ;
        RECT 362.955 2098.765 363.235 2099.045 ;
        RECT 363.665 2098.765 363.945 2099.045 ;
        RECT 364.375 2098.765 364.655 2099.045 ;
        RECT 365.085 2098.765 365.365 2099.045 ;
        RECT 365.795 2098.765 366.075 2099.045 ;
        RECT 366.505 2098.765 366.785 2099.045 ;
        RECT 357.275 2098.055 357.555 2098.335 ;
        RECT 357.985 2098.055 358.265 2098.335 ;
        RECT 358.695 2098.055 358.975 2098.335 ;
        RECT 359.405 2098.055 359.685 2098.335 ;
        RECT 360.115 2098.055 360.395 2098.335 ;
        RECT 360.825 2098.055 361.105 2098.335 ;
        RECT 361.535 2098.055 361.815 2098.335 ;
        RECT 362.245 2098.055 362.525 2098.335 ;
        RECT 362.955 2098.055 363.235 2098.335 ;
        RECT 363.665 2098.055 363.945 2098.335 ;
        RECT 364.375 2098.055 364.655 2098.335 ;
        RECT 365.085 2098.055 365.365 2098.335 ;
        RECT 365.795 2098.055 366.075 2098.335 ;
        RECT 366.505 2098.055 366.785 2098.335 ;
        RECT 357.275 2097.345 357.555 2097.625 ;
        RECT 357.985 2097.345 358.265 2097.625 ;
        RECT 358.695 2097.345 358.975 2097.625 ;
        RECT 359.405 2097.345 359.685 2097.625 ;
        RECT 360.115 2097.345 360.395 2097.625 ;
        RECT 360.825 2097.345 361.105 2097.625 ;
        RECT 361.535 2097.345 361.815 2097.625 ;
        RECT 362.245 2097.345 362.525 2097.625 ;
        RECT 362.955 2097.345 363.235 2097.625 ;
        RECT 363.665 2097.345 363.945 2097.625 ;
        RECT 364.375 2097.345 364.655 2097.625 ;
        RECT 365.085 2097.345 365.365 2097.625 ;
        RECT 365.795 2097.345 366.075 2097.625 ;
        RECT 366.505 2097.345 366.785 2097.625 ;
        RECT 357.275 2096.635 357.555 2096.915 ;
        RECT 357.985 2096.635 358.265 2096.915 ;
        RECT 358.695 2096.635 358.975 2096.915 ;
        RECT 359.405 2096.635 359.685 2096.915 ;
        RECT 360.115 2096.635 360.395 2096.915 ;
        RECT 360.825 2096.635 361.105 2096.915 ;
        RECT 361.535 2096.635 361.815 2096.915 ;
        RECT 362.245 2096.635 362.525 2096.915 ;
        RECT 362.955 2096.635 363.235 2096.915 ;
        RECT 363.665 2096.635 363.945 2096.915 ;
        RECT 364.375 2096.635 364.655 2096.915 ;
        RECT 365.085 2096.635 365.365 2096.915 ;
        RECT 365.795 2096.635 366.075 2096.915 ;
        RECT 366.505 2096.635 366.785 2096.915 ;
        RECT 357.275 2095.925 357.555 2096.205 ;
        RECT 357.985 2095.925 358.265 2096.205 ;
        RECT 358.695 2095.925 358.975 2096.205 ;
        RECT 359.405 2095.925 359.685 2096.205 ;
        RECT 360.115 2095.925 360.395 2096.205 ;
        RECT 360.825 2095.925 361.105 2096.205 ;
        RECT 361.535 2095.925 361.815 2096.205 ;
        RECT 362.245 2095.925 362.525 2096.205 ;
        RECT 362.955 2095.925 363.235 2096.205 ;
        RECT 363.665 2095.925 363.945 2096.205 ;
        RECT 364.375 2095.925 364.655 2096.205 ;
        RECT 365.085 2095.925 365.365 2096.205 ;
        RECT 365.795 2095.925 366.075 2096.205 ;
        RECT 366.505 2095.925 366.785 2096.205 ;
        RECT 357.275 2095.215 357.555 2095.495 ;
        RECT 357.985 2095.215 358.265 2095.495 ;
        RECT 358.695 2095.215 358.975 2095.495 ;
        RECT 359.405 2095.215 359.685 2095.495 ;
        RECT 360.115 2095.215 360.395 2095.495 ;
        RECT 360.825 2095.215 361.105 2095.495 ;
        RECT 361.535 2095.215 361.815 2095.495 ;
        RECT 362.245 2095.215 362.525 2095.495 ;
        RECT 362.955 2095.215 363.235 2095.495 ;
        RECT 363.665 2095.215 363.945 2095.495 ;
        RECT 364.375 2095.215 364.655 2095.495 ;
        RECT 365.085 2095.215 365.365 2095.495 ;
        RECT 365.795 2095.215 366.075 2095.495 ;
        RECT 366.505 2095.215 366.785 2095.495 ;
        RECT 357.275 2094.505 357.555 2094.785 ;
        RECT 357.985 2094.505 358.265 2094.785 ;
        RECT 358.695 2094.505 358.975 2094.785 ;
        RECT 359.405 2094.505 359.685 2094.785 ;
        RECT 360.115 2094.505 360.395 2094.785 ;
        RECT 360.825 2094.505 361.105 2094.785 ;
        RECT 361.535 2094.505 361.815 2094.785 ;
        RECT 362.245 2094.505 362.525 2094.785 ;
        RECT 362.955 2094.505 363.235 2094.785 ;
        RECT 363.665 2094.505 363.945 2094.785 ;
        RECT 364.375 2094.505 364.655 2094.785 ;
        RECT 365.085 2094.505 365.365 2094.785 ;
        RECT 365.795 2094.505 366.075 2094.785 ;
        RECT 366.505 2094.505 366.785 2094.785 ;
        RECT 357.275 2093.795 357.555 2094.075 ;
        RECT 357.985 2093.795 358.265 2094.075 ;
        RECT 358.695 2093.795 358.975 2094.075 ;
        RECT 359.405 2093.795 359.685 2094.075 ;
        RECT 360.115 2093.795 360.395 2094.075 ;
        RECT 360.825 2093.795 361.105 2094.075 ;
        RECT 361.535 2093.795 361.815 2094.075 ;
        RECT 362.245 2093.795 362.525 2094.075 ;
        RECT 362.955 2093.795 363.235 2094.075 ;
        RECT 363.665 2093.795 363.945 2094.075 ;
        RECT 364.375 2093.795 364.655 2094.075 ;
        RECT 365.085 2093.795 365.365 2094.075 ;
        RECT 365.795 2093.795 366.075 2094.075 ;
        RECT 366.505 2093.795 366.785 2094.075 ;
        RECT 357.275 2093.085 357.555 2093.365 ;
        RECT 357.985 2093.085 358.265 2093.365 ;
        RECT 358.695 2093.085 358.975 2093.365 ;
        RECT 359.405 2093.085 359.685 2093.365 ;
        RECT 360.115 2093.085 360.395 2093.365 ;
        RECT 360.825 2093.085 361.105 2093.365 ;
        RECT 361.535 2093.085 361.815 2093.365 ;
        RECT 362.245 2093.085 362.525 2093.365 ;
        RECT 362.955 2093.085 363.235 2093.365 ;
        RECT 363.665 2093.085 363.945 2093.365 ;
        RECT 364.375 2093.085 364.655 2093.365 ;
        RECT 365.085 2093.085 365.365 2093.365 ;
        RECT 365.795 2093.085 366.075 2093.365 ;
        RECT 366.505 2093.085 366.785 2093.365 ;
        RECT 357.275 2092.375 357.555 2092.655 ;
        RECT 357.985 2092.375 358.265 2092.655 ;
        RECT 358.695 2092.375 358.975 2092.655 ;
        RECT 359.405 2092.375 359.685 2092.655 ;
        RECT 360.115 2092.375 360.395 2092.655 ;
        RECT 360.825 2092.375 361.105 2092.655 ;
        RECT 361.535 2092.375 361.815 2092.655 ;
        RECT 362.245 2092.375 362.525 2092.655 ;
        RECT 362.955 2092.375 363.235 2092.655 ;
        RECT 363.665 2092.375 363.945 2092.655 ;
        RECT 364.375 2092.375 364.655 2092.655 ;
        RECT 365.085 2092.375 365.365 2092.655 ;
        RECT 365.795 2092.375 366.075 2092.655 ;
        RECT 366.505 2092.375 366.785 2092.655 ;
        RECT 357.275 2091.665 357.555 2091.945 ;
        RECT 357.985 2091.665 358.265 2091.945 ;
        RECT 358.695 2091.665 358.975 2091.945 ;
        RECT 359.405 2091.665 359.685 2091.945 ;
        RECT 360.115 2091.665 360.395 2091.945 ;
        RECT 360.825 2091.665 361.105 2091.945 ;
        RECT 361.535 2091.665 361.815 2091.945 ;
        RECT 362.245 2091.665 362.525 2091.945 ;
        RECT 362.955 2091.665 363.235 2091.945 ;
        RECT 363.665 2091.665 363.945 2091.945 ;
        RECT 364.375 2091.665 364.655 2091.945 ;
        RECT 365.085 2091.665 365.365 2091.945 ;
        RECT 365.795 2091.665 366.075 2091.945 ;
        RECT 366.505 2091.665 366.785 2091.945 ;
        RECT 357.275 2090.955 357.555 2091.235 ;
        RECT 357.985 2090.955 358.265 2091.235 ;
        RECT 358.695 2090.955 358.975 2091.235 ;
        RECT 359.405 2090.955 359.685 2091.235 ;
        RECT 360.115 2090.955 360.395 2091.235 ;
        RECT 360.825 2090.955 361.105 2091.235 ;
        RECT 361.535 2090.955 361.815 2091.235 ;
        RECT 362.245 2090.955 362.525 2091.235 ;
        RECT 362.955 2090.955 363.235 2091.235 ;
        RECT 363.665 2090.955 363.945 2091.235 ;
        RECT 364.375 2090.955 364.655 2091.235 ;
        RECT 365.085 2090.955 365.365 2091.235 ;
        RECT 365.795 2090.955 366.075 2091.235 ;
        RECT 366.505 2090.955 366.785 2091.235 ;
        RECT 357.275 2088.335 357.555 2088.615 ;
        RECT 357.985 2088.335 358.265 2088.615 ;
        RECT 358.695 2088.335 358.975 2088.615 ;
        RECT 359.405 2088.335 359.685 2088.615 ;
        RECT 360.115 2088.335 360.395 2088.615 ;
        RECT 360.825 2088.335 361.105 2088.615 ;
        RECT 361.535 2088.335 361.815 2088.615 ;
        RECT 362.245 2088.335 362.525 2088.615 ;
        RECT 362.955 2088.335 363.235 2088.615 ;
        RECT 363.665 2088.335 363.945 2088.615 ;
        RECT 364.375 2088.335 364.655 2088.615 ;
        RECT 365.085 2088.335 365.365 2088.615 ;
        RECT 365.795 2088.335 366.075 2088.615 ;
        RECT 366.505 2088.335 366.785 2088.615 ;
        RECT 357.275 2087.625 357.555 2087.905 ;
        RECT 357.985 2087.625 358.265 2087.905 ;
        RECT 358.695 2087.625 358.975 2087.905 ;
        RECT 359.405 2087.625 359.685 2087.905 ;
        RECT 360.115 2087.625 360.395 2087.905 ;
        RECT 360.825 2087.625 361.105 2087.905 ;
        RECT 361.535 2087.625 361.815 2087.905 ;
        RECT 362.245 2087.625 362.525 2087.905 ;
        RECT 362.955 2087.625 363.235 2087.905 ;
        RECT 363.665 2087.625 363.945 2087.905 ;
        RECT 364.375 2087.625 364.655 2087.905 ;
        RECT 365.085 2087.625 365.365 2087.905 ;
        RECT 365.795 2087.625 366.075 2087.905 ;
        RECT 366.505 2087.625 366.785 2087.905 ;
        RECT 357.275 2086.915 357.555 2087.195 ;
        RECT 357.985 2086.915 358.265 2087.195 ;
        RECT 358.695 2086.915 358.975 2087.195 ;
        RECT 359.405 2086.915 359.685 2087.195 ;
        RECT 360.115 2086.915 360.395 2087.195 ;
        RECT 360.825 2086.915 361.105 2087.195 ;
        RECT 361.535 2086.915 361.815 2087.195 ;
        RECT 362.245 2086.915 362.525 2087.195 ;
        RECT 362.955 2086.915 363.235 2087.195 ;
        RECT 363.665 2086.915 363.945 2087.195 ;
        RECT 364.375 2086.915 364.655 2087.195 ;
        RECT 365.085 2086.915 365.365 2087.195 ;
        RECT 365.795 2086.915 366.075 2087.195 ;
        RECT 366.505 2086.915 366.785 2087.195 ;
        RECT 357.275 2086.205 357.555 2086.485 ;
        RECT 357.985 2086.205 358.265 2086.485 ;
        RECT 358.695 2086.205 358.975 2086.485 ;
        RECT 359.405 2086.205 359.685 2086.485 ;
        RECT 360.115 2086.205 360.395 2086.485 ;
        RECT 360.825 2086.205 361.105 2086.485 ;
        RECT 361.535 2086.205 361.815 2086.485 ;
        RECT 362.245 2086.205 362.525 2086.485 ;
        RECT 362.955 2086.205 363.235 2086.485 ;
        RECT 363.665 2086.205 363.945 2086.485 ;
        RECT 364.375 2086.205 364.655 2086.485 ;
        RECT 365.085 2086.205 365.365 2086.485 ;
        RECT 365.795 2086.205 366.075 2086.485 ;
        RECT 366.505 2086.205 366.785 2086.485 ;
        RECT 357.275 2085.495 357.555 2085.775 ;
        RECT 357.985 2085.495 358.265 2085.775 ;
        RECT 358.695 2085.495 358.975 2085.775 ;
        RECT 359.405 2085.495 359.685 2085.775 ;
        RECT 360.115 2085.495 360.395 2085.775 ;
        RECT 360.825 2085.495 361.105 2085.775 ;
        RECT 361.535 2085.495 361.815 2085.775 ;
        RECT 362.245 2085.495 362.525 2085.775 ;
        RECT 362.955 2085.495 363.235 2085.775 ;
        RECT 363.665 2085.495 363.945 2085.775 ;
        RECT 364.375 2085.495 364.655 2085.775 ;
        RECT 365.085 2085.495 365.365 2085.775 ;
        RECT 365.795 2085.495 366.075 2085.775 ;
        RECT 366.505 2085.495 366.785 2085.775 ;
        RECT 357.275 2084.785 357.555 2085.065 ;
        RECT 357.985 2084.785 358.265 2085.065 ;
        RECT 358.695 2084.785 358.975 2085.065 ;
        RECT 359.405 2084.785 359.685 2085.065 ;
        RECT 360.115 2084.785 360.395 2085.065 ;
        RECT 360.825 2084.785 361.105 2085.065 ;
        RECT 361.535 2084.785 361.815 2085.065 ;
        RECT 362.245 2084.785 362.525 2085.065 ;
        RECT 362.955 2084.785 363.235 2085.065 ;
        RECT 363.665 2084.785 363.945 2085.065 ;
        RECT 364.375 2084.785 364.655 2085.065 ;
        RECT 365.085 2084.785 365.365 2085.065 ;
        RECT 365.795 2084.785 366.075 2085.065 ;
        RECT 366.505 2084.785 366.785 2085.065 ;
        RECT 357.275 2084.075 357.555 2084.355 ;
        RECT 357.985 2084.075 358.265 2084.355 ;
        RECT 358.695 2084.075 358.975 2084.355 ;
        RECT 359.405 2084.075 359.685 2084.355 ;
        RECT 360.115 2084.075 360.395 2084.355 ;
        RECT 360.825 2084.075 361.105 2084.355 ;
        RECT 361.535 2084.075 361.815 2084.355 ;
        RECT 362.245 2084.075 362.525 2084.355 ;
        RECT 362.955 2084.075 363.235 2084.355 ;
        RECT 363.665 2084.075 363.945 2084.355 ;
        RECT 364.375 2084.075 364.655 2084.355 ;
        RECT 365.085 2084.075 365.365 2084.355 ;
        RECT 365.795 2084.075 366.075 2084.355 ;
        RECT 366.505 2084.075 366.785 2084.355 ;
        RECT 357.275 2083.365 357.555 2083.645 ;
        RECT 357.985 2083.365 358.265 2083.645 ;
        RECT 358.695 2083.365 358.975 2083.645 ;
        RECT 359.405 2083.365 359.685 2083.645 ;
        RECT 360.115 2083.365 360.395 2083.645 ;
        RECT 360.825 2083.365 361.105 2083.645 ;
        RECT 361.535 2083.365 361.815 2083.645 ;
        RECT 362.245 2083.365 362.525 2083.645 ;
        RECT 362.955 2083.365 363.235 2083.645 ;
        RECT 363.665 2083.365 363.945 2083.645 ;
        RECT 364.375 2083.365 364.655 2083.645 ;
        RECT 365.085 2083.365 365.365 2083.645 ;
        RECT 365.795 2083.365 366.075 2083.645 ;
        RECT 366.505 2083.365 366.785 2083.645 ;
        RECT 357.275 2082.655 357.555 2082.935 ;
        RECT 357.985 2082.655 358.265 2082.935 ;
        RECT 358.695 2082.655 358.975 2082.935 ;
        RECT 359.405 2082.655 359.685 2082.935 ;
        RECT 360.115 2082.655 360.395 2082.935 ;
        RECT 360.825 2082.655 361.105 2082.935 ;
        RECT 361.535 2082.655 361.815 2082.935 ;
        RECT 362.245 2082.655 362.525 2082.935 ;
        RECT 362.955 2082.655 363.235 2082.935 ;
        RECT 363.665 2082.655 363.945 2082.935 ;
        RECT 364.375 2082.655 364.655 2082.935 ;
        RECT 365.085 2082.655 365.365 2082.935 ;
        RECT 365.795 2082.655 366.075 2082.935 ;
        RECT 366.505 2082.655 366.785 2082.935 ;
        RECT 357.275 2081.945 357.555 2082.225 ;
        RECT 357.985 2081.945 358.265 2082.225 ;
        RECT 358.695 2081.945 358.975 2082.225 ;
        RECT 359.405 2081.945 359.685 2082.225 ;
        RECT 360.115 2081.945 360.395 2082.225 ;
        RECT 360.825 2081.945 361.105 2082.225 ;
        RECT 361.535 2081.945 361.815 2082.225 ;
        RECT 362.245 2081.945 362.525 2082.225 ;
        RECT 362.955 2081.945 363.235 2082.225 ;
        RECT 363.665 2081.945 363.945 2082.225 ;
        RECT 364.375 2081.945 364.655 2082.225 ;
        RECT 365.085 2081.945 365.365 2082.225 ;
        RECT 365.795 2081.945 366.075 2082.225 ;
        RECT 366.505 2081.945 366.785 2082.225 ;
        RECT 357.275 2081.235 357.555 2081.515 ;
        RECT 357.985 2081.235 358.265 2081.515 ;
        RECT 358.695 2081.235 358.975 2081.515 ;
        RECT 359.405 2081.235 359.685 2081.515 ;
        RECT 360.115 2081.235 360.395 2081.515 ;
        RECT 360.825 2081.235 361.105 2081.515 ;
        RECT 361.535 2081.235 361.815 2081.515 ;
        RECT 362.245 2081.235 362.525 2081.515 ;
        RECT 362.955 2081.235 363.235 2081.515 ;
        RECT 363.665 2081.235 363.945 2081.515 ;
        RECT 364.375 2081.235 364.655 2081.515 ;
        RECT 365.085 2081.235 365.365 2081.515 ;
        RECT 365.795 2081.235 366.075 2081.515 ;
        RECT 366.505 2081.235 366.785 2081.515 ;
        RECT 357.275 2080.525 357.555 2080.805 ;
        RECT 357.985 2080.525 358.265 2080.805 ;
        RECT 358.695 2080.525 358.975 2080.805 ;
        RECT 359.405 2080.525 359.685 2080.805 ;
        RECT 360.115 2080.525 360.395 2080.805 ;
        RECT 360.825 2080.525 361.105 2080.805 ;
        RECT 361.535 2080.525 361.815 2080.805 ;
        RECT 362.245 2080.525 362.525 2080.805 ;
        RECT 362.955 2080.525 363.235 2080.805 ;
        RECT 363.665 2080.525 363.945 2080.805 ;
        RECT 364.375 2080.525 364.655 2080.805 ;
        RECT 365.085 2080.525 365.365 2080.805 ;
        RECT 365.795 2080.525 366.075 2080.805 ;
        RECT 366.505 2080.525 366.785 2080.805 ;
        RECT 357.275 2079.815 357.555 2080.095 ;
        RECT 357.985 2079.815 358.265 2080.095 ;
        RECT 358.695 2079.815 358.975 2080.095 ;
        RECT 359.405 2079.815 359.685 2080.095 ;
        RECT 360.115 2079.815 360.395 2080.095 ;
        RECT 360.825 2079.815 361.105 2080.095 ;
        RECT 361.535 2079.815 361.815 2080.095 ;
        RECT 362.245 2079.815 362.525 2080.095 ;
        RECT 362.955 2079.815 363.235 2080.095 ;
        RECT 363.665 2079.815 363.945 2080.095 ;
        RECT 364.375 2079.815 364.655 2080.095 ;
        RECT 365.085 2079.815 365.365 2080.095 ;
        RECT 365.795 2079.815 366.075 2080.095 ;
        RECT 366.505 2079.815 366.785 2080.095 ;
        RECT 357.275 2079.105 357.555 2079.385 ;
        RECT 357.985 2079.105 358.265 2079.385 ;
        RECT 358.695 2079.105 358.975 2079.385 ;
        RECT 359.405 2079.105 359.685 2079.385 ;
        RECT 360.115 2079.105 360.395 2079.385 ;
        RECT 360.825 2079.105 361.105 2079.385 ;
        RECT 361.535 2079.105 361.815 2079.385 ;
        RECT 362.245 2079.105 362.525 2079.385 ;
        RECT 362.955 2079.105 363.235 2079.385 ;
        RECT 363.665 2079.105 363.945 2079.385 ;
        RECT 364.375 2079.105 364.655 2079.385 ;
        RECT 365.085 2079.105 365.365 2079.385 ;
        RECT 365.795 2079.105 366.075 2079.385 ;
        RECT 366.505 2079.105 366.785 2079.385 ;
        RECT 357.330 2075.190 357.610 2075.470 ;
        RECT 358.040 2075.190 358.320 2075.470 ;
        RECT 358.750 2075.190 359.030 2075.470 ;
        RECT 359.460 2075.190 359.740 2075.470 ;
        RECT 360.170 2075.190 360.450 2075.470 ;
        RECT 360.880 2075.190 361.160 2075.470 ;
        RECT 361.590 2075.190 361.870 2075.470 ;
        RECT 362.300 2075.190 362.580 2075.470 ;
        RECT 363.010 2075.190 363.290 2075.470 ;
        RECT 363.720 2075.190 364.000 2075.470 ;
        RECT 364.430 2075.190 364.710 2075.470 ;
        RECT 365.140 2075.190 365.420 2075.470 ;
        RECT 365.850 2075.190 366.130 2075.470 ;
        RECT 366.560 2075.190 366.840 2075.470 ;
        RECT 357.330 2074.480 357.610 2074.760 ;
        RECT 358.040 2074.480 358.320 2074.760 ;
        RECT 358.750 2074.480 359.030 2074.760 ;
        RECT 359.460 2074.480 359.740 2074.760 ;
        RECT 360.170 2074.480 360.450 2074.760 ;
        RECT 360.880 2074.480 361.160 2074.760 ;
        RECT 361.590 2074.480 361.870 2074.760 ;
        RECT 362.300 2074.480 362.580 2074.760 ;
        RECT 363.010 2074.480 363.290 2074.760 ;
        RECT 363.720 2074.480 364.000 2074.760 ;
        RECT 364.430 2074.480 364.710 2074.760 ;
        RECT 365.140 2074.480 365.420 2074.760 ;
        RECT 365.850 2074.480 366.130 2074.760 ;
        RECT 366.560 2074.480 366.840 2074.760 ;
        RECT 357.330 2073.770 357.610 2074.050 ;
        RECT 358.040 2073.770 358.320 2074.050 ;
        RECT 358.750 2073.770 359.030 2074.050 ;
        RECT 359.460 2073.770 359.740 2074.050 ;
        RECT 360.170 2073.770 360.450 2074.050 ;
        RECT 360.880 2073.770 361.160 2074.050 ;
        RECT 361.590 2073.770 361.870 2074.050 ;
        RECT 362.300 2073.770 362.580 2074.050 ;
        RECT 363.010 2073.770 363.290 2074.050 ;
        RECT 363.720 2073.770 364.000 2074.050 ;
        RECT 364.430 2073.770 364.710 2074.050 ;
        RECT 365.140 2073.770 365.420 2074.050 ;
        RECT 365.850 2073.770 366.130 2074.050 ;
        RECT 366.560 2073.770 366.840 2074.050 ;
        RECT 357.330 2073.060 357.610 2073.340 ;
        RECT 358.040 2073.060 358.320 2073.340 ;
        RECT 358.750 2073.060 359.030 2073.340 ;
        RECT 359.460 2073.060 359.740 2073.340 ;
        RECT 360.170 2073.060 360.450 2073.340 ;
        RECT 360.880 2073.060 361.160 2073.340 ;
        RECT 361.590 2073.060 361.870 2073.340 ;
        RECT 362.300 2073.060 362.580 2073.340 ;
        RECT 363.010 2073.060 363.290 2073.340 ;
        RECT 363.720 2073.060 364.000 2073.340 ;
        RECT 364.430 2073.060 364.710 2073.340 ;
        RECT 365.140 2073.060 365.420 2073.340 ;
        RECT 365.850 2073.060 366.130 2073.340 ;
        RECT 366.560 2073.060 366.840 2073.340 ;
        RECT 357.330 2072.350 357.610 2072.630 ;
        RECT 358.040 2072.350 358.320 2072.630 ;
        RECT 358.750 2072.350 359.030 2072.630 ;
        RECT 359.460 2072.350 359.740 2072.630 ;
        RECT 360.170 2072.350 360.450 2072.630 ;
        RECT 360.880 2072.350 361.160 2072.630 ;
        RECT 361.590 2072.350 361.870 2072.630 ;
        RECT 362.300 2072.350 362.580 2072.630 ;
        RECT 363.010 2072.350 363.290 2072.630 ;
        RECT 363.720 2072.350 364.000 2072.630 ;
        RECT 364.430 2072.350 364.710 2072.630 ;
        RECT 365.140 2072.350 365.420 2072.630 ;
        RECT 365.850 2072.350 366.130 2072.630 ;
        RECT 366.560 2072.350 366.840 2072.630 ;
        RECT 357.330 2071.640 357.610 2071.920 ;
        RECT 358.040 2071.640 358.320 2071.920 ;
        RECT 358.750 2071.640 359.030 2071.920 ;
        RECT 359.460 2071.640 359.740 2071.920 ;
        RECT 360.170 2071.640 360.450 2071.920 ;
        RECT 360.880 2071.640 361.160 2071.920 ;
        RECT 361.590 2071.640 361.870 2071.920 ;
        RECT 362.300 2071.640 362.580 2071.920 ;
        RECT 363.010 2071.640 363.290 2071.920 ;
        RECT 363.720 2071.640 364.000 2071.920 ;
        RECT 364.430 2071.640 364.710 2071.920 ;
        RECT 365.140 2071.640 365.420 2071.920 ;
        RECT 365.850 2071.640 366.130 2071.920 ;
        RECT 366.560 2071.640 366.840 2071.920 ;
        RECT 357.330 2070.930 357.610 2071.210 ;
        RECT 358.040 2070.930 358.320 2071.210 ;
        RECT 358.750 2070.930 359.030 2071.210 ;
        RECT 359.460 2070.930 359.740 2071.210 ;
        RECT 360.170 2070.930 360.450 2071.210 ;
        RECT 360.880 2070.930 361.160 2071.210 ;
        RECT 361.590 2070.930 361.870 2071.210 ;
        RECT 362.300 2070.930 362.580 2071.210 ;
        RECT 363.010 2070.930 363.290 2071.210 ;
        RECT 363.720 2070.930 364.000 2071.210 ;
        RECT 364.430 2070.930 364.710 2071.210 ;
        RECT 365.140 2070.930 365.420 2071.210 ;
        RECT 365.850 2070.930 366.130 2071.210 ;
        RECT 366.560 2070.930 366.840 2071.210 ;
        RECT 357.330 2070.220 357.610 2070.500 ;
        RECT 358.040 2070.220 358.320 2070.500 ;
        RECT 358.750 2070.220 359.030 2070.500 ;
        RECT 359.460 2070.220 359.740 2070.500 ;
        RECT 360.170 2070.220 360.450 2070.500 ;
        RECT 360.880 2070.220 361.160 2070.500 ;
        RECT 361.590 2070.220 361.870 2070.500 ;
        RECT 362.300 2070.220 362.580 2070.500 ;
        RECT 363.010 2070.220 363.290 2070.500 ;
        RECT 363.720 2070.220 364.000 2070.500 ;
        RECT 364.430 2070.220 364.710 2070.500 ;
        RECT 365.140 2070.220 365.420 2070.500 ;
        RECT 365.850 2070.220 366.130 2070.500 ;
        RECT 366.560 2070.220 366.840 2070.500 ;
        RECT 357.330 2069.510 357.610 2069.790 ;
        RECT 358.040 2069.510 358.320 2069.790 ;
        RECT 358.750 2069.510 359.030 2069.790 ;
        RECT 359.460 2069.510 359.740 2069.790 ;
        RECT 360.170 2069.510 360.450 2069.790 ;
        RECT 360.880 2069.510 361.160 2069.790 ;
        RECT 361.590 2069.510 361.870 2069.790 ;
        RECT 362.300 2069.510 362.580 2069.790 ;
        RECT 363.010 2069.510 363.290 2069.790 ;
        RECT 363.720 2069.510 364.000 2069.790 ;
        RECT 364.430 2069.510 364.710 2069.790 ;
        RECT 365.140 2069.510 365.420 2069.790 ;
        RECT 365.850 2069.510 366.130 2069.790 ;
        RECT 366.560 2069.510 366.840 2069.790 ;
        RECT 357.330 2068.800 357.610 2069.080 ;
        RECT 358.040 2068.800 358.320 2069.080 ;
        RECT 358.750 2068.800 359.030 2069.080 ;
        RECT 359.460 2068.800 359.740 2069.080 ;
        RECT 360.170 2068.800 360.450 2069.080 ;
        RECT 360.880 2068.800 361.160 2069.080 ;
        RECT 361.590 2068.800 361.870 2069.080 ;
        RECT 362.300 2068.800 362.580 2069.080 ;
        RECT 363.010 2068.800 363.290 2069.080 ;
        RECT 363.720 2068.800 364.000 2069.080 ;
        RECT 364.430 2068.800 364.710 2069.080 ;
        RECT 365.140 2068.800 365.420 2069.080 ;
        RECT 365.850 2068.800 366.130 2069.080 ;
        RECT 366.560 2068.800 366.840 2069.080 ;
        RECT 357.330 2068.090 357.610 2068.370 ;
        RECT 358.040 2068.090 358.320 2068.370 ;
        RECT 358.750 2068.090 359.030 2068.370 ;
        RECT 359.460 2068.090 359.740 2068.370 ;
        RECT 360.170 2068.090 360.450 2068.370 ;
        RECT 360.880 2068.090 361.160 2068.370 ;
        RECT 361.590 2068.090 361.870 2068.370 ;
        RECT 362.300 2068.090 362.580 2068.370 ;
        RECT 363.010 2068.090 363.290 2068.370 ;
        RECT 363.720 2068.090 364.000 2068.370 ;
        RECT 364.430 2068.090 364.710 2068.370 ;
        RECT 365.140 2068.090 365.420 2068.370 ;
        RECT 365.850 2068.090 366.130 2068.370 ;
        RECT 366.560 2068.090 366.840 2068.370 ;
        RECT 357.330 2067.380 357.610 2067.660 ;
        RECT 358.040 2067.380 358.320 2067.660 ;
        RECT 358.750 2067.380 359.030 2067.660 ;
        RECT 359.460 2067.380 359.740 2067.660 ;
        RECT 360.170 2067.380 360.450 2067.660 ;
        RECT 360.880 2067.380 361.160 2067.660 ;
        RECT 361.590 2067.380 361.870 2067.660 ;
        RECT 362.300 2067.380 362.580 2067.660 ;
        RECT 363.010 2067.380 363.290 2067.660 ;
        RECT 363.720 2067.380 364.000 2067.660 ;
        RECT 364.430 2067.380 364.710 2067.660 ;
        RECT 365.140 2067.380 365.420 2067.660 ;
        RECT 365.850 2067.380 366.130 2067.660 ;
        RECT 366.560 2067.380 366.840 2067.660 ;
        RECT 357.330 2066.670 357.610 2066.950 ;
        RECT 358.040 2066.670 358.320 2066.950 ;
        RECT 358.750 2066.670 359.030 2066.950 ;
        RECT 359.460 2066.670 359.740 2066.950 ;
        RECT 360.170 2066.670 360.450 2066.950 ;
        RECT 360.880 2066.670 361.160 2066.950 ;
        RECT 361.590 2066.670 361.870 2066.950 ;
        RECT 362.300 2066.670 362.580 2066.950 ;
        RECT 363.010 2066.670 363.290 2066.950 ;
        RECT 363.720 2066.670 364.000 2066.950 ;
        RECT 364.430 2066.670 364.710 2066.950 ;
        RECT 365.140 2066.670 365.420 2066.950 ;
        RECT 365.850 2066.670 366.130 2066.950 ;
        RECT 366.560 2066.670 366.840 2066.950 ;
        RECT 3512.200 2023.050 3512.480 2023.330 ;
        RECT 3512.910 2023.050 3513.190 2023.330 ;
        RECT 3513.620 2023.050 3513.900 2023.330 ;
        RECT 3514.330 2023.050 3514.610 2023.330 ;
        RECT 3515.040 2023.050 3515.320 2023.330 ;
        RECT 3515.750 2023.050 3516.030 2023.330 ;
        RECT 3516.460 2023.050 3516.740 2023.330 ;
        RECT 3517.170 2023.050 3517.450 2023.330 ;
        RECT 3517.880 2023.050 3518.160 2023.330 ;
        RECT 3518.590 2023.050 3518.870 2023.330 ;
        RECT 3519.300 2023.050 3519.580 2023.330 ;
        RECT 3520.010 2023.050 3520.290 2023.330 ;
        RECT 3520.720 2023.050 3521.000 2023.330 ;
        RECT 3521.430 2023.050 3521.710 2023.330 ;
        RECT 3512.200 2022.340 3512.480 2022.620 ;
        RECT 3512.910 2022.340 3513.190 2022.620 ;
        RECT 3513.620 2022.340 3513.900 2022.620 ;
        RECT 3514.330 2022.340 3514.610 2022.620 ;
        RECT 3515.040 2022.340 3515.320 2022.620 ;
        RECT 3515.750 2022.340 3516.030 2022.620 ;
        RECT 3516.460 2022.340 3516.740 2022.620 ;
        RECT 3517.170 2022.340 3517.450 2022.620 ;
        RECT 3517.880 2022.340 3518.160 2022.620 ;
        RECT 3518.590 2022.340 3518.870 2022.620 ;
        RECT 3519.300 2022.340 3519.580 2022.620 ;
        RECT 3520.010 2022.340 3520.290 2022.620 ;
        RECT 3520.720 2022.340 3521.000 2022.620 ;
        RECT 3521.430 2022.340 3521.710 2022.620 ;
        RECT 3512.200 2021.630 3512.480 2021.910 ;
        RECT 3512.910 2021.630 3513.190 2021.910 ;
        RECT 3513.620 2021.630 3513.900 2021.910 ;
        RECT 3514.330 2021.630 3514.610 2021.910 ;
        RECT 3515.040 2021.630 3515.320 2021.910 ;
        RECT 3515.750 2021.630 3516.030 2021.910 ;
        RECT 3516.460 2021.630 3516.740 2021.910 ;
        RECT 3517.170 2021.630 3517.450 2021.910 ;
        RECT 3517.880 2021.630 3518.160 2021.910 ;
        RECT 3518.590 2021.630 3518.870 2021.910 ;
        RECT 3519.300 2021.630 3519.580 2021.910 ;
        RECT 3520.010 2021.630 3520.290 2021.910 ;
        RECT 3520.720 2021.630 3521.000 2021.910 ;
        RECT 3521.430 2021.630 3521.710 2021.910 ;
        RECT 3512.200 2020.920 3512.480 2021.200 ;
        RECT 3512.910 2020.920 3513.190 2021.200 ;
        RECT 3513.620 2020.920 3513.900 2021.200 ;
        RECT 3514.330 2020.920 3514.610 2021.200 ;
        RECT 3515.040 2020.920 3515.320 2021.200 ;
        RECT 3515.750 2020.920 3516.030 2021.200 ;
        RECT 3516.460 2020.920 3516.740 2021.200 ;
        RECT 3517.170 2020.920 3517.450 2021.200 ;
        RECT 3517.880 2020.920 3518.160 2021.200 ;
        RECT 3518.590 2020.920 3518.870 2021.200 ;
        RECT 3519.300 2020.920 3519.580 2021.200 ;
        RECT 3520.010 2020.920 3520.290 2021.200 ;
        RECT 3520.720 2020.920 3521.000 2021.200 ;
        RECT 3521.430 2020.920 3521.710 2021.200 ;
        RECT 3512.200 2020.210 3512.480 2020.490 ;
        RECT 3512.910 2020.210 3513.190 2020.490 ;
        RECT 3513.620 2020.210 3513.900 2020.490 ;
        RECT 3514.330 2020.210 3514.610 2020.490 ;
        RECT 3515.040 2020.210 3515.320 2020.490 ;
        RECT 3515.750 2020.210 3516.030 2020.490 ;
        RECT 3516.460 2020.210 3516.740 2020.490 ;
        RECT 3517.170 2020.210 3517.450 2020.490 ;
        RECT 3517.880 2020.210 3518.160 2020.490 ;
        RECT 3518.590 2020.210 3518.870 2020.490 ;
        RECT 3519.300 2020.210 3519.580 2020.490 ;
        RECT 3520.010 2020.210 3520.290 2020.490 ;
        RECT 3520.720 2020.210 3521.000 2020.490 ;
        RECT 3521.430 2020.210 3521.710 2020.490 ;
        RECT 3512.200 2019.500 3512.480 2019.780 ;
        RECT 3512.910 2019.500 3513.190 2019.780 ;
        RECT 3513.620 2019.500 3513.900 2019.780 ;
        RECT 3514.330 2019.500 3514.610 2019.780 ;
        RECT 3515.040 2019.500 3515.320 2019.780 ;
        RECT 3515.750 2019.500 3516.030 2019.780 ;
        RECT 3516.460 2019.500 3516.740 2019.780 ;
        RECT 3517.170 2019.500 3517.450 2019.780 ;
        RECT 3517.880 2019.500 3518.160 2019.780 ;
        RECT 3518.590 2019.500 3518.870 2019.780 ;
        RECT 3519.300 2019.500 3519.580 2019.780 ;
        RECT 3520.010 2019.500 3520.290 2019.780 ;
        RECT 3520.720 2019.500 3521.000 2019.780 ;
        RECT 3521.430 2019.500 3521.710 2019.780 ;
        RECT 3512.200 2018.790 3512.480 2019.070 ;
        RECT 3512.910 2018.790 3513.190 2019.070 ;
        RECT 3513.620 2018.790 3513.900 2019.070 ;
        RECT 3514.330 2018.790 3514.610 2019.070 ;
        RECT 3515.040 2018.790 3515.320 2019.070 ;
        RECT 3515.750 2018.790 3516.030 2019.070 ;
        RECT 3516.460 2018.790 3516.740 2019.070 ;
        RECT 3517.170 2018.790 3517.450 2019.070 ;
        RECT 3517.880 2018.790 3518.160 2019.070 ;
        RECT 3518.590 2018.790 3518.870 2019.070 ;
        RECT 3519.300 2018.790 3519.580 2019.070 ;
        RECT 3520.010 2018.790 3520.290 2019.070 ;
        RECT 3520.720 2018.790 3521.000 2019.070 ;
        RECT 3521.430 2018.790 3521.710 2019.070 ;
        RECT 3512.200 2018.080 3512.480 2018.360 ;
        RECT 3512.910 2018.080 3513.190 2018.360 ;
        RECT 3513.620 2018.080 3513.900 2018.360 ;
        RECT 3514.330 2018.080 3514.610 2018.360 ;
        RECT 3515.040 2018.080 3515.320 2018.360 ;
        RECT 3515.750 2018.080 3516.030 2018.360 ;
        RECT 3516.460 2018.080 3516.740 2018.360 ;
        RECT 3517.170 2018.080 3517.450 2018.360 ;
        RECT 3517.880 2018.080 3518.160 2018.360 ;
        RECT 3518.590 2018.080 3518.870 2018.360 ;
        RECT 3519.300 2018.080 3519.580 2018.360 ;
        RECT 3520.010 2018.080 3520.290 2018.360 ;
        RECT 3520.720 2018.080 3521.000 2018.360 ;
        RECT 3521.430 2018.080 3521.710 2018.360 ;
        RECT 3512.200 2017.370 3512.480 2017.650 ;
        RECT 3512.910 2017.370 3513.190 2017.650 ;
        RECT 3513.620 2017.370 3513.900 2017.650 ;
        RECT 3514.330 2017.370 3514.610 2017.650 ;
        RECT 3515.040 2017.370 3515.320 2017.650 ;
        RECT 3515.750 2017.370 3516.030 2017.650 ;
        RECT 3516.460 2017.370 3516.740 2017.650 ;
        RECT 3517.170 2017.370 3517.450 2017.650 ;
        RECT 3517.880 2017.370 3518.160 2017.650 ;
        RECT 3518.590 2017.370 3518.870 2017.650 ;
        RECT 3519.300 2017.370 3519.580 2017.650 ;
        RECT 3520.010 2017.370 3520.290 2017.650 ;
        RECT 3520.720 2017.370 3521.000 2017.650 ;
        RECT 3521.430 2017.370 3521.710 2017.650 ;
        RECT 3512.200 2016.660 3512.480 2016.940 ;
        RECT 3512.910 2016.660 3513.190 2016.940 ;
        RECT 3513.620 2016.660 3513.900 2016.940 ;
        RECT 3514.330 2016.660 3514.610 2016.940 ;
        RECT 3515.040 2016.660 3515.320 2016.940 ;
        RECT 3515.750 2016.660 3516.030 2016.940 ;
        RECT 3516.460 2016.660 3516.740 2016.940 ;
        RECT 3517.170 2016.660 3517.450 2016.940 ;
        RECT 3517.880 2016.660 3518.160 2016.940 ;
        RECT 3518.590 2016.660 3518.870 2016.940 ;
        RECT 3519.300 2016.660 3519.580 2016.940 ;
        RECT 3520.010 2016.660 3520.290 2016.940 ;
        RECT 3520.720 2016.660 3521.000 2016.940 ;
        RECT 3521.430 2016.660 3521.710 2016.940 ;
        RECT 3512.200 2015.950 3512.480 2016.230 ;
        RECT 3512.910 2015.950 3513.190 2016.230 ;
        RECT 3513.620 2015.950 3513.900 2016.230 ;
        RECT 3514.330 2015.950 3514.610 2016.230 ;
        RECT 3515.040 2015.950 3515.320 2016.230 ;
        RECT 3515.750 2015.950 3516.030 2016.230 ;
        RECT 3516.460 2015.950 3516.740 2016.230 ;
        RECT 3517.170 2015.950 3517.450 2016.230 ;
        RECT 3517.880 2015.950 3518.160 2016.230 ;
        RECT 3518.590 2015.950 3518.870 2016.230 ;
        RECT 3519.300 2015.950 3519.580 2016.230 ;
        RECT 3520.010 2015.950 3520.290 2016.230 ;
        RECT 3520.720 2015.950 3521.000 2016.230 ;
        RECT 3521.430 2015.950 3521.710 2016.230 ;
        RECT 3512.200 2015.240 3512.480 2015.520 ;
        RECT 3512.910 2015.240 3513.190 2015.520 ;
        RECT 3513.620 2015.240 3513.900 2015.520 ;
        RECT 3514.330 2015.240 3514.610 2015.520 ;
        RECT 3515.040 2015.240 3515.320 2015.520 ;
        RECT 3515.750 2015.240 3516.030 2015.520 ;
        RECT 3516.460 2015.240 3516.740 2015.520 ;
        RECT 3517.170 2015.240 3517.450 2015.520 ;
        RECT 3517.880 2015.240 3518.160 2015.520 ;
        RECT 3518.590 2015.240 3518.870 2015.520 ;
        RECT 3519.300 2015.240 3519.580 2015.520 ;
        RECT 3520.010 2015.240 3520.290 2015.520 ;
        RECT 3520.720 2015.240 3521.000 2015.520 ;
        RECT 3521.430 2015.240 3521.710 2015.520 ;
        RECT 3512.200 2014.530 3512.480 2014.810 ;
        RECT 3512.910 2014.530 3513.190 2014.810 ;
        RECT 3513.620 2014.530 3513.900 2014.810 ;
        RECT 3514.330 2014.530 3514.610 2014.810 ;
        RECT 3515.040 2014.530 3515.320 2014.810 ;
        RECT 3515.750 2014.530 3516.030 2014.810 ;
        RECT 3516.460 2014.530 3516.740 2014.810 ;
        RECT 3517.170 2014.530 3517.450 2014.810 ;
        RECT 3517.880 2014.530 3518.160 2014.810 ;
        RECT 3518.590 2014.530 3518.870 2014.810 ;
        RECT 3519.300 2014.530 3519.580 2014.810 ;
        RECT 3520.010 2014.530 3520.290 2014.810 ;
        RECT 3520.720 2014.530 3521.000 2014.810 ;
        RECT 3521.430 2014.530 3521.710 2014.810 ;
        RECT 3512.255 2010.615 3512.535 2010.895 ;
        RECT 3512.965 2010.615 3513.245 2010.895 ;
        RECT 3513.675 2010.615 3513.955 2010.895 ;
        RECT 3514.385 2010.615 3514.665 2010.895 ;
        RECT 3515.095 2010.615 3515.375 2010.895 ;
        RECT 3515.805 2010.615 3516.085 2010.895 ;
        RECT 3516.515 2010.615 3516.795 2010.895 ;
        RECT 3517.225 2010.615 3517.505 2010.895 ;
        RECT 3517.935 2010.615 3518.215 2010.895 ;
        RECT 3518.645 2010.615 3518.925 2010.895 ;
        RECT 3519.355 2010.615 3519.635 2010.895 ;
        RECT 3520.065 2010.615 3520.345 2010.895 ;
        RECT 3520.775 2010.615 3521.055 2010.895 ;
        RECT 3521.485 2010.615 3521.765 2010.895 ;
        RECT 3512.255 2009.905 3512.535 2010.185 ;
        RECT 3512.965 2009.905 3513.245 2010.185 ;
        RECT 3513.675 2009.905 3513.955 2010.185 ;
        RECT 3514.385 2009.905 3514.665 2010.185 ;
        RECT 3515.095 2009.905 3515.375 2010.185 ;
        RECT 3515.805 2009.905 3516.085 2010.185 ;
        RECT 3516.515 2009.905 3516.795 2010.185 ;
        RECT 3517.225 2009.905 3517.505 2010.185 ;
        RECT 3517.935 2009.905 3518.215 2010.185 ;
        RECT 3518.645 2009.905 3518.925 2010.185 ;
        RECT 3519.355 2009.905 3519.635 2010.185 ;
        RECT 3520.065 2009.905 3520.345 2010.185 ;
        RECT 3520.775 2009.905 3521.055 2010.185 ;
        RECT 3521.485 2009.905 3521.765 2010.185 ;
        RECT 3512.255 2009.195 3512.535 2009.475 ;
        RECT 3512.965 2009.195 3513.245 2009.475 ;
        RECT 3513.675 2009.195 3513.955 2009.475 ;
        RECT 3514.385 2009.195 3514.665 2009.475 ;
        RECT 3515.095 2009.195 3515.375 2009.475 ;
        RECT 3515.805 2009.195 3516.085 2009.475 ;
        RECT 3516.515 2009.195 3516.795 2009.475 ;
        RECT 3517.225 2009.195 3517.505 2009.475 ;
        RECT 3517.935 2009.195 3518.215 2009.475 ;
        RECT 3518.645 2009.195 3518.925 2009.475 ;
        RECT 3519.355 2009.195 3519.635 2009.475 ;
        RECT 3520.065 2009.195 3520.345 2009.475 ;
        RECT 3520.775 2009.195 3521.055 2009.475 ;
        RECT 3521.485 2009.195 3521.765 2009.475 ;
        RECT 3512.255 2008.485 3512.535 2008.765 ;
        RECT 3512.965 2008.485 3513.245 2008.765 ;
        RECT 3513.675 2008.485 3513.955 2008.765 ;
        RECT 3514.385 2008.485 3514.665 2008.765 ;
        RECT 3515.095 2008.485 3515.375 2008.765 ;
        RECT 3515.805 2008.485 3516.085 2008.765 ;
        RECT 3516.515 2008.485 3516.795 2008.765 ;
        RECT 3517.225 2008.485 3517.505 2008.765 ;
        RECT 3517.935 2008.485 3518.215 2008.765 ;
        RECT 3518.645 2008.485 3518.925 2008.765 ;
        RECT 3519.355 2008.485 3519.635 2008.765 ;
        RECT 3520.065 2008.485 3520.345 2008.765 ;
        RECT 3520.775 2008.485 3521.055 2008.765 ;
        RECT 3521.485 2008.485 3521.765 2008.765 ;
        RECT 3512.255 2007.775 3512.535 2008.055 ;
        RECT 3512.965 2007.775 3513.245 2008.055 ;
        RECT 3513.675 2007.775 3513.955 2008.055 ;
        RECT 3514.385 2007.775 3514.665 2008.055 ;
        RECT 3515.095 2007.775 3515.375 2008.055 ;
        RECT 3515.805 2007.775 3516.085 2008.055 ;
        RECT 3516.515 2007.775 3516.795 2008.055 ;
        RECT 3517.225 2007.775 3517.505 2008.055 ;
        RECT 3517.935 2007.775 3518.215 2008.055 ;
        RECT 3518.645 2007.775 3518.925 2008.055 ;
        RECT 3519.355 2007.775 3519.635 2008.055 ;
        RECT 3520.065 2007.775 3520.345 2008.055 ;
        RECT 3520.775 2007.775 3521.055 2008.055 ;
        RECT 3521.485 2007.775 3521.765 2008.055 ;
        RECT 3512.255 2007.065 3512.535 2007.345 ;
        RECT 3512.965 2007.065 3513.245 2007.345 ;
        RECT 3513.675 2007.065 3513.955 2007.345 ;
        RECT 3514.385 2007.065 3514.665 2007.345 ;
        RECT 3515.095 2007.065 3515.375 2007.345 ;
        RECT 3515.805 2007.065 3516.085 2007.345 ;
        RECT 3516.515 2007.065 3516.795 2007.345 ;
        RECT 3517.225 2007.065 3517.505 2007.345 ;
        RECT 3517.935 2007.065 3518.215 2007.345 ;
        RECT 3518.645 2007.065 3518.925 2007.345 ;
        RECT 3519.355 2007.065 3519.635 2007.345 ;
        RECT 3520.065 2007.065 3520.345 2007.345 ;
        RECT 3520.775 2007.065 3521.055 2007.345 ;
        RECT 3521.485 2007.065 3521.765 2007.345 ;
        RECT 3512.255 2006.355 3512.535 2006.635 ;
        RECT 3512.965 2006.355 3513.245 2006.635 ;
        RECT 3513.675 2006.355 3513.955 2006.635 ;
        RECT 3514.385 2006.355 3514.665 2006.635 ;
        RECT 3515.095 2006.355 3515.375 2006.635 ;
        RECT 3515.805 2006.355 3516.085 2006.635 ;
        RECT 3516.515 2006.355 3516.795 2006.635 ;
        RECT 3517.225 2006.355 3517.505 2006.635 ;
        RECT 3517.935 2006.355 3518.215 2006.635 ;
        RECT 3518.645 2006.355 3518.925 2006.635 ;
        RECT 3519.355 2006.355 3519.635 2006.635 ;
        RECT 3520.065 2006.355 3520.345 2006.635 ;
        RECT 3520.775 2006.355 3521.055 2006.635 ;
        RECT 3521.485 2006.355 3521.765 2006.635 ;
        RECT 3512.255 2005.645 3512.535 2005.925 ;
        RECT 3512.965 2005.645 3513.245 2005.925 ;
        RECT 3513.675 2005.645 3513.955 2005.925 ;
        RECT 3514.385 2005.645 3514.665 2005.925 ;
        RECT 3515.095 2005.645 3515.375 2005.925 ;
        RECT 3515.805 2005.645 3516.085 2005.925 ;
        RECT 3516.515 2005.645 3516.795 2005.925 ;
        RECT 3517.225 2005.645 3517.505 2005.925 ;
        RECT 3517.935 2005.645 3518.215 2005.925 ;
        RECT 3518.645 2005.645 3518.925 2005.925 ;
        RECT 3519.355 2005.645 3519.635 2005.925 ;
        RECT 3520.065 2005.645 3520.345 2005.925 ;
        RECT 3520.775 2005.645 3521.055 2005.925 ;
        RECT 3521.485 2005.645 3521.765 2005.925 ;
        RECT 3512.255 2004.935 3512.535 2005.215 ;
        RECT 3512.965 2004.935 3513.245 2005.215 ;
        RECT 3513.675 2004.935 3513.955 2005.215 ;
        RECT 3514.385 2004.935 3514.665 2005.215 ;
        RECT 3515.095 2004.935 3515.375 2005.215 ;
        RECT 3515.805 2004.935 3516.085 2005.215 ;
        RECT 3516.515 2004.935 3516.795 2005.215 ;
        RECT 3517.225 2004.935 3517.505 2005.215 ;
        RECT 3517.935 2004.935 3518.215 2005.215 ;
        RECT 3518.645 2004.935 3518.925 2005.215 ;
        RECT 3519.355 2004.935 3519.635 2005.215 ;
        RECT 3520.065 2004.935 3520.345 2005.215 ;
        RECT 3520.775 2004.935 3521.055 2005.215 ;
        RECT 3521.485 2004.935 3521.765 2005.215 ;
        RECT 3512.255 2004.225 3512.535 2004.505 ;
        RECT 3512.965 2004.225 3513.245 2004.505 ;
        RECT 3513.675 2004.225 3513.955 2004.505 ;
        RECT 3514.385 2004.225 3514.665 2004.505 ;
        RECT 3515.095 2004.225 3515.375 2004.505 ;
        RECT 3515.805 2004.225 3516.085 2004.505 ;
        RECT 3516.515 2004.225 3516.795 2004.505 ;
        RECT 3517.225 2004.225 3517.505 2004.505 ;
        RECT 3517.935 2004.225 3518.215 2004.505 ;
        RECT 3518.645 2004.225 3518.925 2004.505 ;
        RECT 3519.355 2004.225 3519.635 2004.505 ;
        RECT 3520.065 2004.225 3520.345 2004.505 ;
        RECT 3520.775 2004.225 3521.055 2004.505 ;
        RECT 3521.485 2004.225 3521.765 2004.505 ;
        RECT 3512.255 2003.515 3512.535 2003.795 ;
        RECT 3512.965 2003.515 3513.245 2003.795 ;
        RECT 3513.675 2003.515 3513.955 2003.795 ;
        RECT 3514.385 2003.515 3514.665 2003.795 ;
        RECT 3515.095 2003.515 3515.375 2003.795 ;
        RECT 3515.805 2003.515 3516.085 2003.795 ;
        RECT 3516.515 2003.515 3516.795 2003.795 ;
        RECT 3517.225 2003.515 3517.505 2003.795 ;
        RECT 3517.935 2003.515 3518.215 2003.795 ;
        RECT 3518.645 2003.515 3518.925 2003.795 ;
        RECT 3519.355 2003.515 3519.635 2003.795 ;
        RECT 3520.065 2003.515 3520.345 2003.795 ;
        RECT 3520.775 2003.515 3521.055 2003.795 ;
        RECT 3521.485 2003.515 3521.765 2003.795 ;
        RECT 3512.255 2002.805 3512.535 2003.085 ;
        RECT 3512.965 2002.805 3513.245 2003.085 ;
        RECT 3513.675 2002.805 3513.955 2003.085 ;
        RECT 3514.385 2002.805 3514.665 2003.085 ;
        RECT 3515.095 2002.805 3515.375 2003.085 ;
        RECT 3515.805 2002.805 3516.085 2003.085 ;
        RECT 3516.515 2002.805 3516.795 2003.085 ;
        RECT 3517.225 2002.805 3517.505 2003.085 ;
        RECT 3517.935 2002.805 3518.215 2003.085 ;
        RECT 3518.645 2002.805 3518.925 2003.085 ;
        RECT 3519.355 2002.805 3519.635 2003.085 ;
        RECT 3520.065 2002.805 3520.345 2003.085 ;
        RECT 3520.775 2002.805 3521.055 2003.085 ;
        RECT 3521.485 2002.805 3521.765 2003.085 ;
        RECT 3512.255 2002.095 3512.535 2002.375 ;
        RECT 3512.965 2002.095 3513.245 2002.375 ;
        RECT 3513.675 2002.095 3513.955 2002.375 ;
        RECT 3514.385 2002.095 3514.665 2002.375 ;
        RECT 3515.095 2002.095 3515.375 2002.375 ;
        RECT 3515.805 2002.095 3516.085 2002.375 ;
        RECT 3516.515 2002.095 3516.795 2002.375 ;
        RECT 3517.225 2002.095 3517.505 2002.375 ;
        RECT 3517.935 2002.095 3518.215 2002.375 ;
        RECT 3518.645 2002.095 3518.925 2002.375 ;
        RECT 3519.355 2002.095 3519.635 2002.375 ;
        RECT 3520.065 2002.095 3520.345 2002.375 ;
        RECT 3520.775 2002.095 3521.055 2002.375 ;
        RECT 3521.485 2002.095 3521.765 2002.375 ;
        RECT 3512.255 2001.385 3512.535 2001.665 ;
        RECT 3512.965 2001.385 3513.245 2001.665 ;
        RECT 3513.675 2001.385 3513.955 2001.665 ;
        RECT 3514.385 2001.385 3514.665 2001.665 ;
        RECT 3515.095 2001.385 3515.375 2001.665 ;
        RECT 3515.805 2001.385 3516.085 2001.665 ;
        RECT 3516.515 2001.385 3516.795 2001.665 ;
        RECT 3517.225 2001.385 3517.505 2001.665 ;
        RECT 3517.935 2001.385 3518.215 2001.665 ;
        RECT 3518.645 2001.385 3518.925 2001.665 ;
        RECT 3519.355 2001.385 3519.635 2001.665 ;
        RECT 3520.065 2001.385 3520.345 2001.665 ;
        RECT 3520.775 2001.385 3521.055 2001.665 ;
        RECT 3521.485 2001.385 3521.765 2001.665 ;
        RECT 3512.255 1998.765 3512.535 1999.045 ;
        RECT 3512.965 1998.765 3513.245 1999.045 ;
        RECT 3513.675 1998.765 3513.955 1999.045 ;
        RECT 3514.385 1998.765 3514.665 1999.045 ;
        RECT 3515.095 1998.765 3515.375 1999.045 ;
        RECT 3515.805 1998.765 3516.085 1999.045 ;
        RECT 3516.515 1998.765 3516.795 1999.045 ;
        RECT 3517.225 1998.765 3517.505 1999.045 ;
        RECT 3517.935 1998.765 3518.215 1999.045 ;
        RECT 3518.645 1998.765 3518.925 1999.045 ;
        RECT 3519.355 1998.765 3519.635 1999.045 ;
        RECT 3520.065 1998.765 3520.345 1999.045 ;
        RECT 3520.775 1998.765 3521.055 1999.045 ;
        RECT 3521.485 1998.765 3521.765 1999.045 ;
        RECT 3512.255 1998.055 3512.535 1998.335 ;
        RECT 3512.965 1998.055 3513.245 1998.335 ;
        RECT 3513.675 1998.055 3513.955 1998.335 ;
        RECT 3514.385 1998.055 3514.665 1998.335 ;
        RECT 3515.095 1998.055 3515.375 1998.335 ;
        RECT 3515.805 1998.055 3516.085 1998.335 ;
        RECT 3516.515 1998.055 3516.795 1998.335 ;
        RECT 3517.225 1998.055 3517.505 1998.335 ;
        RECT 3517.935 1998.055 3518.215 1998.335 ;
        RECT 3518.645 1998.055 3518.925 1998.335 ;
        RECT 3519.355 1998.055 3519.635 1998.335 ;
        RECT 3520.065 1998.055 3520.345 1998.335 ;
        RECT 3520.775 1998.055 3521.055 1998.335 ;
        RECT 3521.485 1998.055 3521.765 1998.335 ;
        RECT 3512.255 1997.345 3512.535 1997.625 ;
        RECT 3512.965 1997.345 3513.245 1997.625 ;
        RECT 3513.675 1997.345 3513.955 1997.625 ;
        RECT 3514.385 1997.345 3514.665 1997.625 ;
        RECT 3515.095 1997.345 3515.375 1997.625 ;
        RECT 3515.805 1997.345 3516.085 1997.625 ;
        RECT 3516.515 1997.345 3516.795 1997.625 ;
        RECT 3517.225 1997.345 3517.505 1997.625 ;
        RECT 3517.935 1997.345 3518.215 1997.625 ;
        RECT 3518.645 1997.345 3518.925 1997.625 ;
        RECT 3519.355 1997.345 3519.635 1997.625 ;
        RECT 3520.065 1997.345 3520.345 1997.625 ;
        RECT 3520.775 1997.345 3521.055 1997.625 ;
        RECT 3521.485 1997.345 3521.765 1997.625 ;
        RECT 3512.255 1996.635 3512.535 1996.915 ;
        RECT 3512.965 1996.635 3513.245 1996.915 ;
        RECT 3513.675 1996.635 3513.955 1996.915 ;
        RECT 3514.385 1996.635 3514.665 1996.915 ;
        RECT 3515.095 1996.635 3515.375 1996.915 ;
        RECT 3515.805 1996.635 3516.085 1996.915 ;
        RECT 3516.515 1996.635 3516.795 1996.915 ;
        RECT 3517.225 1996.635 3517.505 1996.915 ;
        RECT 3517.935 1996.635 3518.215 1996.915 ;
        RECT 3518.645 1996.635 3518.925 1996.915 ;
        RECT 3519.355 1996.635 3519.635 1996.915 ;
        RECT 3520.065 1996.635 3520.345 1996.915 ;
        RECT 3520.775 1996.635 3521.055 1996.915 ;
        RECT 3521.485 1996.635 3521.765 1996.915 ;
        RECT 3512.255 1995.925 3512.535 1996.205 ;
        RECT 3512.965 1995.925 3513.245 1996.205 ;
        RECT 3513.675 1995.925 3513.955 1996.205 ;
        RECT 3514.385 1995.925 3514.665 1996.205 ;
        RECT 3515.095 1995.925 3515.375 1996.205 ;
        RECT 3515.805 1995.925 3516.085 1996.205 ;
        RECT 3516.515 1995.925 3516.795 1996.205 ;
        RECT 3517.225 1995.925 3517.505 1996.205 ;
        RECT 3517.935 1995.925 3518.215 1996.205 ;
        RECT 3518.645 1995.925 3518.925 1996.205 ;
        RECT 3519.355 1995.925 3519.635 1996.205 ;
        RECT 3520.065 1995.925 3520.345 1996.205 ;
        RECT 3520.775 1995.925 3521.055 1996.205 ;
        RECT 3521.485 1995.925 3521.765 1996.205 ;
        RECT 3512.255 1995.215 3512.535 1995.495 ;
        RECT 3512.965 1995.215 3513.245 1995.495 ;
        RECT 3513.675 1995.215 3513.955 1995.495 ;
        RECT 3514.385 1995.215 3514.665 1995.495 ;
        RECT 3515.095 1995.215 3515.375 1995.495 ;
        RECT 3515.805 1995.215 3516.085 1995.495 ;
        RECT 3516.515 1995.215 3516.795 1995.495 ;
        RECT 3517.225 1995.215 3517.505 1995.495 ;
        RECT 3517.935 1995.215 3518.215 1995.495 ;
        RECT 3518.645 1995.215 3518.925 1995.495 ;
        RECT 3519.355 1995.215 3519.635 1995.495 ;
        RECT 3520.065 1995.215 3520.345 1995.495 ;
        RECT 3520.775 1995.215 3521.055 1995.495 ;
        RECT 3521.485 1995.215 3521.765 1995.495 ;
        RECT 3512.255 1994.505 3512.535 1994.785 ;
        RECT 3512.965 1994.505 3513.245 1994.785 ;
        RECT 3513.675 1994.505 3513.955 1994.785 ;
        RECT 3514.385 1994.505 3514.665 1994.785 ;
        RECT 3515.095 1994.505 3515.375 1994.785 ;
        RECT 3515.805 1994.505 3516.085 1994.785 ;
        RECT 3516.515 1994.505 3516.795 1994.785 ;
        RECT 3517.225 1994.505 3517.505 1994.785 ;
        RECT 3517.935 1994.505 3518.215 1994.785 ;
        RECT 3518.645 1994.505 3518.925 1994.785 ;
        RECT 3519.355 1994.505 3519.635 1994.785 ;
        RECT 3520.065 1994.505 3520.345 1994.785 ;
        RECT 3520.775 1994.505 3521.055 1994.785 ;
        RECT 3521.485 1994.505 3521.765 1994.785 ;
        RECT 3512.255 1993.795 3512.535 1994.075 ;
        RECT 3512.965 1993.795 3513.245 1994.075 ;
        RECT 3513.675 1993.795 3513.955 1994.075 ;
        RECT 3514.385 1993.795 3514.665 1994.075 ;
        RECT 3515.095 1993.795 3515.375 1994.075 ;
        RECT 3515.805 1993.795 3516.085 1994.075 ;
        RECT 3516.515 1993.795 3516.795 1994.075 ;
        RECT 3517.225 1993.795 3517.505 1994.075 ;
        RECT 3517.935 1993.795 3518.215 1994.075 ;
        RECT 3518.645 1993.795 3518.925 1994.075 ;
        RECT 3519.355 1993.795 3519.635 1994.075 ;
        RECT 3520.065 1993.795 3520.345 1994.075 ;
        RECT 3520.775 1993.795 3521.055 1994.075 ;
        RECT 3521.485 1993.795 3521.765 1994.075 ;
        RECT 3512.255 1993.085 3512.535 1993.365 ;
        RECT 3512.965 1993.085 3513.245 1993.365 ;
        RECT 3513.675 1993.085 3513.955 1993.365 ;
        RECT 3514.385 1993.085 3514.665 1993.365 ;
        RECT 3515.095 1993.085 3515.375 1993.365 ;
        RECT 3515.805 1993.085 3516.085 1993.365 ;
        RECT 3516.515 1993.085 3516.795 1993.365 ;
        RECT 3517.225 1993.085 3517.505 1993.365 ;
        RECT 3517.935 1993.085 3518.215 1993.365 ;
        RECT 3518.645 1993.085 3518.925 1993.365 ;
        RECT 3519.355 1993.085 3519.635 1993.365 ;
        RECT 3520.065 1993.085 3520.345 1993.365 ;
        RECT 3520.775 1993.085 3521.055 1993.365 ;
        RECT 3521.485 1993.085 3521.765 1993.365 ;
        RECT 3512.255 1992.375 3512.535 1992.655 ;
        RECT 3512.965 1992.375 3513.245 1992.655 ;
        RECT 3513.675 1992.375 3513.955 1992.655 ;
        RECT 3514.385 1992.375 3514.665 1992.655 ;
        RECT 3515.095 1992.375 3515.375 1992.655 ;
        RECT 3515.805 1992.375 3516.085 1992.655 ;
        RECT 3516.515 1992.375 3516.795 1992.655 ;
        RECT 3517.225 1992.375 3517.505 1992.655 ;
        RECT 3517.935 1992.375 3518.215 1992.655 ;
        RECT 3518.645 1992.375 3518.925 1992.655 ;
        RECT 3519.355 1992.375 3519.635 1992.655 ;
        RECT 3520.065 1992.375 3520.345 1992.655 ;
        RECT 3520.775 1992.375 3521.055 1992.655 ;
        RECT 3521.485 1992.375 3521.765 1992.655 ;
        RECT 3512.255 1991.665 3512.535 1991.945 ;
        RECT 3512.965 1991.665 3513.245 1991.945 ;
        RECT 3513.675 1991.665 3513.955 1991.945 ;
        RECT 3514.385 1991.665 3514.665 1991.945 ;
        RECT 3515.095 1991.665 3515.375 1991.945 ;
        RECT 3515.805 1991.665 3516.085 1991.945 ;
        RECT 3516.515 1991.665 3516.795 1991.945 ;
        RECT 3517.225 1991.665 3517.505 1991.945 ;
        RECT 3517.935 1991.665 3518.215 1991.945 ;
        RECT 3518.645 1991.665 3518.925 1991.945 ;
        RECT 3519.355 1991.665 3519.635 1991.945 ;
        RECT 3520.065 1991.665 3520.345 1991.945 ;
        RECT 3520.775 1991.665 3521.055 1991.945 ;
        RECT 3521.485 1991.665 3521.765 1991.945 ;
        RECT 3512.255 1990.955 3512.535 1991.235 ;
        RECT 3512.965 1990.955 3513.245 1991.235 ;
        RECT 3513.675 1990.955 3513.955 1991.235 ;
        RECT 3514.385 1990.955 3514.665 1991.235 ;
        RECT 3515.095 1990.955 3515.375 1991.235 ;
        RECT 3515.805 1990.955 3516.085 1991.235 ;
        RECT 3516.515 1990.955 3516.795 1991.235 ;
        RECT 3517.225 1990.955 3517.505 1991.235 ;
        RECT 3517.935 1990.955 3518.215 1991.235 ;
        RECT 3518.645 1990.955 3518.925 1991.235 ;
        RECT 3519.355 1990.955 3519.635 1991.235 ;
        RECT 3520.065 1990.955 3520.345 1991.235 ;
        RECT 3520.775 1990.955 3521.055 1991.235 ;
        RECT 3521.485 1990.955 3521.765 1991.235 ;
        RECT 3512.255 1990.245 3512.535 1990.525 ;
        RECT 3512.965 1990.245 3513.245 1990.525 ;
        RECT 3513.675 1990.245 3513.955 1990.525 ;
        RECT 3514.385 1990.245 3514.665 1990.525 ;
        RECT 3515.095 1990.245 3515.375 1990.525 ;
        RECT 3515.805 1990.245 3516.085 1990.525 ;
        RECT 3516.515 1990.245 3516.795 1990.525 ;
        RECT 3517.225 1990.245 3517.505 1990.525 ;
        RECT 3517.935 1990.245 3518.215 1990.525 ;
        RECT 3518.645 1990.245 3518.925 1990.525 ;
        RECT 3519.355 1990.245 3519.635 1990.525 ;
        RECT 3520.065 1990.245 3520.345 1990.525 ;
        RECT 3520.775 1990.245 3521.055 1990.525 ;
        RECT 3521.485 1990.245 3521.765 1990.525 ;
        RECT 3512.255 1989.535 3512.535 1989.815 ;
        RECT 3512.965 1989.535 3513.245 1989.815 ;
        RECT 3513.675 1989.535 3513.955 1989.815 ;
        RECT 3514.385 1989.535 3514.665 1989.815 ;
        RECT 3515.095 1989.535 3515.375 1989.815 ;
        RECT 3515.805 1989.535 3516.085 1989.815 ;
        RECT 3516.515 1989.535 3516.795 1989.815 ;
        RECT 3517.225 1989.535 3517.505 1989.815 ;
        RECT 3517.935 1989.535 3518.215 1989.815 ;
        RECT 3518.645 1989.535 3518.925 1989.815 ;
        RECT 3519.355 1989.535 3519.635 1989.815 ;
        RECT 3520.065 1989.535 3520.345 1989.815 ;
        RECT 3520.775 1989.535 3521.055 1989.815 ;
        RECT 3521.485 1989.535 3521.765 1989.815 ;
        RECT 3512.255 1985.235 3512.535 1985.515 ;
        RECT 3512.965 1985.235 3513.245 1985.515 ;
        RECT 3513.675 1985.235 3513.955 1985.515 ;
        RECT 3514.385 1985.235 3514.665 1985.515 ;
        RECT 3515.095 1985.235 3515.375 1985.515 ;
        RECT 3515.805 1985.235 3516.085 1985.515 ;
        RECT 3516.515 1985.235 3516.795 1985.515 ;
        RECT 3517.225 1985.235 3517.505 1985.515 ;
        RECT 3517.935 1985.235 3518.215 1985.515 ;
        RECT 3518.645 1985.235 3518.925 1985.515 ;
        RECT 3519.355 1985.235 3519.635 1985.515 ;
        RECT 3520.065 1985.235 3520.345 1985.515 ;
        RECT 3520.775 1985.235 3521.055 1985.515 ;
        RECT 3521.485 1985.235 3521.765 1985.515 ;
        RECT 3512.255 1984.525 3512.535 1984.805 ;
        RECT 3512.965 1984.525 3513.245 1984.805 ;
        RECT 3513.675 1984.525 3513.955 1984.805 ;
        RECT 3514.385 1984.525 3514.665 1984.805 ;
        RECT 3515.095 1984.525 3515.375 1984.805 ;
        RECT 3515.805 1984.525 3516.085 1984.805 ;
        RECT 3516.515 1984.525 3516.795 1984.805 ;
        RECT 3517.225 1984.525 3517.505 1984.805 ;
        RECT 3517.935 1984.525 3518.215 1984.805 ;
        RECT 3518.645 1984.525 3518.925 1984.805 ;
        RECT 3519.355 1984.525 3519.635 1984.805 ;
        RECT 3520.065 1984.525 3520.345 1984.805 ;
        RECT 3520.775 1984.525 3521.055 1984.805 ;
        RECT 3521.485 1984.525 3521.765 1984.805 ;
        RECT 3512.255 1983.815 3512.535 1984.095 ;
        RECT 3512.965 1983.815 3513.245 1984.095 ;
        RECT 3513.675 1983.815 3513.955 1984.095 ;
        RECT 3514.385 1983.815 3514.665 1984.095 ;
        RECT 3515.095 1983.815 3515.375 1984.095 ;
        RECT 3515.805 1983.815 3516.085 1984.095 ;
        RECT 3516.515 1983.815 3516.795 1984.095 ;
        RECT 3517.225 1983.815 3517.505 1984.095 ;
        RECT 3517.935 1983.815 3518.215 1984.095 ;
        RECT 3518.645 1983.815 3518.925 1984.095 ;
        RECT 3519.355 1983.815 3519.635 1984.095 ;
        RECT 3520.065 1983.815 3520.345 1984.095 ;
        RECT 3520.775 1983.815 3521.055 1984.095 ;
        RECT 3521.485 1983.815 3521.765 1984.095 ;
        RECT 3512.255 1983.105 3512.535 1983.385 ;
        RECT 3512.965 1983.105 3513.245 1983.385 ;
        RECT 3513.675 1983.105 3513.955 1983.385 ;
        RECT 3514.385 1983.105 3514.665 1983.385 ;
        RECT 3515.095 1983.105 3515.375 1983.385 ;
        RECT 3515.805 1983.105 3516.085 1983.385 ;
        RECT 3516.515 1983.105 3516.795 1983.385 ;
        RECT 3517.225 1983.105 3517.505 1983.385 ;
        RECT 3517.935 1983.105 3518.215 1983.385 ;
        RECT 3518.645 1983.105 3518.925 1983.385 ;
        RECT 3519.355 1983.105 3519.635 1983.385 ;
        RECT 3520.065 1983.105 3520.345 1983.385 ;
        RECT 3520.775 1983.105 3521.055 1983.385 ;
        RECT 3521.485 1983.105 3521.765 1983.385 ;
        RECT 3512.255 1982.395 3512.535 1982.675 ;
        RECT 3512.965 1982.395 3513.245 1982.675 ;
        RECT 3513.675 1982.395 3513.955 1982.675 ;
        RECT 3514.385 1982.395 3514.665 1982.675 ;
        RECT 3515.095 1982.395 3515.375 1982.675 ;
        RECT 3515.805 1982.395 3516.085 1982.675 ;
        RECT 3516.515 1982.395 3516.795 1982.675 ;
        RECT 3517.225 1982.395 3517.505 1982.675 ;
        RECT 3517.935 1982.395 3518.215 1982.675 ;
        RECT 3518.645 1982.395 3518.925 1982.675 ;
        RECT 3519.355 1982.395 3519.635 1982.675 ;
        RECT 3520.065 1982.395 3520.345 1982.675 ;
        RECT 3520.775 1982.395 3521.055 1982.675 ;
        RECT 3521.485 1982.395 3521.765 1982.675 ;
        RECT 3512.255 1981.685 3512.535 1981.965 ;
        RECT 3512.965 1981.685 3513.245 1981.965 ;
        RECT 3513.675 1981.685 3513.955 1981.965 ;
        RECT 3514.385 1981.685 3514.665 1981.965 ;
        RECT 3515.095 1981.685 3515.375 1981.965 ;
        RECT 3515.805 1981.685 3516.085 1981.965 ;
        RECT 3516.515 1981.685 3516.795 1981.965 ;
        RECT 3517.225 1981.685 3517.505 1981.965 ;
        RECT 3517.935 1981.685 3518.215 1981.965 ;
        RECT 3518.645 1981.685 3518.925 1981.965 ;
        RECT 3519.355 1981.685 3519.635 1981.965 ;
        RECT 3520.065 1981.685 3520.345 1981.965 ;
        RECT 3520.775 1981.685 3521.055 1981.965 ;
        RECT 3521.485 1981.685 3521.765 1981.965 ;
        RECT 3512.255 1980.975 3512.535 1981.255 ;
        RECT 3512.965 1980.975 3513.245 1981.255 ;
        RECT 3513.675 1980.975 3513.955 1981.255 ;
        RECT 3514.385 1980.975 3514.665 1981.255 ;
        RECT 3515.095 1980.975 3515.375 1981.255 ;
        RECT 3515.805 1980.975 3516.085 1981.255 ;
        RECT 3516.515 1980.975 3516.795 1981.255 ;
        RECT 3517.225 1980.975 3517.505 1981.255 ;
        RECT 3517.935 1980.975 3518.215 1981.255 ;
        RECT 3518.645 1980.975 3518.925 1981.255 ;
        RECT 3519.355 1980.975 3519.635 1981.255 ;
        RECT 3520.065 1980.975 3520.345 1981.255 ;
        RECT 3520.775 1980.975 3521.055 1981.255 ;
        RECT 3521.485 1980.975 3521.765 1981.255 ;
        RECT 3512.255 1980.265 3512.535 1980.545 ;
        RECT 3512.965 1980.265 3513.245 1980.545 ;
        RECT 3513.675 1980.265 3513.955 1980.545 ;
        RECT 3514.385 1980.265 3514.665 1980.545 ;
        RECT 3515.095 1980.265 3515.375 1980.545 ;
        RECT 3515.805 1980.265 3516.085 1980.545 ;
        RECT 3516.515 1980.265 3516.795 1980.545 ;
        RECT 3517.225 1980.265 3517.505 1980.545 ;
        RECT 3517.935 1980.265 3518.215 1980.545 ;
        RECT 3518.645 1980.265 3518.925 1980.545 ;
        RECT 3519.355 1980.265 3519.635 1980.545 ;
        RECT 3520.065 1980.265 3520.345 1980.545 ;
        RECT 3520.775 1980.265 3521.055 1980.545 ;
        RECT 3521.485 1980.265 3521.765 1980.545 ;
        RECT 3512.255 1979.555 3512.535 1979.835 ;
        RECT 3512.965 1979.555 3513.245 1979.835 ;
        RECT 3513.675 1979.555 3513.955 1979.835 ;
        RECT 3514.385 1979.555 3514.665 1979.835 ;
        RECT 3515.095 1979.555 3515.375 1979.835 ;
        RECT 3515.805 1979.555 3516.085 1979.835 ;
        RECT 3516.515 1979.555 3516.795 1979.835 ;
        RECT 3517.225 1979.555 3517.505 1979.835 ;
        RECT 3517.935 1979.555 3518.215 1979.835 ;
        RECT 3518.645 1979.555 3518.925 1979.835 ;
        RECT 3519.355 1979.555 3519.635 1979.835 ;
        RECT 3520.065 1979.555 3520.345 1979.835 ;
        RECT 3520.775 1979.555 3521.055 1979.835 ;
        RECT 3521.485 1979.555 3521.765 1979.835 ;
        RECT 3512.255 1978.845 3512.535 1979.125 ;
        RECT 3512.965 1978.845 3513.245 1979.125 ;
        RECT 3513.675 1978.845 3513.955 1979.125 ;
        RECT 3514.385 1978.845 3514.665 1979.125 ;
        RECT 3515.095 1978.845 3515.375 1979.125 ;
        RECT 3515.805 1978.845 3516.085 1979.125 ;
        RECT 3516.515 1978.845 3516.795 1979.125 ;
        RECT 3517.225 1978.845 3517.505 1979.125 ;
        RECT 3517.935 1978.845 3518.215 1979.125 ;
        RECT 3518.645 1978.845 3518.925 1979.125 ;
        RECT 3519.355 1978.845 3519.635 1979.125 ;
        RECT 3520.065 1978.845 3520.345 1979.125 ;
        RECT 3520.775 1978.845 3521.055 1979.125 ;
        RECT 3521.485 1978.845 3521.765 1979.125 ;
        RECT 3512.255 1978.135 3512.535 1978.415 ;
        RECT 3512.965 1978.135 3513.245 1978.415 ;
        RECT 3513.675 1978.135 3513.955 1978.415 ;
        RECT 3514.385 1978.135 3514.665 1978.415 ;
        RECT 3515.095 1978.135 3515.375 1978.415 ;
        RECT 3515.805 1978.135 3516.085 1978.415 ;
        RECT 3516.515 1978.135 3516.795 1978.415 ;
        RECT 3517.225 1978.135 3517.505 1978.415 ;
        RECT 3517.935 1978.135 3518.215 1978.415 ;
        RECT 3518.645 1978.135 3518.925 1978.415 ;
        RECT 3519.355 1978.135 3519.635 1978.415 ;
        RECT 3520.065 1978.135 3520.345 1978.415 ;
        RECT 3520.775 1978.135 3521.055 1978.415 ;
        RECT 3521.485 1978.135 3521.765 1978.415 ;
        RECT 3512.255 1977.425 3512.535 1977.705 ;
        RECT 3512.965 1977.425 3513.245 1977.705 ;
        RECT 3513.675 1977.425 3513.955 1977.705 ;
        RECT 3514.385 1977.425 3514.665 1977.705 ;
        RECT 3515.095 1977.425 3515.375 1977.705 ;
        RECT 3515.805 1977.425 3516.085 1977.705 ;
        RECT 3516.515 1977.425 3516.795 1977.705 ;
        RECT 3517.225 1977.425 3517.505 1977.705 ;
        RECT 3517.935 1977.425 3518.215 1977.705 ;
        RECT 3518.645 1977.425 3518.925 1977.705 ;
        RECT 3519.355 1977.425 3519.635 1977.705 ;
        RECT 3520.065 1977.425 3520.345 1977.705 ;
        RECT 3520.775 1977.425 3521.055 1977.705 ;
        RECT 3521.485 1977.425 3521.765 1977.705 ;
        RECT 3512.255 1976.715 3512.535 1976.995 ;
        RECT 3512.965 1976.715 3513.245 1976.995 ;
        RECT 3513.675 1976.715 3513.955 1976.995 ;
        RECT 3514.385 1976.715 3514.665 1976.995 ;
        RECT 3515.095 1976.715 3515.375 1976.995 ;
        RECT 3515.805 1976.715 3516.085 1976.995 ;
        RECT 3516.515 1976.715 3516.795 1976.995 ;
        RECT 3517.225 1976.715 3517.505 1976.995 ;
        RECT 3517.935 1976.715 3518.215 1976.995 ;
        RECT 3518.645 1976.715 3518.925 1976.995 ;
        RECT 3519.355 1976.715 3519.635 1976.995 ;
        RECT 3520.065 1976.715 3520.345 1976.995 ;
        RECT 3520.775 1976.715 3521.055 1976.995 ;
        RECT 3521.485 1976.715 3521.765 1976.995 ;
        RECT 3512.255 1976.005 3512.535 1976.285 ;
        RECT 3512.965 1976.005 3513.245 1976.285 ;
        RECT 3513.675 1976.005 3513.955 1976.285 ;
        RECT 3514.385 1976.005 3514.665 1976.285 ;
        RECT 3515.095 1976.005 3515.375 1976.285 ;
        RECT 3515.805 1976.005 3516.085 1976.285 ;
        RECT 3516.515 1976.005 3516.795 1976.285 ;
        RECT 3517.225 1976.005 3517.505 1976.285 ;
        RECT 3517.935 1976.005 3518.215 1976.285 ;
        RECT 3518.645 1976.005 3518.925 1976.285 ;
        RECT 3519.355 1976.005 3519.635 1976.285 ;
        RECT 3520.065 1976.005 3520.345 1976.285 ;
        RECT 3520.775 1976.005 3521.055 1976.285 ;
        RECT 3521.485 1976.005 3521.765 1976.285 ;
        RECT 3512.255 1973.385 3512.535 1973.665 ;
        RECT 3512.965 1973.385 3513.245 1973.665 ;
        RECT 3513.675 1973.385 3513.955 1973.665 ;
        RECT 3514.385 1973.385 3514.665 1973.665 ;
        RECT 3515.095 1973.385 3515.375 1973.665 ;
        RECT 3515.805 1973.385 3516.085 1973.665 ;
        RECT 3516.515 1973.385 3516.795 1973.665 ;
        RECT 3517.225 1973.385 3517.505 1973.665 ;
        RECT 3517.935 1973.385 3518.215 1973.665 ;
        RECT 3518.645 1973.385 3518.925 1973.665 ;
        RECT 3519.355 1973.385 3519.635 1973.665 ;
        RECT 3520.065 1973.385 3520.345 1973.665 ;
        RECT 3520.775 1973.385 3521.055 1973.665 ;
        RECT 3521.485 1973.385 3521.765 1973.665 ;
        RECT 3512.255 1972.675 3512.535 1972.955 ;
        RECT 3512.965 1972.675 3513.245 1972.955 ;
        RECT 3513.675 1972.675 3513.955 1972.955 ;
        RECT 3514.385 1972.675 3514.665 1972.955 ;
        RECT 3515.095 1972.675 3515.375 1972.955 ;
        RECT 3515.805 1972.675 3516.085 1972.955 ;
        RECT 3516.515 1972.675 3516.795 1972.955 ;
        RECT 3517.225 1972.675 3517.505 1972.955 ;
        RECT 3517.935 1972.675 3518.215 1972.955 ;
        RECT 3518.645 1972.675 3518.925 1972.955 ;
        RECT 3519.355 1972.675 3519.635 1972.955 ;
        RECT 3520.065 1972.675 3520.345 1972.955 ;
        RECT 3520.775 1972.675 3521.055 1972.955 ;
        RECT 3521.485 1972.675 3521.765 1972.955 ;
        RECT 3512.255 1971.965 3512.535 1972.245 ;
        RECT 3512.965 1971.965 3513.245 1972.245 ;
        RECT 3513.675 1971.965 3513.955 1972.245 ;
        RECT 3514.385 1971.965 3514.665 1972.245 ;
        RECT 3515.095 1971.965 3515.375 1972.245 ;
        RECT 3515.805 1971.965 3516.085 1972.245 ;
        RECT 3516.515 1971.965 3516.795 1972.245 ;
        RECT 3517.225 1971.965 3517.505 1972.245 ;
        RECT 3517.935 1971.965 3518.215 1972.245 ;
        RECT 3518.645 1971.965 3518.925 1972.245 ;
        RECT 3519.355 1971.965 3519.635 1972.245 ;
        RECT 3520.065 1971.965 3520.345 1972.245 ;
        RECT 3520.775 1971.965 3521.055 1972.245 ;
        RECT 3521.485 1971.965 3521.765 1972.245 ;
        RECT 3512.255 1971.255 3512.535 1971.535 ;
        RECT 3512.965 1971.255 3513.245 1971.535 ;
        RECT 3513.675 1971.255 3513.955 1971.535 ;
        RECT 3514.385 1971.255 3514.665 1971.535 ;
        RECT 3515.095 1971.255 3515.375 1971.535 ;
        RECT 3515.805 1971.255 3516.085 1971.535 ;
        RECT 3516.515 1971.255 3516.795 1971.535 ;
        RECT 3517.225 1971.255 3517.505 1971.535 ;
        RECT 3517.935 1971.255 3518.215 1971.535 ;
        RECT 3518.645 1971.255 3518.925 1971.535 ;
        RECT 3519.355 1971.255 3519.635 1971.535 ;
        RECT 3520.065 1971.255 3520.345 1971.535 ;
        RECT 3520.775 1971.255 3521.055 1971.535 ;
        RECT 3521.485 1971.255 3521.765 1971.535 ;
        RECT 3512.255 1970.545 3512.535 1970.825 ;
        RECT 3512.965 1970.545 3513.245 1970.825 ;
        RECT 3513.675 1970.545 3513.955 1970.825 ;
        RECT 3514.385 1970.545 3514.665 1970.825 ;
        RECT 3515.095 1970.545 3515.375 1970.825 ;
        RECT 3515.805 1970.545 3516.085 1970.825 ;
        RECT 3516.515 1970.545 3516.795 1970.825 ;
        RECT 3517.225 1970.545 3517.505 1970.825 ;
        RECT 3517.935 1970.545 3518.215 1970.825 ;
        RECT 3518.645 1970.545 3518.925 1970.825 ;
        RECT 3519.355 1970.545 3519.635 1970.825 ;
        RECT 3520.065 1970.545 3520.345 1970.825 ;
        RECT 3520.775 1970.545 3521.055 1970.825 ;
        RECT 3521.485 1970.545 3521.765 1970.825 ;
        RECT 3512.255 1969.835 3512.535 1970.115 ;
        RECT 3512.965 1969.835 3513.245 1970.115 ;
        RECT 3513.675 1969.835 3513.955 1970.115 ;
        RECT 3514.385 1969.835 3514.665 1970.115 ;
        RECT 3515.095 1969.835 3515.375 1970.115 ;
        RECT 3515.805 1969.835 3516.085 1970.115 ;
        RECT 3516.515 1969.835 3516.795 1970.115 ;
        RECT 3517.225 1969.835 3517.505 1970.115 ;
        RECT 3517.935 1969.835 3518.215 1970.115 ;
        RECT 3518.645 1969.835 3518.925 1970.115 ;
        RECT 3519.355 1969.835 3519.635 1970.115 ;
        RECT 3520.065 1969.835 3520.345 1970.115 ;
        RECT 3520.775 1969.835 3521.055 1970.115 ;
        RECT 3521.485 1969.835 3521.765 1970.115 ;
        RECT 3512.255 1969.125 3512.535 1969.405 ;
        RECT 3512.965 1969.125 3513.245 1969.405 ;
        RECT 3513.675 1969.125 3513.955 1969.405 ;
        RECT 3514.385 1969.125 3514.665 1969.405 ;
        RECT 3515.095 1969.125 3515.375 1969.405 ;
        RECT 3515.805 1969.125 3516.085 1969.405 ;
        RECT 3516.515 1969.125 3516.795 1969.405 ;
        RECT 3517.225 1969.125 3517.505 1969.405 ;
        RECT 3517.935 1969.125 3518.215 1969.405 ;
        RECT 3518.645 1969.125 3518.925 1969.405 ;
        RECT 3519.355 1969.125 3519.635 1969.405 ;
        RECT 3520.065 1969.125 3520.345 1969.405 ;
        RECT 3520.775 1969.125 3521.055 1969.405 ;
        RECT 3521.485 1969.125 3521.765 1969.405 ;
        RECT 3512.255 1968.415 3512.535 1968.695 ;
        RECT 3512.965 1968.415 3513.245 1968.695 ;
        RECT 3513.675 1968.415 3513.955 1968.695 ;
        RECT 3514.385 1968.415 3514.665 1968.695 ;
        RECT 3515.095 1968.415 3515.375 1968.695 ;
        RECT 3515.805 1968.415 3516.085 1968.695 ;
        RECT 3516.515 1968.415 3516.795 1968.695 ;
        RECT 3517.225 1968.415 3517.505 1968.695 ;
        RECT 3517.935 1968.415 3518.215 1968.695 ;
        RECT 3518.645 1968.415 3518.925 1968.695 ;
        RECT 3519.355 1968.415 3519.635 1968.695 ;
        RECT 3520.065 1968.415 3520.345 1968.695 ;
        RECT 3520.775 1968.415 3521.055 1968.695 ;
        RECT 3521.485 1968.415 3521.765 1968.695 ;
        RECT 3512.255 1967.705 3512.535 1967.985 ;
        RECT 3512.965 1967.705 3513.245 1967.985 ;
        RECT 3513.675 1967.705 3513.955 1967.985 ;
        RECT 3514.385 1967.705 3514.665 1967.985 ;
        RECT 3515.095 1967.705 3515.375 1967.985 ;
        RECT 3515.805 1967.705 3516.085 1967.985 ;
        RECT 3516.515 1967.705 3516.795 1967.985 ;
        RECT 3517.225 1967.705 3517.505 1967.985 ;
        RECT 3517.935 1967.705 3518.215 1967.985 ;
        RECT 3518.645 1967.705 3518.925 1967.985 ;
        RECT 3519.355 1967.705 3519.635 1967.985 ;
        RECT 3520.065 1967.705 3520.345 1967.985 ;
        RECT 3520.775 1967.705 3521.055 1967.985 ;
        RECT 3521.485 1967.705 3521.765 1967.985 ;
        RECT 3512.255 1966.995 3512.535 1967.275 ;
        RECT 3512.965 1966.995 3513.245 1967.275 ;
        RECT 3513.675 1966.995 3513.955 1967.275 ;
        RECT 3514.385 1966.995 3514.665 1967.275 ;
        RECT 3515.095 1966.995 3515.375 1967.275 ;
        RECT 3515.805 1966.995 3516.085 1967.275 ;
        RECT 3516.515 1966.995 3516.795 1967.275 ;
        RECT 3517.225 1966.995 3517.505 1967.275 ;
        RECT 3517.935 1966.995 3518.215 1967.275 ;
        RECT 3518.645 1966.995 3518.925 1967.275 ;
        RECT 3519.355 1966.995 3519.635 1967.275 ;
        RECT 3520.065 1966.995 3520.345 1967.275 ;
        RECT 3520.775 1966.995 3521.055 1967.275 ;
        RECT 3521.485 1966.995 3521.765 1967.275 ;
        RECT 3512.255 1966.285 3512.535 1966.565 ;
        RECT 3512.965 1966.285 3513.245 1966.565 ;
        RECT 3513.675 1966.285 3513.955 1966.565 ;
        RECT 3514.385 1966.285 3514.665 1966.565 ;
        RECT 3515.095 1966.285 3515.375 1966.565 ;
        RECT 3515.805 1966.285 3516.085 1966.565 ;
        RECT 3516.515 1966.285 3516.795 1966.565 ;
        RECT 3517.225 1966.285 3517.505 1966.565 ;
        RECT 3517.935 1966.285 3518.215 1966.565 ;
        RECT 3518.645 1966.285 3518.925 1966.565 ;
        RECT 3519.355 1966.285 3519.635 1966.565 ;
        RECT 3520.065 1966.285 3520.345 1966.565 ;
        RECT 3520.775 1966.285 3521.055 1966.565 ;
        RECT 3521.485 1966.285 3521.765 1966.565 ;
        RECT 3512.255 1965.575 3512.535 1965.855 ;
        RECT 3512.965 1965.575 3513.245 1965.855 ;
        RECT 3513.675 1965.575 3513.955 1965.855 ;
        RECT 3514.385 1965.575 3514.665 1965.855 ;
        RECT 3515.095 1965.575 3515.375 1965.855 ;
        RECT 3515.805 1965.575 3516.085 1965.855 ;
        RECT 3516.515 1965.575 3516.795 1965.855 ;
        RECT 3517.225 1965.575 3517.505 1965.855 ;
        RECT 3517.935 1965.575 3518.215 1965.855 ;
        RECT 3518.645 1965.575 3518.925 1965.855 ;
        RECT 3519.355 1965.575 3519.635 1965.855 ;
        RECT 3520.065 1965.575 3520.345 1965.855 ;
        RECT 3520.775 1965.575 3521.055 1965.855 ;
        RECT 3521.485 1965.575 3521.765 1965.855 ;
        RECT 3512.255 1964.865 3512.535 1965.145 ;
        RECT 3512.965 1964.865 3513.245 1965.145 ;
        RECT 3513.675 1964.865 3513.955 1965.145 ;
        RECT 3514.385 1964.865 3514.665 1965.145 ;
        RECT 3515.095 1964.865 3515.375 1965.145 ;
        RECT 3515.805 1964.865 3516.085 1965.145 ;
        RECT 3516.515 1964.865 3516.795 1965.145 ;
        RECT 3517.225 1964.865 3517.505 1965.145 ;
        RECT 3517.935 1964.865 3518.215 1965.145 ;
        RECT 3518.645 1964.865 3518.925 1965.145 ;
        RECT 3519.355 1964.865 3519.635 1965.145 ;
        RECT 3520.065 1964.865 3520.345 1965.145 ;
        RECT 3520.775 1964.865 3521.055 1965.145 ;
        RECT 3521.485 1964.865 3521.765 1965.145 ;
        RECT 3512.255 1964.155 3512.535 1964.435 ;
        RECT 3512.965 1964.155 3513.245 1964.435 ;
        RECT 3513.675 1964.155 3513.955 1964.435 ;
        RECT 3514.385 1964.155 3514.665 1964.435 ;
        RECT 3515.095 1964.155 3515.375 1964.435 ;
        RECT 3515.805 1964.155 3516.085 1964.435 ;
        RECT 3516.515 1964.155 3516.795 1964.435 ;
        RECT 3517.225 1964.155 3517.505 1964.435 ;
        RECT 3517.935 1964.155 3518.215 1964.435 ;
        RECT 3518.645 1964.155 3518.925 1964.435 ;
        RECT 3519.355 1964.155 3519.635 1964.435 ;
        RECT 3520.065 1964.155 3520.345 1964.435 ;
        RECT 3520.775 1964.155 3521.055 1964.435 ;
        RECT 3521.485 1964.155 3521.765 1964.435 ;
        RECT 3512.200 1960.270 3512.480 1960.550 ;
        RECT 3512.910 1960.270 3513.190 1960.550 ;
        RECT 3513.620 1960.270 3513.900 1960.550 ;
        RECT 3514.330 1960.270 3514.610 1960.550 ;
        RECT 3515.040 1960.270 3515.320 1960.550 ;
        RECT 3515.750 1960.270 3516.030 1960.550 ;
        RECT 3516.460 1960.270 3516.740 1960.550 ;
        RECT 3517.170 1960.270 3517.450 1960.550 ;
        RECT 3517.880 1960.270 3518.160 1960.550 ;
        RECT 3518.590 1960.270 3518.870 1960.550 ;
        RECT 3519.300 1960.270 3519.580 1960.550 ;
        RECT 3520.010 1960.270 3520.290 1960.550 ;
        RECT 3520.720 1960.270 3521.000 1960.550 ;
        RECT 3521.430 1960.270 3521.710 1960.550 ;
        RECT 3512.200 1959.560 3512.480 1959.840 ;
        RECT 3512.910 1959.560 3513.190 1959.840 ;
        RECT 3513.620 1959.560 3513.900 1959.840 ;
        RECT 3514.330 1959.560 3514.610 1959.840 ;
        RECT 3515.040 1959.560 3515.320 1959.840 ;
        RECT 3515.750 1959.560 3516.030 1959.840 ;
        RECT 3516.460 1959.560 3516.740 1959.840 ;
        RECT 3517.170 1959.560 3517.450 1959.840 ;
        RECT 3517.880 1959.560 3518.160 1959.840 ;
        RECT 3518.590 1959.560 3518.870 1959.840 ;
        RECT 3519.300 1959.560 3519.580 1959.840 ;
        RECT 3520.010 1959.560 3520.290 1959.840 ;
        RECT 3520.720 1959.560 3521.000 1959.840 ;
        RECT 3521.430 1959.560 3521.710 1959.840 ;
        RECT 3512.200 1958.850 3512.480 1959.130 ;
        RECT 3512.910 1958.850 3513.190 1959.130 ;
        RECT 3513.620 1958.850 3513.900 1959.130 ;
        RECT 3514.330 1958.850 3514.610 1959.130 ;
        RECT 3515.040 1958.850 3515.320 1959.130 ;
        RECT 3515.750 1958.850 3516.030 1959.130 ;
        RECT 3516.460 1958.850 3516.740 1959.130 ;
        RECT 3517.170 1958.850 3517.450 1959.130 ;
        RECT 3517.880 1958.850 3518.160 1959.130 ;
        RECT 3518.590 1958.850 3518.870 1959.130 ;
        RECT 3519.300 1958.850 3519.580 1959.130 ;
        RECT 3520.010 1958.850 3520.290 1959.130 ;
        RECT 3520.720 1958.850 3521.000 1959.130 ;
        RECT 3521.430 1958.850 3521.710 1959.130 ;
        RECT 3512.200 1958.140 3512.480 1958.420 ;
        RECT 3512.910 1958.140 3513.190 1958.420 ;
        RECT 3513.620 1958.140 3513.900 1958.420 ;
        RECT 3514.330 1958.140 3514.610 1958.420 ;
        RECT 3515.040 1958.140 3515.320 1958.420 ;
        RECT 3515.750 1958.140 3516.030 1958.420 ;
        RECT 3516.460 1958.140 3516.740 1958.420 ;
        RECT 3517.170 1958.140 3517.450 1958.420 ;
        RECT 3517.880 1958.140 3518.160 1958.420 ;
        RECT 3518.590 1958.140 3518.870 1958.420 ;
        RECT 3519.300 1958.140 3519.580 1958.420 ;
        RECT 3520.010 1958.140 3520.290 1958.420 ;
        RECT 3520.720 1958.140 3521.000 1958.420 ;
        RECT 3521.430 1958.140 3521.710 1958.420 ;
        RECT 3512.200 1957.430 3512.480 1957.710 ;
        RECT 3512.910 1957.430 3513.190 1957.710 ;
        RECT 3513.620 1957.430 3513.900 1957.710 ;
        RECT 3514.330 1957.430 3514.610 1957.710 ;
        RECT 3515.040 1957.430 3515.320 1957.710 ;
        RECT 3515.750 1957.430 3516.030 1957.710 ;
        RECT 3516.460 1957.430 3516.740 1957.710 ;
        RECT 3517.170 1957.430 3517.450 1957.710 ;
        RECT 3517.880 1957.430 3518.160 1957.710 ;
        RECT 3518.590 1957.430 3518.870 1957.710 ;
        RECT 3519.300 1957.430 3519.580 1957.710 ;
        RECT 3520.010 1957.430 3520.290 1957.710 ;
        RECT 3520.720 1957.430 3521.000 1957.710 ;
        RECT 3521.430 1957.430 3521.710 1957.710 ;
        RECT 3512.200 1956.720 3512.480 1957.000 ;
        RECT 3512.910 1956.720 3513.190 1957.000 ;
        RECT 3513.620 1956.720 3513.900 1957.000 ;
        RECT 3514.330 1956.720 3514.610 1957.000 ;
        RECT 3515.040 1956.720 3515.320 1957.000 ;
        RECT 3515.750 1956.720 3516.030 1957.000 ;
        RECT 3516.460 1956.720 3516.740 1957.000 ;
        RECT 3517.170 1956.720 3517.450 1957.000 ;
        RECT 3517.880 1956.720 3518.160 1957.000 ;
        RECT 3518.590 1956.720 3518.870 1957.000 ;
        RECT 3519.300 1956.720 3519.580 1957.000 ;
        RECT 3520.010 1956.720 3520.290 1957.000 ;
        RECT 3520.720 1956.720 3521.000 1957.000 ;
        RECT 3521.430 1956.720 3521.710 1957.000 ;
        RECT 3512.200 1956.010 3512.480 1956.290 ;
        RECT 3512.910 1956.010 3513.190 1956.290 ;
        RECT 3513.620 1956.010 3513.900 1956.290 ;
        RECT 3514.330 1956.010 3514.610 1956.290 ;
        RECT 3515.040 1956.010 3515.320 1956.290 ;
        RECT 3515.750 1956.010 3516.030 1956.290 ;
        RECT 3516.460 1956.010 3516.740 1956.290 ;
        RECT 3517.170 1956.010 3517.450 1956.290 ;
        RECT 3517.880 1956.010 3518.160 1956.290 ;
        RECT 3518.590 1956.010 3518.870 1956.290 ;
        RECT 3519.300 1956.010 3519.580 1956.290 ;
        RECT 3520.010 1956.010 3520.290 1956.290 ;
        RECT 3520.720 1956.010 3521.000 1956.290 ;
        RECT 3521.430 1956.010 3521.710 1956.290 ;
        RECT 3512.200 1955.300 3512.480 1955.580 ;
        RECT 3512.910 1955.300 3513.190 1955.580 ;
        RECT 3513.620 1955.300 3513.900 1955.580 ;
        RECT 3514.330 1955.300 3514.610 1955.580 ;
        RECT 3515.040 1955.300 3515.320 1955.580 ;
        RECT 3515.750 1955.300 3516.030 1955.580 ;
        RECT 3516.460 1955.300 3516.740 1955.580 ;
        RECT 3517.170 1955.300 3517.450 1955.580 ;
        RECT 3517.880 1955.300 3518.160 1955.580 ;
        RECT 3518.590 1955.300 3518.870 1955.580 ;
        RECT 3519.300 1955.300 3519.580 1955.580 ;
        RECT 3520.010 1955.300 3520.290 1955.580 ;
        RECT 3520.720 1955.300 3521.000 1955.580 ;
        RECT 3521.430 1955.300 3521.710 1955.580 ;
        RECT 3512.200 1954.590 3512.480 1954.870 ;
        RECT 3512.910 1954.590 3513.190 1954.870 ;
        RECT 3513.620 1954.590 3513.900 1954.870 ;
        RECT 3514.330 1954.590 3514.610 1954.870 ;
        RECT 3515.040 1954.590 3515.320 1954.870 ;
        RECT 3515.750 1954.590 3516.030 1954.870 ;
        RECT 3516.460 1954.590 3516.740 1954.870 ;
        RECT 3517.170 1954.590 3517.450 1954.870 ;
        RECT 3517.880 1954.590 3518.160 1954.870 ;
        RECT 3518.590 1954.590 3518.870 1954.870 ;
        RECT 3519.300 1954.590 3519.580 1954.870 ;
        RECT 3520.010 1954.590 3520.290 1954.870 ;
        RECT 3520.720 1954.590 3521.000 1954.870 ;
        RECT 3521.430 1954.590 3521.710 1954.870 ;
        RECT 3512.200 1953.880 3512.480 1954.160 ;
        RECT 3512.910 1953.880 3513.190 1954.160 ;
        RECT 3513.620 1953.880 3513.900 1954.160 ;
        RECT 3514.330 1953.880 3514.610 1954.160 ;
        RECT 3515.040 1953.880 3515.320 1954.160 ;
        RECT 3515.750 1953.880 3516.030 1954.160 ;
        RECT 3516.460 1953.880 3516.740 1954.160 ;
        RECT 3517.170 1953.880 3517.450 1954.160 ;
        RECT 3517.880 1953.880 3518.160 1954.160 ;
        RECT 3518.590 1953.880 3518.870 1954.160 ;
        RECT 3519.300 1953.880 3519.580 1954.160 ;
        RECT 3520.010 1953.880 3520.290 1954.160 ;
        RECT 3520.720 1953.880 3521.000 1954.160 ;
        RECT 3521.430 1953.880 3521.710 1954.160 ;
        RECT 3512.200 1953.170 3512.480 1953.450 ;
        RECT 3512.910 1953.170 3513.190 1953.450 ;
        RECT 3513.620 1953.170 3513.900 1953.450 ;
        RECT 3514.330 1953.170 3514.610 1953.450 ;
        RECT 3515.040 1953.170 3515.320 1953.450 ;
        RECT 3515.750 1953.170 3516.030 1953.450 ;
        RECT 3516.460 1953.170 3516.740 1953.450 ;
        RECT 3517.170 1953.170 3517.450 1953.450 ;
        RECT 3517.880 1953.170 3518.160 1953.450 ;
        RECT 3518.590 1953.170 3518.870 1953.450 ;
        RECT 3519.300 1953.170 3519.580 1953.450 ;
        RECT 3520.010 1953.170 3520.290 1953.450 ;
        RECT 3520.720 1953.170 3521.000 1953.450 ;
        RECT 3521.430 1953.170 3521.710 1953.450 ;
        RECT 3512.200 1952.460 3512.480 1952.740 ;
        RECT 3512.910 1952.460 3513.190 1952.740 ;
        RECT 3513.620 1952.460 3513.900 1952.740 ;
        RECT 3514.330 1952.460 3514.610 1952.740 ;
        RECT 3515.040 1952.460 3515.320 1952.740 ;
        RECT 3515.750 1952.460 3516.030 1952.740 ;
        RECT 3516.460 1952.460 3516.740 1952.740 ;
        RECT 3517.170 1952.460 3517.450 1952.740 ;
        RECT 3517.880 1952.460 3518.160 1952.740 ;
        RECT 3518.590 1952.460 3518.870 1952.740 ;
        RECT 3519.300 1952.460 3519.580 1952.740 ;
        RECT 3520.010 1952.460 3520.290 1952.740 ;
        RECT 3520.720 1952.460 3521.000 1952.740 ;
        RECT 3521.430 1952.460 3521.710 1952.740 ;
        RECT 3512.200 1951.750 3512.480 1952.030 ;
        RECT 3512.910 1951.750 3513.190 1952.030 ;
        RECT 3513.620 1951.750 3513.900 1952.030 ;
        RECT 3514.330 1951.750 3514.610 1952.030 ;
        RECT 3515.040 1951.750 3515.320 1952.030 ;
        RECT 3515.750 1951.750 3516.030 1952.030 ;
        RECT 3516.460 1951.750 3516.740 1952.030 ;
        RECT 3517.170 1951.750 3517.450 1952.030 ;
        RECT 3517.880 1951.750 3518.160 1952.030 ;
        RECT 3518.590 1951.750 3518.870 1952.030 ;
        RECT 3519.300 1951.750 3519.580 1952.030 ;
        RECT 3520.010 1951.750 3520.290 1952.030 ;
        RECT 3520.720 1951.750 3521.000 1952.030 ;
        RECT 3521.430 1951.750 3521.710 1952.030 ;
        RECT 369.330 702.970 369.610 703.250 ;
        RECT 370.040 702.970 370.320 703.250 ;
        RECT 370.750 702.970 371.030 703.250 ;
        RECT 371.460 702.970 371.740 703.250 ;
        RECT 372.170 702.970 372.450 703.250 ;
        RECT 372.880 702.970 373.160 703.250 ;
        RECT 373.590 702.970 373.870 703.250 ;
        RECT 374.300 702.970 374.580 703.250 ;
        RECT 375.010 702.970 375.290 703.250 ;
        RECT 375.720 702.970 376.000 703.250 ;
        RECT 376.430 702.970 376.710 703.250 ;
        RECT 369.330 702.260 369.610 702.540 ;
        RECT 370.040 702.260 370.320 702.540 ;
        RECT 370.750 702.260 371.030 702.540 ;
        RECT 371.460 702.260 371.740 702.540 ;
        RECT 372.170 702.260 372.450 702.540 ;
        RECT 372.880 702.260 373.160 702.540 ;
        RECT 373.590 702.260 373.870 702.540 ;
        RECT 374.300 702.260 374.580 702.540 ;
        RECT 375.010 702.260 375.290 702.540 ;
        RECT 375.720 702.260 376.000 702.540 ;
        RECT 376.430 702.260 376.710 702.540 ;
        RECT 369.330 701.550 369.610 701.830 ;
        RECT 370.040 701.550 370.320 701.830 ;
        RECT 370.750 701.550 371.030 701.830 ;
        RECT 371.460 701.550 371.740 701.830 ;
        RECT 372.170 701.550 372.450 701.830 ;
        RECT 372.880 701.550 373.160 701.830 ;
        RECT 373.590 701.550 373.870 701.830 ;
        RECT 374.300 701.550 374.580 701.830 ;
        RECT 375.010 701.550 375.290 701.830 ;
        RECT 375.720 701.550 376.000 701.830 ;
        RECT 376.430 701.550 376.710 701.830 ;
        RECT 369.330 700.840 369.610 701.120 ;
        RECT 370.040 700.840 370.320 701.120 ;
        RECT 370.750 700.840 371.030 701.120 ;
        RECT 371.460 700.840 371.740 701.120 ;
        RECT 372.170 700.840 372.450 701.120 ;
        RECT 372.880 700.840 373.160 701.120 ;
        RECT 373.590 700.840 373.870 701.120 ;
        RECT 374.300 700.840 374.580 701.120 ;
        RECT 375.010 700.840 375.290 701.120 ;
        RECT 375.720 700.840 376.000 701.120 ;
        RECT 376.430 700.840 376.710 701.120 ;
        RECT 369.330 700.130 369.610 700.410 ;
        RECT 370.040 700.130 370.320 700.410 ;
        RECT 370.750 700.130 371.030 700.410 ;
        RECT 371.460 700.130 371.740 700.410 ;
        RECT 372.170 700.130 372.450 700.410 ;
        RECT 372.880 700.130 373.160 700.410 ;
        RECT 373.590 700.130 373.870 700.410 ;
        RECT 374.300 700.130 374.580 700.410 ;
        RECT 375.010 700.130 375.290 700.410 ;
        RECT 375.720 700.130 376.000 700.410 ;
        RECT 376.430 700.130 376.710 700.410 ;
        RECT 369.330 699.420 369.610 699.700 ;
        RECT 370.040 699.420 370.320 699.700 ;
        RECT 370.750 699.420 371.030 699.700 ;
        RECT 371.460 699.420 371.740 699.700 ;
        RECT 372.170 699.420 372.450 699.700 ;
        RECT 372.880 699.420 373.160 699.700 ;
        RECT 373.590 699.420 373.870 699.700 ;
        RECT 374.300 699.420 374.580 699.700 ;
        RECT 375.010 699.420 375.290 699.700 ;
        RECT 375.720 699.420 376.000 699.700 ;
        RECT 376.430 699.420 376.710 699.700 ;
        RECT 369.330 698.710 369.610 698.990 ;
        RECT 370.040 698.710 370.320 698.990 ;
        RECT 370.750 698.710 371.030 698.990 ;
        RECT 371.460 698.710 371.740 698.990 ;
        RECT 372.170 698.710 372.450 698.990 ;
        RECT 372.880 698.710 373.160 698.990 ;
        RECT 373.590 698.710 373.870 698.990 ;
        RECT 374.300 698.710 374.580 698.990 ;
        RECT 375.010 698.710 375.290 698.990 ;
        RECT 375.720 698.710 376.000 698.990 ;
        RECT 376.430 698.710 376.710 698.990 ;
        RECT 369.330 698.000 369.610 698.280 ;
        RECT 370.040 698.000 370.320 698.280 ;
        RECT 370.750 698.000 371.030 698.280 ;
        RECT 371.460 698.000 371.740 698.280 ;
        RECT 372.170 698.000 372.450 698.280 ;
        RECT 372.880 698.000 373.160 698.280 ;
        RECT 373.590 698.000 373.870 698.280 ;
        RECT 374.300 698.000 374.580 698.280 ;
        RECT 375.010 698.000 375.290 698.280 ;
        RECT 375.720 698.000 376.000 698.280 ;
        RECT 376.430 698.000 376.710 698.280 ;
        RECT 369.330 697.290 369.610 697.570 ;
        RECT 370.040 697.290 370.320 697.570 ;
        RECT 370.750 697.290 371.030 697.570 ;
        RECT 371.460 697.290 371.740 697.570 ;
        RECT 372.170 697.290 372.450 697.570 ;
        RECT 372.880 697.290 373.160 697.570 ;
        RECT 373.590 697.290 373.870 697.570 ;
        RECT 374.300 697.290 374.580 697.570 ;
        RECT 375.010 697.290 375.290 697.570 ;
        RECT 375.720 697.290 376.000 697.570 ;
        RECT 376.430 697.290 376.710 697.570 ;
        RECT 369.330 696.580 369.610 696.860 ;
        RECT 370.040 696.580 370.320 696.860 ;
        RECT 370.750 696.580 371.030 696.860 ;
        RECT 371.460 696.580 371.740 696.860 ;
        RECT 372.170 696.580 372.450 696.860 ;
        RECT 372.880 696.580 373.160 696.860 ;
        RECT 373.590 696.580 373.870 696.860 ;
        RECT 374.300 696.580 374.580 696.860 ;
        RECT 375.010 696.580 375.290 696.860 ;
        RECT 375.720 696.580 376.000 696.860 ;
        RECT 376.430 696.580 376.710 696.860 ;
        RECT 369.330 695.870 369.610 696.150 ;
        RECT 370.040 695.870 370.320 696.150 ;
        RECT 370.750 695.870 371.030 696.150 ;
        RECT 371.460 695.870 371.740 696.150 ;
        RECT 372.170 695.870 372.450 696.150 ;
        RECT 372.880 695.870 373.160 696.150 ;
        RECT 373.590 695.870 373.870 696.150 ;
        RECT 374.300 695.870 374.580 696.150 ;
        RECT 375.010 695.870 375.290 696.150 ;
        RECT 375.720 695.870 376.000 696.150 ;
        RECT 376.430 695.870 376.710 696.150 ;
        RECT 369.330 695.160 369.610 695.440 ;
        RECT 370.040 695.160 370.320 695.440 ;
        RECT 370.750 695.160 371.030 695.440 ;
        RECT 371.460 695.160 371.740 695.440 ;
        RECT 372.170 695.160 372.450 695.440 ;
        RECT 372.880 695.160 373.160 695.440 ;
        RECT 373.590 695.160 373.870 695.440 ;
        RECT 374.300 695.160 374.580 695.440 ;
        RECT 375.010 695.160 375.290 695.440 ;
        RECT 375.720 695.160 376.000 695.440 ;
        RECT 376.430 695.160 376.710 695.440 ;
        RECT 369.330 694.450 369.610 694.730 ;
        RECT 370.040 694.450 370.320 694.730 ;
        RECT 370.750 694.450 371.030 694.730 ;
        RECT 371.460 694.450 371.740 694.730 ;
        RECT 372.170 694.450 372.450 694.730 ;
        RECT 372.880 694.450 373.160 694.730 ;
        RECT 373.590 694.450 373.870 694.730 ;
        RECT 374.300 694.450 374.580 694.730 ;
        RECT 375.010 694.450 375.290 694.730 ;
        RECT 375.720 694.450 376.000 694.730 ;
        RECT 376.430 694.450 376.710 694.730 ;
        RECT 369.275 690.565 369.555 690.845 ;
        RECT 369.985 690.565 370.265 690.845 ;
        RECT 370.695 690.565 370.975 690.845 ;
        RECT 371.405 690.565 371.685 690.845 ;
        RECT 372.115 690.565 372.395 690.845 ;
        RECT 372.825 690.565 373.105 690.845 ;
        RECT 373.535 690.565 373.815 690.845 ;
        RECT 374.245 690.565 374.525 690.845 ;
        RECT 374.955 690.565 375.235 690.845 ;
        RECT 375.665 690.565 375.945 690.845 ;
        RECT 376.375 690.565 376.655 690.845 ;
        RECT 369.275 689.855 369.555 690.135 ;
        RECT 369.985 689.855 370.265 690.135 ;
        RECT 370.695 689.855 370.975 690.135 ;
        RECT 371.405 689.855 371.685 690.135 ;
        RECT 372.115 689.855 372.395 690.135 ;
        RECT 372.825 689.855 373.105 690.135 ;
        RECT 373.535 689.855 373.815 690.135 ;
        RECT 374.245 689.855 374.525 690.135 ;
        RECT 374.955 689.855 375.235 690.135 ;
        RECT 375.665 689.855 375.945 690.135 ;
        RECT 376.375 689.855 376.655 690.135 ;
        RECT 369.275 689.145 369.555 689.425 ;
        RECT 369.985 689.145 370.265 689.425 ;
        RECT 370.695 689.145 370.975 689.425 ;
        RECT 371.405 689.145 371.685 689.425 ;
        RECT 372.115 689.145 372.395 689.425 ;
        RECT 372.825 689.145 373.105 689.425 ;
        RECT 373.535 689.145 373.815 689.425 ;
        RECT 374.245 689.145 374.525 689.425 ;
        RECT 374.955 689.145 375.235 689.425 ;
        RECT 375.665 689.145 375.945 689.425 ;
        RECT 376.375 689.145 376.655 689.425 ;
        RECT 369.275 688.435 369.555 688.715 ;
        RECT 369.985 688.435 370.265 688.715 ;
        RECT 370.695 688.435 370.975 688.715 ;
        RECT 371.405 688.435 371.685 688.715 ;
        RECT 372.115 688.435 372.395 688.715 ;
        RECT 372.825 688.435 373.105 688.715 ;
        RECT 373.535 688.435 373.815 688.715 ;
        RECT 374.245 688.435 374.525 688.715 ;
        RECT 374.955 688.435 375.235 688.715 ;
        RECT 375.665 688.435 375.945 688.715 ;
        RECT 376.375 688.435 376.655 688.715 ;
        RECT 369.275 687.725 369.555 688.005 ;
        RECT 369.985 687.725 370.265 688.005 ;
        RECT 370.695 687.725 370.975 688.005 ;
        RECT 371.405 687.725 371.685 688.005 ;
        RECT 372.115 687.725 372.395 688.005 ;
        RECT 372.825 687.725 373.105 688.005 ;
        RECT 373.535 687.725 373.815 688.005 ;
        RECT 374.245 687.725 374.525 688.005 ;
        RECT 374.955 687.725 375.235 688.005 ;
        RECT 375.665 687.725 375.945 688.005 ;
        RECT 376.375 687.725 376.655 688.005 ;
        RECT 369.275 687.015 369.555 687.295 ;
        RECT 369.985 687.015 370.265 687.295 ;
        RECT 370.695 687.015 370.975 687.295 ;
        RECT 371.405 687.015 371.685 687.295 ;
        RECT 372.115 687.015 372.395 687.295 ;
        RECT 372.825 687.015 373.105 687.295 ;
        RECT 373.535 687.015 373.815 687.295 ;
        RECT 374.245 687.015 374.525 687.295 ;
        RECT 374.955 687.015 375.235 687.295 ;
        RECT 375.665 687.015 375.945 687.295 ;
        RECT 376.375 687.015 376.655 687.295 ;
        RECT 369.275 686.305 369.555 686.585 ;
        RECT 369.985 686.305 370.265 686.585 ;
        RECT 370.695 686.305 370.975 686.585 ;
        RECT 371.405 686.305 371.685 686.585 ;
        RECT 372.115 686.305 372.395 686.585 ;
        RECT 372.825 686.305 373.105 686.585 ;
        RECT 373.535 686.305 373.815 686.585 ;
        RECT 374.245 686.305 374.525 686.585 ;
        RECT 374.955 686.305 375.235 686.585 ;
        RECT 375.665 686.305 375.945 686.585 ;
        RECT 376.375 686.305 376.655 686.585 ;
        RECT 369.275 685.595 369.555 685.875 ;
        RECT 369.985 685.595 370.265 685.875 ;
        RECT 370.695 685.595 370.975 685.875 ;
        RECT 371.405 685.595 371.685 685.875 ;
        RECT 372.115 685.595 372.395 685.875 ;
        RECT 372.825 685.595 373.105 685.875 ;
        RECT 373.535 685.595 373.815 685.875 ;
        RECT 374.245 685.595 374.525 685.875 ;
        RECT 374.955 685.595 375.235 685.875 ;
        RECT 375.665 685.595 375.945 685.875 ;
        RECT 376.375 685.595 376.655 685.875 ;
        RECT 369.275 684.885 369.555 685.165 ;
        RECT 369.985 684.885 370.265 685.165 ;
        RECT 370.695 684.885 370.975 685.165 ;
        RECT 371.405 684.885 371.685 685.165 ;
        RECT 372.115 684.885 372.395 685.165 ;
        RECT 372.825 684.885 373.105 685.165 ;
        RECT 373.535 684.885 373.815 685.165 ;
        RECT 374.245 684.885 374.525 685.165 ;
        RECT 374.955 684.885 375.235 685.165 ;
        RECT 375.665 684.885 375.945 685.165 ;
        RECT 376.375 684.885 376.655 685.165 ;
        RECT 369.275 684.175 369.555 684.455 ;
        RECT 369.985 684.175 370.265 684.455 ;
        RECT 370.695 684.175 370.975 684.455 ;
        RECT 371.405 684.175 371.685 684.455 ;
        RECT 372.115 684.175 372.395 684.455 ;
        RECT 372.825 684.175 373.105 684.455 ;
        RECT 373.535 684.175 373.815 684.455 ;
        RECT 374.245 684.175 374.525 684.455 ;
        RECT 374.955 684.175 375.235 684.455 ;
        RECT 375.665 684.175 375.945 684.455 ;
        RECT 376.375 684.175 376.655 684.455 ;
        RECT 369.275 683.465 369.555 683.745 ;
        RECT 369.985 683.465 370.265 683.745 ;
        RECT 370.695 683.465 370.975 683.745 ;
        RECT 371.405 683.465 371.685 683.745 ;
        RECT 372.115 683.465 372.395 683.745 ;
        RECT 372.825 683.465 373.105 683.745 ;
        RECT 373.535 683.465 373.815 683.745 ;
        RECT 374.245 683.465 374.525 683.745 ;
        RECT 374.955 683.465 375.235 683.745 ;
        RECT 375.665 683.465 375.945 683.745 ;
        RECT 376.375 683.465 376.655 683.745 ;
        RECT 369.275 682.755 369.555 683.035 ;
        RECT 369.985 682.755 370.265 683.035 ;
        RECT 370.695 682.755 370.975 683.035 ;
        RECT 371.405 682.755 371.685 683.035 ;
        RECT 372.115 682.755 372.395 683.035 ;
        RECT 372.825 682.755 373.105 683.035 ;
        RECT 373.535 682.755 373.815 683.035 ;
        RECT 374.245 682.755 374.525 683.035 ;
        RECT 374.955 682.755 375.235 683.035 ;
        RECT 375.665 682.755 375.945 683.035 ;
        RECT 376.375 682.755 376.655 683.035 ;
        RECT 369.275 682.045 369.555 682.325 ;
        RECT 369.985 682.045 370.265 682.325 ;
        RECT 370.695 682.045 370.975 682.325 ;
        RECT 371.405 682.045 371.685 682.325 ;
        RECT 372.115 682.045 372.395 682.325 ;
        RECT 372.825 682.045 373.105 682.325 ;
        RECT 373.535 682.045 373.815 682.325 ;
        RECT 374.245 682.045 374.525 682.325 ;
        RECT 374.955 682.045 375.235 682.325 ;
        RECT 375.665 682.045 375.945 682.325 ;
        RECT 376.375 682.045 376.655 682.325 ;
        RECT 369.275 681.335 369.555 681.615 ;
        RECT 369.985 681.335 370.265 681.615 ;
        RECT 370.695 681.335 370.975 681.615 ;
        RECT 371.405 681.335 371.685 681.615 ;
        RECT 372.115 681.335 372.395 681.615 ;
        RECT 372.825 681.335 373.105 681.615 ;
        RECT 373.535 681.335 373.815 681.615 ;
        RECT 374.245 681.335 374.525 681.615 ;
        RECT 374.955 681.335 375.235 681.615 ;
        RECT 375.665 681.335 375.945 681.615 ;
        RECT 376.375 681.335 376.655 681.615 ;
        RECT 369.275 678.715 369.555 678.995 ;
        RECT 369.985 678.715 370.265 678.995 ;
        RECT 370.695 678.715 370.975 678.995 ;
        RECT 371.405 678.715 371.685 678.995 ;
        RECT 372.115 678.715 372.395 678.995 ;
        RECT 372.825 678.715 373.105 678.995 ;
        RECT 373.535 678.715 373.815 678.995 ;
        RECT 374.245 678.715 374.525 678.995 ;
        RECT 374.955 678.715 375.235 678.995 ;
        RECT 375.665 678.715 375.945 678.995 ;
        RECT 376.375 678.715 376.655 678.995 ;
        RECT 369.275 678.005 369.555 678.285 ;
        RECT 369.985 678.005 370.265 678.285 ;
        RECT 370.695 678.005 370.975 678.285 ;
        RECT 371.405 678.005 371.685 678.285 ;
        RECT 372.115 678.005 372.395 678.285 ;
        RECT 372.825 678.005 373.105 678.285 ;
        RECT 373.535 678.005 373.815 678.285 ;
        RECT 374.245 678.005 374.525 678.285 ;
        RECT 374.955 678.005 375.235 678.285 ;
        RECT 375.665 678.005 375.945 678.285 ;
        RECT 376.375 678.005 376.655 678.285 ;
        RECT 369.275 677.295 369.555 677.575 ;
        RECT 369.985 677.295 370.265 677.575 ;
        RECT 370.695 677.295 370.975 677.575 ;
        RECT 371.405 677.295 371.685 677.575 ;
        RECT 372.115 677.295 372.395 677.575 ;
        RECT 372.825 677.295 373.105 677.575 ;
        RECT 373.535 677.295 373.815 677.575 ;
        RECT 374.245 677.295 374.525 677.575 ;
        RECT 374.955 677.295 375.235 677.575 ;
        RECT 375.665 677.295 375.945 677.575 ;
        RECT 376.375 677.295 376.655 677.575 ;
        RECT 369.275 676.585 369.555 676.865 ;
        RECT 369.985 676.585 370.265 676.865 ;
        RECT 370.695 676.585 370.975 676.865 ;
        RECT 371.405 676.585 371.685 676.865 ;
        RECT 372.115 676.585 372.395 676.865 ;
        RECT 372.825 676.585 373.105 676.865 ;
        RECT 373.535 676.585 373.815 676.865 ;
        RECT 374.245 676.585 374.525 676.865 ;
        RECT 374.955 676.585 375.235 676.865 ;
        RECT 375.665 676.585 375.945 676.865 ;
        RECT 376.375 676.585 376.655 676.865 ;
        RECT 369.275 675.875 369.555 676.155 ;
        RECT 369.985 675.875 370.265 676.155 ;
        RECT 370.695 675.875 370.975 676.155 ;
        RECT 371.405 675.875 371.685 676.155 ;
        RECT 372.115 675.875 372.395 676.155 ;
        RECT 372.825 675.875 373.105 676.155 ;
        RECT 373.535 675.875 373.815 676.155 ;
        RECT 374.245 675.875 374.525 676.155 ;
        RECT 374.955 675.875 375.235 676.155 ;
        RECT 375.665 675.875 375.945 676.155 ;
        RECT 376.375 675.875 376.655 676.155 ;
        RECT 369.275 675.165 369.555 675.445 ;
        RECT 369.985 675.165 370.265 675.445 ;
        RECT 370.695 675.165 370.975 675.445 ;
        RECT 371.405 675.165 371.685 675.445 ;
        RECT 372.115 675.165 372.395 675.445 ;
        RECT 372.825 675.165 373.105 675.445 ;
        RECT 373.535 675.165 373.815 675.445 ;
        RECT 374.245 675.165 374.525 675.445 ;
        RECT 374.955 675.165 375.235 675.445 ;
        RECT 375.665 675.165 375.945 675.445 ;
        RECT 376.375 675.165 376.655 675.445 ;
        RECT 369.275 674.455 369.555 674.735 ;
        RECT 369.985 674.455 370.265 674.735 ;
        RECT 370.695 674.455 370.975 674.735 ;
        RECT 371.405 674.455 371.685 674.735 ;
        RECT 372.115 674.455 372.395 674.735 ;
        RECT 372.825 674.455 373.105 674.735 ;
        RECT 373.535 674.455 373.815 674.735 ;
        RECT 374.245 674.455 374.525 674.735 ;
        RECT 374.955 674.455 375.235 674.735 ;
        RECT 375.665 674.455 375.945 674.735 ;
        RECT 376.375 674.455 376.655 674.735 ;
        RECT 369.275 673.745 369.555 674.025 ;
        RECT 369.985 673.745 370.265 674.025 ;
        RECT 370.695 673.745 370.975 674.025 ;
        RECT 371.405 673.745 371.685 674.025 ;
        RECT 372.115 673.745 372.395 674.025 ;
        RECT 372.825 673.745 373.105 674.025 ;
        RECT 373.535 673.745 373.815 674.025 ;
        RECT 374.245 673.745 374.525 674.025 ;
        RECT 374.955 673.745 375.235 674.025 ;
        RECT 375.665 673.745 375.945 674.025 ;
        RECT 376.375 673.745 376.655 674.025 ;
        RECT 369.275 673.035 369.555 673.315 ;
        RECT 369.985 673.035 370.265 673.315 ;
        RECT 370.695 673.035 370.975 673.315 ;
        RECT 371.405 673.035 371.685 673.315 ;
        RECT 372.115 673.035 372.395 673.315 ;
        RECT 372.825 673.035 373.105 673.315 ;
        RECT 373.535 673.035 373.815 673.315 ;
        RECT 374.245 673.035 374.525 673.315 ;
        RECT 374.955 673.035 375.235 673.315 ;
        RECT 375.665 673.035 375.945 673.315 ;
        RECT 376.375 673.035 376.655 673.315 ;
        RECT 369.275 672.325 369.555 672.605 ;
        RECT 369.985 672.325 370.265 672.605 ;
        RECT 370.695 672.325 370.975 672.605 ;
        RECT 371.405 672.325 371.685 672.605 ;
        RECT 372.115 672.325 372.395 672.605 ;
        RECT 372.825 672.325 373.105 672.605 ;
        RECT 373.535 672.325 373.815 672.605 ;
        RECT 374.245 672.325 374.525 672.605 ;
        RECT 374.955 672.325 375.235 672.605 ;
        RECT 375.665 672.325 375.945 672.605 ;
        RECT 376.375 672.325 376.655 672.605 ;
        RECT 369.275 671.615 369.555 671.895 ;
        RECT 369.985 671.615 370.265 671.895 ;
        RECT 370.695 671.615 370.975 671.895 ;
        RECT 371.405 671.615 371.685 671.895 ;
        RECT 372.115 671.615 372.395 671.895 ;
        RECT 372.825 671.615 373.105 671.895 ;
        RECT 373.535 671.615 373.815 671.895 ;
        RECT 374.245 671.615 374.525 671.895 ;
        RECT 374.955 671.615 375.235 671.895 ;
        RECT 375.665 671.615 375.945 671.895 ;
        RECT 376.375 671.615 376.655 671.895 ;
        RECT 369.275 670.905 369.555 671.185 ;
        RECT 369.985 670.905 370.265 671.185 ;
        RECT 370.695 670.905 370.975 671.185 ;
        RECT 371.405 670.905 371.685 671.185 ;
        RECT 372.115 670.905 372.395 671.185 ;
        RECT 372.825 670.905 373.105 671.185 ;
        RECT 373.535 670.905 373.815 671.185 ;
        RECT 374.245 670.905 374.525 671.185 ;
        RECT 374.955 670.905 375.235 671.185 ;
        RECT 375.665 670.905 375.945 671.185 ;
        RECT 376.375 670.905 376.655 671.185 ;
        RECT 369.275 670.195 369.555 670.475 ;
        RECT 369.985 670.195 370.265 670.475 ;
        RECT 370.695 670.195 370.975 670.475 ;
        RECT 371.405 670.195 371.685 670.475 ;
        RECT 372.115 670.195 372.395 670.475 ;
        RECT 372.825 670.195 373.105 670.475 ;
        RECT 373.535 670.195 373.815 670.475 ;
        RECT 374.245 670.195 374.525 670.475 ;
        RECT 374.955 670.195 375.235 670.475 ;
        RECT 375.665 670.195 375.945 670.475 ;
        RECT 376.375 670.195 376.655 670.475 ;
        RECT 369.275 669.485 369.555 669.765 ;
        RECT 369.985 669.485 370.265 669.765 ;
        RECT 370.695 669.485 370.975 669.765 ;
        RECT 371.405 669.485 371.685 669.765 ;
        RECT 372.115 669.485 372.395 669.765 ;
        RECT 372.825 669.485 373.105 669.765 ;
        RECT 373.535 669.485 373.815 669.765 ;
        RECT 374.245 669.485 374.525 669.765 ;
        RECT 374.955 669.485 375.235 669.765 ;
        RECT 375.665 669.485 375.945 669.765 ;
        RECT 376.375 669.485 376.655 669.765 ;
        RECT 369.275 665.185 369.555 665.465 ;
        RECT 369.985 665.185 370.265 665.465 ;
        RECT 370.695 665.185 370.975 665.465 ;
        RECT 371.405 665.185 371.685 665.465 ;
        RECT 372.115 665.185 372.395 665.465 ;
        RECT 372.825 665.185 373.105 665.465 ;
        RECT 373.535 665.185 373.815 665.465 ;
        RECT 374.245 665.185 374.525 665.465 ;
        RECT 374.955 665.185 375.235 665.465 ;
        RECT 375.665 665.185 375.945 665.465 ;
        RECT 376.375 665.185 376.655 665.465 ;
        RECT 369.275 664.475 369.555 664.755 ;
        RECT 369.985 664.475 370.265 664.755 ;
        RECT 370.695 664.475 370.975 664.755 ;
        RECT 371.405 664.475 371.685 664.755 ;
        RECT 372.115 664.475 372.395 664.755 ;
        RECT 372.825 664.475 373.105 664.755 ;
        RECT 373.535 664.475 373.815 664.755 ;
        RECT 374.245 664.475 374.525 664.755 ;
        RECT 374.955 664.475 375.235 664.755 ;
        RECT 375.665 664.475 375.945 664.755 ;
        RECT 376.375 664.475 376.655 664.755 ;
        RECT 369.275 663.765 369.555 664.045 ;
        RECT 369.985 663.765 370.265 664.045 ;
        RECT 370.695 663.765 370.975 664.045 ;
        RECT 371.405 663.765 371.685 664.045 ;
        RECT 372.115 663.765 372.395 664.045 ;
        RECT 372.825 663.765 373.105 664.045 ;
        RECT 373.535 663.765 373.815 664.045 ;
        RECT 374.245 663.765 374.525 664.045 ;
        RECT 374.955 663.765 375.235 664.045 ;
        RECT 375.665 663.765 375.945 664.045 ;
        RECT 376.375 663.765 376.655 664.045 ;
        RECT 369.275 663.055 369.555 663.335 ;
        RECT 369.985 663.055 370.265 663.335 ;
        RECT 370.695 663.055 370.975 663.335 ;
        RECT 371.405 663.055 371.685 663.335 ;
        RECT 372.115 663.055 372.395 663.335 ;
        RECT 372.825 663.055 373.105 663.335 ;
        RECT 373.535 663.055 373.815 663.335 ;
        RECT 374.245 663.055 374.525 663.335 ;
        RECT 374.955 663.055 375.235 663.335 ;
        RECT 375.665 663.055 375.945 663.335 ;
        RECT 376.375 663.055 376.655 663.335 ;
        RECT 369.275 662.345 369.555 662.625 ;
        RECT 369.985 662.345 370.265 662.625 ;
        RECT 370.695 662.345 370.975 662.625 ;
        RECT 371.405 662.345 371.685 662.625 ;
        RECT 372.115 662.345 372.395 662.625 ;
        RECT 372.825 662.345 373.105 662.625 ;
        RECT 373.535 662.345 373.815 662.625 ;
        RECT 374.245 662.345 374.525 662.625 ;
        RECT 374.955 662.345 375.235 662.625 ;
        RECT 375.665 662.345 375.945 662.625 ;
        RECT 376.375 662.345 376.655 662.625 ;
        RECT 369.275 661.635 369.555 661.915 ;
        RECT 369.985 661.635 370.265 661.915 ;
        RECT 370.695 661.635 370.975 661.915 ;
        RECT 371.405 661.635 371.685 661.915 ;
        RECT 372.115 661.635 372.395 661.915 ;
        RECT 372.825 661.635 373.105 661.915 ;
        RECT 373.535 661.635 373.815 661.915 ;
        RECT 374.245 661.635 374.525 661.915 ;
        RECT 374.955 661.635 375.235 661.915 ;
        RECT 375.665 661.635 375.945 661.915 ;
        RECT 376.375 661.635 376.655 661.915 ;
        RECT 369.275 660.925 369.555 661.205 ;
        RECT 369.985 660.925 370.265 661.205 ;
        RECT 370.695 660.925 370.975 661.205 ;
        RECT 371.405 660.925 371.685 661.205 ;
        RECT 372.115 660.925 372.395 661.205 ;
        RECT 372.825 660.925 373.105 661.205 ;
        RECT 373.535 660.925 373.815 661.205 ;
        RECT 374.245 660.925 374.525 661.205 ;
        RECT 374.955 660.925 375.235 661.205 ;
        RECT 375.665 660.925 375.945 661.205 ;
        RECT 376.375 660.925 376.655 661.205 ;
        RECT 369.275 660.215 369.555 660.495 ;
        RECT 369.985 660.215 370.265 660.495 ;
        RECT 370.695 660.215 370.975 660.495 ;
        RECT 371.405 660.215 371.685 660.495 ;
        RECT 372.115 660.215 372.395 660.495 ;
        RECT 372.825 660.215 373.105 660.495 ;
        RECT 373.535 660.215 373.815 660.495 ;
        RECT 374.245 660.215 374.525 660.495 ;
        RECT 374.955 660.215 375.235 660.495 ;
        RECT 375.665 660.215 375.945 660.495 ;
        RECT 376.375 660.215 376.655 660.495 ;
        RECT 369.275 659.505 369.555 659.785 ;
        RECT 369.985 659.505 370.265 659.785 ;
        RECT 370.695 659.505 370.975 659.785 ;
        RECT 371.405 659.505 371.685 659.785 ;
        RECT 372.115 659.505 372.395 659.785 ;
        RECT 372.825 659.505 373.105 659.785 ;
        RECT 373.535 659.505 373.815 659.785 ;
        RECT 374.245 659.505 374.525 659.785 ;
        RECT 374.955 659.505 375.235 659.785 ;
        RECT 375.665 659.505 375.945 659.785 ;
        RECT 376.375 659.505 376.655 659.785 ;
        RECT 369.275 658.795 369.555 659.075 ;
        RECT 369.985 658.795 370.265 659.075 ;
        RECT 370.695 658.795 370.975 659.075 ;
        RECT 371.405 658.795 371.685 659.075 ;
        RECT 372.115 658.795 372.395 659.075 ;
        RECT 372.825 658.795 373.105 659.075 ;
        RECT 373.535 658.795 373.815 659.075 ;
        RECT 374.245 658.795 374.525 659.075 ;
        RECT 374.955 658.795 375.235 659.075 ;
        RECT 375.665 658.795 375.945 659.075 ;
        RECT 376.375 658.795 376.655 659.075 ;
        RECT 369.275 658.085 369.555 658.365 ;
        RECT 369.985 658.085 370.265 658.365 ;
        RECT 370.695 658.085 370.975 658.365 ;
        RECT 371.405 658.085 371.685 658.365 ;
        RECT 372.115 658.085 372.395 658.365 ;
        RECT 372.825 658.085 373.105 658.365 ;
        RECT 373.535 658.085 373.815 658.365 ;
        RECT 374.245 658.085 374.525 658.365 ;
        RECT 374.955 658.085 375.235 658.365 ;
        RECT 375.665 658.085 375.945 658.365 ;
        RECT 376.375 658.085 376.655 658.365 ;
        RECT 369.275 657.375 369.555 657.655 ;
        RECT 369.985 657.375 370.265 657.655 ;
        RECT 370.695 657.375 370.975 657.655 ;
        RECT 371.405 657.375 371.685 657.655 ;
        RECT 372.115 657.375 372.395 657.655 ;
        RECT 372.825 657.375 373.105 657.655 ;
        RECT 373.535 657.375 373.815 657.655 ;
        RECT 374.245 657.375 374.525 657.655 ;
        RECT 374.955 657.375 375.235 657.655 ;
        RECT 375.665 657.375 375.945 657.655 ;
        RECT 376.375 657.375 376.655 657.655 ;
        RECT 369.275 656.665 369.555 656.945 ;
        RECT 369.985 656.665 370.265 656.945 ;
        RECT 370.695 656.665 370.975 656.945 ;
        RECT 371.405 656.665 371.685 656.945 ;
        RECT 372.115 656.665 372.395 656.945 ;
        RECT 372.825 656.665 373.105 656.945 ;
        RECT 373.535 656.665 373.815 656.945 ;
        RECT 374.245 656.665 374.525 656.945 ;
        RECT 374.955 656.665 375.235 656.945 ;
        RECT 375.665 656.665 375.945 656.945 ;
        RECT 376.375 656.665 376.655 656.945 ;
        RECT 369.275 655.955 369.555 656.235 ;
        RECT 369.985 655.955 370.265 656.235 ;
        RECT 370.695 655.955 370.975 656.235 ;
        RECT 371.405 655.955 371.685 656.235 ;
        RECT 372.115 655.955 372.395 656.235 ;
        RECT 372.825 655.955 373.105 656.235 ;
        RECT 373.535 655.955 373.815 656.235 ;
        RECT 374.245 655.955 374.525 656.235 ;
        RECT 374.955 655.955 375.235 656.235 ;
        RECT 375.665 655.955 375.945 656.235 ;
        RECT 376.375 655.955 376.655 656.235 ;
        RECT 369.275 653.335 369.555 653.615 ;
        RECT 369.985 653.335 370.265 653.615 ;
        RECT 370.695 653.335 370.975 653.615 ;
        RECT 371.405 653.335 371.685 653.615 ;
        RECT 372.115 653.335 372.395 653.615 ;
        RECT 372.825 653.335 373.105 653.615 ;
        RECT 373.535 653.335 373.815 653.615 ;
        RECT 374.245 653.335 374.525 653.615 ;
        RECT 374.955 653.335 375.235 653.615 ;
        RECT 375.665 653.335 375.945 653.615 ;
        RECT 376.375 653.335 376.655 653.615 ;
        RECT 369.275 652.625 369.555 652.905 ;
        RECT 369.985 652.625 370.265 652.905 ;
        RECT 370.695 652.625 370.975 652.905 ;
        RECT 371.405 652.625 371.685 652.905 ;
        RECT 372.115 652.625 372.395 652.905 ;
        RECT 372.825 652.625 373.105 652.905 ;
        RECT 373.535 652.625 373.815 652.905 ;
        RECT 374.245 652.625 374.525 652.905 ;
        RECT 374.955 652.625 375.235 652.905 ;
        RECT 375.665 652.625 375.945 652.905 ;
        RECT 376.375 652.625 376.655 652.905 ;
        RECT 369.275 651.915 369.555 652.195 ;
        RECT 369.985 651.915 370.265 652.195 ;
        RECT 370.695 651.915 370.975 652.195 ;
        RECT 371.405 651.915 371.685 652.195 ;
        RECT 372.115 651.915 372.395 652.195 ;
        RECT 372.825 651.915 373.105 652.195 ;
        RECT 373.535 651.915 373.815 652.195 ;
        RECT 374.245 651.915 374.525 652.195 ;
        RECT 374.955 651.915 375.235 652.195 ;
        RECT 375.665 651.915 375.945 652.195 ;
        RECT 376.375 651.915 376.655 652.195 ;
        RECT 369.275 651.205 369.555 651.485 ;
        RECT 369.985 651.205 370.265 651.485 ;
        RECT 370.695 651.205 370.975 651.485 ;
        RECT 371.405 651.205 371.685 651.485 ;
        RECT 372.115 651.205 372.395 651.485 ;
        RECT 372.825 651.205 373.105 651.485 ;
        RECT 373.535 651.205 373.815 651.485 ;
        RECT 374.245 651.205 374.525 651.485 ;
        RECT 374.955 651.205 375.235 651.485 ;
        RECT 375.665 651.205 375.945 651.485 ;
        RECT 376.375 651.205 376.655 651.485 ;
        RECT 369.275 650.495 369.555 650.775 ;
        RECT 369.985 650.495 370.265 650.775 ;
        RECT 370.695 650.495 370.975 650.775 ;
        RECT 371.405 650.495 371.685 650.775 ;
        RECT 372.115 650.495 372.395 650.775 ;
        RECT 372.825 650.495 373.105 650.775 ;
        RECT 373.535 650.495 373.815 650.775 ;
        RECT 374.245 650.495 374.525 650.775 ;
        RECT 374.955 650.495 375.235 650.775 ;
        RECT 375.665 650.495 375.945 650.775 ;
        RECT 376.375 650.495 376.655 650.775 ;
        RECT 369.275 649.785 369.555 650.065 ;
        RECT 369.985 649.785 370.265 650.065 ;
        RECT 370.695 649.785 370.975 650.065 ;
        RECT 371.405 649.785 371.685 650.065 ;
        RECT 372.115 649.785 372.395 650.065 ;
        RECT 372.825 649.785 373.105 650.065 ;
        RECT 373.535 649.785 373.815 650.065 ;
        RECT 374.245 649.785 374.525 650.065 ;
        RECT 374.955 649.785 375.235 650.065 ;
        RECT 375.665 649.785 375.945 650.065 ;
        RECT 376.375 649.785 376.655 650.065 ;
        RECT 369.275 649.075 369.555 649.355 ;
        RECT 369.985 649.075 370.265 649.355 ;
        RECT 370.695 649.075 370.975 649.355 ;
        RECT 371.405 649.075 371.685 649.355 ;
        RECT 372.115 649.075 372.395 649.355 ;
        RECT 372.825 649.075 373.105 649.355 ;
        RECT 373.535 649.075 373.815 649.355 ;
        RECT 374.245 649.075 374.525 649.355 ;
        RECT 374.955 649.075 375.235 649.355 ;
        RECT 375.665 649.075 375.945 649.355 ;
        RECT 376.375 649.075 376.655 649.355 ;
        RECT 369.275 648.365 369.555 648.645 ;
        RECT 369.985 648.365 370.265 648.645 ;
        RECT 370.695 648.365 370.975 648.645 ;
        RECT 371.405 648.365 371.685 648.645 ;
        RECT 372.115 648.365 372.395 648.645 ;
        RECT 372.825 648.365 373.105 648.645 ;
        RECT 373.535 648.365 373.815 648.645 ;
        RECT 374.245 648.365 374.525 648.645 ;
        RECT 374.955 648.365 375.235 648.645 ;
        RECT 375.665 648.365 375.945 648.645 ;
        RECT 376.375 648.365 376.655 648.645 ;
        RECT 369.275 647.655 369.555 647.935 ;
        RECT 369.985 647.655 370.265 647.935 ;
        RECT 370.695 647.655 370.975 647.935 ;
        RECT 371.405 647.655 371.685 647.935 ;
        RECT 372.115 647.655 372.395 647.935 ;
        RECT 372.825 647.655 373.105 647.935 ;
        RECT 373.535 647.655 373.815 647.935 ;
        RECT 374.245 647.655 374.525 647.935 ;
        RECT 374.955 647.655 375.235 647.935 ;
        RECT 375.665 647.655 375.945 647.935 ;
        RECT 376.375 647.655 376.655 647.935 ;
        RECT 369.275 646.945 369.555 647.225 ;
        RECT 369.985 646.945 370.265 647.225 ;
        RECT 370.695 646.945 370.975 647.225 ;
        RECT 371.405 646.945 371.685 647.225 ;
        RECT 372.115 646.945 372.395 647.225 ;
        RECT 372.825 646.945 373.105 647.225 ;
        RECT 373.535 646.945 373.815 647.225 ;
        RECT 374.245 646.945 374.525 647.225 ;
        RECT 374.955 646.945 375.235 647.225 ;
        RECT 375.665 646.945 375.945 647.225 ;
        RECT 376.375 646.945 376.655 647.225 ;
        RECT 369.275 646.235 369.555 646.515 ;
        RECT 369.985 646.235 370.265 646.515 ;
        RECT 370.695 646.235 370.975 646.515 ;
        RECT 371.405 646.235 371.685 646.515 ;
        RECT 372.115 646.235 372.395 646.515 ;
        RECT 372.825 646.235 373.105 646.515 ;
        RECT 373.535 646.235 373.815 646.515 ;
        RECT 374.245 646.235 374.525 646.515 ;
        RECT 374.955 646.235 375.235 646.515 ;
        RECT 375.665 646.235 375.945 646.515 ;
        RECT 376.375 646.235 376.655 646.515 ;
        RECT 369.275 645.525 369.555 645.805 ;
        RECT 369.985 645.525 370.265 645.805 ;
        RECT 370.695 645.525 370.975 645.805 ;
        RECT 371.405 645.525 371.685 645.805 ;
        RECT 372.115 645.525 372.395 645.805 ;
        RECT 372.825 645.525 373.105 645.805 ;
        RECT 373.535 645.525 373.815 645.805 ;
        RECT 374.245 645.525 374.525 645.805 ;
        RECT 374.955 645.525 375.235 645.805 ;
        RECT 375.665 645.525 375.945 645.805 ;
        RECT 376.375 645.525 376.655 645.805 ;
        RECT 369.275 644.815 369.555 645.095 ;
        RECT 369.985 644.815 370.265 645.095 ;
        RECT 370.695 644.815 370.975 645.095 ;
        RECT 371.405 644.815 371.685 645.095 ;
        RECT 372.115 644.815 372.395 645.095 ;
        RECT 372.825 644.815 373.105 645.095 ;
        RECT 373.535 644.815 373.815 645.095 ;
        RECT 374.245 644.815 374.525 645.095 ;
        RECT 374.955 644.815 375.235 645.095 ;
        RECT 375.665 644.815 375.945 645.095 ;
        RECT 376.375 644.815 376.655 645.095 ;
        RECT 369.275 644.105 369.555 644.385 ;
        RECT 369.985 644.105 370.265 644.385 ;
        RECT 370.695 644.105 370.975 644.385 ;
        RECT 371.405 644.105 371.685 644.385 ;
        RECT 372.115 644.105 372.395 644.385 ;
        RECT 372.825 644.105 373.105 644.385 ;
        RECT 373.535 644.105 373.815 644.385 ;
        RECT 374.245 644.105 374.525 644.385 ;
        RECT 374.955 644.105 375.235 644.385 ;
        RECT 375.665 644.105 375.945 644.385 ;
        RECT 376.375 644.105 376.655 644.385 ;
        RECT 369.330 640.190 369.610 640.470 ;
        RECT 370.040 640.190 370.320 640.470 ;
        RECT 370.750 640.190 371.030 640.470 ;
        RECT 371.460 640.190 371.740 640.470 ;
        RECT 372.170 640.190 372.450 640.470 ;
        RECT 372.880 640.190 373.160 640.470 ;
        RECT 373.590 640.190 373.870 640.470 ;
        RECT 374.300 640.190 374.580 640.470 ;
        RECT 375.010 640.190 375.290 640.470 ;
        RECT 375.720 640.190 376.000 640.470 ;
        RECT 376.430 640.190 376.710 640.470 ;
        RECT 369.330 639.480 369.610 639.760 ;
        RECT 370.040 639.480 370.320 639.760 ;
        RECT 370.750 639.480 371.030 639.760 ;
        RECT 371.460 639.480 371.740 639.760 ;
        RECT 372.170 639.480 372.450 639.760 ;
        RECT 372.880 639.480 373.160 639.760 ;
        RECT 373.590 639.480 373.870 639.760 ;
        RECT 374.300 639.480 374.580 639.760 ;
        RECT 375.010 639.480 375.290 639.760 ;
        RECT 375.720 639.480 376.000 639.760 ;
        RECT 376.430 639.480 376.710 639.760 ;
        RECT 369.330 638.770 369.610 639.050 ;
        RECT 370.040 638.770 370.320 639.050 ;
        RECT 370.750 638.770 371.030 639.050 ;
        RECT 371.460 638.770 371.740 639.050 ;
        RECT 372.170 638.770 372.450 639.050 ;
        RECT 372.880 638.770 373.160 639.050 ;
        RECT 373.590 638.770 373.870 639.050 ;
        RECT 374.300 638.770 374.580 639.050 ;
        RECT 375.010 638.770 375.290 639.050 ;
        RECT 375.720 638.770 376.000 639.050 ;
        RECT 376.430 638.770 376.710 639.050 ;
        RECT 369.330 638.060 369.610 638.340 ;
        RECT 370.040 638.060 370.320 638.340 ;
        RECT 370.750 638.060 371.030 638.340 ;
        RECT 371.460 638.060 371.740 638.340 ;
        RECT 372.170 638.060 372.450 638.340 ;
        RECT 372.880 638.060 373.160 638.340 ;
        RECT 373.590 638.060 373.870 638.340 ;
        RECT 374.300 638.060 374.580 638.340 ;
        RECT 375.010 638.060 375.290 638.340 ;
        RECT 375.720 638.060 376.000 638.340 ;
        RECT 376.430 638.060 376.710 638.340 ;
        RECT 369.330 637.350 369.610 637.630 ;
        RECT 370.040 637.350 370.320 637.630 ;
        RECT 370.750 637.350 371.030 637.630 ;
        RECT 371.460 637.350 371.740 637.630 ;
        RECT 372.170 637.350 372.450 637.630 ;
        RECT 372.880 637.350 373.160 637.630 ;
        RECT 373.590 637.350 373.870 637.630 ;
        RECT 374.300 637.350 374.580 637.630 ;
        RECT 375.010 637.350 375.290 637.630 ;
        RECT 375.720 637.350 376.000 637.630 ;
        RECT 376.430 637.350 376.710 637.630 ;
        RECT 369.330 636.640 369.610 636.920 ;
        RECT 370.040 636.640 370.320 636.920 ;
        RECT 370.750 636.640 371.030 636.920 ;
        RECT 371.460 636.640 371.740 636.920 ;
        RECT 372.170 636.640 372.450 636.920 ;
        RECT 372.880 636.640 373.160 636.920 ;
        RECT 373.590 636.640 373.870 636.920 ;
        RECT 374.300 636.640 374.580 636.920 ;
        RECT 375.010 636.640 375.290 636.920 ;
        RECT 375.720 636.640 376.000 636.920 ;
        RECT 376.430 636.640 376.710 636.920 ;
        RECT 369.330 635.930 369.610 636.210 ;
        RECT 370.040 635.930 370.320 636.210 ;
        RECT 370.750 635.930 371.030 636.210 ;
        RECT 371.460 635.930 371.740 636.210 ;
        RECT 372.170 635.930 372.450 636.210 ;
        RECT 372.880 635.930 373.160 636.210 ;
        RECT 373.590 635.930 373.870 636.210 ;
        RECT 374.300 635.930 374.580 636.210 ;
        RECT 375.010 635.930 375.290 636.210 ;
        RECT 375.720 635.930 376.000 636.210 ;
        RECT 376.430 635.930 376.710 636.210 ;
        RECT 369.330 635.220 369.610 635.500 ;
        RECT 370.040 635.220 370.320 635.500 ;
        RECT 370.750 635.220 371.030 635.500 ;
        RECT 371.460 635.220 371.740 635.500 ;
        RECT 372.170 635.220 372.450 635.500 ;
        RECT 372.880 635.220 373.160 635.500 ;
        RECT 373.590 635.220 373.870 635.500 ;
        RECT 374.300 635.220 374.580 635.500 ;
        RECT 375.010 635.220 375.290 635.500 ;
        RECT 375.720 635.220 376.000 635.500 ;
        RECT 376.430 635.220 376.710 635.500 ;
        RECT 369.330 634.510 369.610 634.790 ;
        RECT 370.040 634.510 370.320 634.790 ;
        RECT 370.750 634.510 371.030 634.790 ;
        RECT 371.460 634.510 371.740 634.790 ;
        RECT 372.170 634.510 372.450 634.790 ;
        RECT 372.880 634.510 373.160 634.790 ;
        RECT 373.590 634.510 373.870 634.790 ;
        RECT 374.300 634.510 374.580 634.790 ;
        RECT 375.010 634.510 375.290 634.790 ;
        RECT 375.720 634.510 376.000 634.790 ;
        RECT 376.430 634.510 376.710 634.790 ;
        RECT 369.330 633.800 369.610 634.080 ;
        RECT 370.040 633.800 370.320 634.080 ;
        RECT 370.750 633.800 371.030 634.080 ;
        RECT 371.460 633.800 371.740 634.080 ;
        RECT 372.170 633.800 372.450 634.080 ;
        RECT 372.880 633.800 373.160 634.080 ;
        RECT 373.590 633.800 373.870 634.080 ;
        RECT 374.300 633.800 374.580 634.080 ;
        RECT 375.010 633.800 375.290 634.080 ;
        RECT 375.720 633.800 376.000 634.080 ;
        RECT 376.430 633.800 376.710 634.080 ;
        RECT 369.330 633.090 369.610 633.370 ;
        RECT 370.040 633.090 370.320 633.370 ;
        RECT 370.750 633.090 371.030 633.370 ;
        RECT 371.460 633.090 371.740 633.370 ;
        RECT 372.170 633.090 372.450 633.370 ;
        RECT 372.880 633.090 373.160 633.370 ;
        RECT 373.590 633.090 373.870 633.370 ;
        RECT 374.300 633.090 374.580 633.370 ;
        RECT 375.010 633.090 375.290 633.370 ;
        RECT 375.720 633.090 376.000 633.370 ;
        RECT 376.430 633.090 376.710 633.370 ;
        RECT 369.330 632.380 369.610 632.660 ;
        RECT 370.040 632.380 370.320 632.660 ;
        RECT 370.750 632.380 371.030 632.660 ;
        RECT 371.460 632.380 371.740 632.660 ;
        RECT 372.170 632.380 372.450 632.660 ;
        RECT 372.880 632.380 373.160 632.660 ;
        RECT 373.590 632.380 373.870 632.660 ;
        RECT 374.300 632.380 374.580 632.660 ;
        RECT 375.010 632.380 375.290 632.660 ;
        RECT 375.720 632.380 376.000 632.660 ;
        RECT 376.430 632.380 376.710 632.660 ;
        RECT 369.330 631.670 369.610 631.950 ;
        RECT 370.040 631.670 370.320 631.950 ;
        RECT 370.750 631.670 371.030 631.950 ;
        RECT 371.460 631.670 371.740 631.950 ;
        RECT 372.170 631.670 372.450 631.950 ;
        RECT 372.880 631.670 373.160 631.950 ;
        RECT 373.590 631.670 373.870 631.950 ;
        RECT 374.300 631.670 374.580 631.950 ;
        RECT 375.010 631.670 375.290 631.950 ;
        RECT 375.720 631.670 376.000 631.950 ;
        RECT 376.430 631.670 376.710 631.950 ;
        RECT 369.330 497.970 369.610 498.250 ;
        RECT 370.040 497.970 370.320 498.250 ;
        RECT 370.750 497.970 371.030 498.250 ;
        RECT 371.460 497.970 371.740 498.250 ;
        RECT 372.170 497.970 372.450 498.250 ;
        RECT 372.880 497.970 373.160 498.250 ;
        RECT 373.590 497.970 373.870 498.250 ;
        RECT 374.300 497.970 374.580 498.250 ;
        RECT 375.010 497.970 375.290 498.250 ;
        RECT 375.720 497.970 376.000 498.250 ;
        RECT 376.430 497.970 376.710 498.250 ;
        RECT 369.330 497.260 369.610 497.540 ;
        RECT 370.040 497.260 370.320 497.540 ;
        RECT 370.750 497.260 371.030 497.540 ;
        RECT 371.460 497.260 371.740 497.540 ;
        RECT 372.170 497.260 372.450 497.540 ;
        RECT 372.880 497.260 373.160 497.540 ;
        RECT 373.590 497.260 373.870 497.540 ;
        RECT 374.300 497.260 374.580 497.540 ;
        RECT 375.010 497.260 375.290 497.540 ;
        RECT 375.720 497.260 376.000 497.540 ;
        RECT 376.430 497.260 376.710 497.540 ;
        RECT 369.330 496.550 369.610 496.830 ;
        RECT 370.040 496.550 370.320 496.830 ;
        RECT 370.750 496.550 371.030 496.830 ;
        RECT 371.460 496.550 371.740 496.830 ;
        RECT 372.170 496.550 372.450 496.830 ;
        RECT 372.880 496.550 373.160 496.830 ;
        RECT 373.590 496.550 373.870 496.830 ;
        RECT 374.300 496.550 374.580 496.830 ;
        RECT 375.010 496.550 375.290 496.830 ;
        RECT 375.720 496.550 376.000 496.830 ;
        RECT 376.430 496.550 376.710 496.830 ;
        RECT 369.330 495.840 369.610 496.120 ;
        RECT 370.040 495.840 370.320 496.120 ;
        RECT 370.750 495.840 371.030 496.120 ;
        RECT 371.460 495.840 371.740 496.120 ;
        RECT 372.170 495.840 372.450 496.120 ;
        RECT 372.880 495.840 373.160 496.120 ;
        RECT 373.590 495.840 373.870 496.120 ;
        RECT 374.300 495.840 374.580 496.120 ;
        RECT 375.010 495.840 375.290 496.120 ;
        RECT 375.720 495.840 376.000 496.120 ;
        RECT 376.430 495.840 376.710 496.120 ;
        RECT 369.330 495.130 369.610 495.410 ;
        RECT 370.040 495.130 370.320 495.410 ;
        RECT 370.750 495.130 371.030 495.410 ;
        RECT 371.460 495.130 371.740 495.410 ;
        RECT 372.170 495.130 372.450 495.410 ;
        RECT 372.880 495.130 373.160 495.410 ;
        RECT 373.590 495.130 373.870 495.410 ;
        RECT 374.300 495.130 374.580 495.410 ;
        RECT 375.010 495.130 375.290 495.410 ;
        RECT 375.720 495.130 376.000 495.410 ;
        RECT 376.430 495.130 376.710 495.410 ;
        RECT 369.330 494.420 369.610 494.700 ;
        RECT 370.040 494.420 370.320 494.700 ;
        RECT 370.750 494.420 371.030 494.700 ;
        RECT 371.460 494.420 371.740 494.700 ;
        RECT 372.170 494.420 372.450 494.700 ;
        RECT 372.880 494.420 373.160 494.700 ;
        RECT 373.590 494.420 373.870 494.700 ;
        RECT 374.300 494.420 374.580 494.700 ;
        RECT 375.010 494.420 375.290 494.700 ;
        RECT 375.720 494.420 376.000 494.700 ;
        RECT 376.430 494.420 376.710 494.700 ;
        RECT 369.330 493.710 369.610 493.990 ;
        RECT 370.040 493.710 370.320 493.990 ;
        RECT 370.750 493.710 371.030 493.990 ;
        RECT 371.460 493.710 371.740 493.990 ;
        RECT 372.170 493.710 372.450 493.990 ;
        RECT 372.880 493.710 373.160 493.990 ;
        RECT 373.590 493.710 373.870 493.990 ;
        RECT 374.300 493.710 374.580 493.990 ;
        RECT 375.010 493.710 375.290 493.990 ;
        RECT 375.720 493.710 376.000 493.990 ;
        RECT 376.430 493.710 376.710 493.990 ;
        RECT 369.330 493.000 369.610 493.280 ;
        RECT 370.040 493.000 370.320 493.280 ;
        RECT 370.750 493.000 371.030 493.280 ;
        RECT 371.460 493.000 371.740 493.280 ;
        RECT 372.170 493.000 372.450 493.280 ;
        RECT 372.880 493.000 373.160 493.280 ;
        RECT 373.590 493.000 373.870 493.280 ;
        RECT 374.300 493.000 374.580 493.280 ;
        RECT 375.010 493.000 375.290 493.280 ;
        RECT 375.720 493.000 376.000 493.280 ;
        RECT 376.430 493.000 376.710 493.280 ;
        RECT 369.330 492.290 369.610 492.570 ;
        RECT 370.040 492.290 370.320 492.570 ;
        RECT 370.750 492.290 371.030 492.570 ;
        RECT 371.460 492.290 371.740 492.570 ;
        RECT 372.170 492.290 372.450 492.570 ;
        RECT 372.880 492.290 373.160 492.570 ;
        RECT 373.590 492.290 373.870 492.570 ;
        RECT 374.300 492.290 374.580 492.570 ;
        RECT 375.010 492.290 375.290 492.570 ;
        RECT 375.720 492.290 376.000 492.570 ;
        RECT 376.430 492.290 376.710 492.570 ;
        RECT 369.330 491.580 369.610 491.860 ;
        RECT 370.040 491.580 370.320 491.860 ;
        RECT 370.750 491.580 371.030 491.860 ;
        RECT 371.460 491.580 371.740 491.860 ;
        RECT 372.170 491.580 372.450 491.860 ;
        RECT 372.880 491.580 373.160 491.860 ;
        RECT 373.590 491.580 373.870 491.860 ;
        RECT 374.300 491.580 374.580 491.860 ;
        RECT 375.010 491.580 375.290 491.860 ;
        RECT 375.720 491.580 376.000 491.860 ;
        RECT 376.430 491.580 376.710 491.860 ;
        RECT 369.330 490.870 369.610 491.150 ;
        RECT 370.040 490.870 370.320 491.150 ;
        RECT 370.750 490.870 371.030 491.150 ;
        RECT 371.460 490.870 371.740 491.150 ;
        RECT 372.170 490.870 372.450 491.150 ;
        RECT 372.880 490.870 373.160 491.150 ;
        RECT 373.590 490.870 373.870 491.150 ;
        RECT 374.300 490.870 374.580 491.150 ;
        RECT 375.010 490.870 375.290 491.150 ;
        RECT 375.720 490.870 376.000 491.150 ;
        RECT 376.430 490.870 376.710 491.150 ;
        RECT 369.330 490.160 369.610 490.440 ;
        RECT 370.040 490.160 370.320 490.440 ;
        RECT 370.750 490.160 371.030 490.440 ;
        RECT 371.460 490.160 371.740 490.440 ;
        RECT 372.170 490.160 372.450 490.440 ;
        RECT 372.880 490.160 373.160 490.440 ;
        RECT 373.590 490.160 373.870 490.440 ;
        RECT 374.300 490.160 374.580 490.440 ;
        RECT 375.010 490.160 375.290 490.440 ;
        RECT 375.720 490.160 376.000 490.440 ;
        RECT 376.430 490.160 376.710 490.440 ;
        RECT 369.330 489.450 369.610 489.730 ;
        RECT 370.040 489.450 370.320 489.730 ;
        RECT 370.750 489.450 371.030 489.730 ;
        RECT 371.460 489.450 371.740 489.730 ;
        RECT 372.170 489.450 372.450 489.730 ;
        RECT 372.880 489.450 373.160 489.730 ;
        RECT 373.590 489.450 373.870 489.730 ;
        RECT 374.300 489.450 374.580 489.730 ;
        RECT 375.010 489.450 375.290 489.730 ;
        RECT 375.720 489.450 376.000 489.730 ;
        RECT 376.430 489.450 376.710 489.730 ;
        RECT 369.275 485.565 369.555 485.845 ;
        RECT 369.985 485.565 370.265 485.845 ;
        RECT 370.695 485.565 370.975 485.845 ;
        RECT 371.405 485.565 371.685 485.845 ;
        RECT 372.115 485.565 372.395 485.845 ;
        RECT 372.825 485.565 373.105 485.845 ;
        RECT 373.535 485.565 373.815 485.845 ;
        RECT 374.245 485.565 374.525 485.845 ;
        RECT 374.955 485.565 375.235 485.845 ;
        RECT 375.665 485.565 375.945 485.845 ;
        RECT 376.375 485.565 376.655 485.845 ;
        RECT 369.275 484.855 369.555 485.135 ;
        RECT 369.985 484.855 370.265 485.135 ;
        RECT 370.695 484.855 370.975 485.135 ;
        RECT 371.405 484.855 371.685 485.135 ;
        RECT 372.115 484.855 372.395 485.135 ;
        RECT 372.825 484.855 373.105 485.135 ;
        RECT 373.535 484.855 373.815 485.135 ;
        RECT 374.245 484.855 374.525 485.135 ;
        RECT 374.955 484.855 375.235 485.135 ;
        RECT 375.665 484.855 375.945 485.135 ;
        RECT 376.375 484.855 376.655 485.135 ;
        RECT 369.275 484.145 369.555 484.425 ;
        RECT 369.985 484.145 370.265 484.425 ;
        RECT 370.695 484.145 370.975 484.425 ;
        RECT 371.405 484.145 371.685 484.425 ;
        RECT 372.115 484.145 372.395 484.425 ;
        RECT 372.825 484.145 373.105 484.425 ;
        RECT 373.535 484.145 373.815 484.425 ;
        RECT 374.245 484.145 374.525 484.425 ;
        RECT 374.955 484.145 375.235 484.425 ;
        RECT 375.665 484.145 375.945 484.425 ;
        RECT 376.375 484.145 376.655 484.425 ;
        RECT 369.275 483.435 369.555 483.715 ;
        RECT 369.985 483.435 370.265 483.715 ;
        RECT 370.695 483.435 370.975 483.715 ;
        RECT 371.405 483.435 371.685 483.715 ;
        RECT 372.115 483.435 372.395 483.715 ;
        RECT 372.825 483.435 373.105 483.715 ;
        RECT 373.535 483.435 373.815 483.715 ;
        RECT 374.245 483.435 374.525 483.715 ;
        RECT 374.955 483.435 375.235 483.715 ;
        RECT 375.665 483.435 375.945 483.715 ;
        RECT 376.375 483.435 376.655 483.715 ;
        RECT 369.275 482.725 369.555 483.005 ;
        RECT 369.985 482.725 370.265 483.005 ;
        RECT 370.695 482.725 370.975 483.005 ;
        RECT 371.405 482.725 371.685 483.005 ;
        RECT 372.115 482.725 372.395 483.005 ;
        RECT 372.825 482.725 373.105 483.005 ;
        RECT 373.535 482.725 373.815 483.005 ;
        RECT 374.245 482.725 374.525 483.005 ;
        RECT 374.955 482.725 375.235 483.005 ;
        RECT 375.665 482.725 375.945 483.005 ;
        RECT 376.375 482.725 376.655 483.005 ;
        RECT 369.275 482.015 369.555 482.295 ;
        RECT 369.985 482.015 370.265 482.295 ;
        RECT 370.695 482.015 370.975 482.295 ;
        RECT 371.405 482.015 371.685 482.295 ;
        RECT 372.115 482.015 372.395 482.295 ;
        RECT 372.825 482.015 373.105 482.295 ;
        RECT 373.535 482.015 373.815 482.295 ;
        RECT 374.245 482.015 374.525 482.295 ;
        RECT 374.955 482.015 375.235 482.295 ;
        RECT 375.665 482.015 375.945 482.295 ;
        RECT 376.375 482.015 376.655 482.295 ;
        RECT 369.275 481.305 369.555 481.585 ;
        RECT 369.985 481.305 370.265 481.585 ;
        RECT 370.695 481.305 370.975 481.585 ;
        RECT 371.405 481.305 371.685 481.585 ;
        RECT 372.115 481.305 372.395 481.585 ;
        RECT 372.825 481.305 373.105 481.585 ;
        RECT 373.535 481.305 373.815 481.585 ;
        RECT 374.245 481.305 374.525 481.585 ;
        RECT 374.955 481.305 375.235 481.585 ;
        RECT 375.665 481.305 375.945 481.585 ;
        RECT 376.375 481.305 376.655 481.585 ;
        RECT 369.275 480.595 369.555 480.875 ;
        RECT 369.985 480.595 370.265 480.875 ;
        RECT 370.695 480.595 370.975 480.875 ;
        RECT 371.405 480.595 371.685 480.875 ;
        RECT 372.115 480.595 372.395 480.875 ;
        RECT 372.825 480.595 373.105 480.875 ;
        RECT 373.535 480.595 373.815 480.875 ;
        RECT 374.245 480.595 374.525 480.875 ;
        RECT 374.955 480.595 375.235 480.875 ;
        RECT 375.665 480.595 375.945 480.875 ;
        RECT 376.375 480.595 376.655 480.875 ;
        RECT 369.275 479.885 369.555 480.165 ;
        RECT 369.985 479.885 370.265 480.165 ;
        RECT 370.695 479.885 370.975 480.165 ;
        RECT 371.405 479.885 371.685 480.165 ;
        RECT 372.115 479.885 372.395 480.165 ;
        RECT 372.825 479.885 373.105 480.165 ;
        RECT 373.535 479.885 373.815 480.165 ;
        RECT 374.245 479.885 374.525 480.165 ;
        RECT 374.955 479.885 375.235 480.165 ;
        RECT 375.665 479.885 375.945 480.165 ;
        RECT 376.375 479.885 376.655 480.165 ;
        RECT 369.275 479.175 369.555 479.455 ;
        RECT 369.985 479.175 370.265 479.455 ;
        RECT 370.695 479.175 370.975 479.455 ;
        RECT 371.405 479.175 371.685 479.455 ;
        RECT 372.115 479.175 372.395 479.455 ;
        RECT 372.825 479.175 373.105 479.455 ;
        RECT 373.535 479.175 373.815 479.455 ;
        RECT 374.245 479.175 374.525 479.455 ;
        RECT 374.955 479.175 375.235 479.455 ;
        RECT 375.665 479.175 375.945 479.455 ;
        RECT 376.375 479.175 376.655 479.455 ;
        RECT 369.275 478.465 369.555 478.745 ;
        RECT 369.985 478.465 370.265 478.745 ;
        RECT 370.695 478.465 370.975 478.745 ;
        RECT 371.405 478.465 371.685 478.745 ;
        RECT 372.115 478.465 372.395 478.745 ;
        RECT 372.825 478.465 373.105 478.745 ;
        RECT 373.535 478.465 373.815 478.745 ;
        RECT 374.245 478.465 374.525 478.745 ;
        RECT 374.955 478.465 375.235 478.745 ;
        RECT 375.665 478.465 375.945 478.745 ;
        RECT 376.375 478.465 376.655 478.745 ;
        RECT 369.275 477.755 369.555 478.035 ;
        RECT 369.985 477.755 370.265 478.035 ;
        RECT 370.695 477.755 370.975 478.035 ;
        RECT 371.405 477.755 371.685 478.035 ;
        RECT 372.115 477.755 372.395 478.035 ;
        RECT 372.825 477.755 373.105 478.035 ;
        RECT 373.535 477.755 373.815 478.035 ;
        RECT 374.245 477.755 374.525 478.035 ;
        RECT 374.955 477.755 375.235 478.035 ;
        RECT 375.665 477.755 375.945 478.035 ;
        RECT 376.375 477.755 376.655 478.035 ;
        RECT 369.275 477.045 369.555 477.325 ;
        RECT 369.985 477.045 370.265 477.325 ;
        RECT 370.695 477.045 370.975 477.325 ;
        RECT 371.405 477.045 371.685 477.325 ;
        RECT 372.115 477.045 372.395 477.325 ;
        RECT 372.825 477.045 373.105 477.325 ;
        RECT 373.535 477.045 373.815 477.325 ;
        RECT 374.245 477.045 374.525 477.325 ;
        RECT 374.955 477.045 375.235 477.325 ;
        RECT 375.665 477.045 375.945 477.325 ;
        RECT 376.375 477.045 376.655 477.325 ;
        RECT 369.275 476.335 369.555 476.615 ;
        RECT 369.985 476.335 370.265 476.615 ;
        RECT 370.695 476.335 370.975 476.615 ;
        RECT 371.405 476.335 371.685 476.615 ;
        RECT 372.115 476.335 372.395 476.615 ;
        RECT 372.825 476.335 373.105 476.615 ;
        RECT 373.535 476.335 373.815 476.615 ;
        RECT 374.245 476.335 374.525 476.615 ;
        RECT 374.955 476.335 375.235 476.615 ;
        RECT 375.665 476.335 375.945 476.615 ;
        RECT 376.375 476.335 376.655 476.615 ;
        RECT 369.275 473.715 369.555 473.995 ;
        RECT 369.985 473.715 370.265 473.995 ;
        RECT 370.695 473.715 370.975 473.995 ;
        RECT 371.405 473.715 371.685 473.995 ;
        RECT 372.115 473.715 372.395 473.995 ;
        RECT 372.825 473.715 373.105 473.995 ;
        RECT 373.535 473.715 373.815 473.995 ;
        RECT 374.245 473.715 374.525 473.995 ;
        RECT 374.955 473.715 375.235 473.995 ;
        RECT 375.665 473.715 375.945 473.995 ;
        RECT 376.375 473.715 376.655 473.995 ;
        RECT 369.275 473.005 369.555 473.285 ;
        RECT 369.985 473.005 370.265 473.285 ;
        RECT 370.695 473.005 370.975 473.285 ;
        RECT 371.405 473.005 371.685 473.285 ;
        RECT 372.115 473.005 372.395 473.285 ;
        RECT 372.825 473.005 373.105 473.285 ;
        RECT 373.535 473.005 373.815 473.285 ;
        RECT 374.245 473.005 374.525 473.285 ;
        RECT 374.955 473.005 375.235 473.285 ;
        RECT 375.665 473.005 375.945 473.285 ;
        RECT 376.375 473.005 376.655 473.285 ;
        RECT 369.275 472.295 369.555 472.575 ;
        RECT 369.985 472.295 370.265 472.575 ;
        RECT 370.695 472.295 370.975 472.575 ;
        RECT 371.405 472.295 371.685 472.575 ;
        RECT 372.115 472.295 372.395 472.575 ;
        RECT 372.825 472.295 373.105 472.575 ;
        RECT 373.535 472.295 373.815 472.575 ;
        RECT 374.245 472.295 374.525 472.575 ;
        RECT 374.955 472.295 375.235 472.575 ;
        RECT 375.665 472.295 375.945 472.575 ;
        RECT 376.375 472.295 376.655 472.575 ;
        RECT 369.275 471.585 369.555 471.865 ;
        RECT 369.985 471.585 370.265 471.865 ;
        RECT 370.695 471.585 370.975 471.865 ;
        RECT 371.405 471.585 371.685 471.865 ;
        RECT 372.115 471.585 372.395 471.865 ;
        RECT 372.825 471.585 373.105 471.865 ;
        RECT 373.535 471.585 373.815 471.865 ;
        RECT 374.245 471.585 374.525 471.865 ;
        RECT 374.955 471.585 375.235 471.865 ;
        RECT 375.665 471.585 375.945 471.865 ;
        RECT 376.375 471.585 376.655 471.865 ;
        RECT 369.275 470.875 369.555 471.155 ;
        RECT 369.985 470.875 370.265 471.155 ;
        RECT 370.695 470.875 370.975 471.155 ;
        RECT 371.405 470.875 371.685 471.155 ;
        RECT 372.115 470.875 372.395 471.155 ;
        RECT 372.825 470.875 373.105 471.155 ;
        RECT 373.535 470.875 373.815 471.155 ;
        RECT 374.245 470.875 374.525 471.155 ;
        RECT 374.955 470.875 375.235 471.155 ;
        RECT 375.665 470.875 375.945 471.155 ;
        RECT 376.375 470.875 376.655 471.155 ;
        RECT 369.275 470.165 369.555 470.445 ;
        RECT 369.985 470.165 370.265 470.445 ;
        RECT 370.695 470.165 370.975 470.445 ;
        RECT 371.405 470.165 371.685 470.445 ;
        RECT 372.115 470.165 372.395 470.445 ;
        RECT 372.825 470.165 373.105 470.445 ;
        RECT 373.535 470.165 373.815 470.445 ;
        RECT 374.245 470.165 374.525 470.445 ;
        RECT 374.955 470.165 375.235 470.445 ;
        RECT 375.665 470.165 375.945 470.445 ;
        RECT 376.375 470.165 376.655 470.445 ;
        RECT 369.275 469.455 369.555 469.735 ;
        RECT 369.985 469.455 370.265 469.735 ;
        RECT 370.695 469.455 370.975 469.735 ;
        RECT 371.405 469.455 371.685 469.735 ;
        RECT 372.115 469.455 372.395 469.735 ;
        RECT 372.825 469.455 373.105 469.735 ;
        RECT 373.535 469.455 373.815 469.735 ;
        RECT 374.245 469.455 374.525 469.735 ;
        RECT 374.955 469.455 375.235 469.735 ;
        RECT 375.665 469.455 375.945 469.735 ;
        RECT 376.375 469.455 376.655 469.735 ;
        RECT 369.275 468.745 369.555 469.025 ;
        RECT 369.985 468.745 370.265 469.025 ;
        RECT 370.695 468.745 370.975 469.025 ;
        RECT 371.405 468.745 371.685 469.025 ;
        RECT 372.115 468.745 372.395 469.025 ;
        RECT 372.825 468.745 373.105 469.025 ;
        RECT 373.535 468.745 373.815 469.025 ;
        RECT 374.245 468.745 374.525 469.025 ;
        RECT 374.955 468.745 375.235 469.025 ;
        RECT 375.665 468.745 375.945 469.025 ;
        RECT 376.375 468.745 376.655 469.025 ;
        RECT 369.275 468.035 369.555 468.315 ;
        RECT 369.985 468.035 370.265 468.315 ;
        RECT 370.695 468.035 370.975 468.315 ;
        RECT 371.405 468.035 371.685 468.315 ;
        RECT 372.115 468.035 372.395 468.315 ;
        RECT 372.825 468.035 373.105 468.315 ;
        RECT 373.535 468.035 373.815 468.315 ;
        RECT 374.245 468.035 374.525 468.315 ;
        RECT 374.955 468.035 375.235 468.315 ;
        RECT 375.665 468.035 375.945 468.315 ;
        RECT 376.375 468.035 376.655 468.315 ;
        RECT 369.275 467.325 369.555 467.605 ;
        RECT 369.985 467.325 370.265 467.605 ;
        RECT 370.695 467.325 370.975 467.605 ;
        RECT 371.405 467.325 371.685 467.605 ;
        RECT 372.115 467.325 372.395 467.605 ;
        RECT 372.825 467.325 373.105 467.605 ;
        RECT 373.535 467.325 373.815 467.605 ;
        RECT 374.245 467.325 374.525 467.605 ;
        RECT 374.955 467.325 375.235 467.605 ;
        RECT 375.665 467.325 375.945 467.605 ;
        RECT 376.375 467.325 376.655 467.605 ;
        RECT 369.275 466.615 369.555 466.895 ;
        RECT 369.985 466.615 370.265 466.895 ;
        RECT 370.695 466.615 370.975 466.895 ;
        RECT 371.405 466.615 371.685 466.895 ;
        RECT 372.115 466.615 372.395 466.895 ;
        RECT 372.825 466.615 373.105 466.895 ;
        RECT 373.535 466.615 373.815 466.895 ;
        RECT 374.245 466.615 374.525 466.895 ;
        RECT 374.955 466.615 375.235 466.895 ;
        RECT 375.665 466.615 375.945 466.895 ;
        RECT 376.375 466.615 376.655 466.895 ;
        RECT 369.275 465.905 369.555 466.185 ;
        RECT 369.985 465.905 370.265 466.185 ;
        RECT 370.695 465.905 370.975 466.185 ;
        RECT 371.405 465.905 371.685 466.185 ;
        RECT 372.115 465.905 372.395 466.185 ;
        RECT 372.825 465.905 373.105 466.185 ;
        RECT 373.535 465.905 373.815 466.185 ;
        RECT 374.245 465.905 374.525 466.185 ;
        RECT 374.955 465.905 375.235 466.185 ;
        RECT 375.665 465.905 375.945 466.185 ;
        RECT 376.375 465.905 376.655 466.185 ;
        RECT 369.275 465.195 369.555 465.475 ;
        RECT 369.985 465.195 370.265 465.475 ;
        RECT 370.695 465.195 370.975 465.475 ;
        RECT 371.405 465.195 371.685 465.475 ;
        RECT 372.115 465.195 372.395 465.475 ;
        RECT 372.825 465.195 373.105 465.475 ;
        RECT 373.535 465.195 373.815 465.475 ;
        RECT 374.245 465.195 374.525 465.475 ;
        RECT 374.955 465.195 375.235 465.475 ;
        RECT 375.665 465.195 375.945 465.475 ;
        RECT 376.375 465.195 376.655 465.475 ;
        RECT 369.275 464.485 369.555 464.765 ;
        RECT 369.985 464.485 370.265 464.765 ;
        RECT 370.695 464.485 370.975 464.765 ;
        RECT 371.405 464.485 371.685 464.765 ;
        RECT 372.115 464.485 372.395 464.765 ;
        RECT 372.825 464.485 373.105 464.765 ;
        RECT 373.535 464.485 373.815 464.765 ;
        RECT 374.245 464.485 374.525 464.765 ;
        RECT 374.955 464.485 375.235 464.765 ;
        RECT 375.665 464.485 375.945 464.765 ;
        RECT 376.375 464.485 376.655 464.765 ;
        RECT 369.275 460.185 369.555 460.465 ;
        RECT 369.985 460.185 370.265 460.465 ;
        RECT 370.695 460.185 370.975 460.465 ;
        RECT 371.405 460.185 371.685 460.465 ;
        RECT 372.115 460.185 372.395 460.465 ;
        RECT 372.825 460.185 373.105 460.465 ;
        RECT 373.535 460.185 373.815 460.465 ;
        RECT 374.245 460.185 374.525 460.465 ;
        RECT 374.955 460.185 375.235 460.465 ;
        RECT 375.665 460.185 375.945 460.465 ;
        RECT 376.375 460.185 376.655 460.465 ;
        RECT 369.275 459.475 369.555 459.755 ;
        RECT 369.985 459.475 370.265 459.755 ;
        RECT 370.695 459.475 370.975 459.755 ;
        RECT 371.405 459.475 371.685 459.755 ;
        RECT 372.115 459.475 372.395 459.755 ;
        RECT 372.825 459.475 373.105 459.755 ;
        RECT 373.535 459.475 373.815 459.755 ;
        RECT 374.245 459.475 374.525 459.755 ;
        RECT 374.955 459.475 375.235 459.755 ;
        RECT 375.665 459.475 375.945 459.755 ;
        RECT 376.375 459.475 376.655 459.755 ;
        RECT 369.275 458.765 369.555 459.045 ;
        RECT 369.985 458.765 370.265 459.045 ;
        RECT 370.695 458.765 370.975 459.045 ;
        RECT 371.405 458.765 371.685 459.045 ;
        RECT 372.115 458.765 372.395 459.045 ;
        RECT 372.825 458.765 373.105 459.045 ;
        RECT 373.535 458.765 373.815 459.045 ;
        RECT 374.245 458.765 374.525 459.045 ;
        RECT 374.955 458.765 375.235 459.045 ;
        RECT 375.665 458.765 375.945 459.045 ;
        RECT 376.375 458.765 376.655 459.045 ;
        RECT 369.275 458.055 369.555 458.335 ;
        RECT 369.985 458.055 370.265 458.335 ;
        RECT 370.695 458.055 370.975 458.335 ;
        RECT 371.405 458.055 371.685 458.335 ;
        RECT 372.115 458.055 372.395 458.335 ;
        RECT 372.825 458.055 373.105 458.335 ;
        RECT 373.535 458.055 373.815 458.335 ;
        RECT 374.245 458.055 374.525 458.335 ;
        RECT 374.955 458.055 375.235 458.335 ;
        RECT 375.665 458.055 375.945 458.335 ;
        RECT 376.375 458.055 376.655 458.335 ;
        RECT 369.275 457.345 369.555 457.625 ;
        RECT 369.985 457.345 370.265 457.625 ;
        RECT 370.695 457.345 370.975 457.625 ;
        RECT 371.405 457.345 371.685 457.625 ;
        RECT 372.115 457.345 372.395 457.625 ;
        RECT 372.825 457.345 373.105 457.625 ;
        RECT 373.535 457.345 373.815 457.625 ;
        RECT 374.245 457.345 374.525 457.625 ;
        RECT 374.955 457.345 375.235 457.625 ;
        RECT 375.665 457.345 375.945 457.625 ;
        RECT 376.375 457.345 376.655 457.625 ;
        RECT 369.275 456.635 369.555 456.915 ;
        RECT 369.985 456.635 370.265 456.915 ;
        RECT 370.695 456.635 370.975 456.915 ;
        RECT 371.405 456.635 371.685 456.915 ;
        RECT 372.115 456.635 372.395 456.915 ;
        RECT 372.825 456.635 373.105 456.915 ;
        RECT 373.535 456.635 373.815 456.915 ;
        RECT 374.245 456.635 374.525 456.915 ;
        RECT 374.955 456.635 375.235 456.915 ;
        RECT 375.665 456.635 375.945 456.915 ;
        RECT 376.375 456.635 376.655 456.915 ;
        RECT 369.275 455.925 369.555 456.205 ;
        RECT 369.985 455.925 370.265 456.205 ;
        RECT 370.695 455.925 370.975 456.205 ;
        RECT 371.405 455.925 371.685 456.205 ;
        RECT 372.115 455.925 372.395 456.205 ;
        RECT 372.825 455.925 373.105 456.205 ;
        RECT 373.535 455.925 373.815 456.205 ;
        RECT 374.245 455.925 374.525 456.205 ;
        RECT 374.955 455.925 375.235 456.205 ;
        RECT 375.665 455.925 375.945 456.205 ;
        RECT 376.375 455.925 376.655 456.205 ;
        RECT 369.275 455.215 369.555 455.495 ;
        RECT 369.985 455.215 370.265 455.495 ;
        RECT 370.695 455.215 370.975 455.495 ;
        RECT 371.405 455.215 371.685 455.495 ;
        RECT 372.115 455.215 372.395 455.495 ;
        RECT 372.825 455.215 373.105 455.495 ;
        RECT 373.535 455.215 373.815 455.495 ;
        RECT 374.245 455.215 374.525 455.495 ;
        RECT 374.955 455.215 375.235 455.495 ;
        RECT 375.665 455.215 375.945 455.495 ;
        RECT 376.375 455.215 376.655 455.495 ;
        RECT 369.275 454.505 369.555 454.785 ;
        RECT 369.985 454.505 370.265 454.785 ;
        RECT 370.695 454.505 370.975 454.785 ;
        RECT 371.405 454.505 371.685 454.785 ;
        RECT 372.115 454.505 372.395 454.785 ;
        RECT 372.825 454.505 373.105 454.785 ;
        RECT 373.535 454.505 373.815 454.785 ;
        RECT 374.245 454.505 374.525 454.785 ;
        RECT 374.955 454.505 375.235 454.785 ;
        RECT 375.665 454.505 375.945 454.785 ;
        RECT 376.375 454.505 376.655 454.785 ;
        RECT 369.275 453.795 369.555 454.075 ;
        RECT 369.985 453.795 370.265 454.075 ;
        RECT 370.695 453.795 370.975 454.075 ;
        RECT 371.405 453.795 371.685 454.075 ;
        RECT 372.115 453.795 372.395 454.075 ;
        RECT 372.825 453.795 373.105 454.075 ;
        RECT 373.535 453.795 373.815 454.075 ;
        RECT 374.245 453.795 374.525 454.075 ;
        RECT 374.955 453.795 375.235 454.075 ;
        RECT 375.665 453.795 375.945 454.075 ;
        RECT 376.375 453.795 376.655 454.075 ;
        RECT 369.275 453.085 369.555 453.365 ;
        RECT 369.985 453.085 370.265 453.365 ;
        RECT 370.695 453.085 370.975 453.365 ;
        RECT 371.405 453.085 371.685 453.365 ;
        RECT 372.115 453.085 372.395 453.365 ;
        RECT 372.825 453.085 373.105 453.365 ;
        RECT 373.535 453.085 373.815 453.365 ;
        RECT 374.245 453.085 374.525 453.365 ;
        RECT 374.955 453.085 375.235 453.365 ;
        RECT 375.665 453.085 375.945 453.365 ;
        RECT 376.375 453.085 376.655 453.365 ;
        RECT 369.275 452.375 369.555 452.655 ;
        RECT 369.985 452.375 370.265 452.655 ;
        RECT 370.695 452.375 370.975 452.655 ;
        RECT 371.405 452.375 371.685 452.655 ;
        RECT 372.115 452.375 372.395 452.655 ;
        RECT 372.825 452.375 373.105 452.655 ;
        RECT 373.535 452.375 373.815 452.655 ;
        RECT 374.245 452.375 374.525 452.655 ;
        RECT 374.955 452.375 375.235 452.655 ;
        RECT 375.665 452.375 375.945 452.655 ;
        RECT 376.375 452.375 376.655 452.655 ;
        RECT 369.275 451.665 369.555 451.945 ;
        RECT 369.985 451.665 370.265 451.945 ;
        RECT 370.695 451.665 370.975 451.945 ;
        RECT 371.405 451.665 371.685 451.945 ;
        RECT 372.115 451.665 372.395 451.945 ;
        RECT 372.825 451.665 373.105 451.945 ;
        RECT 373.535 451.665 373.815 451.945 ;
        RECT 374.245 451.665 374.525 451.945 ;
        RECT 374.955 451.665 375.235 451.945 ;
        RECT 375.665 451.665 375.945 451.945 ;
        RECT 376.375 451.665 376.655 451.945 ;
        RECT 369.275 450.955 369.555 451.235 ;
        RECT 369.985 450.955 370.265 451.235 ;
        RECT 370.695 450.955 370.975 451.235 ;
        RECT 371.405 450.955 371.685 451.235 ;
        RECT 372.115 450.955 372.395 451.235 ;
        RECT 372.825 450.955 373.105 451.235 ;
        RECT 373.535 450.955 373.815 451.235 ;
        RECT 374.245 450.955 374.525 451.235 ;
        RECT 374.955 450.955 375.235 451.235 ;
        RECT 375.665 450.955 375.945 451.235 ;
        RECT 376.375 450.955 376.655 451.235 ;
        RECT 369.275 448.335 369.555 448.615 ;
        RECT 369.985 448.335 370.265 448.615 ;
        RECT 370.695 448.335 370.975 448.615 ;
        RECT 371.405 448.335 371.685 448.615 ;
        RECT 372.115 448.335 372.395 448.615 ;
        RECT 372.825 448.335 373.105 448.615 ;
        RECT 373.535 448.335 373.815 448.615 ;
        RECT 374.245 448.335 374.525 448.615 ;
        RECT 374.955 448.335 375.235 448.615 ;
        RECT 375.665 448.335 375.945 448.615 ;
        RECT 376.375 448.335 376.655 448.615 ;
        RECT 369.275 447.625 369.555 447.905 ;
        RECT 369.985 447.625 370.265 447.905 ;
        RECT 370.695 447.625 370.975 447.905 ;
        RECT 371.405 447.625 371.685 447.905 ;
        RECT 372.115 447.625 372.395 447.905 ;
        RECT 372.825 447.625 373.105 447.905 ;
        RECT 373.535 447.625 373.815 447.905 ;
        RECT 374.245 447.625 374.525 447.905 ;
        RECT 374.955 447.625 375.235 447.905 ;
        RECT 375.665 447.625 375.945 447.905 ;
        RECT 376.375 447.625 376.655 447.905 ;
        RECT 369.275 446.915 369.555 447.195 ;
        RECT 369.985 446.915 370.265 447.195 ;
        RECT 370.695 446.915 370.975 447.195 ;
        RECT 371.405 446.915 371.685 447.195 ;
        RECT 372.115 446.915 372.395 447.195 ;
        RECT 372.825 446.915 373.105 447.195 ;
        RECT 373.535 446.915 373.815 447.195 ;
        RECT 374.245 446.915 374.525 447.195 ;
        RECT 374.955 446.915 375.235 447.195 ;
        RECT 375.665 446.915 375.945 447.195 ;
        RECT 376.375 446.915 376.655 447.195 ;
        RECT 369.275 446.205 369.555 446.485 ;
        RECT 369.985 446.205 370.265 446.485 ;
        RECT 370.695 446.205 370.975 446.485 ;
        RECT 371.405 446.205 371.685 446.485 ;
        RECT 372.115 446.205 372.395 446.485 ;
        RECT 372.825 446.205 373.105 446.485 ;
        RECT 373.535 446.205 373.815 446.485 ;
        RECT 374.245 446.205 374.525 446.485 ;
        RECT 374.955 446.205 375.235 446.485 ;
        RECT 375.665 446.205 375.945 446.485 ;
        RECT 376.375 446.205 376.655 446.485 ;
        RECT 369.275 445.495 369.555 445.775 ;
        RECT 369.985 445.495 370.265 445.775 ;
        RECT 370.695 445.495 370.975 445.775 ;
        RECT 371.405 445.495 371.685 445.775 ;
        RECT 372.115 445.495 372.395 445.775 ;
        RECT 372.825 445.495 373.105 445.775 ;
        RECT 373.535 445.495 373.815 445.775 ;
        RECT 374.245 445.495 374.525 445.775 ;
        RECT 374.955 445.495 375.235 445.775 ;
        RECT 375.665 445.495 375.945 445.775 ;
        RECT 376.375 445.495 376.655 445.775 ;
        RECT 369.275 444.785 369.555 445.065 ;
        RECT 369.985 444.785 370.265 445.065 ;
        RECT 370.695 444.785 370.975 445.065 ;
        RECT 371.405 444.785 371.685 445.065 ;
        RECT 372.115 444.785 372.395 445.065 ;
        RECT 372.825 444.785 373.105 445.065 ;
        RECT 373.535 444.785 373.815 445.065 ;
        RECT 374.245 444.785 374.525 445.065 ;
        RECT 374.955 444.785 375.235 445.065 ;
        RECT 375.665 444.785 375.945 445.065 ;
        RECT 376.375 444.785 376.655 445.065 ;
        RECT 369.275 444.075 369.555 444.355 ;
        RECT 369.985 444.075 370.265 444.355 ;
        RECT 370.695 444.075 370.975 444.355 ;
        RECT 371.405 444.075 371.685 444.355 ;
        RECT 372.115 444.075 372.395 444.355 ;
        RECT 372.825 444.075 373.105 444.355 ;
        RECT 373.535 444.075 373.815 444.355 ;
        RECT 374.245 444.075 374.525 444.355 ;
        RECT 374.955 444.075 375.235 444.355 ;
        RECT 375.665 444.075 375.945 444.355 ;
        RECT 376.375 444.075 376.655 444.355 ;
        RECT 369.275 443.365 369.555 443.645 ;
        RECT 369.985 443.365 370.265 443.645 ;
        RECT 370.695 443.365 370.975 443.645 ;
        RECT 371.405 443.365 371.685 443.645 ;
        RECT 372.115 443.365 372.395 443.645 ;
        RECT 372.825 443.365 373.105 443.645 ;
        RECT 373.535 443.365 373.815 443.645 ;
        RECT 374.245 443.365 374.525 443.645 ;
        RECT 374.955 443.365 375.235 443.645 ;
        RECT 375.665 443.365 375.945 443.645 ;
        RECT 376.375 443.365 376.655 443.645 ;
        RECT 369.275 442.655 369.555 442.935 ;
        RECT 369.985 442.655 370.265 442.935 ;
        RECT 370.695 442.655 370.975 442.935 ;
        RECT 371.405 442.655 371.685 442.935 ;
        RECT 372.115 442.655 372.395 442.935 ;
        RECT 372.825 442.655 373.105 442.935 ;
        RECT 373.535 442.655 373.815 442.935 ;
        RECT 374.245 442.655 374.525 442.935 ;
        RECT 374.955 442.655 375.235 442.935 ;
        RECT 375.665 442.655 375.945 442.935 ;
        RECT 376.375 442.655 376.655 442.935 ;
        RECT 369.275 441.945 369.555 442.225 ;
        RECT 369.985 441.945 370.265 442.225 ;
        RECT 370.695 441.945 370.975 442.225 ;
        RECT 371.405 441.945 371.685 442.225 ;
        RECT 372.115 441.945 372.395 442.225 ;
        RECT 372.825 441.945 373.105 442.225 ;
        RECT 373.535 441.945 373.815 442.225 ;
        RECT 374.245 441.945 374.525 442.225 ;
        RECT 374.955 441.945 375.235 442.225 ;
        RECT 375.665 441.945 375.945 442.225 ;
        RECT 376.375 441.945 376.655 442.225 ;
        RECT 369.275 441.235 369.555 441.515 ;
        RECT 369.985 441.235 370.265 441.515 ;
        RECT 370.695 441.235 370.975 441.515 ;
        RECT 371.405 441.235 371.685 441.515 ;
        RECT 372.115 441.235 372.395 441.515 ;
        RECT 372.825 441.235 373.105 441.515 ;
        RECT 373.535 441.235 373.815 441.515 ;
        RECT 374.245 441.235 374.525 441.515 ;
        RECT 374.955 441.235 375.235 441.515 ;
        RECT 375.665 441.235 375.945 441.515 ;
        RECT 376.375 441.235 376.655 441.515 ;
        RECT 369.275 440.525 369.555 440.805 ;
        RECT 369.985 440.525 370.265 440.805 ;
        RECT 370.695 440.525 370.975 440.805 ;
        RECT 371.405 440.525 371.685 440.805 ;
        RECT 372.115 440.525 372.395 440.805 ;
        RECT 372.825 440.525 373.105 440.805 ;
        RECT 373.535 440.525 373.815 440.805 ;
        RECT 374.245 440.525 374.525 440.805 ;
        RECT 374.955 440.525 375.235 440.805 ;
        RECT 375.665 440.525 375.945 440.805 ;
        RECT 376.375 440.525 376.655 440.805 ;
        RECT 369.275 439.815 369.555 440.095 ;
        RECT 369.985 439.815 370.265 440.095 ;
        RECT 370.695 439.815 370.975 440.095 ;
        RECT 371.405 439.815 371.685 440.095 ;
        RECT 372.115 439.815 372.395 440.095 ;
        RECT 372.825 439.815 373.105 440.095 ;
        RECT 373.535 439.815 373.815 440.095 ;
        RECT 374.245 439.815 374.525 440.095 ;
        RECT 374.955 439.815 375.235 440.095 ;
        RECT 375.665 439.815 375.945 440.095 ;
        RECT 376.375 439.815 376.655 440.095 ;
        RECT 369.275 439.105 369.555 439.385 ;
        RECT 369.985 439.105 370.265 439.385 ;
        RECT 370.695 439.105 370.975 439.385 ;
        RECT 371.405 439.105 371.685 439.385 ;
        RECT 372.115 439.105 372.395 439.385 ;
        RECT 372.825 439.105 373.105 439.385 ;
        RECT 373.535 439.105 373.815 439.385 ;
        RECT 374.245 439.105 374.525 439.385 ;
        RECT 374.955 439.105 375.235 439.385 ;
        RECT 375.665 439.105 375.945 439.385 ;
        RECT 376.375 439.105 376.655 439.385 ;
        RECT 369.330 435.190 369.610 435.470 ;
        RECT 370.040 435.190 370.320 435.470 ;
        RECT 370.750 435.190 371.030 435.470 ;
        RECT 371.460 435.190 371.740 435.470 ;
        RECT 372.170 435.190 372.450 435.470 ;
        RECT 372.880 435.190 373.160 435.470 ;
        RECT 373.590 435.190 373.870 435.470 ;
        RECT 374.300 435.190 374.580 435.470 ;
        RECT 375.010 435.190 375.290 435.470 ;
        RECT 375.720 435.190 376.000 435.470 ;
        RECT 376.430 435.190 376.710 435.470 ;
        RECT 369.330 434.480 369.610 434.760 ;
        RECT 370.040 434.480 370.320 434.760 ;
        RECT 370.750 434.480 371.030 434.760 ;
        RECT 371.460 434.480 371.740 434.760 ;
        RECT 372.170 434.480 372.450 434.760 ;
        RECT 372.880 434.480 373.160 434.760 ;
        RECT 373.590 434.480 373.870 434.760 ;
        RECT 374.300 434.480 374.580 434.760 ;
        RECT 375.010 434.480 375.290 434.760 ;
        RECT 375.720 434.480 376.000 434.760 ;
        RECT 376.430 434.480 376.710 434.760 ;
        RECT 369.330 433.770 369.610 434.050 ;
        RECT 370.040 433.770 370.320 434.050 ;
        RECT 370.750 433.770 371.030 434.050 ;
        RECT 371.460 433.770 371.740 434.050 ;
        RECT 372.170 433.770 372.450 434.050 ;
        RECT 372.880 433.770 373.160 434.050 ;
        RECT 373.590 433.770 373.870 434.050 ;
        RECT 374.300 433.770 374.580 434.050 ;
        RECT 375.010 433.770 375.290 434.050 ;
        RECT 375.720 433.770 376.000 434.050 ;
        RECT 376.430 433.770 376.710 434.050 ;
        RECT 369.330 433.060 369.610 433.340 ;
        RECT 370.040 433.060 370.320 433.340 ;
        RECT 370.750 433.060 371.030 433.340 ;
        RECT 371.460 433.060 371.740 433.340 ;
        RECT 372.170 433.060 372.450 433.340 ;
        RECT 372.880 433.060 373.160 433.340 ;
        RECT 373.590 433.060 373.870 433.340 ;
        RECT 374.300 433.060 374.580 433.340 ;
        RECT 375.010 433.060 375.290 433.340 ;
        RECT 375.720 433.060 376.000 433.340 ;
        RECT 376.430 433.060 376.710 433.340 ;
        RECT 369.330 432.350 369.610 432.630 ;
        RECT 370.040 432.350 370.320 432.630 ;
        RECT 370.750 432.350 371.030 432.630 ;
        RECT 371.460 432.350 371.740 432.630 ;
        RECT 372.170 432.350 372.450 432.630 ;
        RECT 372.880 432.350 373.160 432.630 ;
        RECT 373.590 432.350 373.870 432.630 ;
        RECT 374.300 432.350 374.580 432.630 ;
        RECT 375.010 432.350 375.290 432.630 ;
        RECT 375.720 432.350 376.000 432.630 ;
        RECT 376.430 432.350 376.710 432.630 ;
        RECT 369.330 431.640 369.610 431.920 ;
        RECT 370.040 431.640 370.320 431.920 ;
        RECT 370.750 431.640 371.030 431.920 ;
        RECT 371.460 431.640 371.740 431.920 ;
        RECT 372.170 431.640 372.450 431.920 ;
        RECT 372.880 431.640 373.160 431.920 ;
        RECT 373.590 431.640 373.870 431.920 ;
        RECT 374.300 431.640 374.580 431.920 ;
        RECT 375.010 431.640 375.290 431.920 ;
        RECT 375.720 431.640 376.000 431.920 ;
        RECT 376.430 431.640 376.710 431.920 ;
        RECT 369.330 430.930 369.610 431.210 ;
        RECT 370.040 430.930 370.320 431.210 ;
        RECT 370.750 430.930 371.030 431.210 ;
        RECT 371.460 430.930 371.740 431.210 ;
        RECT 372.170 430.930 372.450 431.210 ;
        RECT 372.880 430.930 373.160 431.210 ;
        RECT 373.590 430.930 373.870 431.210 ;
        RECT 374.300 430.930 374.580 431.210 ;
        RECT 375.010 430.930 375.290 431.210 ;
        RECT 375.720 430.930 376.000 431.210 ;
        RECT 376.430 430.930 376.710 431.210 ;
        RECT 369.330 430.220 369.610 430.500 ;
        RECT 370.040 430.220 370.320 430.500 ;
        RECT 370.750 430.220 371.030 430.500 ;
        RECT 371.460 430.220 371.740 430.500 ;
        RECT 372.170 430.220 372.450 430.500 ;
        RECT 372.880 430.220 373.160 430.500 ;
        RECT 373.590 430.220 373.870 430.500 ;
        RECT 374.300 430.220 374.580 430.500 ;
        RECT 375.010 430.220 375.290 430.500 ;
        RECT 375.720 430.220 376.000 430.500 ;
        RECT 376.430 430.220 376.710 430.500 ;
        RECT 369.330 429.510 369.610 429.790 ;
        RECT 370.040 429.510 370.320 429.790 ;
        RECT 370.750 429.510 371.030 429.790 ;
        RECT 371.460 429.510 371.740 429.790 ;
        RECT 372.170 429.510 372.450 429.790 ;
        RECT 372.880 429.510 373.160 429.790 ;
        RECT 373.590 429.510 373.870 429.790 ;
        RECT 374.300 429.510 374.580 429.790 ;
        RECT 375.010 429.510 375.290 429.790 ;
        RECT 375.720 429.510 376.000 429.790 ;
        RECT 376.430 429.510 376.710 429.790 ;
        RECT 369.330 428.800 369.610 429.080 ;
        RECT 370.040 428.800 370.320 429.080 ;
        RECT 370.750 428.800 371.030 429.080 ;
        RECT 371.460 428.800 371.740 429.080 ;
        RECT 372.170 428.800 372.450 429.080 ;
        RECT 372.880 428.800 373.160 429.080 ;
        RECT 373.590 428.800 373.870 429.080 ;
        RECT 374.300 428.800 374.580 429.080 ;
        RECT 375.010 428.800 375.290 429.080 ;
        RECT 375.720 428.800 376.000 429.080 ;
        RECT 376.430 428.800 376.710 429.080 ;
        RECT 369.330 428.090 369.610 428.370 ;
        RECT 370.040 428.090 370.320 428.370 ;
        RECT 370.750 428.090 371.030 428.370 ;
        RECT 371.460 428.090 371.740 428.370 ;
        RECT 372.170 428.090 372.450 428.370 ;
        RECT 372.880 428.090 373.160 428.370 ;
        RECT 373.590 428.090 373.870 428.370 ;
        RECT 374.300 428.090 374.580 428.370 ;
        RECT 375.010 428.090 375.290 428.370 ;
        RECT 375.720 428.090 376.000 428.370 ;
        RECT 376.430 428.090 376.710 428.370 ;
        RECT 369.330 427.380 369.610 427.660 ;
        RECT 370.040 427.380 370.320 427.660 ;
        RECT 370.750 427.380 371.030 427.660 ;
        RECT 371.460 427.380 371.740 427.660 ;
        RECT 372.170 427.380 372.450 427.660 ;
        RECT 372.880 427.380 373.160 427.660 ;
        RECT 373.590 427.380 373.870 427.660 ;
        RECT 374.300 427.380 374.580 427.660 ;
        RECT 375.010 427.380 375.290 427.660 ;
        RECT 375.720 427.380 376.000 427.660 ;
        RECT 376.430 427.380 376.710 427.660 ;
        RECT 369.330 426.670 369.610 426.950 ;
        RECT 370.040 426.670 370.320 426.950 ;
        RECT 370.750 426.670 371.030 426.950 ;
        RECT 371.460 426.670 371.740 426.950 ;
        RECT 372.170 426.670 372.450 426.950 ;
        RECT 372.880 426.670 373.160 426.950 ;
        RECT 373.590 426.670 373.870 426.950 ;
        RECT 374.300 426.670 374.580 426.950 ;
        RECT 375.010 426.670 375.290 426.950 ;
        RECT 375.720 426.670 376.000 426.950 ;
        RECT 376.430 426.670 376.710 426.950 ;
        RECT 3276.715 379.895 3276.995 380.175 ;
        RECT 3277.425 379.895 3277.705 380.175 ;
        RECT 3278.135 379.895 3278.415 380.175 ;
        RECT 3278.845 379.895 3279.125 380.175 ;
        RECT 3279.555 379.895 3279.835 380.175 ;
        RECT 3280.265 379.895 3280.545 380.175 ;
        RECT 3280.975 379.895 3281.255 380.175 ;
        RECT 3281.685 379.895 3281.965 380.175 ;
        RECT 3276.715 379.185 3276.995 379.465 ;
        RECT 3277.425 379.185 3277.705 379.465 ;
        RECT 3278.135 379.185 3278.415 379.465 ;
        RECT 3278.845 379.185 3279.125 379.465 ;
        RECT 3279.555 379.185 3279.835 379.465 ;
        RECT 3280.265 379.185 3280.545 379.465 ;
        RECT 3280.975 379.185 3281.255 379.465 ;
        RECT 3281.685 379.185 3281.965 379.465 ;
        RECT 3276.715 378.475 3276.995 378.755 ;
        RECT 3277.425 378.475 3277.705 378.755 ;
        RECT 3278.135 378.475 3278.415 378.755 ;
        RECT 3278.845 378.475 3279.125 378.755 ;
        RECT 3279.555 378.475 3279.835 378.755 ;
        RECT 3280.265 378.475 3280.545 378.755 ;
        RECT 3280.975 378.475 3281.255 378.755 ;
        RECT 3281.685 378.475 3281.965 378.755 ;
        RECT 3276.715 377.765 3276.995 378.045 ;
        RECT 3277.425 377.765 3277.705 378.045 ;
        RECT 3278.135 377.765 3278.415 378.045 ;
        RECT 3278.845 377.765 3279.125 378.045 ;
        RECT 3279.555 377.765 3279.835 378.045 ;
        RECT 3280.265 377.765 3280.545 378.045 ;
        RECT 3280.975 377.765 3281.255 378.045 ;
        RECT 3281.685 377.765 3281.965 378.045 ;
        RECT 3276.715 377.055 3276.995 377.335 ;
        RECT 3277.425 377.055 3277.705 377.335 ;
        RECT 3278.135 377.055 3278.415 377.335 ;
        RECT 3278.845 377.055 3279.125 377.335 ;
        RECT 3279.555 377.055 3279.835 377.335 ;
        RECT 3280.265 377.055 3280.545 377.335 ;
        RECT 3280.975 377.055 3281.255 377.335 ;
        RECT 3281.685 377.055 3281.965 377.335 ;
        RECT 3276.715 376.345 3276.995 376.625 ;
        RECT 3277.425 376.345 3277.705 376.625 ;
        RECT 3278.135 376.345 3278.415 376.625 ;
        RECT 3278.845 376.345 3279.125 376.625 ;
        RECT 3279.555 376.345 3279.835 376.625 ;
        RECT 3280.265 376.345 3280.545 376.625 ;
        RECT 3280.975 376.345 3281.255 376.625 ;
        RECT 3281.685 376.345 3281.965 376.625 ;
        RECT 3276.715 375.635 3276.995 375.915 ;
        RECT 3277.425 375.635 3277.705 375.915 ;
        RECT 3278.135 375.635 3278.415 375.915 ;
        RECT 3278.845 375.635 3279.125 375.915 ;
        RECT 3279.555 375.635 3279.835 375.915 ;
        RECT 3280.265 375.635 3280.545 375.915 ;
        RECT 3280.975 375.635 3281.255 375.915 ;
        RECT 3281.685 375.635 3281.965 375.915 ;
        RECT 3276.715 374.925 3276.995 375.205 ;
        RECT 3277.425 374.925 3277.705 375.205 ;
        RECT 3278.135 374.925 3278.415 375.205 ;
        RECT 3278.845 374.925 3279.125 375.205 ;
        RECT 3279.555 374.925 3279.835 375.205 ;
        RECT 3280.265 374.925 3280.545 375.205 ;
        RECT 3280.975 374.925 3281.255 375.205 ;
        RECT 3281.685 374.925 3281.965 375.205 ;
        RECT 3276.715 374.215 3276.995 374.495 ;
        RECT 3277.425 374.215 3277.705 374.495 ;
        RECT 3278.135 374.215 3278.415 374.495 ;
        RECT 3278.845 374.215 3279.125 374.495 ;
        RECT 3279.555 374.215 3279.835 374.495 ;
        RECT 3280.265 374.215 3280.545 374.495 ;
        RECT 3280.975 374.215 3281.255 374.495 ;
        RECT 3281.685 374.215 3281.965 374.495 ;
        RECT 3276.715 373.505 3276.995 373.785 ;
        RECT 3277.425 373.505 3277.705 373.785 ;
        RECT 3278.135 373.505 3278.415 373.785 ;
        RECT 3278.845 373.505 3279.125 373.785 ;
        RECT 3279.555 373.505 3279.835 373.785 ;
        RECT 3280.265 373.505 3280.545 373.785 ;
        RECT 3280.975 373.505 3281.255 373.785 ;
        RECT 3281.685 373.505 3281.965 373.785 ;
        RECT 3276.715 372.795 3276.995 373.075 ;
        RECT 3277.425 372.795 3277.705 373.075 ;
        RECT 3278.135 372.795 3278.415 373.075 ;
        RECT 3278.845 372.795 3279.125 373.075 ;
        RECT 3279.555 372.795 3279.835 373.075 ;
        RECT 3280.265 372.795 3280.545 373.075 ;
        RECT 3280.975 372.795 3281.255 373.075 ;
        RECT 3281.685 372.795 3281.965 373.075 ;
        RECT 3289.115 379.895 3289.395 380.175 ;
        RECT 3289.825 379.895 3290.105 380.175 ;
        RECT 3290.535 379.895 3290.815 380.175 ;
        RECT 3291.245 379.895 3291.525 380.175 ;
        RECT 3291.955 379.895 3292.235 380.175 ;
        RECT 3292.665 379.895 3292.945 380.175 ;
        RECT 3293.375 379.895 3293.655 380.175 ;
        RECT 3294.085 379.895 3294.365 380.175 ;
        RECT 3294.795 379.895 3295.075 380.175 ;
        RECT 3295.505 379.895 3295.785 380.175 ;
        RECT 3296.215 379.895 3296.495 380.175 ;
        RECT 3296.925 379.895 3297.205 380.175 ;
        RECT 3297.635 379.895 3297.915 380.175 ;
        RECT 3298.345 379.895 3298.625 380.175 ;
        RECT 3289.115 379.185 3289.395 379.465 ;
        RECT 3289.825 379.185 3290.105 379.465 ;
        RECT 3290.535 379.185 3290.815 379.465 ;
        RECT 3291.245 379.185 3291.525 379.465 ;
        RECT 3291.955 379.185 3292.235 379.465 ;
        RECT 3292.665 379.185 3292.945 379.465 ;
        RECT 3293.375 379.185 3293.655 379.465 ;
        RECT 3294.085 379.185 3294.365 379.465 ;
        RECT 3294.795 379.185 3295.075 379.465 ;
        RECT 3295.505 379.185 3295.785 379.465 ;
        RECT 3296.215 379.185 3296.495 379.465 ;
        RECT 3296.925 379.185 3297.205 379.465 ;
        RECT 3297.635 379.185 3297.915 379.465 ;
        RECT 3298.345 379.185 3298.625 379.465 ;
        RECT 3289.115 378.475 3289.395 378.755 ;
        RECT 3289.825 378.475 3290.105 378.755 ;
        RECT 3290.535 378.475 3290.815 378.755 ;
        RECT 3291.245 378.475 3291.525 378.755 ;
        RECT 3291.955 378.475 3292.235 378.755 ;
        RECT 3292.665 378.475 3292.945 378.755 ;
        RECT 3293.375 378.475 3293.655 378.755 ;
        RECT 3294.085 378.475 3294.365 378.755 ;
        RECT 3294.795 378.475 3295.075 378.755 ;
        RECT 3295.505 378.475 3295.785 378.755 ;
        RECT 3296.215 378.475 3296.495 378.755 ;
        RECT 3296.925 378.475 3297.205 378.755 ;
        RECT 3297.635 378.475 3297.915 378.755 ;
        RECT 3298.345 378.475 3298.625 378.755 ;
        RECT 3289.115 377.765 3289.395 378.045 ;
        RECT 3289.825 377.765 3290.105 378.045 ;
        RECT 3290.535 377.765 3290.815 378.045 ;
        RECT 3291.245 377.765 3291.525 378.045 ;
        RECT 3291.955 377.765 3292.235 378.045 ;
        RECT 3292.665 377.765 3292.945 378.045 ;
        RECT 3293.375 377.765 3293.655 378.045 ;
        RECT 3294.085 377.765 3294.365 378.045 ;
        RECT 3294.795 377.765 3295.075 378.045 ;
        RECT 3295.505 377.765 3295.785 378.045 ;
        RECT 3296.215 377.765 3296.495 378.045 ;
        RECT 3296.925 377.765 3297.205 378.045 ;
        RECT 3297.635 377.765 3297.915 378.045 ;
        RECT 3298.345 377.765 3298.625 378.045 ;
        RECT 3289.115 377.055 3289.395 377.335 ;
        RECT 3289.825 377.055 3290.105 377.335 ;
        RECT 3290.535 377.055 3290.815 377.335 ;
        RECT 3291.245 377.055 3291.525 377.335 ;
        RECT 3291.955 377.055 3292.235 377.335 ;
        RECT 3292.665 377.055 3292.945 377.335 ;
        RECT 3293.375 377.055 3293.655 377.335 ;
        RECT 3294.085 377.055 3294.365 377.335 ;
        RECT 3294.795 377.055 3295.075 377.335 ;
        RECT 3295.505 377.055 3295.785 377.335 ;
        RECT 3296.215 377.055 3296.495 377.335 ;
        RECT 3296.925 377.055 3297.205 377.335 ;
        RECT 3297.635 377.055 3297.915 377.335 ;
        RECT 3298.345 377.055 3298.625 377.335 ;
        RECT 3289.115 376.345 3289.395 376.625 ;
        RECT 3289.825 376.345 3290.105 376.625 ;
        RECT 3290.535 376.345 3290.815 376.625 ;
        RECT 3291.245 376.345 3291.525 376.625 ;
        RECT 3291.955 376.345 3292.235 376.625 ;
        RECT 3292.665 376.345 3292.945 376.625 ;
        RECT 3293.375 376.345 3293.655 376.625 ;
        RECT 3294.085 376.345 3294.365 376.625 ;
        RECT 3294.795 376.345 3295.075 376.625 ;
        RECT 3295.505 376.345 3295.785 376.625 ;
        RECT 3296.215 376.345 3296.495 376.625 ;
        RECT 3296.925 376.345 3297.205 376.625 ;
        RECT 3297.635 376.345 3297.915 376.625 ;
        RECT 3298.345 376.345 3298.625 376.625 ;
        RECT 3289.115 375.635 3289.395 375.915 ;
        RECT 3289.825 375.635 3290.105 375.915 ;
        RECT 3290.535 375.635 3290.815 375.915 ;
        RECT 3291.245 375.635 3291.525 375.915 ;
        RECT 3291.955 375.635 3292.235 375.915 ;
        RECT 3292.665 375.635 3292.945 375.915 ;
        RECT 3293.375 375.635 3293.655 375.915 ;
        RECT 3294.085 375.635 3294.365 375.915 ;
        RECT 3294.795 375.635 3295.075 375.915 ;
        RECT 3295.505 375.635 3295.785 375.915 ;
        RECT 3296.215 375.635 3296.495 375.915 ;
        RECT 3296.925 375.635 3297.205 375.915 ;
        RECT 3297.635 375.635 3297.915 375.915 ;
        RECT 3298.345 375.635 3298.625 375.915 ;
        RECT 3289.115 374.925 3289.395 375.205 ;
        RECT 3289.825 374.925 3290.105 375.205 ;
        RECT 3290.535 374.925 3290.815 375.205 ;
        RECT 3291.245 374.925 3291.525 375.205 ;
        RECT 3291.955 374.925 3292.235 375.205 ;
        RECT 3292.665 374.925 3292.945 375.205 ;
        RECT 3293.375 374.925 3293.655 375.205 ;
        RECT 3294.085 374.925 3294.365 375.205 ;
        RECT 3294.795 374.925 3295.075 375.205 ;
        RECT 3295.505 374.925 3295.785 375.205 ;
        RECT 3296.215 374.925 3296.495 375.205 ;
        RECT 3296.925 374.925 3297.205 375.205 ;
        RECT 3297.635 374.925 3297.915 375.205 ;
        RECT 3298.345 374.925 3298.625 375.205 ;
        RECT 3289.115 374.215 3289.395 374.495 ;
        RECT 3289.825 374.215 3290.105 374.495 ;
        RECT 3290.535 374.215 3290.815 374.495 ;
        RECT 3291.245 374.215 3291.525 374.495 ;
        RECT 3291.955 374.215 3292.235 374.495 ;
        RECT 3292.665 374.215 3292.945 374.495 ;
        RECT 3293.375 374.215 3293.655 374.495 ;
        RECT 3294.085 374.215 3294.365 374.495 ;
        RECT 3294.795 374.215 3295.075 374.495 ;
        RECT 3295.505 374.215 3295.785 374.495 ;
        RECT 3296.215 374.215 3296.495 374.495 ;
        RECT 3296.925 374.215 3297.205 374.495 ;
        RECT 3297.635 374.215 3297.915 374.495 ;
        RECT 3298.345 374.215 3298.625 374.495 ;
        RECT 3289.115 373.505 3289.395 373.785 ;
        RECT 3289.825 373.505 3290.105 373.785 ;
        RECT 3290.535 373.505 3290.815 373.785 ;
        RECT 3291.245 373.505 3291.525 373.785 ;
        RECT 3291.955 373.505 3292.235 373.785 ;
        RECT 3292.665 373.505 3292.945 373.785 ;
        RECT 3293.375 373.505 3293.655 373.785 ;
        RECT 3294.085 373.505 3294.365 373.785 ;
        RECT 3294.795 373.505 3295.075 373.785 ;
        RECT 3295.505 373.505 3295.785 373.785 ;
        RECT 3296.215 373.505 3296.495 373.785 ;
        RECT 3296.925 373.505 3297.205 373.785 ;
        RECT 3297.635 373.505 3297.915 373.785 ;
        RECT 3298.345 373.505 3298.625 373.785 ;
        RECT 3289.115 372.795 3289.395 373.075 ;
        RECT 3289.825 372.795 3290.105 373.075 ;
        RECT 3290.535 372.795 3290.815 373.075 ;
        RECT 3291.245 372.795 3291.525 373.075 ;
        RECT 3291.955 372.795 3292.235 373.075 ;
        RECT 3292.665 372.795 3292.945 373.075 ;
        RECT 3293.375 372.795 3293.655 373.075 ;
        RECT 3294.085 372.795 3294.365 373.075 ;
        RECT 3294.795 372.795 3295.075 373.075 ;
        RECT 3295.505 372.795 3295.785 373.075 ;
        RECT 3296.215 372.795 3296.495 373.075 ;
        RECT 3296.925 372.795 3297.205 373.075 ;
        RECT 3297.635 372.795 3297.915 373.075 ;
        RECT 3298.345 372.795 3298.625 373.075 ;
        RECT 3300.965 379.895 3301.245 380.175 ;
        RECT 3301.675 379.895 3301.955 380.175 ;
        RECT 3302.385 379.895 3302.665 380.175 ;
        RECT 3303.095 379.895 3303.375 380.175 ;
        RECT 3303.805 379.895 3304.085 380.175 ;
        RECT 3304.515 379.895 3304.795 380.175 ;
        RECT 3305.225 379.895 3305.505 380.175 ;
        RECT 3305.935 379.895 3306.215 380.175 ;
        RECT 3306.645 379.895 3306.925 380.175 ;
        RECT 3307.355 379.895 3307.635 380.175 ;
        RECT 3308.065 379.895 3308.345 380.175 ;
        RECT 3308.775 379.895 3309.055 380.175 ;
        RECT 3309.485 379.895 3309.765 380.175 ;
        RECT 3310.195 379.895 3310.475 380.175 ;
        RECT 3300.965 379.185 3301.245 379.465 ;
        RECT 3301.675 379.185 3301.955 379.465 ;
        RECT 3302.385 379.185 3302.665 379.465 ;
        RECT 3303.095 379.185 3303.375 379.465 ;
        RECT 3303.805 379.185 3304.085 379.465 ;
        RECT 3304.515 379.185 3304.795 379.465 ;
        RECT 3305.225 379.185 3305.505 379.465 ;
        RECT 3305.935 379.185 3306.215 379.465 ;
        RECT 3306.645 379.185 3306.925 379.465 ;
        RECT 3307.355 379.185 3307.635 379.465 ;
        RECT 3308.065 379.185 3308.345 379.465 ;
        RECT 3308.775 379.185 3309.055 379.465 ;
        RECT 3309.485 379.185 3309.765 379.465 ;
        RECT 3310.195 379.185 3310.475 379.465 ;
        RECT 3300.965 378.475 3301.245 378.755 ;
        RECT 3301.675 378.475 3301.955 378.755 ;
        RECT 3302.385 378.475 3302.665 378.755 ;
        RECT 3303.095 378.475 3303.375 378.755 ;
        RECT 3303.805 378.475 3304.085 378.755 ;
        RECT 3304.515 378.475 3304.795 378.755 ;
        RECT 3305.225 378.475 3305.505 378.755 ;
        RECT 3305.935 378.475 3306.215 378.755 ;
        RECT 3306.645 378.475 3306.925 378.755 ;
        RECT 3307.355 378.475 3307.635 378.755 ;
        RECT 3308.065 378.475 3308.345 378.755 ;
        RECT 3308.775 378.475 3309.055 378.755 ;
        RECT 3309.485 378.475 3309.765 378.755 ;
        RECT 3310.195 378.475 3310.475 378.755 ;
        RECT 3300.965 377.765 3301.245 378.045 ;
        RECT 3301.675 377.765 3301.955 378.045 ;
        RECT 3302.385 377.765 3302.665 378.045 ;
        RECT 3303.095 377.765 3303.375 378.045 ;
        RECT 3303.805 377.765 3304.085 378.045 ;
        RECT 3304.515 377.765 3304.795 378.045 ;
        RECT 3305.225 377.765 3305.505 378.045 ;
        RECT 3305.935 377.765 3306.215 378.045 ;
        RECT 3306.645 377.765 3306.925 378.045 ;
        RECT 3307.355 377.765 3307.635 378.045 ;
        RECT 3308.065 377.765 3308.345 378.045 ;
        RECT 3308.775 377.765 3309.055 378.045 ;
        RECT 3309.485 377.765 3309.765 378.045 ;
        RECT 3310.195 377.765 3310.475 378.045 ;
        RECT 3300.965 377.055 3301.245 377.335 ;
        RECT 3301.675 377.055 3301.955 377.335 ;
        RECT 3302.385 377.055 3302.665 377.335 ;
        RECT 3303.095 377.055 3303.375 377.335 ;
        RECT 3303.805 377.055 3304.085 377.335 ;
        RECT 3304.515 377.055 3304.795 377.335 ;
        RECT 3305.225 377.055 3305.505 377.335 ;
        RECT 3305.935 377.055 3306.215 377.335 ;
        RECT 3306.645 377.055 3306.925 377.335 ;
        RECT 3307.355 377.055 3307.635 377.335 ;
        RECT 3308.065 377.055 3308.345 377.335 ;
        RECT 3308.775 377.055 3309.055 377.335 ;
        RECT 3309.485 377.055 3309.765 377.335 ;
        RECT 3310.195 377.055 3310.475 377.335 ;
        RECT 3300.965 376.345 3301.245 376.625 ;
        RECT 3301.675 376.345 3301.955 376.625 ;
        RECT 3302.385 376.345 3302.665 376.625 ;
        RECT 3303.095 376.345 3303.375 376.625 ;
        RECT 3303.805 376.345 3304.085 376.625 ;
        RECT 3304.515 376.345 3304.795 376.625 ;
        RECT 3305.225 376.345 3305.505 376.625 ;
        RECT 3305.935 376.345 3306.215 376.625 ;
        RECT 3306.645 376.345 3306.925 376.625 ;
        RECT 3307.355 376.345 3307.635 376.625 ;
        RECT 3308.065 376.345 3308.345 376.625 ;
        RECT 3308.775 376.345 3309.055 376.625 ;
        RECT 3309.485 376.345 3309.765 376.625 ;
        RECT 3310.195 376.345 3310.475 376.625 ;
        RECT 3300.965 375.635 3301.245 375.915 ;
        RECT 3301.675 375.635 3301.955 375.915 ;
        RECT 3302.385 375.635 3302.665 375.915 ;
        RECT 3303.095 375.635 3303.375 375.915 ;
        RECT 3303.805 375.635 3304.085 375.915 ;
        RECT 3304.515 375.635 3304.795 375.915 ;
        RECT 3305.225 375.635 3305.505 375.915 ;
        RECT 3305.935 375.635 3306.215 375.915 ;
        RECT 3306.645 375.635 3306.925 375.915 ;
        RECT 3307.355 375.635 3307.635 375.915 ;
        RECT 3308.065 375.635 3308.345 375.915 ;
        RECT 3308.775 375.635 3309.055 375.915 ;
        RECT 3309.485 375.635 3309.765 375.915 ;
        RECT 3310.195 375.635 3310.475 375.915 ;
        RECT 3300.965 374.925 3301.245 375.205 ;
        RECT 3301.675 374.925 3301.955 375.205 ;
        RECT 3302.385 374.925 3302.665 375.205 ;
        RECT 3303.095 374.925 3303.375 375.205 ;
        RECT 3303.805 374.925 3304.085 375.205 ;
        RECT 3304.515 374.925 3304.795 375.205 ;
        RECT 3305.225 374.925 3305.505 375.205 ;
        RECT 3305.935 374.925 3306.215 375.205 ;
        RECT 3306.645 374.925 3306.925 375.205 ;
        RECT 3307.355 374.925 3307.635 375.205 ;
        RECT 3308.065 374.925 3308.345 375.205 ;
        RECT 3308.775 374.925 3309.055 375.205 ;
        RECT 3309.485 374.925 3309.765 375.205 ;
        RECT 3310.195 374.925 3310.475 375.205 ;
        RECT 3300.965 374.215 3301.245 374.495 ;
        RECT 3301.675 374.215 3301.955 374.495 ;
        RECT 3302.385 374.215 3302.665 374.495 ;
        RECT 3303.095 374.215 3303.375 374.495 ;
        RECT 3303.805 374.215 3304.085 374.495 ;
        RECT 3304.515 374.215 3304.795 374.495 ;
        RECT 3305.225 374.215 3305.505 374.495 ;
        RECT 3305.935 374.215 3306.215 374.495 ;
        RECT 3306.645 374.215 3306.925 374.495 ;
        RECT 3307.355 374.215 3307.635 374.495 ;
        RECT 3308.065 374.215 3308.345 374.495 ;
        RECT 3308.775 374.215 3309.055 374.495 ;
        RECT 3309.485 374.215 3309.765 374.495 ;
        RECT 3310.195 374.215 3310.475 374.495 ;
        RECT 3300.965 373.505 3301.245 373.785 ;
        RECT 3301.675 373.505 3301.955 373.785 ;
        RECT 3302.385 373.505 3302.665 373.785 ;
        RECT 3303.095 373.505 3303.375 373.785 ;
        RECT 3303.805 373.505 3304.085 373.785 ;
        RECT 3304.515 373.505 3304.795 373.785 ;
        RECT 3305.225 373.505 3305.505 373.785 ;
        RECT 3305.935 373.505 3306.215 373.785 ;
        RECT 3306.645 373.505 3306.925 373.785 ;
        RECT 3307.355 373.505 3307.635 373.785 ;
        RECT 3308.065 373.505 3308.345 373.785 ;
        RECT 3308.775 373.505 3309.055 373.785 ;
        RECT 3309.485 373.505 3309.765 373.785 ;
        RECT 3310.195 373.505 3310.475 373.785 ;
        RECT 3300.965 372.795 3301.245 373.075 ;
        RECT 3301.675 372.795 3301.955 373.075 ;
        RECT 3302.385 372.795 3302.665 373.075 ;
        RECT 3303.095 372.795 3303.375 373.075 ;
        RECT 3303.805 372.795 3304.085 373.075 ;
        RECT 3304.515 372.795 3304.795 373.075 ;
        RECT 3305.225 372.795 3305.505 373.075 ;
        RECT 3305.935 372.795 3306.215 373.075 ;
        RECT 3306.645 372.795 3306.925 373.075 ;
        RECT 3307.355 372.795 3307.635 373.075 ;
        RECT 3308.065 372.795 3308.345 373.075 ;
        RECT 3308.775 372.795 3309.055 373.075 ;
        RECT 3309.485 372.795 3309.765 373.075 ;
        RECT 3310.195 372.795 3310.475 373.075 ;
        RECT 3314.495 379.895 3314.775 380.175 ;
        RECT 3315.205 379.895 3315.485 380.175 ;
        RECT 3315.915 379.895 3316.195 380.175 ;
        RECT 3316.625 379.895 3316.905 380.175 ;
        RECT 3317.335 379.895 3317.615 380.175 ;
        RECT 3318.045 379.895 3318.325 380.175 ;
        RECT 3318.755 379.895 3319.035 380.175 ;
        RECT 3319.465 379.895 3319.745 380.175 ;
        RECT 3320.175 379.895 3320.455 380.175 ;
        RECT 3320.885 379.895 3321.165 380.175 ;
        RECT 3321.595 379.895 3321.875 380.175 ;
        RECT 3322.305 379.895 3322.585 380.175 ;
        RECT 3323.015 379.895 3323.295 380.175 ;
        RECT 3323.725 379.895 3324.005 380.175 ;
        RECT 3314.495 379.185 3314.775 379.465 ;
        RECT 3315.205 379.185 3315.485 379.465 ;
        RECT 3315.915 379.185 3316.195 379.465 ;
        RECT 3316.625 379.185 3316.905 379.465 ;
        RECT 3317.335 379.185 3317.615 379.465 ;
        RECT 3318.045 379.185 3318.325 379.465 ;
        RECT 3318.755 379.185 3319.035 379.465 ;
        RECT 3319.465 379.185 3319.745 379.465 ;
        RECT 3320.175 379.185 3320.455 379.465 ;
        RECT 3320.885 379.185 3321.165 379.465 ;
        RECT 3321.595 379.185 3321.875 379.465 ;
        RECT 3322.305 379.185 3322.585 379.465 ;
        RECT 3323.015 379.185 3323.295 379.465 ;
        RECT 3323.725 379.185 3324.005 379.465 ;
        RECT 3314.495 378.475 3314.775 378.755 ;
        RECT 3315.205 378.475 3315.485 378.755 ;
        RECT 3315.915 378.475 3316.195 378.755 ;
        RECT 3316.625 378.475 3316.905 378.755 ;
        RECT 3317.335 378.475 3317.615 378.755 ;
        RECT 3318.045 378.475 3318.325 378.755 ;
        RECT 3318.755 378.475 3319.035 378.755 ;
        RECT 3319.465 378.475 3319.745 378.755 ;
        RECT 3320.175 378.475 3320.455 378.755 ;
        RECT 3320.885 378.475 3321.165 378.755 ;
        RECT 3321.595 378.475 3321.875 378.755 ;
        RECT 3322.305 378.475 3322.585 378.755 ;
        RECT 3323.015 378.475 3323.295 378.755 ;
        RECT 3323.725 378.475 3324.005 378.755 ;
        RECT 3314.495 377.765 3314.775 378.045 ;
        RECT 3315.205 377.765 3315.485 378.045 ;
        RECT 3315.915 377.765 3316.195 378.045 ;
        RECT 3316.625 377.765 3316.905 378.045 ;
        RECT 3317.335 377.765 3317.615 378.045 ;
        RECT 3318.045 377.765 3318.325 378.045 ;
        RECT 3318.755 377.765 3319.035 378.045 ;
        RECT 3319.465 377.765 3319.745 378.045 ;
        RECT 3320.175 377.765 3320.455 378.045 ;
        RECT 3320.885 377.765 3321.165 378.045 ;
        RECT 3321.595 377.765 3321.875 378.045 ;
        RECT 3322.305 377.765 3322.585 378.045 ;
        RECT 3323.015 377.765 3323.295 378.045 ;
        RECT 3323.725 377.765 3324.005 378.045 ;
        RECT 3314.495 377.055 3314.775 377.335 ;
        RECT 3315.205 377.055 3315.485 377.335 ;
        RECT 3315.915 377.055 3316.195 377.335 ;
        RECT 3316.625 377.055 3316.905 377.335 ;
        RECT 3317.335 377.055 3317.615 377.335 ;
        RECT 3318.045 377.055 3318.325 377.335 ;
        RECT 3318.755 377.055 3319.035 377.335 ;
        RECT 3319.465 377.055 3319.745 377.335 ;
        RECT 3320.175 377.055 3320.455 377.335 ;
        RECT 3320.885 377.055 3321.165 377.335 ;
        RECT 3321.595 377.055 3321.875 377.335 ;
        RECT 3322.305 377.055 3322.585 377.335 ;
        RECT 3323.015 377.055 3323.295 377.335 ;
        RECT 3323.725 377.055 3324.005 377.335 ;
        RECT 3314.495 376.345 3314.775 376.625 ;
        RECT 3315.205 376.345 3315.485 376.625 ;
        RECT 3315.915 376.345 3316.195 376.625 ;
        RECT 3316.625 376.345 3316.905 376.625 ;
        RECT 3317.335 376.345 3317.615 376.625 ;
        RECT 3318.045 376.345 3318.325 376.625 ;
        RECT 3318.755 376.345 3319.035 376.625 ;
        RECT 3319.465 376.345 3319.745 376.625 ;
        RECT 3320.175 376.345 3320.455 376.625 ;
        RECT 3320.885 376.345 3321.165 376.625 ;
        RECT 3321.595 376.345 3321.875 376.625 ;
        RECT 3322.305 376.345 3322.585 376.625 ;
        RECT 3323.015 376.345 3323.295 376.625 ;
        RECT 3323.725 376.345 3324.005 376.625 ;
        RECT 3314.495 375.635 3314.775 375.915 ;
        RECT 3315.205 375.635 3315.485 375.915 ;
        RECT 3315.915 375.635 3316.195 375.915 ;
        RECT 3316.625 375.635 3316.905 375.915 ;
        RECT 3317.335 375.635 3317.615 375.915 ;
        RECT 3318.045 375.635 3318.325 375.915 ;
        RECT 3318.755 375.635 3319.035 375.915 ;
        RECT 3319.465 375.635 3319.745 375.915 ;
        RECT 3320.175 375.635 3320.455 375.915 ;
        RECT 3320.885 375.635 3321.165 375.915 ;
        RECT 3321.595 375.635 3321.875 375.915 ;
        RECT 3322.305 375.635 3322.585 375.915 ;
        RECT 3323.015 375.635 3323.295 375.915 ;
        RECT 3323.725 375.635 3324.005 375.915 ;
        RECT 3314.495 374.925 3314.775 375.205 ;
        RECT 3315.205 374.925 3315.485 375.205 ;
        RECT 3315.915 374.925 3316.195 375.205 ;
        RECT 3316.625 374.925 3316.905 375.205 ;
        RECT 3317.335 374.925 3317.615 375.205 ;
        RECT 3318.045 374.925 3318.325 375.205 ;
        RECT 3318.755 374.925 3319.035 375.205 ;
        RECT 3319.465 374.925 3319.745 375.205 ;
        RECT 3320.175 374.925 3320.455 375.205 ;
        RECT 3320.885 374.925 3321.165 375.205 ;
        RECT 3321.595 374.925 3321.875 375.205 ;
        RECT 3322.305 374.925 3322.585 375.205 ;
        RECT 3323.015 374.925 3323.295 375.205 ;
        RECT 3323.725 374.925 3324.005 375.205 ;
        RECT 3314.495 374.215 3314.775 374.495 ;
        RECT 3315.205 374.215 3315.485 374.495 ;
        RECT 3315.915 374.215 3316.195 374.495 ;
        RECT 3316.625 374.215 3316.905 374.495 ;
        RECT 3317.335 374.215 3317.615 374.495 ;
        RECT 3318.045 374.215 3318.325 374.495 ;
        RECT 3318.755 374.215 3319.035 374.495 ;
        RECT 3319.465 374.215 3319.745 374.495 ;
        RECT 3320.175 374.215 3320.455 374.495 ;
        RECT 3320.885 374.215 3321.165 374.495 ;
        RECT 3321.595 374.215 3321.875 374.495 ;
        RECT 3322.305 374.215 3322.585 374.495 ;
        RECT 3323.015 374.215 3323.295 374.495 ;
        RECT 3323.725 374.215 3324.005 374.495 ;
        RECT 3314.495 373.505 3314.775 373.785 ;
        RECT 3315.205 373.505 3315.485 373.785 ;
        RECT 3315.915 373.505 3316.195 373.785 ;
        RECT 3316.625 373.505 3316.905 373.785 ;
        RECT 3317.335 373.505 3317.615 373.785 ;
        RECT 3318.045 373.505 3318.325 373.785 ;
        RECT 3318.755 373.505 3319.035 373.785 ;
        RECT 3319.465 373.505 3319.745 373.785 ;
        RECT 3320.175 373.505 3320.455 373.785 ;
        RECT 3320.885 373.505 3321.165 373.785 ;
        RECT 3321.595 373.505 3321.875 373.785 ;
        RECT 3322.305 373.505 3322.585 373.785 ;
        RECT 3323.015 373.505 3323.295 373.785 ;
        RECT 3323.725 373.505 3324.005 373.785 ;
        RECT 3314.495 372.795 3314.775 373.075 ;
        RECT 3315.205 372.795 3315.485 373.075 ;
        RECT 3315.915 372.795 3316.195 373.075 ;
        RECT 3316.625 372.795 3316.905 373.075 ;
        RECT 3317.335 372.795 3317.615 373.075 ;
        RECT 3318.045 372.795 3318.325 373.075 ;
        RECT 3318.755 372.795 3319.035 373.075 ;
        RECT 3319.465 372.795 3319.745 373.075 ;
        RECT 3320.175 372.795 3320.455 373.075 ;
        RECT 3320.885 372.795 3321.165 373.075 ;
        RECT 3321.595 372.795 3321.875 373.075 ;
        RECT 3322.305 372.795 3322.585 373.075 ;
        RECT 3323.015 372.795 3323.295 373.075 ;
        RECT 3323.725 372.795 3324.005 373.075 ;
        RECT 3326.345 379.895 3326.625 380.175 ;
        RECT 3327.055 379.895 3327.335 380.175 ;
        RECT 3327.765 379.895 3328.045 380.175 ;
        RECT 3328.475 379.895 3328.755 380.175 ;
        RECT 3329.185 379.895 3329.465 380.175 ;
        RECT 3329.895 379.895 3330.175 380.175 ;
        RECT 3330.605 379.895 3330.885 380.175 ;
        RECT 3331.315 379.895 3331.595 380.175 ;
        RECT 3332.025 379.895 3332.305 380.175 ;
        RECT 3332.735 379.895 3333.015 380.175 ;
        RECT 3333.445 379.895 3333.725 380.175 ;
        RECT 3334.155 379.895 3334.435 380.175 ;
        RECT 3334.865 379.895 3335.145 380.175 ;
        RECT 3335.575 379.895 3335.855 380.175 ;
        RECT 3326.345 379.185 3326.625 379.465 ;
        RECT 3327.055 379.185 3327.335 379.465 ;
        RECT 3327.765 379.185 3328.045 379.465 ;
        RECT 3328.475 379.185 3328.755 379.465 ;
        RECT 3329.185 379.185 3329.465 379.465 ;
        RECT 3329.895 379.185 3330.175 379.465 ;
        RECT 3330.605 379.185 3330.885 379.465 ;
        RECT 3331.315 379.185 3331.595 379.465 ;
        RECT 3332.025 379.185 3332.305 379.465 ;
        RECT 3332.735 379.185 3333.015 379.465 ;
        RECT 3333.445 379.185 3333.725 379.465 ;
        RECT 3334.155 379.185 3334.435 379.465 ;
        RECT 3334.865 379.185 3335.145 379.465 ;
        RECT 3335.575 379.185 3335.855 379.465 ;
        RECT 3326.345 378.475 3326.625 378.755 ;
        RECT 3327.055 378.475 3327.335 378.755 ;
        RECT 3327.765 378.475 3328.045 378.755 ;
        RECT 3328.475 378.475 3328.755 378.755 ;
        RECT 3329.185 378.475 3329.465 378.755 ;
        RECT 3329.895 378.475 3330.175 378.755 ;
        RECT 3330.605 378.475 3330.885 378.755 ;
        RECT 3331.315 378.475 3331.595 378.755 ;
        RECT 3332.025 378.475 3332.305 378.755 ;
        RECT 3332.735 378.475 3333.015 378.755 ;
        RECT 3333.445 378.475 3333.725 378.755 ;
        RECT 3334.155 378.475 3334.435 378.755 ;
        RECT 3334.865 378.475 3335.145 378.755 ;
        RECT 3335.575 378.475 3335.855 378.755 ;
        RECT 3326.345 377.765 3326.625 378.045 ;
        RECT 3327.055 377.765 3327.335 378.045 ;
        RECT 3327.765 377.765 3328.045 378.045 ;
        RECT 3328.475 377.765 3328.755 378.045 ;
        RECT 3329.185 377.765 3329.465 378.045 ;
        RECT 3329.895 377.765 3330.175 378.045 ;
        RECT 3330.605 377.765 3330.885 378.045 ;
        RECT 3331.315 377.765 3331.595 378.045 ;
        RECT 3332.025 377.765 3332.305 378.045 ;
        RECT 3332.735 377.765 3333.015 378.045 ;
        RECT 3333.445 377.765 3333.725 378.045 ;
        RECT 3334.155 377.765 3334.435 378.045 ;
        RECT 3334.865 377.765 3335.145 378.045 ;
        RECT 3335.575 377.765 3335.855 378.045 ;
        RECT 3326.345 377.055 3326.625 377.335 ;
        RECT 3327.055 377.055 3327.335 377.335 ;
        RECT 3327.765 377.055 3328.045 377.335 ;
        RECT 3328.475 377.055 3328.755 377.335 ;
        RECT 3329.185 377.055 3329.465 377.335 ;
        RECT 3329.895 377.055 3330.175 377.335 ;
        RECT 3330.605 377.055 3330.885 377.335 ;
        RECT 3331.315 377.055 3331.595 377.335 ;
        RECT 3332.025 377.055 3332.305 377.335 ;
        RECT 3332.735 377.055 3333.015 377.335 ;
        RECT 3333.445 377.055 3333.725 377.335 ;
        RECT 3334.155 377.055 3334.435 377.335 ;
        RECT 3334.865 377.055 3335.145 377.335 ;
        RECT 3335.575 377.055 3335.855 377.335 ;
        RECT 3326.345 376.345 3326.625 376.625 ;
        RECT 3327.055 376.345 3327.335 376.625 ;
        RECT 3327.765 376.345 3328.045 376.625 ;
        RECT 3328.475 376.345 3328.755 376.625 ;
        RECT 3329.185 376.345 3329.465 376.625 ;
        RECT 3329.895 376.345 3330.175 376.625 ;
        RECT 3330.605 376.345 3330.885 376.625 ;
        RECT 3331.315 376.345 3331.595 376.625 ;
        RECT 3332.025 376.345 3332.305 376.625 ;
        RECT 3332.735 376.345 3333.015 376.625 ;
        RECT 3333.445 376.345 3333.725 376.625 ;
        RECT 3334.155 376.345 3334.435 376.625 ;
        RECT 3334.865 376.345 3335.145 376.625 ;
        RECT 3335.575 376.345 3335.855 376.625 ;
        RECT 3326.345 375.635 3326.625 375.915 ;
        RECT 3327.055 375.635 3327.335 375.915 ;
        RECT 3327.765 375.635 3328.045 375.915 ;
        RECT 3328.475 375.635 3328.755 375.915 ;
        RECT 3329.185 375.635 3329.465 375.915 ;
        RECT 3329.895 375.635 3330.175 375.915 ;
        RECT 3330.605 375.635 3330.885 375.915 ;
        RECT 3331.315 375.635 3331.595 375.915 ;
        RECT 3332.025 375.635 3332.305 375.915 ;
        RECT 3332.735 375.635 3333.015 375.915 ;
        RECT 3333.445 375.635 3333.725 375.915 ;
        RECT 3334.155 375.635 3334.435 375.915 ;
        RECT 3334.865 375.635 3335.145 375.915 ;
        RECT 3335.575 375.635 3335.855 375.915 ;
        RECT 3326.345 374.925 3326.625 375.205 ;
        RECT 3327.055 374.925 3327.335 375.205 ;
        RECT 3327.765 374.925 3328.045 375.205 ;
        RECT 3328.475 374.925 3328.755 375.205 ;
        RECT 3329.185 374.925 3329.465 375.205 ;
        RECT 3329.895 374.925 3330.175 375.205 ;
        RECT 3330.605 374.925 3330.885 375.205 ;
        RECT 3331.315 374.925 3331.595 375.205 ;
        RECT 3332.025 374.925 3332.305 375.205 ;
        RECT 3332.735 374.925 3333.015 375.205 ;
        RECT 3333.445 374.925 3333.725 375.205 ;
        RECT 3334.155 374.925 3334.435 375.205 ;
        RECT 3334.865 374.925 3335.145 375.205 ;
        RECT 3335.575 374.925 3335.855 375.205 ;
        RECT 3326.345 374.215 3326.625 374.495 ;
        RECT 3327.055 374.215 3327.335 374.495 ;
        RECT 3327.765 374.215 3328.045 374.495 ;
        RECT 3328.475 374.215 3328.755 374.495 ;
        RECT 3329.185 374.215 3329.465 374.495 ;
        RECT 3329.895 374.215 3330.175 374.495 ;
        RECT 3330.605 374.215 3330.885 374.495 ;
        RECT 3331.315 374.215 3331.595 374.495 ;
        RECT 3332.025 374.215 3332.305 374.495 ;
        RECT 3332.735 374.215 3333.015 374.495 ;
        RECT 3333.445 374.215 3333.725 374.495 ;
        RECT 3334.155 374.215 3334.435 374.495 ;
        RECT 3334.865 374.215 3335.145 374.495 ;
        RECT 3335.575 374.215 3335.855 374.495 ;
        RECT 3326.345 373.505 3326.625 373.785 ;
        RECT 3327.055 373.505 3327.335 373.785 ;
        RECT 3327.765 373.505 3328.045 373.785 ;
        RECT 3328.475 373.505 3328.755 373.785 ;
        RECT 3329.185 373.505 3329.465 373.785 ;
        RECT 3329.895 373.505 3330.175 373.785 ;
        RECT 3330.605 373.505 3330.885 373.785 ;
        RECT 3331.315 373.505 3331.595 373.785 ;
        RECT 3332.025 373.505 3332.305 373.785 ;
        RECT 3332.735 373.505 3333.015 373.785 ;
        RECT 3333.445 373.505 3333.725 373.785 ;
        RECT 3334.155 373.505 3334.435 373.785 ;
        RECT 3334.865 373.505 3335.145 373.785 ;
        RECT 3335.575 373.505 3335.855 373.785 ;
        RECT 3326.345 372.795 3326.625 373.075 ;
        RECT 3327.055 372.795 3327.335 373.075 ;
        RECT 3327.765 372.795 3328.045 373.075 ;
        RECT 3328.475 372.795 3328.755 373.075 ;
        RECT 3329.185 372.795 3329.465 373.075 ;
        RECT 3329.895 372.795 3330.175 373.075 ;
        RECT 3330.605 372.795 3330.885 373.075 ;
        RECT 3331.315 372.795 3331.595 373.075 ;
        RECT 3332.025 372.795 3332.305 373.075 ;
        RECT 3332.735 372.795 3333.015 373.075 ;
        RECT 3333.445 372.795 3333.725 373.075 ;
        RECT 3334.155 372.795 3334.435 373.075 ;
        RECT 3334.865 372.795 3335.145 373.075 ;
        RECT 3335.575 372.795 3335.855 373.075 ;
        RECT 3339.495 379.895 3339.775 380.175 ;
        RECT 3340.205 379.895 3340.485 380.175 ;
        RECT 3340.915 379.895 3341.195 380.175 ;
        RECT 3341.625 379.895 3341.905 380.175 ;
        RECT 3342.335 379.895 3342.615 380.175 ;
        RECT 3343.045 379.895 3343.325 380.175 ;
        RECT 3343.755 379.895 3344.035 380.175 ;
        RECT 3344.465 379.895 3344.745 380.175 ;
        RECT 3345.175 379.895 3345.455 380.175 ;
        RECT 3345.885 379.895 3346.165 380.175 ;
        RECT 3346.595 379.895 3346.875 380.175 ;
        RECT 3347.305 379.895 3347.585 380.175 ;
        RECT 3348.015 379.895 3348.295 380.175 ;
        RECT 3339.495 379.185 3339.775 379.465 ;
        RECT 3340.205 379.185 3340.485 379.465 ;
        RECT 3340.915 379.185 3341.195 379.465 ;
        RECT 3341.625 379.185 3341.905 379.465 ;
        RECT 3342.335 379.185 3342.615 379.465 ;
        RECT 3343.045 379.185 3343.325 379.465 ;
        RECT 3343.755 379.185 3344.035 379.465 ;
        RECT 3344.465 379.185 3344.745 379.465 ;
        RECT 3345.175 379.185 3345.455 379.465 ;
        RECT 3345.885 379.185 3346.165 379.465 ;
        RECT 3346.595 379.185 3346.875 379.465 ;
        RECT 3347.305 379.185 3347.585 379.465 ;
        RECT 3348.015 379.185 3348.295 379.465 ;
        RECT 3339.495 378.475 3339.775 378.755 ;
        RECT 3340.205 378.475 3340.485 378.755 ;
        RECT 3340.915 378.475 3341.195 378.755 ;
        RECT 3341.625 378.475 3341.905 378.755 ;
        RECT 3342.335 378.475 3342.615 378.755 ;
        RECT 3343.045 378.475 3343.325 378.755 ;
        RECT 3343.755 378.475 3344.035 378.755 ;
        RECT 3344.465 378.475 3344.745 378.755 ;
        RECT 3345.175 378.475 3345.455 378.755 ;
        RECT 3345.885 378.475 3346.165 378.755 ;
        RECT 3346.595 378.475 3346.875 378.755 ;
        RECT 3347.305 378.475 3347.585 378.755 ;
        RECT 3348.015 378.475 3348.295 378.755 ;
        RECT 3339.495 377.765 3339.775 378.045 ;
        RECT 3340.205 377.765 3340.485 378.045 ;
        RECT 3340.915 377.765 3341.195 378.045 ;
        RECT 3341.625 377.765 3341.905 378.045 ;
        RECT 3342.335 377.765 3342.615 378.045 ;
        RECT 3343.045 377.765 3343.325 378.045 ;
        RECT 3343.755 377.765 3344.035 378.045 ;
        RECT 3344.465 377.765 3344.745 378.045 ;
        RECT 3345.175 377.765 3345.455 378.045 ;
        RECT 3345.885 377.765 3346.165 378.045 ;
        RECT 3346.595 377.765 3346.875 378.045 ;
        RECT 3347.305 377.765 3347.585 378.045 ;
        RECT 3348.015 377.765 3348.295 378.045 ;
        RECT 3339.495 377.055 3339.775 377.335 ;
        RECT 3340.205 377.055 3340.485 377.335 ;
        RECT 3340.915 377.055 3341.195 377.335 ;
        RECT 3341.625 377.055 3341.905 377.335 ;
        RECT 3342.335 377.055 3342.615 377.335 ;
        RECT 3343.045 377.055 3343.325 377.335 ;
        RECT 3343.755 377.055 3344.035 377.335 ;
        RECT 3344.465 377.055 3344.745 377.335 ;
        RECT 3345.175 377.055 3345.455 377.335 ;
        RECT 3345.885 377.055 3346.165 377.335 ;
        RECT 3346.595 377.055 3346.875 377.335 ;
        RECT 3347.305 377.055 3347.585 377.335 ;
        RECT 3348.015 377.055 3348.295 377.335 ;
        RECT 3339.495 376.345 3339.775 376.625 ;
        RECT 3340.205 376.345 3340.485 376.625 ;
        RECT 3340.915 376.345 3341.195 376.625 ;
        RECT 3341.625 376.345 3341.905 376.625 ;
        RECT 3342.335 376.345 3342.615 376.625 ;
        RECT 3343.045 376.345 3343.325 376.625 ;
        RECT 3343.755 376.345 3344.035 376.625 ;
        RECT 3344.465 376.345 3344.745 376.625 ;
        RECT 3345.175 376.345 3345.455 376.625 ;
        RECT 3345.885 376.345 3346.165 376.625 ;
        RECT 3346.595 376.345 3346.875 376.625 ;
        RECT 3347.305 376.345 3347.585 376.625 ;
        RECT 3348.015 376.345 3348.295 376.625 ;
        RECT 3339.495 375.635 3339.775 375.915 ;
        RECT 3340.205 375.635 3340.485 375.915 ;
        RECT 3340.915 375.635 3341.195 375.915 ;
        RECT 3341.625 375.635 3341.905 375.915 ;
        RECT 3342.335 375.635 3342.615 375.915 ;
        RECT 3343.045 375.635 3343.325 375.915 ;
        RECT 3343.755 375.635 3344.035 375.915 ;
        RECT 3344.465 375.635 3344.745 375.915 ;
        RECT 3345.175 375.635 3345.455 375.915 ;
        RECT 3345.885 375.635 3346.165 375.915 ;
        RECT 3346.595 375.635 3346.875 375.915 ;
        RECT 3347.305 375.635 3347.585 375.915 ;
        RECT 3348.015 375.635 3348.295 375.915 ;
        RECT 3339.495 374.925 3339.775 375.205 ;
        RECT 3340.205 374.925 3340.485 375.205 ;
        RECT 3340.915 374.925 3341.195 375.205 ;
        RECT 3341.625 374.925 3341.905 375.205 ;
        RECT 3342.335 374.925 3342.615 375.205 ;
        RECT 3343.045 374.925 3343.325 375.205 ;
        RECT 3343.755 374.925 3344.035 375.205 ;
        RECT 3344.465 374.925 3344.745 375.205 ;
        RECT 3345.175 374.925 3345.455 375.205 ;
        RECT 3345.885 374.925 3346.165 375.205 ;
        RECT 3346.595 374.925 3346.875 375.205 ;
        RECT 3347.305 374.925 3347.585 375.205 ;
        RECT 3348.015 374.925 3348.295 375.205 ;
        RECT 3339.495 374.215 3339.775 374.495 ;
        RECT 3340.205 374.215 3340.485 374.495 ;
        RECT 3340.915 374.215 3341.195 374.495 ;
        RECT 3341.625 374.215 3341.905 374.495 ;
        RECT 3342.335 374.215 3342.615 374.495 ;
        RECT 3343.045 374.215 3343.325 374.495 ;
        RECT 3343.755 374.215 3344.035 374.495 ;
        RECT 3344.465 374.215 3344.745 374.495 ;
        RECT 3345.175 374.215 3345.455 374.495 ;
        RECT 3345.885 374.215 3346.165 374.495 ;
        RECT 3346.595 374.215 3346.875 374.495 ;
        RECT 3347.305 374.215 3347.585 374.495 ;
        RECT 3348.015 374.215 3348.295 374.495 ;
        RECT 3339.495 373.505 3339.775 373.785 ;
        RECT 3340.205 373.505 3340.485 373.785 ;
        RECT 3340.915 373.505 3341.195 373.785 ;
        RECT 3341.625 373.505 3341.905 373.785 ;
        RECT 3342.335 373.505 3342.615 373.785 ;
        RECT 3343.045 373.505 3343.325 373.785 ;
        RECT 3343.755 373.505 3344.035 373.785 ;
        RECT 3344.465 373.505 3344.745 373.785 ;
        RECT 3345.175 373.505 3345.455 373.785 ;
        RECT 3345.885 373.505 3346.165 373.785 ;
        RECT 3346.595 373.505 3346.875 373.785 ;
        RECT 3347.305 373.505 3347.585 373.785 ;
        RECT 3348.015 373.505 3348.295 373.785 ;
        RECT 3339.495 372.795 3339.775 373.075 ;
        RECT 3340.205 372.795 3340.485 373.075 ;
        RECT 3340.915 372.795 3341.195 373.075 ;
        RECT 3341.625 372.795 3341.905 373.075 ;
        RECT 3342.335 372.795 3342.615 373.075 ;
        RECT 3343.045 372.795 3343.325 373.075 ;
        RECT 3343.755 372.795 3344.035 373.075 ;
        RECT 3344.465 372.795 3344.745 373.075 ;
        RECT 3345.175 372.795 3345.455 373.075 ;
        RECT 3345.885 372.795 3346.165 373.075 ;
        RECT 3346.595 372.795 3346.875 373.075 ;
        RECT 3347.305 372.795 3347.585 373.075 ;
        RECT 3348.015 372.795 3348.295 373.075 ;
        RECT 526.715 369.895 526.995 370.175 ;
        RECT 527.425 369.895 527.705 370.175 ;
        RECT 528.135 369.895 528.415 370.175 ;
        RECT 528.845 369.895 529.125 370.175 ;
        RECT 529.555 369.895 529.835 370.175 ;
        RECT 530.265 369.895 530.545 370.175 ;
        RECT 530.975 369.895 531.255 370.175 ;
        RECT 531.685 369.895 531.965 370.175 ;
        RECT 532.395 369.895 532.675 370.175 ;
        RECT 533.105 369.895 533.385 370.175 ;
        RECT 533.815 369.895 534.095 370.175 ;
        RECT 534.525 369.895 534.805 370.175 ;
        RECT 535.235 369.895 535.515 370.175 ;
        RECT 526.715 369.185 526.995 369.465 ;
        RECT 527.425 369.185 527.705 369.465 ;
        RECT 528.135 369.185 528.415 369.465 ;
        RECT 528.845 369.185 529.125 369.465 ;
        RECT 529.555 369.185 529.835 369.465 ;
        RECT 530.265 369.185 530.545 369.465 ;
        RECT 530.975 369.185 531.255 369.465 ;
        RECT 531.685 369.185 531.965 369.465 ;
        RECT 532.395 369.185 532.675 369.465 ;
        RECT 533.105 369.185 533.385 369.465 ;
        RECT 533.815 369.185 534.095 369.465 ;
        RECT 534.525 369.185 534.805 369.465 ;
        RECT 535.235 369.185 535.515 369.465 ;
        RECT 526.715 368.475 526.995 368.755 ;
        RECT 527.425 368.475 527.705 368.755 ;
        RECT 528.135 368.475 528.415 368.755 ;
        RECT 528.845 368.475 529.125 368.755 ;
        RECT 529.555 368.475 529.835 368.755 ;
        RECT 530.265 368.475 530.545 368.755 ;
        RECT 530.975 368.475 531.255 368.755 ;
        RECT 531.685 368.475 531.965 368.755 ;
        RECT 532.395 368.475 532.675 368.755 ;
        RECT 533.105 368.475 533.385 368.755 ;
        RECT 533.815 368.475 534.095 368.755 ;
        RECT 534.525 368.475 534.805 368.755 ;
        RECT 535.235 368.475 535.515 368.755 ;
        RECT 526.715 367.765 526.995 368.045 ;
        RECT 527.425 367.765 527.705 368.045 ;
        RECT 528.135 367.765 528.415 368.045 ;
        RECT 528.845 367.765 529.125 368.045 ;
        RECT 529.555 367.765 529.835 368.045 ;
        RECT 530.265 367.765 530.545 368.045 ;
        RECT 530.975 367.765 531.255 368.045 ;
        RECT 531.685 367.765 531.965 368.045 ;
        RECT 532.395 367.765 532.675 368.045 ;
        RECT 533.105 367.765 533.385 368.045 ;
        RECT 533.815 367.765 534.095 368.045 ;
        RECT 534.525 367.765 534.805 368.045 ;
        RECT 535.235 367.765 535.515 368.045 ;
        RECT 526.715 367.055 526.995 367.335 ;
        RECT 527.425 367.055 527.705 367.335 ;
        RECT 528.135 367.055 528.415 367.335 ;
        RECT 528.845 367.055 529.125 367.335 ;
        RECT 529.555 367.055 529.835 367.335 ;
        RECT 530.265 367.055 530.545 367.335 ;
        RECT 530.975 367.055 531.255 367.335 ;
        RECT 531.685 367.055 531.965 367.335 ;
        RECT 532.395 367.055 532.675 367.335 ;
        RECT 533.105 367.055 533.385 367.335 ;
        RECT 533.815 367.055 534.095 367.335 ;
        RECT 534.525 367.055 534.805 367.335 ;
        RECT 535.235 367.055 535.515 367.335 ;
        RECT 526.715 366.345 526.995 366.625 ;
        RECT 527.425 366.345 527.705 366.625 ;
        RECT 528.135 366.345 528.415 366.625 ;
        RECT 528.845 366.345 529.125 366.625 ;
        RECT 529.555 366.345 529.835 366.625 ;
        RECT 530.265 366.345 530.545 366.625 ;
        RECT 530.975 366.345 531.255 366.625 ;
        RECT 531.685 366.345 531.965 366.625 ;
        RECT 532.395 366.345 532.675 366.625 ;
        RECT 533.105 366.345 533.385 366.625 ;
        RECT 533.815 366.345 534.095 366.625 ;
        RECT 534.525 366.345 534.805 366.625 ;
        RECT 535.235 366.345 535.515 366.625 ;
        RECT 526.715 365.635 526.995 365.915 ;
        RECT 527.425 365.635 527.705 365.915 ;
        RECT 528.135 365.635 528.415 365.915 ;
        RECT 528.845 365.635 529.125 365.915 ;
        RECT 529.555 365.635 529.835 365.915 ;
        RECT 530.265 365.635 530.545 365.915 ;
        RECT 530.975 365.635 531.255 365.915 ;
        RECT 531.685 365.635 531.965 365.915 ;
        RECT 532.395 365.635 532.675 365.915 ;
        RECT 533.105 365.635 533.385 365.915 ;
        RECT 533.815 365.635 534.095 365.915 ;
        RECT 534.525 365.635 534.805 365.915 ;
        RECT 535.235 365.635 535.515 365.915 ;
        RECT 526.715 364.925 526.995 365.205 ;
        RECT 527.425 364.925 527.705 365.205 ;
        RECT 528.135 364.925 528.415 365.205 ;
        RECT 528.845 364.925 529.125 365.205 ;
        RECT 529.555 364.925 529.835 365.205 ;
        RECT 530.265 364.925 530.545 365.205 ;
        RECT 530.975 364.925 531.255 365.205 ;
        RECT 531.685 364.925 531.965 365.205 ;
        RECT 532.395 364.925 532.675 365.205 ;
        RECT 533.105 364.925 533.385 365.205 ;
        RECT 533.815 364.925 534.095 365.205 ;
        RECT 534.525 364.925 534.805 365.205 ;
        RECT 535.235 364.925 535.515 365.205 ;
        RECT 526.715 364.215 526.995 364.495 ;
        RECT 527.425 364.215 527.705 364.495 ;
        RECT 528.135 364.215 528.415 364.495 ;
        RECT 528.845 364.215 529.125 364.495 ;
        RECT 529.555 364.215 529.835 364.495 ;
        RECT 530.265 364.215 530.545 364.495 ;
        RECT 530.975 364.215 531.255 364.495 ;
        RECT 531.685 364.215 531.965 364.495 ;
        RECT 532.395 364.215 532.675 364.495 ;
        RECT 533.105 364.215 533.385 364.495 ;
        RECT 533.815 364.215 534.095 364.495 ;
        RECT 534.525 364.215 534.805 364.495 ;
        RECT 535.235 364.215 535.515 364.495 ;
        RECT 526.715 363.505 526.995 363.785 ;
        RECT 527.425 363.505 527.705 363.785 ;
        RECT 528.135 363.505 528.415 363.785 ;
        RECT 528.845 363.505 529.125 363.785 ;
        RECT 529.555 363.505 529.835 363.785 ;
        RECT 530.265 363.505 530.545 363.785 ;
        RECT 530.975 363.505 531.255 363.785 ;
        RECT 531.685 363.505 531.965 363.785 ;
        RECT 532.395 363.505 532.675 363.785 ;
        RECT 533.105 363.505 533.385 363.785 ;
        RECT 533.815 363.505 534.095 363.785 ;
        RECT 534.525 363.505 534.805 363.785 ;
        RECT 535.235 363.505 535.515 363.785 ;
        RECT 526.715 362.795 526.995 363.075 ;
        RECT 527.425 362.795 527.705 363.075 ;
        RECT 528.135 362.795 528.415 363.075 ;
        RECT 528.845 362.795 529.125 363.075 ;
        RECT 529.555 362.795 529.835 363.075 ;
        RECT 530.265 362.795 530.545 363.075 ;
        RECT 530.975 362.795 531.255 363.075 ;
        RECT 531.685 362.795 531.965 363.075 ;
        RECT 532.395 362.795 532.675 363.075 ;
        RECT 533.105 362.795 533.385 363.075 ;
        RECT 533.815 362.795 534.095 363.075 ;
        RECT 534.525 362.795 534.805 363.075 ;
        RECT 535.235 362.795 535.515 363.075 ;
        RECT 526.715 362.085 526.995 362.365 ;
        RECT 527.425 362.085 527.705 362.365 ;
        RECT 528.135 362.085 528.415 362.365 ;
        RECT 528.845 362.085 529.125 362.365 ;
        RECT 529.555 362.085 529.835 362.365 ;
        RECT 530.265 362.085 530.545 362.365 ;
        RECT 530.975 362.085 531.255 362.365 ;
        RECT 531.685 362.085 531.965 362.365 ;
        RECT 532.395 362.085 532.675 362.365 ;
        RECT 533.105 362.085 533.385 362.365 ;
        RECT 533.815 362.085 534.095 362.365 ;
        RECT 534.525 362.085 534.805 362.365 ;
        RECT 535.235 362.085 535.515 362.365 ;
        RECT 526.715 361.375 526.995 361.655 ;
        RECT 527.425 361.375 527.705 361.655 ;
        RECT 528.135 361.375 528.415 361.655 ;
        RECT 528.845 361.375 529.125 361.655 ;
        RECT 529.555 361.375 529.835 361.655 ;
        RECT 530.265 361.375 530.545 361.655 ;
        RECT 530.975 361.375 531.255 361.655 ;
        RECT 531.685 361.375 531.965 361.655 ;
        RECT 532.395 361.375 532.675 361.655 ;
        RECT 533.105 361.375 533.385 361.655 ;
        RECT 533.815 361.375 534.095 361.655 ;
        RECT 534.525 361.375 534.805 361.655 ;
        RECT 535.235 361.375 535.515 361.655 ;
        RECT 526.715 360.665 526.995 360.945 ;
        RECT 527.425 360.665 527.705 360.945 ;
        RECT 528.135 360.665 528.415 360.945 ;
        RECT 528.845 360.665 529.125 360.945 ;
        RECT 529.555 360.665 529.835 360.945 ;
        RECT 530.265 360.665 530.545 360.945 ;
        RECT 530.975 360.665 531.255 360.945 ;
        RECT 531.685 360.665 531.965 360.945 ;
        RECT 532.395 360.665 532.675 360.945 ;
        RECT 533.105 360.665 533.385 360.945 ;
        RECT 533.815 360.665 534.095 360.945 ;
        RECT 534.525 360.665 534.805 360.945 ;
        RECT 535.235 360.665 535.515 360.945 ;
        RECT 544.975 369.895 545.255 370.175 ;
        RECT 545.685 369.895 545.965 370.175 ;
        RECT 546.395 369.895 546.675 370.175 ;
        RECT 547.105 369.895 547.385 370.175 ;
        RECT 547.815 369.895 548.095 370.175 ;
        RECT 548.525 369.895 548.805 370.175 ;
        RECT 544.975 369.185 545.255 369.465 ;
        RECT 545.685 369.185 545.965 369.465 ;
        RECT 546.395 369.185 546.675 369.465 ;
        RECT 547.105 369.185 547.385 369.465 ;
        RECT 547.815 369.185 548.095 369.465 ;
        RECT 548.525 369.185 548.805 369.465 ;
        RECT 544.975 368.475 545.255 368.755 ;
        RECT 545.685 368.475 545.965 368.755 ;
        RECT 546.395 368.475 546.675 368.755 ;
        RECT 547.105 368.475 547.385 368.755 ;
        RECT 547.815 368.475 548.095 368.755 ;
        RECT 548.525 368.475 548.805 368.755 ;
        RECT 544.975 367.765 545.255 368.045 ;
        RECT 545.685 367.765 545.965 368.045 ;
        RECT 546.395 367.765 546.675 368.045 ;
        RECT 547.105 367.765 547.385 368.045 ;
        RECT 547.815 367.765 548.095 368.045 ;
        RECT 548.525 367.765 548.805 368.045 ;
        RECT 544.975 367.055 545.255 367.335 ;
        RECT 545.685 367.055 545.965 367.335 ;
        RECT 546.395 367.055 546.675 367.335 ;
        RECT 547.105 367.055 547.385 367.335 ;
        RECT 547.815 367.055 548.095 367.335 ;
        RECT 548.525 367.055 548.805 367.335 ;
        RECT 544.975 366.345 545.255 366.625 ;
        RECT 545.685 366.345 545.965 366.625 ;
        RECT 546.395 366.345 546.675 366.625 ;
        RECT 547.105 366.345 547.385 366.625 ;
        RECT 547.815 366.345 548.095 366.625 ;
        RECT 548.525 366.345 548.805 366.625 ;
        RECT 544.975 365.635 545.255 365.915 ;
        RECT 545.685 365.635 545.965 365.915 ;
        RECT 546.395 365.635 546.675 365.915 ;
        RECT 547.105 365.635 547.385 365.915 ;
        RECT 547.815 365.635 548.095 365.915 ;
        RECT 548.525 365.635 548.805 365.915 ;
        RECT 544.975 364.925 545.255 365.205 ;
        RECT 545.685 364.925 545.965 365.205 ;
        RECT 546.395 364.925 546.675 365.205 ;
        RECT 547.105 364.925 547.385 365.205 ;
        RECT 547.815 364.925 548.095 365.205 ;
        RECT 548.525 364.925 548.805 365.205 ;
        RECT 544.975 364.215 545.255 364.495 ;
        RECT 545.685 364.215 545.965 364.495 ;
        RECT 546.395 364.215 546.675 364.495 ;
        RECT 547.105 364.215 547.385 364.495 ;
        RECT 547.815 364.215 548.095 364.495 ;
        RECT 548.525 364.215 548.805 364.495 ;
        RECT 544.975 363.505 545.255 363.785 ;
        RECT 545.685 363.505 545.965 363.785 ;
        RECT 546.395 363.505 546.675 363.785 ;
        RECT 547.105 363.505 547.385 363.785 ;
        RECT 547.815 363.505 548.095 363.785 ;
        RECT 548.525 363.505 548.805 363.785 ;
        RECT 544.975 362.795 545.255 363.075 ;
        RECT 545.685 362.795 545.965 363.075 ;
        RECT 546.395 362.795 546.675 363.075 ;
        RECT 547.105 362.795 547.385 363.075 ;
        RECT 547.815 362.795 548.095 363.075 ;
        RECT 548.525 362.795 548.805 363.075 ;
        RECT 544.975 362.085 545.255 362.365 ;
        RECT 545.685 362.085 545.965 362.365 ;
        RECT 546.395 362.085 546.675 362.365 ;
        RECT 547.105 362.085 547.385 362.365 ;
        RECT 547.815 362.085 548.095 362.365 ;
        RECT 548.525 362.085 548.805 362.365 ;
        RECT 544.975 361.375 545.255 361.655 ;
        RECT 545.685 361.375 545.965 361.655 ;
        RECT 546.395 361.375 546.675 361.655 ;
        RECT 547.105 361.375 547.385 361.655 ;
        RECT 547.815 361.375 548.095 361.655 ;
        RECT 548.525 361.375 548.805 361.655 ;
        RECT 544.975 360.665 545.255 360.945 ;
        RECT 545.685 360.665 545.965 360.945 ;
        RECT 546.395 360.665 546.675 360.945 ;
        RECT 547.105 360.665 547.385 360.945 ;
        RECT 547.815 360.665 548.095 360.945 ;
        RECT 548.525 360.665 548.805 360.945 ;
        RECT 550.965 369.895 551.245 370.175 ;
        RECT 551.675 369.895 551.955 370.175 ;
        RECT 552.385 369.895 552.665 370.175 ;
        RECT 553.095 369.895 553.375 370.175 ;
        RECT 553.805 369.895 554.085 370.175 ;
        RECT 554.515 369.895 554.795 370.175 ;
        RECT 555.225 369.895 555.505 370.175 ;
        RECT 555.935 369.895 556.215 370.175 ;
        RECT 556.645 369.895 556.925 370.175 ;
        RECT 557.355 369.895 557.635 370.175 ;
        RECT 558.065 369.895 558.345 370.175 ;
        RECT 558.775 369.895 559.055 370.175 ;
        RECT 559.485 369.895 559.765 370.175 ;
        RECT 560.195 369.895 560.475 370.175 ;
        RECT 550.965 369.185 551.245 369.465 ;
        RECT 551.675 369.185 551.955 369.465 ;
        RECT 552.385 369.185 552.665 369.465 ;
        RECT 553.095 369.185 553.375 369.465 ;
        RECT 553.805 369.185 554.085 369.465 ;
        RECT 554.515 369.185 554.795 369.465 ;
        RECT 555.225 369.185 555.505 369.465 ;
        RECT 555.935 369.185 556.215 369.465 ;
        RECT 556.645 369.185 556.925 369.465 ;
        RECT 557.355 369.185 557.635 369.465 ;
        RECT 558.065 369.185 558.345 369.465 ;
        RECT 558.775 369.185 559.055 369.465 ;
        RECT 559.485 369.185 559.765 369.465 ;
        RECT 560.195 369.185 560.475 369.465 ;
        RECT 550.965 368.475 551.245 368.755 ;
        RECT 551.675 368.475 551.955 368.755 ;
        RECT 552.385 368.475 552.665 368.755 ;
        RECT 553.095 368.475 553.375 368.755 ;
        RECT 553.805 368.475 554.085 368.755 ;
        RECT 554.515 368.475 554.795 368.755 ;
        RECT 555.225 368.475 555.505 368.755 ;
        RECT 555.935 368.475 556.215 368.755 ;
        RECT 556.645 368.475 556.925 368.755 ;
        RECT 557.355 368.475 557.635 368.755 ;
        RECT 558.065 368.475 558.345 368.755 ;
        RECT 558.775 368.475 559.055 368.755 ;
        RECT 559.485 368.475 559.765 368.755 ;
        RECT 560.195 368.475 560.475 368.755 ;
        RECT 550.965 367.765 551.245 368.045 ;
        RECT 551.675 367.765 551.955 368.045 ;
        RECT 552.385 367.765 552.665 368.045 ;
        RECT 553.095 367.765 553.375 368.045 ;
        RECT 553.805 367.765 554.085 368.045 ;
        RECT 554.515 367.765 554.795 368.045 ;
        RECT 555.225 367.765 555.505 368.045 ;
        RECT 555.935 367.765 556.215 368.045 ;
        RECT 556.645 367.765 556.925 368.045 ;
        RECT 557.355 367.765 557.635 368.045 ;
        RECT 558.065 367.765 558.345 368.045 ;
        RECT 558.775 367.765 559.055 368.045 ;
        RECT 559.485 367.765 559.765 368.045 ;
        RECT 560.195 367.765 560.475 368.045 ;
        RECT 550.965 367.055 551.245 367.335 ;
        RECT 551.675 367.055 551.955 367.335 ;
        RECT 552.385 367.055 552.665 367.335 ;
        RECT 553.095 367.055 553.375 367.335 ;
        RECT 553.805 367.055 554.085 367.335 ;
        RECT 554.515 367.055 554.795 367.335 ;
        RECT 555.225 367.055 555.505 367.335 ;
        RECT 555.935 367.055 556.215 367.335 ;
        RECT 556.645 367.055 556.925 367.335 ;
        RECT 557.355 367.055 557.635 367.335 ;
        RECT 558.065 367.055 558.345 367.335 ;
        RECT 558.775 367.055 559.055 367.335 ;
        RECT 559.485 367.055 559.765 367.335 ;
        RECT 560.195 367.055 560.475 367.335 ;
        RECT 550.965 366.345 551.245 366.625 ;
        RECT 551.675 366.345 551.955 366.625 ;
        RECT 552.385 366.345 552.665 366.625 ;
        RECT 553.095 366.345 553.375 366.625 ;
        RECT 553.805 366.345 554.085 366.625 ;
        RECT 554.515 366.345 554.795 366.625 ;
        RECT 555.225 366.345 555.505 366.625 ;
        RECT 555.935 366.345 556.215 366.625 ;
        RECT 556.645 366.345 556.925 366.625 ;
        RECT 557.355 366.345 557.635 366.625 ;
        RECT 558.065 366.345 558.345 366.625 ;
        RECT 558.775 366.345 559.055 366.625 ;
        RECT 559.485 366.345 559.765 366.625 ;
        RECT 560.195 366.345 560.475 366.625 ;
        RECT 550.965 365.635 551.245 365.915 ;
        RECT 551.675 365.635 551.955 365.915 ;
        RECT 552.385 365.635 552.665 365.915 ;
        RECT 553.095 365.635 553.375 365.915 ;
        RECT 553.805 365.635 554.085 365.915 ;
        RECT 554.515 365.635 554.795 365.915 ;
        RECT 555.225 365.635 555.505 365.915 ;
        RECT 555.935 365.635 556.215 365.915 ;
        RECT 556.645 365.635 556.925 365.915 ;
        RECT 557.355 365.635 557.635 365.915 ;
        RECT 558.065 365.635 558.345 365.915 ;
        RECT 558.775 365.635 559.055 365.915 ;
        RECT 559.485 365.635 559.765 365.915 ;
        RECT 560.195 365.635 560.475 365.915 ;
        RECT 550.965 364.925 551.245 365.205 ;
        RECT 551.675 364.925 551.955 365.205 ;
        RECT 552.385 364.925 552.665 365.205 ;
        RECT 553.095 364.925 553.375 365.205 ;
        RECT 553.805 364.925 554.085 365.205 ;
        RECT 554.515 364.925 554.795 365.205 ;
        RECT 555.225 364.925 555.505 365.205 ;
        RECT 555.935 364.925 556.215 365.205 ;
        RECT 556.645 364.925 556.925 365.205 ;
        RECT 557.355 364.925 557.635 365.205 ;
        RECT 558.065 364.925 558.345 365.205 ;
        RECT 558.775 364.925 559.055 365.205 ;
        RECT 559.485 364.925 559.765 365.205 ;
        RECT 560.195 364.925 560.475 365.205 ;
        RECT 550.965 364.215 551.245 364.495 ;
        RECT 551.675 364.215 551.955 364.495 ;
        RECT 552.385 364.215 552.665 364.495 ;
        RECT 553.095 364.215 553.375 364.495 ;
        RECT 553.805 364.215 554.085 364.495 ;
        RECT 554.515 364.215 554.795 364.495 ;
        RECT 555.225 364.215 555.505 364.495 ;
        RECT 555.935 364.215 556.215 364.495 ;
        RECT 556.645 364.215 556.925 364.495 ;
        RECT 557.355 364.215 557.635 364.495 ;
        RECT 558.065 364.215 558.345 364.495 ;
        RECT 558.775 364.215 559.055 364.495 ;
        RECT 559.485 364.215 559.765 364.495 ;
        RECT 560.195 364.215 560.475 364.495 ;
        RECT 550.965 363.505 551.245 363.785 ;
        RECT 551.675 363.505 551.955 363.785 ;
        RECT 552.385 363.505 552.665 363.785 ;
        RECT 553.095 363.505 553.375 363.785 ;
        RECT 553.805 363.505 554.085 363.785 ;
        RECT 554.515 363.505 554.795 363.785 ;
        RECT 555.225 363.505 555.505 363.785 ;
        RECT 555.935 363.505 556.215 363.785 ;
        RECT 556.645 363.505 556.925 363.785 ;
        RECT 557.355 363.505 557.635 363.785 ;
        RECT 558.065 363.505 558.345 363.785 ;
        RECT 558.775 363.505 559.055 363.785 ;
        RECT 559.485 363.505 559.765 363.785 ;
        RECT 560.195 363.505 560.475 363.785 ;
        RECT 550.965 362.795 551.245 363.075 ;
        RECT 551.675 362.795 551.955 363.075 ;
        RECT 552.385 362.795 552.665 363.075 ;
        RECT 553.095 362.795 553.375 363.075 ;
        RECT 553.805 362.795 554.085 363.075 ;
        RECT 554.515 362.795 554.795 363.075 ;
        RECT 555.225 362.795 555.505 363.075 ;
        RECT 555.935 362.795 556.215 363.075 ;
        RECT 556.645 362.795 556.925 363.075 ;
        RECT 557.355 362.795 557.635 363.075 ;
        RECT 558.065 362.795 558.345 363.075 ;
        RECT 558.775 362.795 559.055 363.075 ;
        RECT 559.485 362.795 559.765 363.075 ;
        RECT 560.195 362.795 560.475 363.075 ;
        RECT 550.965 362.085 551.245 362.365 ;
        RECT 551.675 362.085 551.955 362.365 ;
        RECT 552.385 362.085 552.665 362.365 ;
        RECT 553.095 362.085 553.375 362.365 ;
        RECT 553.805 362.085 554.085 362.365 ;
        RECT 554.515 362.085 554.795 362.365 ;
        RECT 555.225 362.085 555.505 362.365 ;
        RECT 555.935 362.085 556.215 362.365 ;
        RECT 556.645 362.085 556.925 362.365 ;
        RECT 557.355 362.085 557.635 362.365 ;
        RECT 558.065 362.085 558.345 362.365 ;
        RECT 558.775 362.085 559.055 362.365 ;
        RECT 559.485 362.085 559.765 362.365 ;
        RECT 560.195 362.085 560.475 362.365 ;
        RECT 550.965 361.375 551.245 361.655 ;
        RECT 551.675 361.375 551.955 361.655 ;
        RECT 552.385 361.375 552.665 361.655 ;
        RECT 553.095 361.375 553.375 361.655 ;
        RECT 553.805 361.375 554.085 361.655 ;
        RECT 554.515 361.375 554.795 361.655 ;
        RECT 555.225 361.375 555.505 361.655 ;
        RECT 555.935 361.375 556.215 361.655 ;
        RECT 556.645 361.375 556.925 361.655 ;
        RECT 557.355 361.375 557.635 361.655 ;
        RECT 558.065 361.375 558.345 361.655 ;
        RECT 558.775 361.375 559.055 361.655 ;
        RECT 559.485 361.375 559.765 361.655 ;
        RECT 560.195 361.375 560.475 361.655 ;
        RECT 550.965 360.665 551.245 360.945 ;
        RECT 551.675 360.665 551.955 360.945 ;
        RECT 552.385 360.665 552.665 360.945 ;
        RECT 553.095 360.665 553.375 360.945 ;
        RECT 553.805 360.665 554.085 360.945 ;
        RECT 554.515 360.665 554.795 360.945 ;
        RECT 555.225 360.665 555.505 360.945 ;
        RECT 555.935 360.665 556.215 360.945 ;
        RECT 556.645 360.665 556.925 360.945 ;
        RECT 557.355 360.665 557.635 360.945 ;
        RECT 558.065 360.665 558.345 360.945 ;
        RECT 558.775 360.665 559.055 360.945 ;
        RECT 559.485 360.665 559.765 360.945 ;
        RECT 560.195 360.665 560.475 360.945 ;
        RECT 566.625 369.895 566.905 370.175 ;
        RECT 567.335 369.895 567.615 370.175 ;
        RECT 568.045 369.895 568.325 370.175 ;
        RECT 568.755 369.895 569.035 370.175 ;
        RECT 569.465 369.895 569.745 370.175 ;
        RECT 570.175 369.895 570.455 370.175 ;
        RECT 570.885 369.895 571.165 370.175 ;
        RECT 571.595 369.895 571.875 370.175 ;
        RECT 572.305 369.895 572.585 370.175 ;
        RECT 573.015 369.895 573.295 370.175 ;
        RECT 573.725 369.895 574.005 370.175 ;
        RECT 566.625 369.185 566.905 369.465 ;
        RECT 567.335 369.185 567.615 369.465 ;
        RECT 568.045 369.185 568.325 369.465 ;
        RECT 568.755 369.185 569.035 369.465 ;
        RECT 569.465 369.185 569.745 369.465 ;
        RECT 570.175 369.185 570.455 369.465 ;
        RECT 570.885 369.185 571.165 369.465 ;
        RECT 571.595 369.185 571.875 369.465 ;
        RECT 572.305 369.185 572.585 369.465 ;
        RECT 573.015 369.185 573.295 369.465 ;
        RECT 573.725 369.185 574.005 369.465 ;
        RECT 566.625 368.475 566.905 368.755 ;
        RECT 567.335 368.475 567.615 368.755 ;
        RECT 568.045 368.475 568.325 368.755 ;
        RECT 568.755 368.475 569.035 368.755 ;
        RECT 569.465 368.475 569.745 368.755 ;
        RECT 570.175 368.475 570.455 368.755 ;
        RECT 570.885 368.475 571.165 368.755 ;
        RECT 571.595 368.475 571.875 368.755 ;
        RECT 572.305 368.475 572.585 368.755 ;
        RECT 573.015 368.475 573.295 368.755 ;
        RECT 573.725 368.475 574.005 368.755 ;
        RECT 566.625 367.765 566.905 368.045 ;
        RECT 567.335 367.765 567.615 368.045 ;
        RECT 568.045 367.765 568.325 368.045 ;
        RECT 568.755 367.765 569.035 368.045 ;
        RECT 569.465 367.765 569.745 368.045 ;
        RECT 570.175 367.765 570.455 368.045 ;
        RECT 570.885 367.765 571.165 368.045 ;
        RECT 571.595 367.765 571.875 368.045 ;
        RECT 572.305 367.765 572.585 368.045 ;
        RECT 573.015 367.765 573.295 368.045 ;
        RECT 573.725 367.765 574.005 368.045 ;
        RECT 566.625 367.055 566.905 367.335 ;
        RECT 567.335 367.055 567.615 367.335 ;
        RECT 568.045 367.055 568.325 367.335 ;
        RECT 568.755 367.055 569.035 367.335 ;
        RECT 569.465 367.055 569.745 367.335 ;
        RECT 570.175 367.055 570.455 367.335 ;
        RECT 570.885 367.055 571.165 367.335 ;
        RECT 571.595 367.055 571.875 367.335 ;
        RECT 572.305 367.055 572.585 367.335 ;
        RECT 573.015 367.055 573.295 367.335 ;
        RECT 573.725 367.055 574.005 367.335 ;
        RECT 566.625 366.345 566.905 366.625 ;
        RECT 567.335 366.345 567.615 366.625 ;
        RECT 568.045 366.345 568.325 366.625 ;
        RECT 568.755 366.345 569.035 366.625 ;
        RECT 569.465 366.345 569.745 366.625 ;
        RECT 570.175 366.345 570.455 366.625 ;
        RECT 570.885 366.345 571.165 366.625 ;
        RECT 571.595 366.345 571.875 366.625 ;
        RECT 572.305 366.345 572.585 366.625 ;
        RECT 573.015 366.345 573.295 366.625 ;
        RECT 573.725 366.345 574.005 366.625 ;
        RECT 566.625 365.635 566.905 365.915 ;
        RECT 567.335 365.635 567.615 365.915 ;
        RECT 568.045 365.635 568.325 365.915 ;
        RECT 568.755 365.635 569.035 365.915 ;
        RECT 569.465 365.635 569.745 365.915 ;
        RECT 570.175 365.635 570.455 365.915 ;
        RECT 570.885 365.635 571.165 365.915 ;
        RECT 571.595 365.635 571.875 365.915 ;
        RECT 572.305 365.635 572.585 365.915 ;
        RECT 573.015 365.635 573.295 365.915 ;
        RECT 573.725 365.635 574.005 365.915 ;
        RECT 566.625 364.925 566.905 365.205 ;
        RECT 567.335 364.925 567.615 365.205 ;
        RECT 568.045 364.925 568.325 365.205 ;
        RECT 568.755 364.925 569.035 365.205 ;
        RECT 569.465 364.925 569.745 365.205 ;
        RECT 570.175 364.925 570.455 365.205 ;
        RECT 570.885 364.925 571.165 365.205 ;
        RECT 571.595 364.925 571.875 365.205 ;
        RECT 572.305 364.925 572.585 365.205 ;
        RECT 573.015 364.925 573.295 365.205 ;
        RECT 573.725 364.925 574.005 365.205 ;
        RECT 566.625 364.215 566.905 364.495 ;
        RECT 567.335 364.215 567.615 364.495 ;
        RECT 568.045 364.215 568.325 364.495 ;
        RECT 568.755 364.215 569.035 364.495 ;
        RECT 569.465 364.215 569.745 364.495 ;
        RECT 570.175 364.215 570.455 364.495 ;
        RECT 570.885 364.215 571.165 364.495 ;
        RECT 571.595 364.215 571.875 364.495 ;
        RECT 572.305 364.215 572.585 364.495 ;
        RECT 573.015 364.215 573.295 364.495 ;
        RECT 573.725 364.215 574.005 364.495 ;
        RECT 566.625 363.505 566.905 363.785 ;
        RECT 567.335 363.505 567.615 363.785 ;
        RECT 568.045 363.505 568.325 363.785 ;
        RECT 568.755 363.505 569.035 363.785 ;
        RECT 569.465 363.505 569.745 363.785 ;
        RECT 570.175 363.505 570.455 363.785 ;
        RECT 570.885 363.505 571.165 363.785 ;
        RECT 571.595 363.505 571.875 363.785 ;
        RECT 572.305 363.505 572.585 363.785 ;
        RECT 573.015 363.505 573.295 363.785 ;
        RECT 573.725 363.505 574.005 363.785 ;
        RECT 566.625 362.795 566.905 363.075 ;
        RECT 567.335 362.795 567.615 363.075 ;
        RECT 568.045 362.795 568.325 363.075 ;
        RECT 568.755 362.795 569.035 363.075 ;
        RECT 569.465 362.795 569.745 363.075 ;
        RECT 570.175 362.795 570.455 363.075 ;
        RECT 570.885 362.795 571.165 363.075 ;
        RECT 571.595 362.795 571.875 363.075 ;
        RECT 572.305 362.795 572.585 363.075 ;
        RECT 573.015 362.795 573.295 363.075 ;
        RECT 573.725 362.795 574.005 363.075 ;
        RECT 566.625 362.085 566.905 362.365 ;
        RECT 567.335 362.085 567.615 362.365 ;
        RECT 568.045 362.085 568.325 362.365 ;
        RECT 568.755 362.085 569.035 362.365 ;
        RECT 569.465 362.085 569.745 362.365 ;
        RECT 570.175 362.085 570.455 362.365 ;
        RECT 570.885 362.085 571.165 362.365 ;
        RECT 571.595 362.085 571.875 362.365 ;
        RECT 572.305 362.085 572.585 362.365 ;
        RECT 573.015 362.085 573.295 362.365 ;
        RECT 573.725 362.085 574.005 362.365 ;
        RECT 566.625 361.375 566.905 361.655 ;
        RECT 567.335 361.375 567.615 361.655 ;
        RECT 568.045 361.375 568.325 361.655 ;
        RECT 568.755 361.375 569.035 361.655 ;
        RECT 569.465 361.375 569.745 361.655 ;
        RECT 570.175 361.375 570.455 361.655 ;
        RECT 570.885 361.375 571.165 361.655 ;
        RECT 571.595 361.375 571.875 361.655 ;
        RECT 572.305 361.375 572.585 361.655 ;
        RECT 573.015 361.375 573.295 361.655 ;
        RECT 573.725 361.375 574.005 361.655 ;
        RECT 566.625 360.665 566.905 360.945 ;
        RECT 567.335 360.665 567.615 360.945 ;
        RECT 568.045 360.665 568.325 360.945 ;
        RECT 568.755 360.665 569.035 360.945 ;
        RECT 569.465 360.665 569.745 360.945 ;
        RECT 570.175 360.665 570.455 360.945 ;
        RECT 570.885 360.665 571.165 360.945 ;
        RECT 571.595 360.665 571.875 360.945 ;
        RECT 572.305 360.665 572.585 360.945 ;
        RECT 573.015 360.665 573.295 360.945 ;
        RECT 573.725 360.665 574.005 360.945 ;
        RECT 576.345 369.895 576.625 370.175 ;
        RECT 577.055 369.895 577.335 370.175 ;
        RECT 577.765 369.895 578.045 370.175 ;
        RECT 578.475 369.895 578.755 370.175 ;
        RECT 579.185 369.895 579.465 370.175 ;
        RECT 579.895 369.895 580.175 370.175 ;
        RECT 580.605 369.895 580.885 370.175 ;
        RECT 581.315 369.895 581.595 370.175 ;
        RECT 582.025 369.895 582.305 370.175 ;
        RECT 582.735 369.895 583.015 370.175 ;
        RECT 583.445 369.895 583.725 370.175 ;
        RECT 584.155 369.895 584.435 370.175 ;
        RECT 584.865 369.895 585.145 370.175 ;
        RECT 585.575 369.895 585.855 370.175 ;
        RECT 576.345 369.185 576.625 369.465 ;
        RECT 577.055 369.185 577.335 369.465 ;
        RECT 577.765 369.185 578.045 369.465 ;
        RECT 578.475 369.185 578.755 369.465 ;
        RECT 579.185 369.185 579.465 369.465 ;
        RECT 579.895 369.185 580.175 369.465 ;
        RECT 580.605 369.185 580.885 369.465 ;
        RECT 581.315 369.185 581.595 369.465 ;
        RECT 582.025 369.185 582.305 369.465 ;
        RECT 582.735 369.185 583.015 369.465 ;
        RECT 583.445 369.185 583.725 369.465 ;
        RECT 584.155 369.185 584.435 369.465 ;
        RECT 584.865 369.185 585.145 369.465 ;
        RECT 585.575 369.185 585.855 369.465 ;
        RECT 576.345 368.475 576.625 368.755 ;
        RECT 577.055 368.475 577.335 368.755 ;
        RECT 577.765 368.475 578.045 368.755 ;
        RECT 578.475 368.475 578.755 368.755 ;
        RECT 579.185 368.475 579.465 368.755 ;
        RECT 579.895 368.475 580.175 368.755 ;
        RECT 580.605 368.475 580.885 368.755 ;
        RECT 581.315 368.475 581.595 368.755 ;
        RECT 582.025 368.475 582.305 368.755 ;
        RECT 582.735 368.475 583.015 368.755 ;
        RECT 583.445 368.475 583.725 368.755 ;
        RECT 584.155 368.475 584.435 368.755 ;
        RECT 584.865 368.475 585.145 368.755 ;
        RECT 585.575 368.475 585.855 368.755 ;
        RECT 576.345 367.765 576.625 368.045 ;
        RECT 577.055 367.765 577.335 368.045 ;
        RECT 577.765 367.765 578.045 368.045 ;
        RECT 578.475 367.765 578.755 368.045 ;
        RECT 579.185 367.765 579.465 368.045 ;
        RECT 579.895 367.765 580.175 368.045 ;
        RECT 580.605 367.765 580.885 368.045 ;
        RECT 581.315 367.765 581.595 368.045 ;
        RECT 582.025 367.765 582.305 368.045 ;
        RECT 582.735 367.765 583.015 368.045 ;
        RECT 583.445 367.765 583.725 368.045 ;
        RECT 584.155 367.765 584.435 368.045 ;
        RECT 584.865 367.765 585.145 368.045 ;
        RECT 585.575 367.765 585.855 368.045 ;
        RECT 576.345 367.055 576.625 367.335 ;
        RECT 577.055 367.055 577.335 367.335 ;
        RECT 577.765 367.055 578.045 367.335 ;
        RECT 578.475 367.055 578.755 367.335 ;
        RECT 579.185 367.055 579.465 367.335 ;
        RECT 579.895 367.055 580.175 367.335 ;
        RECT 580.605 367.055 580.885 367.335 ;
        RECT 581.315 367.055 581.595 367.335 ;
        RECT 582.025 367.055 582.305 367.335 ;
        RECT 582.735 367.055 583.015 367.335 ;
        RECT 583.445 367.055 583.725 367.335 ;
        RECT 584.155 367.055 584.435 367.335 ;
        RECT 584.865 367.055 585.145 367.335 ;
        RECT 585.575 367.055 585.855 367.335 ;
        RECT 576.345 366.345 576.625 366.625 ;
        RECT 577.055 366.345 577.335 366.625 ;
        RECT 577.765 366.345 578.045 366.625 ;
        RECT 578.475 366.345 578.755 366.625 ;
        RECT 579.185 366.345 579.465 366.625 ;
        RECT 579.895 366.345 580.175 366.625 ;
        RECT 580.605 366.345 580.885 366.625 ;
        RECT 581.315 366.345 581.595 366.625 ;
        RECT 582.025 366.345 582.305 366.625 ;
        RECT 582.735 366.345 583.015 366.625 ;
        RECT 583.445 366.345 583.725 366.625 ;
        RECT 584.155 366.345 584.435 366.625 ;
        RECT 584.865 366.345 585.145 366.625 ;
        RECT 585.575 366.345 585.855 366.625 ;
        RECT 576.345 365.635 576.625 365.915 ;
        RECT 577.055 365.635 577.335 365.915 ;
        RECT 577.765 365.635 578.045 365.915 ;
        RECT 578.475 365.635 578.755 365.915 ;
        RECT 579.185 365.635 579.465 365.915 ;
        RECT 579.895 365.635 580.175 365.915 ;
        RECT 580.605 365.635 580.885 365.915 ;
        RECT 581.315 365.635 581.595 365.915 ;
        RECT 582.025 365.635 582.305 365.915 ;
        RECT 582.735 365.635 583.015 365.915 ;
        RECT 583.445 365.635 583.725 365.915 ;
        RECT 584.155 365.635 584.435 365.915 ;
        RECT 584.865 365.635 585.145 365.915 ;
        RECT 585.575 365.635 585.855 365.915 ;
        RECT 576.345 364.925 576.625 365.205 ;
        RECT 577.055 364.925 577.335 365.205 ;
        RECT 577.765 364.925 578.045 365.205 ;
        RECT 578.475 364.925 578.755 365.205 ;
        RECT 579.185 364.925 579.465 365.205 ;
        RECT 579.895 364.925 580.175 365.205 ;
        RECT 580.605 364.925 580.885 365.205 ;
        RECT 581.315 364.925 581.595 365.205 ;
        RECT 582.025 364.925 582.305 365.205 ;
        RECT 582.735 364.925 583.015 365.205 ;
        RECT 583.445 364.925 583.725 365.205 ;
        RECT 584.155 364.925 584.435 365.205 ;
        RECT 584.865 364.925 585.145 365.205 ;
        RECT 585.575 364.925 585.855 365.205 ;
        RECT 576.345 364.215 576.625 364.495 ;
        RECT 577.055 364.215 577.335 364.495 ;
        RECT 577.765 364.215 578.045 364.495 ;
        RECT 578.475 364.215 578.755 364.495 ;
        RECT 579.185 364.215 579.465 364.495 ;
        RECT 579.895 364.215 580.175 364.495 ;
        RECT 580.605 364.215 580.885 364.495 ;
        RECT 581.315 364.215 581.595 364.495 ;
        RECT 582.025 364.215 582.305 364.495 ;
        RECT 582.735 364.215 583.015 364.495 ;
        RECT 583.445 364.215 583.725 364.495 ;
        RECT 584.155 364.215 584.435 364.495 ;
        RECT 584.865 364.215 585.145 364.495 ;
        RECT 585.575 364.215 585.855 364.495 ;
        RECT 576.345 363.505 576.625 363.785 ;
        RECT 577.055 363.505 577.335 363.785 ;
        RECT 577.765 363.505 578.045 363.785 ;
        RECT 578.475 363.505 578.755 363.785 ;
        RECT 579.185 363.505 579.465 363.785 ;
        RECT 579.895 363.505 580.175 363.785 ;
        RECT 580.605 363.505 580.885 363.785 ;
        RECT 581.315 363.505 581.595 363.785 ;
        RECT 582.025 363.505 582.305 363.785 ;
        RECT 582.735 363.505 583.015 363.785 ;
        RECT 583.445 363.505 583.725 363.785 ;
        RECT 584.155 363.505 584.435 363.785 ;
        RECT 584.865 363.505 585.145 363.785 ;
        RECT 585.575 363.505 585.855 363.785 ;
        RECT 576.345 362.795 576.625 363.075 ;
        RECT 577.055 362.795 577.335 363.075 ;
        RECT 577.765 362.795 578.045 363.075 ;
        RECT 578.475 362.795 578.755 363.075 ;
        RECT 579.185 362.795 579.465 363.075 ;
        RECT 579.895 362.795 580.175 363.075 ;
        RECT 580.605 362.795 580.885 363.075 ;
        RECT 581.315 362.795 581.595 363.075 ;
        RECT 582.025 362.795 582.305 363.075 ;
        RECT 582.735 362.795 583.015 363.075 ;
        RECT 583.445 362.795 583.725 363.075 ;
        RECT 584.155 362.795 584.435 363.075 ;
        RECT 584.865 362.795 585.145 363.075 ;
        RECT 585.575 362.795 585.855 363.075 ;
        RECT 576.345 362.085 576.625 362.365 ;
        RECT 577.055 362.085 577.335 362.365 ;
        RECT 577.765 362.085 578.045 362.365 ;
        RECT 578.475 362.085 578.755 362.365 ;
        RECT 579.185 362.085 579.465 362.365 ;
        RECT 579.895 362.085 580.175 362.365 ;
        RECT 580.605 362.085 580.885 362.365 ;
        RECT 581.315 362.085 581.595 362.365 ;
        RECT 582.025 362.085 582.305 362.365 ;
        RECT 582.735 362.085 583.015 362.365 ;
        RECT 583.445 362.085 583.725 362.365 ;
        RECT 584.155 362.085 584.435 362.365 ;
        RECT 584.865 362.085 585.145 362.365 ;
        RECT 585.575 362.085 585.855 362.365 ;
        RECT 576.345 361.375 576.625 361.655 ;
        RECT 577.055 361.375 577.335 361.655 ;
        RECT 577.765 361.375 578.045 361.655 ;
        RECT 578.475 361.375 578.755 361.655 ;
        RECT 579.185 361.375 579.465 361.655 ;
        RECT 579.895 361.375 580.175 361.655 ;
        RECT 580.605 361.375 580.885 361.655 ;
        RECT 581.315 361.375 581.595 361.655 ;
        RECT 582.025 361.375 582.305 361.655 ;
        RECT 582.735 361.375 583.015 361.655 ;
        RECT 583.445 361.375 583.725 361.655 ;
        RECT 584.155 361.375 584.435 361.655 ;
        RECT 584.865 361.375 585.145 361.655 ;
        RECT 585.575 361.375 585.855 361.655 ;
        RECT 576.345 360.665 576.625 360.945 ;
        RECT 577.055 360.665 577.335 360.945 ;
        RECT 577.765 360.665 578.045 360.945 ;
        RECT 578.475 360.665 578.755 360.945 ;
        RECT 579.185 360.665 579.465 360.945 ;
        RECT 579.895 360.665 580.175 360.945 ;
        RECT 580.605 360.665 580.885 360.945 ;
        RECT 581.315 360.665 581.595 360.945 ;
        RECT 582.025 360.665 582.305 360.945 ;
        RECT 582.735 360.665 583.015 360.945 ;
        RECT 583.445 360.665 583.725 360.945 ;
        RECT 584.155 360.665 584.435 360.945 ;
        RECT 584.865 360.665 585.145 360.945 ;
        RECT 585.575 360.665 585.855 360.945 ;
        RECT 589.495 369.895 589.775 370.175 ;
        RECT 590.205 369.895 590.485 370.175 ;
        RECT 590.915 369.895 591.195 370.175 ;
        RECT 591.625 369.895 591.905 370.175 ;
        RECT 592.335 369.895 592.615 370.175 ;
        RECT 593.045 369.895 593.325 370.175 ;
        RECT 593.755 369.895 594.035 370.175 ;
        RECT 594.465 369.895 594.745 370.175 ;
        RECT 595.175 369.895 595.455 370.175 ;
        RECT 595.885 369.895 596.165 370.175 ;
        RECT 596.595 369.895 596.875 370.175 ;
        RECT 597.305 369.895 597.585 370.175 ;
        RECT 598.015 369.895 598.295 370.175 ;
        RECT 589.495 369.185 589.775 369.465 ;
        RECT 590.205 369.185 590.485 369.465 ;
        RECT 590.915 369.185 591.195 369.465 ;
        RECT 591.625 369.185 591.905 369.465 ;
        RECT 592.335 369.185 592.615 369.465 ;
        RECT 593.045 369.185 593.325 369.465 ;
        RECT 593.755 369.185 594.035 369.465 ;
        RECT 594.465 369.185 594.745 369.465 ;
        RECT 595.175 369.185 595.455 369.465 ;
        RECT 595.885 369.185 596.165 369.465 ;
        RECT 596.595 369.185 596.875 369.465 ;
        RECT 597.305 369.185 597.585 369.465 ;
        RECT 598.015 369.185 598.295 369.465 ;
        RECT 589.495 368.475 589.775 368.755 ;
        RECT 590.205 368.475 590.485 368.755 ;
        RECT 590.915 368.475 591.195 368.755 ;
        RECT 591.625 368.475 591.905 368.755 ;
        RECT 592.335 368.475 592.615 368.755 ;
        RECT 593.045 368.475 593.325 368.755 ;
        RECT 593.755 368.475 594.035 368.755 ;
        RECT 594.465 368.475 594.745 368.755 ;
        RECT 595.175 368.475 595.455 368.755 ;
        RECT 595.885 368.475 596.165 368.755 ;
        RECT 596.595 368.475 596.875 368.755 ;
        RECT 597.305 368.475 597.585 368.755 ;
        RECT 598.015 368.475 598.295 368.755 ;
        RECT 589.495 367.765 589.775 368.045 ;
        RECT 590.205 367.765 590.485 368.045 ;
        RECT 590.915 367.765 591.195 368.045 ;
        RECT 591.625 367.765 591.905 368.045 ;
        RECT 592.335 367.765 592.615 368.045 ;
        RECT 593.045 367.765 593.325 368.045 ;
        RECT 593.755 367.765 594.035 368.045 ;
        RECT 594.465 367.765 594.745 368.045 ;
        RECT 595.175 367.765 595.455 368.045 ;
        RECT 595.885 367.765 596.165 368.045 ;
        RECT 596.595 367.765 596.875 368.045 ;
        RECT 597.305 367.765 597.585 368.045 ;
        RECT 598.015 367.765 598.295 368.045 ;
        RECT 589.495 367.055 589.775 367.335 ;
        RECT 590.205 367.055 590.485 367.335 ;
        RECT 590.915 367.055 591.195 367.335 ;
        RECT 591.625 367.055 591.905 367.335 ;
        RECT 592.335 367.055 592.615 367.335 ;
        RECT 593.045 367.055 593.325 367.335 ;
        RECT 593.755 367.055 594.035 367.335 ;
        RECT 594.465 367.055 594.745 367.335 ;
        RECT 595.175 367.055 595.455 367.335 ;
        RECT 595.885 367.055 596.165 367.335 ;
        RECT 596.595 367.055 596.875 367.335 ;
        RECT 597.305 367.055 597.585 367.335 ;
        RECT 598.015 367.055 598.295 367.335 ;
        RECT 589.495 366.345 589.775 366.625 ;
        RECT 590.205 366.345 590.485 366.625 ;
        RECT 590.915 366.345 591.195 366.625 ;
        RECT 591.625 366.345 591.905 366.625 ;
        RECT 592.335 366.345 592.615 366.625 ;
        RECT 593.045 366.345 593.325 366.625 ;
        RECT 593.755 366.345 594.035 366.625 ;
        RECT 594.465 366.345 594.745 366.625 ;
        RECT 595.175 366.345 595.455 366.625 ;
        RECT 595.885 366.345 596.165 366.625 ;
        RECT 596.595 366.345 596.875 366.625 ;
        RECT 597.305 366.345 597.585 366.625 ;
        RECT 598.015 366.345 598.295 366.625 ;
        RECT 589.495 365.635 589.775 365.915 ;
        RECT 590.205 365.635 590.485 365.915 ;
        RECT 590.915 365.635 591.195 365.915 ;
        RECT 591.625 365.635 591.905 365.915 ;
        RECT 592.335 365.635 592.615 365.915 ;
        RECT 593.045 365.635 593.325 365.915 ;
        RECT 593.755 365.635 594.035 365.915 ;
        RECT 594.465 365.635 594.745 365.915 ;
        RECT 595.175 365.635 595.455 365.915 ;
        RECT 595.885 365.635 596.165 365.915 ;
        RECT 596.595 365.635 596.875 365.915 ;
        RECT 597.305 365.635 597.585 365.915 ;
        RECT 598.015 365.635 598.295 365.915 ;
        RECT 589.495 364.925 589.775 365.205 ;
        RECT 590.205 364.925 590.485 365.205 ;
        RECT 590.915 364.925 591.195 365.205 ;
        RECT 591.625 364.925 591.905 365.205 ;
        RECT 592.335 364.925 592.615 365.205 ;
        RECT 593.045 364.925 593.325 365.205 ;
        RECT 593.755 364.925 594.035 365.205 ;
        RECT 594.465 364.925 594.745 365.205 ;
        RECT 595.175 364.925 595.455 365.205 ;
        RECT 595.885 364.925 596.165 365.205 ;
        RECT 596.595 364.925 596.875 365.205 ;
        RECT 597.305 364.925 597.585 365.205 ;
        RECT 598.015 364.925 598.295 365.205 ;
        RECT 589.495 364.215 589.775 364.495 ;
        RECT 590.205 364.215 590.485 364.495 ;
        RECT 590.915 364.215 591.195 364.495 ;
        RECT 591.625 364.215 591.905 364.495 ;
        RECT 592.335 364.215 592.615 364.495 ;
        RECT 593.045 364.215 593.325 364.495 ;
        RECT 593.755 364.215 594.035 364.495 ;
        RECT 594.465 364.215 594.745 364.495 ;
        RECT 595.175 364.215 595.455 364.495 ;
        RECT 595.885 364.215 596.165 364.495 ;
        RECT 596.595 364.215 596.875 364.495 ;
        RECT 597.305 364.215 597.585 364.495 ;
        RECT 598.015 364.215 598.295 364.495 ;
        RECT 589.495 363.505 589.775 363.785 ;
        RECT 590.205 363.505 590.485 363.785 ;
        RECT 590.915 363.505 591.195 363.785 ;
        RECT 591.625 363.505 591.905 363.785 ;
        RECT 592.335 363.505 592.615 363.785 ;
        RECT 593.045 363.505 593.325 363.785 ;
        RECT 593.755 363.505 594.035 363.785 ;
        RECT 594.465 363.505 594.745 363.785 ;
        RECT 595.175 363.505 595.455 363.785 ;
        RECT 595.885 363.505 596.165 363.785 ;
        RECT 596.595 363.505 596.875 363.785 ;
        RECT 597.305 363.505 597.585 363.785 ;
        RECT 598.015 363.505 598.295 363.785 ;
        RECT 589.495 362.795 589.775 363.075 ;
        RECT 590.205 362.795 590.485 363.075 ;
        RECT 590.915 362.795 591.195 363.075 ;
        RECT 591.625 362.795 591.905 363.075 ;
        RECT 592.335 362.795 592.615 363.075 ;
        RECT 593.045 362.795 593.325 363.075 ;
        RECT 593.755 362.795 594.035 363.075 ;
        RECT 594.465 362.795 594.745 363.075 ;
        RECT 595.175 362.795 595.455 363.075 ;
        RECT 595.885 362.795 596.165 363.075 ;
        RECT 596.595 362.795 596.875 363.075 ;
        RECT 597.305 362.795 597.585 363.075 ;
        RECT 598.015 362.795 598.295 363.075 ;
        RECT 589.495 362.085 589.775 362.365 ;
        RECT 590.205 362.085 590.485 362.365 ;
        RECT 590.915 362.085 591.195 362.365 ;
        RECT 591.625 362.085 591.905 362.365 ;
        RECT 592.335 362.085 592.615 362.365 ;
        RECT 593.045 362.085 593.325 362.365 ;
        RECT 593.755 362.085 594.035 362.365 ;
        RECT 594.465 362.085 594.745 362.365 ;
        RECT 595.175 362.085 595.455 362.365 ;
        RECT 595.885 362.085 596.165 362.365 ;
        RECT 596.595 362.085 596.875 362.365 ;
        RECT 597.305 362.085 597.585 362.365 ;
        RECT 598.015 362.085 598.295 362.365 ;
        RECT 589.495 361.375 589.775 361.655 ;
        RECT 590.205 361.375 590.485 361.655 ;
        RECT 590.915 361.375 591.195 361.655 ;
        RECT 591.625 361.375 591.905 361.655 ;
        RECT 592.335 361.375 592.615 361.655 ;
        RECT 593.045 361.375 593.325 361.655 ;
        RECT 593.755 361.375 594.035 361.655 ;
        RECT 594.465 361.375 594.745 361.655 ;
        RECT 595.175 361.375 595.455 361.655 ;
        RECT 595.885 361.375 596.165 361.655 ;
        RECT 596.595 361.375 596.875 361.655 ;
        RECT 597.305 361.375 597.585 361.655 ;
        RECT 598.015 361.375 598.295 361.655 ;
        RECT 589.495 360.665 589.775 360.945 ;
        RECT 590.205 360.665 590.485 360.945 ;
        RECT 590.915 360.665 591.195 360.945 ;
        RECT 591.625 360.665 591.905 360.945 ;
        RECT 592.335 360.665 592.615 360.945 ;
        RECT 593.045 360.665 593.325 360.945 ;
        RECT 593.755 360.665 594.035 360.945 ;
        RECT 594.465 360.665 594.745 360.945 ;
        RECT 595.175 360.665 595.455 360.945 ;
        RECT 595.885 360.665 596.165 360.945 ;
        RECT 596.595 360.665 596.875 360.945 ;
        RECT 597.305 360.665 597.585 360.945 ;
        RECT 598.015 360.665 598.295 360.945 ;
        RECT 1351.715 369.895 1351.995 370.175 ;
        RECT 1352.425 369.895 1352.705 370.175 ;
        RECT 1353.135 369.895 1353.415 370.175 ;
        RECT 1353.845 369.895 1354.125 370.175 ;
        RECT 1354.555 369.895 1354.835 370.175 ;
        RECT 1355.265 369.895 1355.545 370.175 ;
        RECT 1355.975 369.895 1356.255 370.175 ;
        RECT 1356.685 369.895 1356.965 370.175 ;
        RECT 1357.395 369.895 1357.675 370.175 ;
        RECT 1358.105 369.895 1358.385 370.175 ;
        RECT 1358.815 369.895 1359.095 370.175 ;
        RECT 1359.525 369.895 1359.805 370.175 ;
        RECT 1360.235 369.895 1360.515 370.175 ;
        RECT 1351.715 369.185 1351.995 369.465 ;
        RECT 1352.425 369.185 1352.705 369.465 ;
        RECT 1353.135 369.185 1353.415 369.465 ;
        RECT 1353.845 369.185 1354.125 369.465 ;
        RECT 1354.555 369.185 1354.835 369.465 ;
        RECT 1355.265 369.185 1355.545 369.465 ;
        RECT 1355.975 369.185 1356.255 369.465 ;
        RECT 1356.685 369.185 1356.965 369.465 ;
        RECT 1357.395 369.185 1357.675 369.465 ;
        RECT 1358.105 369.185 1358.385 369.465 ;
        RECT 1358.815 369.185 1359.095 369.465 ;
        RECT 1359.525 369.185 1359.805 369.465 ;
        RECT 1360.235 369.185 1360.515 369.465 ;
        RECT 1351.715 368.475 1351.995 368.755 ;
        RECT 1352.425 368.475 1352.705 368.755 ;
        RECT 1353.135 368.475 1353.415 368.755 ;
        RECT 1353.845 368.475 1354.125 368.755 ;
        RECT 1354.555 368.475 1354.835 368.755 ;
        RECT 1355.265 368.475 1355.545 368.755 ;
        RECT 1355.975 368.475 1356.255 368.755 ;
        RECT 1356.685 368.475 1356.965 368.755 ;
        RECT 1357.395 368.475 1357.675 368.755 ;
        RECT 1358.105 368.475 1358.385 368.755 ;
        RECT 1358.815 368.475 1359.095 368.755 ;
        RECT 1359.525 368.475 1359.805 368.755 ;
        RECT 1360.235 368.475 1360.515 368.755 ;
        RECT 1351.715 367.765 1351.995 368.045 ;
        RECT 1352.425 367.765 1352.705 368.045 ;
        RECT 1353.135 367.765 1353.415 368.045 ;
        RECT 1353.845 367.765 1354.125 368.045 ;
        RECT 1354.555 367.765 1354.835 368.045 ;
        RECT 1355.265 367.765 1355.545 368.045 ;
        RECT 1355.975 367.765 1356.255 368.045 ;
        RECT 1356.685 367.765 1356.965 368.045 ;
        RECT 1357.395 367.765 1357.675 368.045 ;
        RECT 1358.105 367.765 1358.385 368.045 ;
        RECT 1358.815 367.765 1359.095 368.045 ;
        RECT 1359.525 367.765 1359.805 368.045 ;
        RECT 1360.235 367.765 1360.515 368.045 ;
        RECT 1351.715 367.055 1351.995 367.335 ;
        RECT 1352.425 367.055 1352.705 367.335 ;
        RECT 1353.135 367.055 1353.415 367.335 ;
        RECT 1353.845 367.055 1354.125 367.335 ;
        RECT 1354.555 367.055 1354.835 367.335 ;
        RECT 1355.265 367.055 1355.545 367.335 ;
        RECT 1355.975 367.055 1356.255 367.335 ;
        RECT 1356.685 367.055 1356.965 367.335 ;
        RECT 1357.395 367.055 1357.675 367.335 ;
        RECT 1358.105 367.055 1358.385 367.335 ;
        RECT 1358.815 367.055 1359.095 367.335 ;
        RECT 1359.525 367.055 1359.805 367.335 ;
        RECT 1360.235 367.055 1360.515 367.335 ;
        RECT 1351.715 366.345 1351.995 366.625 ;
        RECT 1352.425 366.345 1352.705 366.625 ;
        RECT 1353.135 366.345 1353.415 366.625 ;
        RECT 1353.845 366.345 1354.125 366.625 ;
        RECT 1354.555 366.345 1354.835 366.625 ;
        RECT 1355.265 366.345 1355.545 366.625 ;
        RECT 1355.975 366.345 1356.255 366.625 ;
        RECT 1356.685 366.345 1356.965 366.625 ;
        RECT 1357.395 366.345 1357.675 366.625 ;
        RECT 1358.105 366.345 1358.385 366.625 ;
        RECT 1358.815 366.345 1359.095 366.625 ;
        RECT 1359.525 366.345 1359.805 366.625 ;
        RECT 1360.235 366.345 1360.515 366.625 ;
        RECT 1351.715 365.635 1351.995 365.915 ;
        RECT 1352.425 365.635 1352.705 365.915 ;
        RECT 1353.135 365.635 1353.415 365.915 ;
        RECT 1353.845 365.635 1354.125 365.915 ;
        RECT 1354.555 365.635 1354.835 365.915 ;
        RECT 1355.265 365.635 1355.545 365.915 ;
        RECT 1355.975 365.635 1356.255 365.915 ;
        RECT 1356.685 365.635 1356.965 365.915 ;
        RECT 1357.395 365.635 1357.675 365.915 ;
        RECT 1358.105 365.635 1358.385 365.915 ;
        RECT 1358.815 365.635 1359.095 365.915 ;
        RECT 1359.525 365.635 1359.805 365.915 ;
        RECT 1360.235 365.635 1360.515 365.915 ;
        RECT 1351.715 364.925 1351.995 365.205 ;
        RECT 1352.425 364.925 1352.705 365.205 ;
        RECT 1353.135 364.925 1353.415 365.205 ;
        RECT 1353.845 364.925 1354.125 365.205 ;
        RECT 1354.555 364.925 1354.835 365.205 ;
        RECT 1355.265 364.925 1355.545 365.205 ;
        RECT 1355.975 364.925 1356.255 365.205 ;
        RECT 1356.685 364.925 1356.965 365.205 ;
        RECT 1357.395 364.925 1357.675 365.205 ;
        RECT 1358.105 364.925 1358.385 365.205 ;
        RECT 1358.815 364.925 1359.095 365.205 ;
        RECT 1359.525 364.925 1359.805 365.205 ;
        RECT 1360.235 364.925 1360.515 365.205 ;
        RECT 1351.715 364.215 1351.995 364.495 ;
        RECT 1352.425 364.215 1352.705 364.495 ;
        RECT 1353.135 364.215 1353.415 364.495 ;
        RECT 1353.845 364.215 1354.125 364.495 ;
        RECT 1354.555 364.215 1354.835 364.495 ;
        RECT 1355.265 364.215 1355.545 364.495 ;
        RECT 1355.975 364.215 1356.255 364.495 ;
        RECT 1356.685 364.215 1356.965 364.495 ;
        RECT 1357.395 364.215 1357.675 364.495 ;
        RECT 1358.105 364.215 1358.385 364.495 ;
        RECT 1358.815 364.215 1359.095 364.495 ;
        RECT 1359.525 364.215 1359.805 364.495 ;
        RECT 1360.235 364.215 1360.515 364.495 ;
        RECT 1351.715 363.505 1351.995 363.785 ;
        RECT 1352.425 363.505 1352.705 363.785 ;
        RECT 1353.135 363.505 1353.415 363.785 ;
        RECT 1353.845 363.505 1354.125 363.785 ;
        RECT 1354.555 363.505 1354.835 363.785 ;
        RECT 1355.265 363.505 1355.545 363.785 ;
        RECT 1355.975 363.505 1356.255 363.785 ;
        RECT 1356.685 363.505 1356.965 363.785 ;
        RECT 1357.395 363.505 1357.675 363.785 ;
        RECT 1358.105 363.505 1358.385 363.785 ;
        RECT 1358.815 363.505 1359.095 363.785 ;
        RECT 1359.525 363.505 1359.805 363.785 ;
        RECT 1360.235 363.505 1360.515 363.785 ;
        RECT 1351.715 362.795 1351.995 363.075 ;
        RECT 1352.425 362.795 1352.705 363.075 ;
        RECT 1353.135 362.795 1353.415 363.075 ;
        RECT 1353.845 362.795 1354.125 363.075 ;
        RECT 1354.555 362.795 1354.835 363.075 ;
        RECT 1355.265 362.795 1355.545 363.075 ;
        RECT 1355.975 362.795 1356.255 363.075 ;
        RECT 1356.685 362.795 1356.965 363.075 ;
        RECT 1357.395 362.795 1357.675 363.075 ;
        RECT 1358.105 362.795 1358.385 363.075 ;
        RECT 1358.815 362.795 1359.095 363.075 ;
        RECT 1359.525 362.795 1359.805 363.075 ;
        RECT 1360.235 362.795 1360.515 363.075 ;
        RECT 1351.715 362.085 1351.995 362.365 ;
        RECT 1352.425 362.085 1352.705 362.365 ;
        RECT 1353.135 362.085 1353.415 362.365 ;
        RECT 1353.845 362.085 1354.125 362.365 ;
        RECT 1354.555 362.085 1354.835 362.365 ;
        RECT 1355.265 362.085 1355.545 362.365 ;
        RECT 1355.975 362.085 1356.255 362.365 ;
        RECT 1356.685 362.085 1356.965 362.365 ;
        RECT 1357.395 362.085 1357.675 362.365 ;
        RECT 1358.105 362.085 1358.385 362.365 ;
        RECT 1358.815 362.085 1359.095 362.365 ;
        RECT 1359.525 362.085 1359.805 362.365 ;
        RECT 1360.235 362.085 1360.515 362.365 ;
        RECT 1351.715 361.375 1351.995 361.655 ;
        RECT 1352.425 361.375 1352.705 361.655 ;
        RECT 1353.135 361.375 1353.415 361.655 ;
        RECT 1353.845 361.375 1354.125 361.655 ;
        RECT 1354.555 361.375 1354.835 361.655 ;
        RECT 1355.265 361.375 1355.545 361.655 ;
        RECT 1355.975 361.375 1356.255 361.655 ;
        RECT 1356.685 361.375 1356.965 361.655 ;
        RECT 1357.395 361.375 1357.675 361.655 ;
        RECT 1358.105 361.375 1358.385 361.655 ;
        RECT 1358.815 361.375 1359.095 361.655 ;
        RECT 1359.525 361.375 1359.805 361.655 ;
        RECT 1360.235 361.375 1360.515 361.655 ;
        RECT 1351.715 360.665 1351.995 360.945 ;
        RECT 1352.425 360.665 1352.705 360.945 ;
        RECT 1353.135 360.665 1353.415 360.945 ;
        RECT 1353.845 360.665 1354.125 360.945 ;
        RECT 1354.555 360.665 1354.835 360.945 ;
        RECT 1355.265 360.665 1355.545 360.945 ;
        RECT 1355.975 360.665 1356.255 360.945 ;
        RECT 1356.685 360.665 1356.965 360.945 ;
        RECT 1357.395 360.665 1357.675 360.945 ;
        RECT 1358.105 360.665 1358.385 360.945 ;
        RECT 1358.815 360.665 1359.095 360.945 ;
        RECT 1359.525 360.665 1359.805 360.945 ;
        RECT 1360.235 360.665 1360.515 360.945 ;
        RECT 1364.115 369.895 1364.395 370.175 ;
        RECT 1364.825 369.895 1365.105 370.175 ;
        RECT 1365.535 369.895 1365.815 370.175 ;
        RECT 1366.245 369.895 1366.525 370.175 ;
        RECT 1366.955 369.895 1367.235 370.175 ;
        RECT 1367.665 369.895 1367.945 370.175 ;
        RECT 1368.375 369.895 1368.655 370.175 ;
        RECT 1369.085 369.895 1369.365 370.175 ;
        RECT 1369.795 369.895 1370.075 370.175 ;
        RECT 1370.505 369.895 1370.785 370.175 ;
        RECT 1371.215 369.895 1371.495 370.175 ;
        RECT 1371.925 369.895 1372.205 370.175 ;
        RECT 1372.635 369.895 1372.915 370.175 ;
        RECT 1373.345 369.895 1373.625 370.175 ;
        RECT 1364.115 369.185 1364.395 369.465 ;
        RECT 1364.825 369.185 1365.105 369.465 ;
        RECT 1365.535 369.185 1365.815 369.465 ;
        RECT 1366.245 369.185 1366.525 369.465 ;
        RECT 1366.955 369.185 1367.235 369.465 ;
        RECT 1367.665 369.185 1367.945 369.465 ;
        RECT 1368.375 369.185 1368.655 369.465 ;
        RECT 1369.085 369.185 1369.365 369.465 ;
        RECT 1369.795 369.185 1370.075 369.465 ;
        RECT 1370.505 369.185 1370.785 369.465 ;
        RECT 1371.215 369.185 1371.495 369.465 ;
        RECT 1371.925 369.185 1372.205 369.465 ;
        RECT 1372.635 369.185 1372.915 369.465 ;
        RECT 1373.345 369.185 1373.625 369.465 ;
        RECT 1364.115 368.475 1364.395 368.755 ;
        RECT 1364.825 368.475 1365.105 368.755 ;
        RECT 1365.535 368.475 1365.815 368.755 ;
        RECT 1366.245 368.475 1366.525 368.755 ;
        RECT 1366.955 368.475 1367.235 368.755 ;
        RECT 1367.665 368.475 1367.945 368.755 ;
        RECT 1368.375 368.475 1368.655 368.755 ;
        RECT 1369.085 368.475 1369.365 368.755 ;
        RECT 1369.795 368.475 1370.075 368.755 ;
        RECT 1370.505 368.475 1370.785 368.755 ;
        RECT 1371.215 368.475 1371.495 368.755 ;
        RECT 1371.925 368.475 1372.205 368.755 ;
        RECT 1372.635 368.475 1372.915 368.755 ;
        RECT 1373.345 368.475 1373.625 368.755 ;
        RECT 1364.115 367.765 1364.395 368.045 ;
        RECT 1364.825 367.765 1365.105 368.045 ;
        RECT 1365.535 367.765 1365.815 368.045 ;
        RECT 1366.245 367.765 1366.525 368.045 ;
        RECT 1366.955 367.765 1367.235 368.045 ;
        RECT 1367.665 367.765 1367.945 368.045 ;
        RECT 1368.375 367.765 1368.655 368.045 ;
        RECT 1369.085 367.765 1369.365 368.045 ;
        RECT 1369.795 367.765 1370.075 368.045 ;
        RECT 1370.505 367.765 1370.785 368.045 ;
        RECT 1371.215 367.765 1371.495 368.045 ;
        RECT 1371.925 367.765 1372.205 368.045 ;
        RECT 1372.635 367.765 1372.915 368.045 ;
        RECT 1373.345 367.765 1373.625 368.045 ;
        RECT 1364.115 367.055 1364.395 367.335 ;
        RECT 1364.825 367.055 1365.105 367.335 ;
        RECT 1365.535 367.055 1365.815 367.335 ;
        RECT 1366.245 367.055 1366.525 367.335 ;
        RECT 1366.955 367.055 1367.235 367.335 ;
        RECT 1367.665 367.055 1367.945 367.335 ;
        RECT 1368.375 367.055 1368.655 367.335 ;
        RECT 1369.085 367.055 1369.365 367.335 ;
        RECT 1369.795 367.055 1370.075 367.335 ;
        RECT 1370.505 367.055 1370.785 367.335 ;
        RECT 1371.215 367.055 1371.495 367.335 ;
        RECT 1371.925 367.055 1372.205 367.335 ;
        RECT 1372.635 367.055 1372.915 367.335 ;
        RECT 1373.345 367.055 1373.625 367.335 ;
        RECT 1364.115 366.345 1364.395 366.625 ;
        RECT 1364.825 366.345 1365.105 366.625 ;
        RECT 1365.535 366.345 1365.815 366.625 ;
        RECT 1366.245 366.345 1366.525 366.625 ;
        RECT 1366.955 366.345 1367.235 366.625 ;
        RECT 1367.665 366.345 1367.945 366.625 ;
        RECT 1368.375 366.345 1368.655 366.625 ;
        RECT 1369.085 366.345 1369.365 366.625 ;
        RECT 1369.795 366.345 1370.075 366.625 ;
        RECT 1370.505 366.345 1370.785 366.625 ;
        RECT 1371.215 366.345 1371.495 366.625 ;
        RECT 1371.925 366.345 1372.205 366.625 ;
        RECT 1372.635 366.345 1372.915 366.625 ;
        RECT 1373.345 366.345 1373.625 366.625 ;
        RECT 1364.115 365.635 1364.395 365.915 ;
        RECT 1364.825 365.635 1365.105 365.915 ;
        RECT 1365.535 365.635 1365.815 365.915 ;
        RECT 1366.245 365.635 1366.525 365.915 ;
        RECT 1366.955 365.635 1367.235 365.915 ;
        RECT 1367.665 365.635 1367.945 365.915 ;
        RECT 1368.375 365.635 1368.655 365.915 ;
        RECT 1369.085 365.635 1369.365 365.915 ;
        RECT 1369.795 365.635 1370.075 365.915 ;
        RECT 1370.505 365.635 1370.785 365.915 ;
        RECT 1371.215 365.635 1371.495 365.915 ;
        RECT 1371.925 365.635 1372.205 365.915 ;
        RECT 1372.635 365.635 1372.915 365.915 ;
        RECT 1373.345 365.635 1373.625 365.915 ;
        RECT 1364.115 364.925 1364.395 365.205 ;
        RECT 1364.825 364.925 1365.105 365.205 ;
        RECT 1365.535 364.925 1365.815 365.205 ;
        RECT 1366.245 364.925 1366.525 365.205 ;
        RECT 1366.955 364.925 1367.235 365.205 ;
        RECT 1367.665 364.925 1367.945 365.205 ;
        RECT 1368.375 364.925 1368.655 365.205 ;
        RECT 1369.085 364.925 1369.365 365.205 ;
        RECT 1369.795 364.925 1370.075 365.205 ;
        RECT 1370.505 364.925 1370.785 365.205 ;
        RECT 1371.215 364.925 1371.495 365.205 ;
        RECT 1371.925 364.925 1372.205 365.205 ;
        RECT 1372.635 364.925 1372.915 365.205 ;
        RECT 1373.345 364.925 1373.625 365.205 ;
        RECT 1364.115 364.215 1364.395 364.495 ;
        RECT 1364.825 364.215 1365.105 364.495 ;
        RECT 1365.535 364.215 1365.815 364.495 ;
        RECT 1366.245 364.215 1366.525 364.495 ;
        RECT 1366.955 364.215 1367.235 364.495 ;
        RECT 1367.665 364.215 1367.945 364.495 ;
        RECT 1368.375 364.215 1368.655 364.495 ;
        RECT 1369.085 364.215 1369.365 364.495 ;
        RECT 1369.795 364.215 1370.075 364.495 ;
        RECT 1370.505 364.215 1370.785 364.495 ;
        RECT 1371.215 364.215 1371.495 364.495 ;
        RECT 1371.925 364.215 1372.205 364.495 ;
        RECT 1372.635 364.215 1372.915 364.495 ;
        RECT 1373.345 364.215 1373.625 364.495 ;
        RECT 1364.115 363.505 1364.395 363.785 ;
        RECT 1364.825 363.505 1365.105 363.785 ;
        RECT 1365.535 363.505 1365.815 363.785 ;
        RECT 1366.245 363.505 1366.525 363.785 ;
        RECT 1366.955 363.505 1367.235 363.785 ;
        RECT 1367.665 363.505 1367.945 363.785 ;
        RECT 1368.375 363.505 1368.655 363.785 ;
        RECT 1369.085 363.505 1369.365 363.785 ;
        RECT 1369.795 363.505 1370.075 363.785 ;
        RECT 1370.505 363.505 1370.785 363.785 ;
        RECT 1371.215 363.505 1371.495 363.785 ;
        RECT 1371.925 363.505 1372.205 363.785 ;
        RECT 1372.635 363.505 1372.915 363.785 ;
        RECT 1373.345 363.505 1373.625 363.785 ;
        RECT 1364.115 362.795 1364.395 363.075 ;
        RECT 1364.825 362.795 1365.105 363.075 ;
        RECT 1365.535 362.795 1365.815 363.075 ;
        RECT 1366.245 362.795 1366.525 363.075 ;
        RECT 1366.955 362.795 1367.235 363.075 ;
        RECT 1367.665 362.795 1367.945 363.075 ;
        RECT 1368.375 362.795 1368.655 363.075 ;
        RECT 1369.085 362.795 1369.365 363.075 ;
        RECT 1369.795 362.795 1370.075 363.075 ;
        RECT 1370.505 362.795 1370.785 363.075 ;
        RECT 1371.215 362.795 1371.495 363.075 ;
        RECT 1371.925 362.795 1372.205 363.075 ;
        RECT 1372.635 362.795 1372.915 363.075 ;
        RECT 1373.345 362.795 1373.625 363.075 ;
        RECT 1364.115 362.085 1364.395 362.365 ;
        RECT 1364.825 362.085 1365.105 362.365 ;
        RECT 1365.535 362.085 1365.815 362.365 ;
        RECT 1366.245 362.085 1366.525 362.365 ;
        RECT 1366.955 362.085 1367.235 362.365 ;
        RECT 1367.665 362.085 1367.945 362.365 ;
        RECT 1368.375 362.085 1368.655 362.365 ;
        RECT 1369.085 362.085 1369.365 362.365 ;
        RECT 1369.795 362.085 1370.075 362.365 ;
        RECT 1370.505 362.085 1370.785 362.365 ;
        RECT 1371.215 362.085 1371.495 362.365 ;
        RECT 1371.925 362.085 1372.205 362.365 ;
        RECT 1372.635 362.085 1372.915 362.365 ;
        RECT 1373.345 362.085 1373.625 362.365 ;
        RECT 1364.115 361.375 1364.395 361.655 ;
        RECT 1364.825 361.375 1365.105 361.655 ;
        RECT 1365.535 361.375 1365.815 361.655 ;
        RECT 1366.245 361.375 1366.525 361.655 ;
        RECT 1366.955 361.375 1367.235 361.655 ;
        RECT 1367.665 361.375 1367.945 361.655 ;
        RECT 1368.375 361.375 1368.655 361.655 ;
        RECT 1369.085 361.375 1369.365 361.655 ;
        RECT 1369.795 361.375 1370.075 361.655 ;
        RECT 1370.505 361.375 1370.785 361.655 ;
        RECT 1371.215 361.375 1371.495 361.655 ;
        RECT 1371.925 361.375 1372.205 361.655 ;
        RECT 1372.635 361.375 1372.915 361.655 ;
        RECT 1373.345 361.375 1373.625 361.655 ;
        RECT 1364.115 360.665 1364.395 360.945 ;
        RECT 1364.825 360.665 1365.105 360.945 ;
        RECT 1365.535 360.665 1365.815 360.945 ;
        RECT 1366.245 360.665 1366.525 360.945 ;
        RECT 1366.955 360.665 1367.235 360.945 ;
        RECT 1367.665 360.665 1367.945 360.945 ;
        RECT 1368.375 360.665 1368.655 360.945 ;
        RECT 1369.085 360.665 1369.365 360.945 ;
        RECT 1369.795 360.665 1370.075 360.945 ;
        RECT 1370.505 360.665 1370.785 360.945 ;
        RECT 1371.215 360.665 1371.495 360.945 ;
        RECT 1371.925 360.665 1372.205 360.945 ;
        RECT 1372.635 360.665 1372.915 360.945 ;
        RECT 1373.345 360.665 1373.625 360.945 ;
        RECT 1375.965 369.895 1376.245 370.175 ;
        RECT 1376.675 369.895 1376.955 370.175 ;
        RECT 1377.385 369.895 1377.665 370.175 ;
        RECT 1378.095 369.895 1378.375 370.175 ;
        RECT 1378.805 369.895 1379.085 370.175 ;
        RECT 1379.515 369.895 1379.795 370.175 ;
        RECT 1380.225 369.895 1380.505 370.175 ;
        RECT 1380.935 369.895 1381.215 370.175 ;
        RECT 1381.645 369.895 1381.925 370.175 ;
        RECT 1382.355 369.895 1382.635 370.175 ;
        RECT 1383.065 369.895 1383.345 370.175 ;
        RECT 1383.775 369.895 1384.055 370.175 ;
        RECT 1384.485 369.895 1384.765 370.175 ;
        RECT 1385.195 369.895 1385.475 370.175 ;
        RECT 1375.965 369.185 1376.245 369.465 ;
        RECT 1376.675 369.185 1376.955 369.465 ;
        RECT 1377.385 369.185 1377.665 369.465 ;
        RECT 1378.095 369.185 1378.375 369.465 ;
        RECT 1378.805 369.185 1379.085 369.465 ;
        RECT 1379.515 369.185 1379.795 369.465 ;
        RECT 1380.225 369.185 1380.505 369.465 ;
        RECT 1380.935 369.185 1381.215 369.465 ;
        RECT 1381.645 369.185 1381.925 369.465 ;
        RECT 1382.355 369.185 1382.635 369.465 ;
        RECT 1383.065 369.185 1383.345 369.465 ;
        RECT 1383.775 369.185 1384.055 369.465 ;
        RECT 1384.485 369.185 1384.765 369.465 ;
        RECT 1385.195 369.185 1385.475 369.465 ;
        RECT 1375.965 368.475 1376.245 368.755 ;
        RECT 1376.675 368.475 1376.955 368.755 ;
        RECT 1377.385 368.475 1377.665 368.755 ;
        RECT 1378.095 368.475 1378.375 368.755 ;
        RECT 1378.805 368.475 1379.085 368.755 ;
        RECT 1379.515 368.475 1379.795 368.755 ;
        RECT 1380.225 368.475 1380.505 368.755 ;
        RECT 1380.935 368.475 1381.215 368.755 ;
        RECT 1381.645 368.475 1381.925 368.755 ;
        RECT 1382.355 368.475 1382.635 368.755 ;
        RECT 1383.065 368.475 1383.345 368.755 ;
        RECT 1383.775 368.475 1384.055 368.755 ;
        RECT 1384.485 368.475 1384.765 368.755 ;
        RECT 1385.195 368.475 1385.475 368.755 ;
        RECT 1375.965 367.765 1376.245 368.045 ;
        RECT 1376.675 367.765 1376.955 368.045 ;
        RECT 1377.385 367.765 1377.665 368.045 ;
        RECT 1378.095 367.765 1378.375 368.045 ;
        RECT 1378.805 367.765 1379.085 368.045 ;
        RECT 1379.515 367.765 1379.795 368.045 ;
        RECT 1380.225 367.765 1380.505 368.045 ;
        RECT 1380.935 367.765 1381.215 368.045 ;
        RECT 1381.645 367.765 1381.925 368.045 ;
        RECT 1382.355 367.765 1382.635 368.045 ;
        RECT 1383.065 367.765 1383.345 368.045 ;
        RECT 1383.775 367.765 1384.055 368.045 ;
        RECT 1384.485 367.765 1384.765 368.045 ;
        RECT 1385.195 367.765 1385.475 368.045 ;
        RECT 1375.965 367.055 1376.245 367.335 ;
        RECT 1376.675 367.055 1376.955 367.335 ;
        RECT 1377.385 367.055 1377.665 367.335 ;
        RECT 1378.095 367.055 1378.375 367.335 ;
        RECT 1378.805 367.055 1379.085 367.335 ;
        RECT 1379.515 367.055 1379.795 367.335 ;
        RECT 1380.225 367.055 1380.505 367.335 ;
        RECT 1380.935 367.055 1381.215 367.335 ;
        RECT 1381.645 367.055 1381.925 367.335 ;
        RECT 1382.355 367.055 1382.635 367.335 ;
        RECT 1383.065 367.055 1383.345 367.335 ;
        RECT 1383.775 367.055 1384.055 367.335 ;
        RECT 1384.485 367.055 1384.765 367.335 ;
        RECT 1385.195 367.055 1385.475 367.335 ;
        RECT 1375.965 366.345 1376.245 366.625 ;
        RECT 1376.675 366.345 1376.955 366.625 ;
        RECT 1377.385 366.345 1377.665 366.625 ;
        RECT 1378.095 366.345 1378.375 366.625 ;
        RECT 1378.805 366.345 1379.085 366.625 ;
        RECT 1379.515 366.345 1379.795 366.625 ;
        RECT 1380.225 366.345 1380.505 366.625 ;
        RECT 1380.935 366.345 1381.215 366.625 ;
        RECT 1381.645 366.345 1381.925 366.625 ;
        RECT 1382.355 366.345 1382.635 366.625 ;
        RECT 1383.065 366.345 1383.345 366.625 ;
        RECT 1383.775 366.345 1384.055 366.625 ;
        RECT 1384.485 366.345 1384.765 366.625 ;
        RECT 1385.195 366.345 1385.475 366.625 ;
        RECT 1375.965 365.635 1376.245 365.915 ;
        RECT 1376.675 365.635 1376.955 365.915 ;
        RECT 1377.385 365.635 1377.665 365.915 ;
        RECT 1378.095 365.635 1378.375 365.915 ;
        RECT 1378.805 365.635 1379.085 365.915 ;
        RECT 1379.515 365.635 1379.795 365.915 ;
        RECT 1380.225 365.635 1380.505 365.915 ;
        RECT 1380.935 365.635 1381.215 365.915 ;
        RECT 1381.645 365.635 1381.925 365.915 ;
        RECT 1382.355 365.635 1382.635 365.915 ;
        RECT 1383.065 365.635 1383.345 365.915 ;
        RECT 1383.775 365.635 1384.055 365.915 ;
        RECT 1384.485 365.635 1384.765 365.915 ;
        RECT 1385.195 365.635 1385.475 365.915 ;
        RECT 1375.965 364.925 1376.245 365.205 ;
        RECT 1376.675 364.925 1376.955 365.205 ;
        RECT 1377.385 364.925 1377.665 365.205 ;
        RECT 1378.095 364.925 1378.375 365.205 ;
        RECT 1378.805 364.925 1379.085 365.205 ;
        RECT 1379.515 364.925 1379.795 365.205 ;
        RECT 1380.225 364.925 1380.505 365.205 ;
        RECT 1380.935 364.925 1381.215 365.205 ;
        RECT 1381.645 364.925 1381.925 365.205 ;
        RECT 1382.355 364.925 1382.635 365.205 ;
        RECT 1383.065 364.925 1383.345 365.205 ;
        RECT 1383.775 364.925 1384.055 365.205 ;
        RECT 1384.485 364.925 1384.765 365.205 ;
        RECT 1385.195 364.925 1385.475 365.205 ;
        RECT 1375.965 364.215 1376.245 364.495 ;
        RECT 1376.675 364.215 1376.955 364.495 ;
        RECT 1377.385 364.215 1377.665 364.495 ;
        RECT 1378.095 364.215 1378.375 364.495 ;
        RECT 1378.805 364.215 1379.085 364.495 ;
        RECT 1379.515 364.215 1379.795 364.495 ;
        RECT 1380.225 364.215 1380.505 364.495 ;
        RECT 1380.935 364.215 1381.215 364.495 ;
        RECT 1381.645 364.215 1381.925 364.495 ;
        RECT 1382.355 364.215 1382.635 364.495 ;
        RECT 1383.065 364.215 1383.345 364.495 ;
        RECT 1383.775 364.215 1384.055 364.495 ;
        RECT 1384.485 364.215 1384.765 364.495 ;
        RECT 1385.195 364.215 1385.475 364.495 ;
        RECT 1375.965 363.505 1376.245 363.785 ;
        RECT 1376.675 363.505 1376.955 363.785 ;
        RECT 1377.385 363.505 1377.665 363.785 ;
        RECT 1378.095 363.505 1378.375 363.785 ;
        RECT 1378.805 363.505 1379.085 363.785 ;
        RECT 1379.515 363.505 1379.795 363.785 ;
        RECT 1380.225 363.505 1380.505 363.785 ;
        RECT 1380.935 363.505 1381.215 363.785 ;
        RECT 1381.645 363.505 1381.925 363.785 ;
        RECT 1382.355 363.505 1382.635 363.785 ;
        RECT 1383.065 363.505 1383.345 363.785 ;
        RECT 1383.775 363.505 1384.055 363.785 ;
        RECT 1384.485 363.505 1384.765 363.785 ;
        RECT 1385.195 363.505 1385.475 363.785 ;
        RECT 1375.965 362.795 1376.245 363.075 ;
        RECT 1376.675 362.795 1376.955 363.075 ;
        RECT 1377.385 362.795 1377.665 363.075 ;
        RECT 1378.095 362.795 1378.375 363.075 ;
        RECT 1378.805 362.795 1379.085 363.075 ;
        RECT 1379.515 362.795 1379.795 363.075 ;
        RECT 1380.225 362.795 1380.505 363.075 ;
        RECT 1380.935 362.795 1381.215 363.075 ;
        RECT 1381.645 362.795 1381.925 363.075 ;
        RECT 1382.355 362.795 1382.635 363.075 ;
        RECT 1383.065 362.795 1383.345 363.075 ;
        RECT 1383.775 362.795 1384.055 363.075 ;
        RECT 1384.485 362.795 1384.765 363.075 ;
        RECT 1385.195 362.795 1385.475 363.075 ;
        RECT 1375.965 362.085 1376.245 362.365 ;
        RECT 1376.675 362.085 1376.955 362.365 ;
        RECT 1377.385 362.085 1377.665 362.365 ;
        RECT 1378.095 362.085 1378.375 362.365 ;
        RECT 1378.805 362.085 1379.085 362.365 ;
        RECT 1379.515 362.085 1379.795 362.365 ;
        RECT 1380.225 362.085 1380.505 362.365 ;
        RECT 1380.935 362.085 1381.215 362.365 ;
        RECT 1381.645 362.085 1381.925 362.365 ;
        RECT 1382.355 362.085 1382.635 362.365 ;
        RECT 1383.065 362.085 1383.345 362.365 ;
        RECT 1383.775 362.085 1384.055 362.365 ;
        RECT 1384.485 362.085 1384.765 362.365 ;
        RECT 1385.195 362.085 1385.475 362.365 ;
        RECT 1375.965 361.375 1376.245 361.655 ;
        RECT 1376.675 361.375 1376.955 361.655 ;
        RECT 1377.385 361.375 1377.665 361.655 ;
        RECT 1378.095 361.375 1378.375 361.655 ;
        RECT 1378.805 361.375 1379.085 361.655 ;
        RECT 1379.515 361.375 1379.795 361.655 ;
        RECT 1380.225 361.375 1380.505 361.655 ;
        RECT 1380.935 361.375 1381.215 361.655 ;
        RECT 1381.645 361.375 1381.925 361.655 ;
        RECT 1382.355 361.375 1382.635 361.655 ;
        RECT 1383.065 361.375 1383.345 361.655 ;
        RECT 1383.775 361.375 1384.055 361.655 ;
        RECT 1384.485 361.375 1384.765 361.655 ;
        RECT 1385.195 361.375 1385.475 361.655 ;
        RECT 1375.965 360.665 1376.245 360.945 ;
        RECT 1376.675 360.665 1376.955 360.945 ;
        RECT 1377.385 360.665 1377.665 360.945 ;
        RECT 1378.095 360.665 1378.375 360.945 ;
        RECT 1378.805 360.665 1379.085 360.945 ;
        RECT 1379.515 360.665 1379.795 360.945 ;
        RECT 1380.225 360.665 1380.505 360.945 ;
        RECT 1380.935 360.665 1381.215 360.945 ;
        RECT 1381.645 360.665 1381.925 360.945 ;
        RECT 1382.355 360.665 1382.635 360.945 ;
        RECT 1383.065 360.665 1383.345 360.945 ;
        RECT 1383.775 360.665 1384.055 360.945 ;
        RECT 1384.485 360.665 1384.765 360.945 ;
        RECT 1385.195 360.665 1385.475 360.945 ;
        RECT 1389.495 369.895 1389.775 370.175 ;
        RECT 1390.205 369.895 1390.485 370.175 ;
        RECT 1390.915 369.895 1391.195 370.175 ;
        RECT 1391.625 369.895 1391.905 370.175 ;
        RECT 1392.335 369.895 1392.615 370.175 ;
        RECT 1393.045 369.895 1393.325 370.175 ;
        RECT 1393.755 369.895 1394.035 370.175 ;
        RECT 1394.465 369.895 1394.745 370.175 ;
        RECT 1395.175 369.895 1395.455 370.175 ;
        RECT 1395.885 369.895 1396.165 370.175 ;
        RECT 1396.595 369.895 1396.875 370.175 ;
        RECT 1397.305 369.895 1397.585 370.175 ;
        RECT 1398.015 369.895 1398.295 370.175 ;
        RECT 1398.725 369.895 1399.005 370.175 ;
        RECT 1389.495 369.185 1389.775 369.465 ;
        RECT 1390.205 369.185 1390.485 369.465 ;
        RECT 1390.915 369.185 1391.195 369.465 ;
        RECT 1391.625 369.185 1391.905 369.465 ;
        RECT 1392.335 369.185 1392.615 369.465 ;
        RECT 1393.045 369.185 1393.325 369.465 ;
        RECT 1393.755 369.185 1394.035 369.465 ;
        RECT 1394.465 369.185 1394.745 369.465 ;
        RECT 1395.175 369.185 1395.455 369.465 ;
        RECT 1395.885 369.185 1396.165 369.465 ;
        RECT 1396.595 369.185 1396.875 369.465 ;
        RECT 1397.305 369.185 1397.585 369.465 ;
        RECT 1398.015 369.185 1398.295 369.465 ;
        RECT 1398.725 369.185 1399.005 369.465 ;
        RECT 1389.495 368.475 1389.775 368.755 ;
        RECT 1390.205 368.475 1390.485 368.755 ;
        RECT 1390.915 368.475 1391.195 368.755 ;
        RECT 1391.625 368.475 1391.905 368.755 ;
        RECT 1392.335 368.475 1392.615 368.755 ;
        RECT 1393.045 368.475 1393.325 368.755 ;
        RECT 1393.755 368.475 1394.035 368.755 ;
        RECT 1394.465 368.475 1394.745 368.755 ;
        RECT 1395.175 368.475 1395.455 368.755 ;
        RECT 1395.885 368.475 1396.165 368.755 ;
        RECT 1396.595 368.475 1396.875 368.755 ;
        RECT 1397.305 368.475 1397.585 368.755 ;
        RECT 1398.015 368.475 1398.295 368.755 ;
        RECT 1398.725 368.475 1399.005 368.755 ;
        RECT 1389.495 367.765 1389.775 368.045 ;
        RECT 1390.205 367.765 1390.485 368.045 ;
        RECT 1390.915 367.765 1391.195 368.045 ;
        RECT 1391.625 367.765 1391.905 368.045 ;
        RECT 1392.335 367.765 1392.615 368.045 ;
        RECT 1393.045 367.765 1393.325 368.045 ;
        RECT 1393.755 367.765 1394.035 368.045 ;
        RECT 1394.465 367.765 1394.745 368.045 ;
        RECT 1395.175 367.765 1395.455 368.045 ;
        RECT 1395.885 367.765 1396.165 368.045 ;
        RECT 1396.595 367.765 1396.875 368.045 ;
        RECT 1397.305 367.765 1397.585 368.045 ;
        RECT 1398.015 367.765 1398.295 368.045 ;
        RECT 1398.725 367.765 1399.005 368.045 ;
        RECT 1389.495 367.055 1389.775 367.335 ;
        RECT 1390.205 367.055 1390.485 367.335 ;
        RECT 1390.915 367.055 1391.195 367.335 ;
        RECT 1391.625 367.055 1391.905 367.335 ;
        RECT 1392.335 367.055 1392.615 367.335 ;
        RECT 1393.045 367.055 1393.325 367.335 ;
        RECT 1393.755 367.055 1394.035 367.335 ;
        RECT 1394.465 367.055 1394.745 367.335 ;
        RECT 1395.175 367.055 1395.455 367.335 ;
        RECT 1395.885 367.055 1396.165 367.335 ;
        RECT 1396.595 367.055 1396.875 367.335 ;
        RECT 1397.305 367.055 1397.585 367.335 ;
        RECT 1398.015 367.055 1398.295 367.335 ;
        RECT 1398.725 367.055 1399.005 367.335 ;
        RECT 1389.495 366.345 1389.775 366.625 ;
        RECT 1390.205 366.345 1390.485 366.625 ;
        RECT 1390.915 366.345 1391.195 366.625 ;
        RECT 1391.625 366.345 1391.905 366.625 ;
        RECT 1392.335 366.345 1392.615 366.625 ;
        RECT 1393.045 366.345 1393.325 366.625 ;
        RECT 1393.755 366.345 1394.035 366.625 ;
        RECT 1394.465 366.345 1394.745 366.625 ;
        RECT 1395.175 366.345 1395.455 366.625 ;
        RECT 1395.885 366.345 1396.165 366.625 ;
        RECT 1396.595 366.345 1396.875 366.625 ;
        RECT 1397.305 366.345 1397.585 366.625 ;
        RECT 1398.015 366.345 1398.295 366.625 ;
        RECT 1398.725 366.345 1399.005 366.625 ;
        RECT 1389.495 365.635 1389.775 365.915 ;
        RECT 1390.205 365.635 1390.485 365.915 ;
        RECT 1390.915 365.635 1391.195 365.915 ;
        RECT 1391.625 365.635 1391.905 365.915 ;
        RECT 1392.335 365.635 1392.615 365.915 ;
        RECT 1393.045 365.635 1393.325 365.915 ;
        RECT 1393.755 365.635 1394.035 365.915 ;
        RECT 1394.465 365.635 1394.745 365.915 ;
        RECT 1395.175 365.635 1395.455 365.915 ;
        RECT 1395.885 365.635 1396.165 365.915 ;
        RECT 1396.595 365.635 1396.875 365.915 ;
        RECT 1397.305 365.635 1397.585 365.915 ;
        RECT 1398.015 365.635 1398.295 365.915 ;
        RECT 1398.725 365.635 1399.005 365.915 ;
        RECT 1389.495 364.925 1389.775 365.205 ;
        RECT 1390.205 364.925 1390.485 365.205 ;
        RECT 1390.915 364.925 1391.195 365.205 ;
        RECT 1391.625 364.925 1391.905 365.205 ;
        RECT 1392.335 364.925 1392.615 365.205 ;
        RECT 1393.045 364.925 1393.325 365.205 ;
        RECT 1393.755 364.925 1394.035 365.205 ;
        RECT 1394.465 364.925 1394.745 365.205 ;
        RECT 1395.175 364.925 1395.455 365.205 ;
        RECT 1395.885 364.925 1396.165 365.205 ;
        RECT 1396.595 364.925 1396.875 365.205 ;
        RECT 1397.305 364.925 1397.585 365.205 ;
        RECT 1398.015 364.925 1398.295 365.205 ;
        RECT 1398.725 364.925 1399.005 365.205 ;
        RECT 1389.495 364.215 1389.775 364.495 ;
        RECT 1390.205 364.215 1390.485 364.495 ;
        RECT 1390.915 364.215 1391.195 364.495 ;
        RECT 1391.625 364.215 1391.905 364.495 ;
        RECT 1392.335 364.215 1392.615 364.495 ;
        RECT 1393.045 364.215 1393.325 364.495 ;
        RECT 1393.755 364.215 1394.035 364.495 ;
        RECT 1394.465 364.215 1394.745 364.495 ;
        RECT 1395.175 364.215 1395.455 364.495 ;
        RECT 1395.885 364.215 1396.165 364.495 ;
        RECT 1396.595 364.215 1396.875 364.495 ;
        RECT 1397.305 364.215 1397.585 364.495 ;
        RECT 1398.015 364.215 1398.295 364.495 ;
        RECT 1398.725 364.215 1399.005 364.495 ;
        RECT 1389.495 363.505 1389.775 363.785 ;
        RECT 1390.205 363.505 1390.485 363.785 ;
        RECT 1390.915 363.505 1391.195 363.785 ;
        RECT 1391.625 363.505 1391.905 363.785 ;
        RECT 1392.335 363.505 1392.615 363.785 ;
        RECT 1393.045 363.505 1393.325 363.785 ;
        RECT 1393.755 363.505 1394.035 363.785 ;
        RECT 1394.465 363.505 1394.745 363.785 ;
        RECT 1395.175 363.505 1395.455 363.785 ;
        RECT 1395.885 363.505 1396.165 363.785 ;
        RECT 1396.595 363.505 1396.875 363.785 ;
        RECT 1397.305 363.505 1397.585 363.785 ;
        RECT 1398.015 363.505 1398.295 363.785 ;
        RECT 1398.725 363.505 1399.005 363.785 ;
        RECT 1389.495 362.795 1389.775 363.075 ;
        RECT 1390.205 362.795 1390.485 363.075 ;
        RECT 1390.915 362.795 1391.195 363.075 ;
        RECT 1391.625 362.795 1391.905 363.075 ;
        RECT 1392.335 362.795 1392.615 363.075 ;
        RECT 1393.045 362.795 1393.325 363.075 ;
        RECT 1393.755 362.795 1394.035 363.075 ;
        RECT 1394.465 362.795 1394.745 363.075 ;
        RECT 1395.175 362.795 1395.455 363.075 ;
        RECT 1395.885 362.795 1396.165 363.075 ;
        RECT 1396.595 362.795 1396.875 363.075 ;
        RECT 1397.305 362.795 1397.585 363.075 ;
        RECT 1398.015 362.795 1398.295 363.075 ;
        RECT 1398.725 362.795 1399.005 363.075 ;
        RECT 1389.495 362.085 1389.775 362.365 ;
        RECT 1390.205 362.085 1390.485 362.365 ;
        RECT 1390.915 362.085 1391.195 362.365 ;
        RECT 1391.625 362.085 1391.905 362.365 ;
        RECT 1392.335 362.085 1392.615 362.365 ;
        RECT 1393.045 362.085 1393.325 362.365 ;
        RECT 1393.755 362.085 1394.035 362.365 ;
        RECT 1394.465 362.085 1394.745 362.365 ;
        RECT 1395.175 362.085 1395.455 362.365 ;
        RECT 1395.885 362.085 1396.165 362.365 ;
        RECT 1396.595 362.085 1396.875 362.365 ;
        RECT 1397.305 362.085 1397.585 362.365 ;
        RECT 1398.015 362.085 1398.295 362.365 ;
        RECT 1398.725 362.085 1399.005 362.365 ;
        RECT 1389.495 361.375 1389.775 361.655 ;
        RECT 1390.205 361.375 1390.485 361.655 ;
        RECT 1390.915 361.375 1391.195 361.655 ;
        RECT 1391.625 361.375 1391.905 361.655 ;
        RECT 1392.335 361.375 1392.615 361.655 ;
        RECT 1393.045 361.375 1393.325 361.655 ;
        RECT 1393.755 361.375 1394.035 361.655 ;
        RECT 1394.465 361.375 1394.745 361.655 ;
        RECT 1395.175 361.375 1395.455 361.655 ;
        RECT 1395.885 361.375 1396.165 361.655 ;
        RECT 1396.595 361.375 1396.875 361.655 ;
        RECT 1397.305 361.375 1397.585 361.655 ;
        RECT 1398.015 361.375 1398.295 361.655 ;
        RECT 1398.725 361.375 1399.005 361.655 ;
        RECT 1389.495 360.665 1389.775 360.945 ;
        RECT 1390.205 360.665 1390.485 360.945 ;
        RECT 1390.915 360.665 1391.195 360.945 ;
        RECT 1391.625 360.665 1391.905 360.945 ;
        RECT 1392.335 360.665 1392.615 360.945 ;
        RECT 1393.045 360.665 1393.325 360.945 ;
        RECT 1393.755 360.665 1394.035 360.945 ;
        RECT 1394.465 360.665 1394.745 360.945 ;
        RECT 1395.175 360.665 1395.455 360.945 ;
        RECT 1395.885 360.665 1396.165 360.945 ;
        RECT 1396.595 360.665 1396.875 360.945 ;
        RECT 1397.305 360.665 1397.585 360.945 ;
        RECT 1398.015 360.665 1398.295 360.945 ;
        RECT 1398.725 360.665 1399.005 360.945 ;
        RECT 1401.345 369.895 1401.625 370.175 ;
        RECT 1402.055 369.895 1402.335 370.175 ;
        RECT 1402.765 369.895 1403.045 370.175 ;
        RECT 1403.475 369.895 1403.755 370.175 ;
        RECT 1404.185 369.895 1404.465 370.175 ;
        RECT 1404.895 369.895 1405.175 370.175 ;
        RECT 1405.605 369.895 1405.885 370.175 ;
        RECT 1406.315 369.895 1406.595 370.175 ;
        RECT 1407.025 369.895 1407.305 370.175 ;
        RECT 1407.735 369.895 1408.015 370.175 ;
        RECT 1408.445 369.895 1408.725 370.175 ;
        RECT 1409.155 369.895 1409.435 370.175 ;
        RECT 1409.865 369.895 1410.145 370.175 ;
        RECT 1410.575 369.895 1410.855 370.175 ;
        RECT 1401.345 369.185 1401.625 369.465 ;
        RECT 1402.055 369.185 1402.335 369.465 ;
        RECT 1402.765 369.185 1403.045 369.465 ;
        RECT 1403.475 369.185 1403.755 369.465 ;
        RECT 1404.185 369.185 1404.465 369.465 ;
        RECT 1404.895 369.185 1405.175 369.465 ;
        RECT 1405.605 369.185 1405.885 369.465 ;
        RECT 1406.315 369.185 1406.595 369.465 ;
        RECT 1407.025 369.185 1407.305 369.465 ;
        RECT 1407.735 369.185 1408.015 369.465 ;
        RECT 1408.445 369.185 1408.725 369.465 ;
        RECT 1409.155 369.185 1409.435 369.465 ;
        RECT 1409.865 369.185 1410.145 369.465 ;
        RECT 1410.575 369.185 1410.855 369.465 ;
        RECT 1401.345 368.475 1401.625 368.755 ;
        RECT 1402.055 368.475 1402.335 368.755 ;
        RECT 1402.765 368.475 1403.045 368.755 ;
        RECT 1403.475 368.475 1403.755 368.755 ;
        RECT 1404.185 368.475 1404.465 368.755 ;
        RECT 1404.895 368.475 1405.175 368.755 ;
        RECT 1405.605 368.475 1405.885 368.755 ;
        RECT 1406.315 368.475 1406.595 368.755 ;
        RECT 1407.025 368.475 1407.305 368.755 ;
        RECT 1407.735 368.475 1408.015 368.755 ;
        RECT 1408.445 368.475 1408.725 368.755 ;
        RECT 1409.155 368.475 1409.435 368.755 ;
        RECT 1409.865 368.475 1410.145 368.755 ;
        RECT 1410.575 368.475 1410.855 368.755 ;
        RECT 1401.345 367.765 1401.625 368.045 ;
        RECT 1402.055 367.765 1402.335 368.045 ;
        RECT 1402.765 367.765 1403.045 368.045 ;
        RECT 1403.475 367.765 1403.755 368.045 ;
        RECT 1404.185 367.765 1404.465 368.045 ;
        RECT 1404.895 367.765 1405.175 368.045 ;
        RECT 1405.605 367.765 1405.885 368.045 ;
        RECT 1406.315 367.765 1406.595 368.045 ;
        RECT 1407.025 367.765 1407.305 368.045 ;
        RECT 1407.735 367.765 1408.015 368.045 ;
        RECT 1408.445 367.765 1408.725 368.045 ;
        RECT 1409.155 367.765 1409.435 368.045 ;
        RECT 1409.865 367.765 1410.145 368.045 ;
        RECT 1410.575 367.765 1410.855 368.045 ;
        RECT 1401.345 367.055 1401.625 367.335 ;
        RECT 1402.055 367.055 1402.335 367.335 ;
        RECT 1402.765 367.055 1403.045 367.335 ;
        RECT 1403.475 367.055 1403.755 367.335 ;
        RECT 1404.185 367.055 1404.465 367.335 ;
        RECT 1404.895 367.055 1405.175 367.335 ;
        RECT 1405.605 367.055 1405.885 367.335 ;
        RECT 1406.315 367.055 1406.595 367.335 ;
        RECT 1407.025 367.055 1407.305 367.335 ;
        RECT 1407.735 367.055 1408.015 367.335 ;
        RECT 1408.445 367.055 1408.725 367.335 ;
        RECT 1409.155 367.055 1409.435 367.335 ;
        RECT 1409.865 367.055 1410.145 367.335 ;
        RECT 1410.575 367.055 1410.855 367.335 ;
        RECT 1401.345 366.345 1401.625 366.625 ;
        RECT 1402.055 366.345 1402.335 366.625 ;
        RECT 1402.765 366.345 1403.045 366.625 ;
        RECT 1403.475 366.345 1403.755 366.625 ;
        RECT 1404.185 366.345 1404.465 366.625 ;
        RECT 1404.895 366.345 1405.175 366.625 ;
        RECT 1405.605 366.345 1405.885 366.625 ;
        RECT 1406.315 366.345 1406.595 366.625 ;
        RECT 1407.025 366.345 1407.305 366.625 ;
        RECT 1407.735 366.345 1408.015 366.625 ;
        RECT 1408.445 366.345 1408.725 366.625 ;
        RECT 1409.155 366.345 1409.435 366.625 ;
        RECT 1409.865 366.345 1410.145 366.625 ;
        RECT 1410.575 366.345 1410.855 366.625 ;
        RECT 1401.345 365.635 1401.625 365.915 ;
        RECT 1402.055 365.635 1402.335 365.915 ;
        RECT 1402.765 365.635 1403.045 365.915 ;
        RECT 1403.475 365.635 1403.755 365.915 ;
        RECT 1404.185 365.635 1404.465 365.915 ;
        RECT 1404.895 365.635 1405.175 365.915 ;
        RECT 1405.605 365.635 1405.885 365.915 ;
        RECT 1406.315 365.635 1406.595 365.915 ;
        RECT 1407.025 365.635 1407.305 365.915 ;
        RECT 1407.735 365.635 1408.015 365.915 ;
        RECT 1408.445 365.635 1408.725 365.915 ;
        RECT 1409.155 365.635 1409.435 365.915 ;
        RECT 1409.865 365.635 1410.145 365.915 ;
        RECT 1410.575 365.635 1410.855 365.915 ;
        RECT 1401.345 364.925 1401.625 365.205 ;
        RECT 1402.055 364.925 1402.335 365.205 ;
        RECT 1402.765 364.925 1403.045 365.205 ;
        RECT 1403.475 364.925 1403.755 365.205 ;
        RECT 1404.185 364.925 1404.465 365.205 ;
        RECT 1404.895 364.925 1405.175 365.205 ;
        RECT 1405.605 364.925 1405.885 365.205 ;
        RECT 1406.315 364.925 1406.595 365.205 ;
        RECT 1407.025 364.925 1407.305 365.205 ;
        RECT 1407.735 364.925 1408.015 365.205 ;
        RECT 1408.445 364.925 1408.725 365.205 ;
        RECT 1409.155 364.925 1409.435 365.205 ;
        RECT 1409.865 364.925 1410.145 365.205 ;
        RECT 1410.575 364.925 1410.855 365.205 ;
        RECT 1401.345 364.215 1401.625 364.495 ;
        RECT 1402.055 364.215 1402.335 364.495 ;
        RECT 1402.765 364.215 1403.045 364.495 ;
        RECT 1403.475 364.215 1403.755 364.495 ;
        RECT 1404.185 364.215 1404.465 364.495 ;
        RECT 1404.895 364.215 1405.175 364.495 ;
        RECT 1405.605 364.215 1405.885 364.495 ;
        RECT 1406.315 364.215 1406.595 364.495 ;
        RECT 1407.025 364.215 1407.305 364.495 ;
        RECT 1407.735 364.215 1408.015 364.495 ;
        RECT 1408.445 364.215 1408.725 364.495 ;
        RECT 1409.155 364.215 1409.435 364.495 ;
        RECT 1409.865 364.215 1410.145 364.495 ;
        RECT 1410.575 364.215 1410.855 364.495 ;
        RECT 1401.345 363.505 1401.625 363.785 ;
        RECT 1402.055 363.505 1402.335 363.785 ;
        RECT 1402.765 363.505 1403.045 363.785 ;
        RECT 1403.475 363.505 1403.755 363.785 ;
        RECT 1404.185 363.505 1404.465 363.785 ;
        RECT 1404.895 363.505 1405.175 363.785 ;
        RECT 1405.605 363.505 1405.885 363.785 ;
        RECT 1406.315 363.505 1406.595 363.785 ;
        RECT 1407.025 363.505 1407.305 363.785 ;
        RECT 1407.735 363.505 1408.015 363.785 ;
        RECT 1408.445 363.505 1408.725 363.785 ;
        RECT 1409.155 363.505 1409.435 363.785 ;
        RECT 1409.865 363.505 1410.145 363.785 ;
        RECT 1410.575 363.505 1410.855 363.785 ;
        RECT 1401.345 362.795 1401.625 363.075 ;
        RECT 1402.055 362.795 1402.335 363.075 ;
        RECT 1402.765 362.795 1403.045 363.075 ;
        RECT 1403.475 362.795 1403.755 363.075 ;
        RECT 1404.185 362.795 1404.465 363.075 ;
        RECT 1404.895 362.795 1405.175 363.075 ;
        RECT 1405.605 362.795 1405.885 363.075 ;
        RECT 1406.315 362.795 1406.595 363.075 ;
        RECT 1407.025 362.795 1407.305 363.075 ;
        RECT 1407.735 362.795 1408.015 363.075 ;
        RECT 1408.445 362.795 1408.725 363.075 ;
        RECT 1409.155 362.795 1409.435 363.075 ;
        RECT 1409.865 362.795 1410.145 363.075 ;
        RECT 1410.575 362.795 1410.855 363.075 ;
        RECT 1401.345 362.085 1401.625 362.365 ;
        RECT 1402.055 362.085 1402.335 362.365 ;
        RECT 1402.765 362.085 1403.045 362.365 ;
        RECT 1403.475 362.085 1403.755 362.365 ;
        RECT 1404.185 362.085 1404.465 362.365 ;
        RECT 1404.895 362.085 1405.175 362.365 ;
        RECT 1405.605 362.085 1405.885 362.365 ;
        RECT 1406.315 362.085 1406.595 362.365 ;
        RECT 1407.025 362.085 1407.305 362.365 ;
        RECT 1407.735 362.085 1408.015 362.365 ;
        RECT 1408.445 362.085 1408.725 362.365 ;
        RECT 1409.155 362.085 1409.435 362.365 ;
        RECT 1409.865 362.085 1410.145 362.365 ;
        RECT 1410.575 362.085 1410.855 362.365 ;
        RECT 1401.345 361.375 1401.625 361.655 ;
        RECT 1402.055 361.375 1402.335 361.655 ;
        RECT 1402.765 361.375 1403.045 361.655 ;
        RECT 1403.475 361.375 1403.755 361.655 ;
        RECT 1404.185 361.375 1404.465 361.655 ;
        RECT 1404.895 361.375 1405.175 361.655 ;
        RECT 1405.605 361.375 1405.885 361.655 ;
        RECT 1406.315 361.375 1406.595 361.655 ;
        RECT 1407.025 361.375 1407.305 361.655 ;
        RECT 1407.735 361.375 1408.015 361.655 ;
        RECT 1408.445 361.375 1408.725 361.655 ;
        RECT 1409.155 361.375 1409.435 361.655 ;
        RECT 1409.865 361.375 1410.145 361.655 ;
        RECT 1410.575 361.375 1410.855 361.655 ;
        RECT 1401.345 360.665 1401.625 360.945 ;
        RECT 1402.055 360.665 1402.335 360.945 ;
        RECT 1402.765 360.665 1403.045 360.945 ;
        RECT 1403.475 360.665 1403.755 360.945 ;
        RECT 1404.185 360.665 1404.465 360.945 ;
        RECT 1404.895 360.665 1405.175 360.945 ;
        RECT 1405.605 360.665 1405.885 360.945 ;
        RECT 1406.315 360.665 1406.595 360.945 ;
        RECT 1407.025 360.665 1407.305 360.945 ;
        RECT 1407.735 360.665 1408.015 360.945 ;
        RECT 1408.445 360.665 1408.725 360.945 ;
        RECT 1409.155 360.665 1409.435 360.945 ;
        RECT 1409.865 360.665 1410.145 360.945 ;
        RECT 1410.575 360.665 1410.855 360.945 ;
        RECT 1414.495 369.895 1414.775 370.175 ;
        RECT 1415.205 369.895 1415.485 370.175 ;
        RECT 1415.915 369.895 1416.195 370.175 ;
        RECT 1416.625 369.895 1416.905 370.175 ;
        RECT 1417.335 369.895 1417.615 370.175 ;
        RECT 1418.045 369.895 1418.325 370.175 ;
        RECT 1418.755 369.895 1419.035 370.175 ;
        RECT 1419.465 369.895 1419.745 370.175 ;
        RECT 1414.495 369.185 1414.775 369.465 ;
        RECT 1415.205 369.185 1415.485 369.465 ;
        RECT 1415.915 369.185 1416.195 369.465 ;
        RECT 1416.625 369.185 1416.905 369.465 ;
        RECT 1417.335 369.185 1417.615 369.465 ;
        RECT 1418.045 369.185 1418.325 369.465 ;
        RECT 1418.755 369.185 1419.035 369.465 ;
        RECT 1419.465 369.185 1419.745 369.465 ;
        RECT 1414.495 368.475 1414.775 368.755 ;
        RECT 1415.205 368.475 1415.485 368.755 ;
        RECT 1415.915 368.475 1416.195 368.755 ;
        RECT 1416.625 368.475 1416.905 368.755 ;
        RECT 1417.335 368.475 1417.615 368.755 ;
        RECT 1418.045 368.475 1418.325 368.755 ;
        RECT 1418.755 368.475 1419.035 368.755 ;
        RECT 1419.465 368.475 1419.745 368.755 ;
        RECT 1414.495 367.765 1414.775 368.045 ;
        RECT 1415.205 367.765 1415.485 368.045 ;
        RECT 1415.915 367.765 1416.195 368.045 ;
        RECT 1416.625 367.765 1416.905 368.045 ;
        RECT 1417.335 367.765 1417.615 368.045 ;
        RECT 1418.045 367.765 1418.325 368.045 ;
        RECT 1418.755 367.765 1419.035 368.045 ;
        RECT 1419.465 367.765 1419.745 368.045 ;
        RECT 1414.495 367.055 1414.775 367.335 ;
        RECT 1415.205 367.055 1415.485 367.335 ;
        RECT 1415.915 367.055 1416.195 367.335 ;
        RECT 1416.625 367.055 1416.905 367.335 ;
        RECT 1417.335 367.055 1417.615 367.335 ;
        RECT 1418.045 367.055 1418.325 367.335 ;
        RECT 1418.755 367.055 1419.035 367.335 ;
        RECT 1419.465 367.055 1419.745 367.335 ;
        RECT 1414.495 366.345 1414.775 366.625 ;
        RECT 1415.205 366.345 1415.485 366.625 ;
        RECT 1415.915 366.345 1416.195 366.625 ;
        RECT 1416.625 366.345 1416.905 366.625 ;
        RECT 1417.335 366.345 1417.615 366.625 ;
        RECT 1418.045 366.345 1418.325 366.625 ;
        RECT 1418.755 366.345 1419.035 366.625 ;
        RECT 1419.465 366.345 1419.745 366.625 ;
        RECT 1414.495 365.635 1414.775 365.915 ;
        RECT 1415.205 365.635 1415.485 365.915 ;
        RECT 1415.915 365.635 1416.195 365.915 ;
        RECT 1416.625 365.635 1416.905 365.915 ;
        RECT 1417.335 365.635 1417.615 365.915 ;
        RECT 1418.045 365.635 1418.325 365.915 ;
        RECT 1418.755 365.635 1419.035 365.915 ;
        RECT 1419.465 365.635 1419.745 365.915 ;
        RECT 1414.495 364.925 1414.775 365.205 ;
        RECT 1415.205 364.925 1415.485 365.205 ;
        RECT 1415.915 364.925 1416.195 365.205 ;
        RECT 1416.625 364.925 1416.905 365.205 ;
        RECT 1417.335 364.925 1417.615 365.205 ;
        RECT 1418.045 364.925 1418.325 365.205 ;
        RECT 1418.755 364.925 1419.035 365.205 ;
        RECT 1419.465 364.925 1419.745 365.205 ;
        RECT 1414.495 364.215 1414.775 364.495 ;
        RECT 1415.205 364.215 1415.485 364.495 ;
        RECT 1415.915 364.215 1416.195 364.495 ;
        RECT 1416.625 364.215 1416.905 364.495 ;
        RECT 1417.335 364.215 1417.615 364.495 ;
        RECT 1418.045 364.215 1418.325 364.495 ;
        RECT 1418.755 364.215 1419.035 364.495 ;
        RECT 1419.465 364.215 1419.745 364.495 ;
        RECT 1414.495 363.505 1414.775 363.785 ;
        RECT 1415.205 363.505 1415.485 363.785 ;
        RECT 1415.915 363.505 1416.195 363.785 ;
        RECT 1416.625 363.505 1416.905 363.785 ;
        RECT 1417.335 363.505 1417.615 363.785 ;
        RECT 1418.045 363.505 1418.325 363.785 ;
        RECT 1418.755 363.505 1419.035 363.785 ;
        RECT 1419.465 363.505 1419.745 363.785 ;
        RECT 1414.495 362.795 1414.775 363.075 ;
        RECT 1415.205 362.795 1415.485 363.075 ;
        RECT 1415.915 362.795 1416.195 363.075 ;
        RECT 1416.625 362.795 1416.905 363.075 ;
        RECT 1417.335 362.795 1417.615 363.075 ;
        RECT 1418.045 362.795 1418.325 363.075 ;
        RECT 1418.755 362.795 1419.035 363.075 ;
        RECT 1419.465 362.795 1419.745 363.075 ;
        RECT 1414.495 362.085 1414.775 362.365 ;
        RECT 1415.205 362.085 1415.485 362.365 ;
        RECT 1415.915 362.085 1416.195 362.365 ;
        RECT 1416.625 362.085 1416.905 362.365 ;
        RECT 1417.335 362.085 1417.615 362.365 ;
        RECT 1418.045 362.085 1418.325 362.365 ;
        RECT 1418.755 362.085 1419.035 362.365 ;
        RECT 1419.465 362.085 1419.745 362.365 ;
        RECT 1414.495 361.375 1414.775 361.655 ;
        RECT 1415.205 361.375 1415.485 361.655 ;
        RECT 1415.915 361.375 1416.195 361.655 ;
        RECT 1416.625 361.375 1416.905 361.655 ;
        RECT 1417.335 361.375 1417.615 361.655 ;
        RECT 1418.045 361.375 1418.325 361.655 ;
        RECT 1418.755 361.375 1419.035 361.655 ;
        RECT 1419.465 361.375 1419.745 361.655 ;
        RECT 1414.495 360.665 1414.775 360.945 ;
        RECT 1415.205 360.665 1415.485 360.945 ;
        RECT 1415.915 360.665 1416.195 360.945 ;
        RECT 1416.625 360.665 1416.905 360.945 ;
        RECT 1417.335 360.665 1417.615 360.945 ;
        RECT 1418.045 360.665 1418.325 360.945 ;
        RECT 1418.755 360.665 1419.035 360.945 ;
        RECT 1419.465 360.665 1419.745 360.945 ;
        RECT 3001.715 369.895 3001.995 370.175 ;
        RECT 3002.425 369.895 3002.705 370.175 ;
        RECT 3003.135 369.895 3003.415 370.175 ;
        RECT 3003.845 369.895 3004.125 370.175 ;
        RECT 3004.555 369.895 3004.835 370.175 ;
        RECT 3005.265 369.895 3005.545 370.175 ;
        RECT 3005.975 369.895 3006.255 370.175 ;
        RECT 3006.685 369.895 3006.965 370.175 ;
        RECT 3007.395 369.895 3007.675 370.175 ;
        RECT 3008.105 369.895 3008.385 370.175 ;
        RECT 3008.815 369.895 3009.095 370.175 ;
        RECT 3009.525 369.895 3009.805 370.175 ;
        RECT 3010.235 369.895 3010.515 370.175 ;
        RECT 3001.715 369.185 3001.995 369.465 ;
        RECT 3002.425 369.185 3002.705 369.465 ;
        RECT 3003.135 369.185 3003.415 369.465 ;
        RECT 3003.845 369.185 3004.125 369.465 ;
        RECT 3004.555 369.185 3004.835 369.465 ;
        RECT 3005.265 369.185 3005.545 369.465 ;
        RECT 3005.975 369.185 3006.255 369.465 ;
        RECT 3006.685 369.185 3006.965 369.465 ;
        RECT 3007.395 369.185 3007.675 369.465 ;
        RECT 3008.105 369.185 3008.385 369.465 ;
        RECT 3008.815 369.185 3009.095 369.465 ;
        RECT 3009.525 369.185 3009.805 369.465 ;
        RECT 3010.235 369.185 3010.515 369.465 ;
        RECT 3001.715 368.475 3001.995 368.755 ;
        RECT 3002.425 368.475 3002.705 368.755 ;
        RECT 3003.135 368.475 3003.415 368.755 ;
        RECT 3003.845 368.475 3004.125 368.755 ;
        RECT 3004.555 368.475 3004.835 368.755 ;
        RECT 3005.265 368.475 3005.545 368.755 ;
        RECT 3005.975 368.475 3006.255 368.755 ;
        RECT 3006.685 368.475 3006.965 368.755 ;
        RECT 3007.395 368.475 3007.675 368.755 ;
        RECT 3008.105 368.475 3008.385 368.755 ;
        RECT 3008.815 368.475 3009.095 368.755 ;
        RECT 3009.525 368.475 3009.805 368.755 ;
        RECT 3010.235 368.475 3010.515 368.755 ;
        RECT 3001.715 367.765 3001.995 368.045 ;
        RECT 3002.425 367.765 3002.705 368.045 ;
        RECT 3003.135 367.765 3003.415 368.045 ;
        RECT 3003.845 367.765 3004.125 368.045 ;
        RECT 3004.555 367.765 3004.835 368.045 ;
        RECT 3005.265 367.765 3005.545 368.045 ;
        RECT 3005.975 367.765 3006.255 368.045 ;
        RECT 3006.685 367.765 3006.965 368.045 ;
        RECT 3007.395 367.765 3007.675 368.045 ;
        RECT 3008.105 367.765 3008.385 368.045 ;
        RECT 3008.815 367.765 3009.095 368.045 ;
        RECT 3009.525 367.765 3009.805 368.045 ;
        RECT 3010.235 367.765 3010.515 368.045 ;
        RECT 3001.715 367.055 3001.995 367.335 ;
        RECT 3002.425 367.055 3002.705 367.335 ;
        RECT 3003.135 367.055 3003.415 367.335 ;
        RECT 3003.845 367.055 3004.125 367.335 ;
        RECT 3004.555 367.055 3004.835 367.335 ;
        RECT 3005.265 367.055 3005.545 367.335 ;
        RECT 3005.975 367.055 3006.255 367.335 ;
        RECT 3006.685 367.055 3006.965 367.335 ;
        RECT 3007.395 367.055 3007.675 367.335 ;
        RECT 3008.105 367.055 3008.385 367.335 ;
        RECT 3008.815 367.055 3009.095 367.335 ;
        RECT 3009.525 367.055 3009.805 367.335 ;
        RECT 3010.235 367.055 3010.515 367.335 ;
        RECT 3001.715 366.345 3001.995 366.625 ;
        RECT 3002.425 366.345 3002.705 366.625 ;
        RECT 3003.135 366.345 3003.415 366.625 ;
        RECT 3003.845 366.345 3004.125 366.625 ;
        RECT 3004.555 366.345 3004.835 366.625 ;
        RECT 3005.265 366.345 3005.545 366.625 ;
        RECT 3005.975 366.345 3006.255 366.625 ;
        RECT 3006.685 366.345 3006.965 366.625 ;
        RECT 3007.395 366.345 3007.675 366.625 ;
        RECT 3008.105 366.345 3008.385 366.625 ;
        RECT 3008.815 366.345 3009.095 366.625 ;
        RECT 3009.525 366.345 3009.805 366.625 ;
        RECT 3010.235 366.345 3010.515 366.625 ;
        RECT 3001.715 365.635 3001.995 365.915 ;
        RECT 3002.425 365.635 3002.705 365.915 ;
        RECT 3003.135 365.635 3003.415 365.915 ;
        RECT 3003.845 365.635 3004.125 365.915 ;
        RECT 3004.555 365.635 3004.835 365.915 ;
        RECT 3005.265 365.635 3005.545 365.915 ;
        RECT 3005.975 365.635 3006.255 365.915 ;
        RECT 3006.685 365.635 3006.965 365.915 ;
        RECT 3007.395 365.635 3007.675 365.915 ;
        RECT 3008.105 365.635 3008.385 365.915 ;
        RECT 3008.815 365.635 3009.095 365.915 ;
        RECT 3009.525 365.635 3009.805 365.915 ;
        RECT 3010.235 365.635 3010.515 365.915 ;
        RECT 3001.715 364.925 3001.995 365.205 ;
        RECT 3002.425 364.925 3002.705 365.205 ;
        RECT 3003.135 364.925 3003.415 365.205 ;
        RECT 3003.845 364.925 3004.125 365.205 ;
        RECT 3004.555 364.925 3004.835 365.205 ;
        RECT 3005.265 364.925 3005.545 365.205 ;
        RECT 3005.975 364.925 3006.255 365.205 ;
        RECT 3006.685 364.925 3006.965 365.205 ;
        RECT 3007.395 364.925 3007.675 365.205 ;
        RECT 3008.105 364.925 3008.385 365.205 ;
        RECT 3008.815 364.925 3009.095 365.205 ;
        RECT 3009.525 364.925 3009.805 365.205 ;
        RECT 3010.235 364.925 3010.515 365.205 ;
        RECT 3001.715 364.215 3001.995 364.495 ;
        RECT 3002.425 364.215 3002.705 364.495 ;
        RECT 3003.135 364.215 3003.415 364.495 ;
        RECT 3003.845 364.215 3004.125 364.495 ;
        RECT 3004.555 364.215 3004.835 364.495 ;
        RECT 3005.265 364.215 3005.545 364.495 ;
        RECT 3005.975 364.215 3006.255 364.495 ;
        RECT 3006.685 364.215 3006.965 364.495 ;
        RECT 3007.395 364.215 3007.675 364.495 ;
        RECT 3008.105 364.215 3008.385 364.495 ;
        RECT 3008.815 364.215 3009.095 364.495 ;
        RECT 3009.525 364.215 3009.805 364.495 ;
        RECT 3010.235 364.215 3010.515 364.495 ;
        RECT 3001.715 363.505 3001.995 363.785 ;
        RECT 3002.425 363.505 3002.705 363.785 ;
        RECT 3003.135 363.505 3003.415 363.785 ;
        RECT 3003.845 363.505 3004.125 363.785 ;
        RECT 3004.555 363.505 3004.835 363.785 ;
        RECT 3005.265 363.505 3005.545 363.785 ;
        RECT 3005.975 363.505 3006.255 363.785 ;
        RECT 3006.685 363.505 3006.965 363.785 ;
        RECT 3007.395 363.505 3007.675 363.785 ;
        RECT 3008.105 363.505 3008.385 363.785 ;
        RECT 3008.815 363.505 3009.095 363.785 ;
        RECT 3009.525 363.505 3009.805 363.785 ;
        RECT 3010.235 363.505 3010.515 363.785 ;
        RECT 3001.715 362.795 3001.995 363.075 ;
        RECT 3002.425 362.795 3002.705 363.075 ;
        RECT 3003.135 362.795 3003.415 363.075 ;
        RECT 3003.845 362.795 3004.125 363.075 ;
        RECT 3004.555 362.795 3004.835 363.075 ;
        RECT 3005.265 362.795 3005.545 363.075 ;
        RECT 3005.975 362.795 3006.255 363.075 ;
        RECT 3006.685 362.795 3006.965 363.075 ;
        RECT 3007.395 362.795 3007.675 363.075 ;
        RECT 3008.105 362.795 3008.385 363.075 ;
        RECT 3008.815 362.795 3009.095 363.075 ;
        RECT 3009.525 362.795 3009.805 363.075 ;
        RECT 3010.235 362.795 3010.515 363.075 ;
        RECT 3001.715 362.085 3001.995 362.365 ;
        RECT 3002.425 362.085 3002.705 362.365 ;
        RECT 3003.135 362.085 3003.415 362.365 ;
        RECT 3003.845 362.085 3004.125 362.365 ;
        RECT 3004.555 362.085 3004.835 362.365 ;
        RECT 3005.265 362.085 3005.545 362.365 ;
        RECT 3005.975 362.085 3006.255 362.365 ;
        RECT 3006.685 362.085 3006.965 362.365 ;
        RECT 3007.395 362.085 3007.675 362.365 ;
        RECT 3008.105 362.085 3008.385 362.365 ;
        RECT 3008.815 362.085 3009.095 362.365 ;
        RECT 3009.525 362.085 3009.805 362.365 ;
        RECT 3010.235 362.085 3010.515 362.365 ;
        RECT 3001.715 361.375 3001.995 361.655 ;
        RECT 3002.425 361.375 3002.705 361.655 ;
        RECT 3003.135 361.375 3003.415 361.655 ;
        RECT 3003.845 361.375 3004.125 361.655 ;
        RECT 3004.555 361.375 3004.835 361.655 ;
        RECT 3005.265 361.375 3005.545 361.655 ;
        RECT 3005.975 361.375 3006.255 361.655 ;
        RECT 3006.685 361.375 3006.965 361.655 ;
        RECT 3007.395 361.375 3007.675 361.655 ;
        RECT 3008.105 361.375 3008.385 361.655 ;
        RECT 3008.815 361.375 3009.095 361.655 ;
        RECT 3009.525 361.375 3009.805 361.655 ;
        RECT 3010.235 361.375 3010.515 361.655 ;
        RECT 3001.715 360.665 3001.995 360.945 ;
        RECT 3002.425 360.665 3002.705 360.945 ;
        RECT 3003.135 360.665 3003.415 360.945 ;
        RECT 3003.845 360.665 3004.125 360.945 ;
        RECT 3004.555 360.665 3004.835 360.945 ;
        RECT 3005.265 360.665 3005.545 360.945 ;
        RECT 3005.975 360.665 3006.255 360.945 ;
        RECT 3006.685 360.665 3006.965 360.945 ;
        RECT 3007.395 360.665 3007.675 360.945 ;
        RECT 3008.105 360.665 3008.385 360.945 ;
        RECT 3008.815 360.665 3009.095 360.945 ;
        RECT 3009.525 360.665 3009.805 360.945 ;
        RECT 3010.235 360.665 3010.515 360.945 ;
        RECT 3014.115 369.895 3014.395 370.175 ;
        RECT 3014.825 369.895 3015.105 370.175 ;
        RECT 3015.535 369.895 3015.815 370.175 ;
        RECT 3016.245 369.895 3016.525 370.175 ;
        RECT 3016.955 369.895 3017.235 370.175 ;
        RECT 3017.665 369.895 3017.945 370.175 ;
        RECT 3018.375 369.895 3018.655 370.175 ;
        RECT 3019.085 369.895 3019.365 370.175 ;
        RECT 3019.795 369.895 3020.075 370.175 ;
        RECT 3014.115 369.185 3014.395 369.465 ;
        RECT 3014.825 369.185 3015.105 369.465 ;
        RECT 3015.535 369.185 3015.815 369.465 ;
        RECT 3016.245 369.185 3016.525 369.465 ;
        RECT 3016.955 369.185 3017.235 369.465 ;
        RECT 3017.665 369.185 3017.945 369.465 ;
        RECT 3018.375 369.185 3018.655 369.465 ;
        RECT 3019.085 369.185 3019.365 369.465 ;
        RECT 3019.795 369.185 3020.075 369.465 ;
        RECT 3014.115 368.475 3014.395 368.755 ;
        RECT 3014.825 368.475 3015.105 368.755 ;
        RECT 3015.535 368.475 3015.815 368.755 ;
        RECT 3016.245 368.475 3016.525 368.755 ;
        RECT 3016.955 368.475 3017.235 368.755 ;
        RECT 3017.665 368.475 3017.945 368.755 ;
        RECT 3018.375 368.475 3018.655 368.755 ;
        RECT 3019.085 368.475 3019.365 368.755 ;
        RECT 3019.795 368.475 3020.075 368.755 ;
        RECT 3014.115 367.765 3014.395 368.045 ;
        RECT 3014.825 367.765 3015.105 368.045 ;
        RECT 3015.535 367.765 3015.815 368.045 ;
        RECT 3016.245 367.765 3016.525 368.045 ;
        RECT 3016.955 367.765 3017.235 368.045 ;
        RECT 3017.665 367.765 3017.945 368.045 ;
        RECT 3018.375 367.765 3018.655 368.045 ;
        RECT 3019.085 367.765 3019.365 368.045 ;
        RECT 3019.795 367.765 3020.075 368.045 ;
        RECT 3014.115 367.055 3014.395 367.335 ;
        RECT 3014.825 367.055 3015.105 367.335 ;
        RECT 3015.535 367.055 3015.815 367.335 ;
        RECT 3016.245 367.055 3016.525 367.335 ;
        RECT 3016.955 367.055 3017.235 367.335 ;
        RECT 3017.665 367.055 3017.945 367.335 ;
        RECT 3018.375 367.055 3018.655 367.335 ;
        RECT 3019.085 367.055 3019.365 367.335 ;
        RECT 3019.795 367.055 3020.075 367.335 ;
        RECT 3014.115 366.345 3014.395 366.625 ;
        RECT 3014.825 366.345 3015.105 366.625 ;
        RECT 3015.535 366.345 3015.815 366.625 ;
        RECT 3016.245 366.345 3016.525 366.625 ;
        RECT 3016.955 366.345 3017.235 366.625 ;
        RECT 3017.665 366.345 3017.945 366.625 ;
        RECT 3018.375 366.345 3018.655 366.625 ;
        RECT 3019.085 366.345 3019.365 366.625 ;
        RECT 3019.795 366.345 3020.075 366.625 ;
        RECT 3014.115 365.635 3014.395 365.915 ;
        RECT 3014.825 365.635 3015.105 365.915 ;
        RECT 3015.535 365.635 3015.815 365.915 ;
        RECT 3016.245 365.635 3016.525 365.915 ;
        RECT 3016.955 365.635 3017.235 365.915 ;
        RECT 3017.665 365.635 3017.945 365.915 ;
        RECT 3018.375 365.635 3018.655 365.915 ;
        RECT 3019.085 365.635 3019.365 365.915 ;
        RECT 3019.795 365.635 3020.075 365.915 ;
        RECT 3014.115 364.925 3014.395 365.205 ;
        RECT 3014.825 364.925 3015.105 365.205 ;
        RECT 3015.535 364.925 3015.815 365.205 ;
        RECT 3016.245 364.925 3016.525 365.205 ;
        RECT 3016.955 364.925 3017.235 365.205 ;
        RECT 3017.665 364.925 3017.945 365.205 ;
        RECT 3018.375 364.925 3018.655 365.205 ;
        RECT 3019.085 364.925 3019.365 365.205 ;
        RECT 3019.795 364.925 3020.075 365.205 ;
        RECT 3014.115 364.215 3014.395 364.495 ;
        RECT 3014.825 364.215 3015.105 364.495 ;
        RECT 3015.535 364.215 3015.815 364.495 ;
        RECT 3016.245 364.215 3016.525 364.495 ;
        RECT 3016.955 364.215 3017.235 364.495 ;
        RECT 3017.665 364.215 3017.945 364.495 ;
        RECT 3018.375 364.215 3018.655 364.495 ;
        RECT 3019.085 364.215 3019.365 364.495 ;
        RECT 3019.795 364.215 3020.075 364.495 ;
        RECT 3014.115 363.505 3014.395 363.785 ;
        RECT 3014.825 363.505 3015.105 363.785 ;
        RECT 3015.535 363.505 3015.815 363.785 ;
        RECT 3016.245 363.505 3016.525 363.785 ;
        RECT 3016.955 363.505 3017.235 363.785 ;
        RECT 3017.665 363.505 3017.945 363.785 ;
        RECT 3018.375 363.505 3018.655 363.785 ;
        RECT 3019.085 363.505 3019.365 363.785 ;
        RECT 3019.795 363.505 3020.075 363.785 ;
        RECT 3014.115 362.795 3014.395 363.075 ;
        RECT 3014.825 362.795 3015.105 363.075 ;
        RECT 3015.535 362.795 3015.815 363.075 ;
        RECT 3016.245 362.795 3016.525 363.075 ;
        RECT 3016.955 362.795 3017.235 363.075 ;
        RECT 3017.665 362.795 3017.945 363.075 ;
        RECT 3018.375 362.795 3018.655 363.075 ;
        RECT 3019.085 362.795 3019.365 363.075 ;
        RECT 3019.795 362.795 3020.075 363.075 ;
        RECT 3014.115 362.085 3014.395 362.365 ;
        RECT 3014.825 362.085 3015.105 362.365 ;
        RECT 3015.535 362.085 3015.815 362.365 ;
        RECT 3016.245 362.085 3016.525 362.365 ;
        RECT 3016.955 362.085 3017.235 362.365 ;
        RECT 3017.665 362.085 3017.945 362.365 ;
        RECT 3018.375 362.085 3018.655 362.365 ;
        RECT 3019.085 362.085 3019.365 362.365 ;
        RECT 3019.795 362.085 3020.075 362.365 ;
        RECT 3014.115 361.375 3014.395 361.655 ;
        RECT 3014.825 361.375 3015.105 361.655 ;
        RECT 3015.535 361.375 3015.815 361.655 ;
        RECT 3016.245 361.375 3016.525 361.655 ;
        RECT 3016.955 361.375 3017.235 361.655 ;
        RECT 3017.665 361.375 3017.945 361.655 ;
        RECT 3018.375 361.375 3018.655 361.655 ;
        RECT 3019.085 361.375 3019.365 361.655 ;
        RECT 3019.795 361.375 3020.075 361.655 ;
        RECT 3014.115 360.665 3014.395 360.945 ;
        RECT 3014.825 360.665 3015.105 360.945 ;
        RECT 3015.535 360.665 3015.815 360.945 ;
        RECT 3016.245 360.665 3016.525 360.945 ;
        RECT 3016.955 360.665 3017.235 360.945 ;
        RECT 3017.665 360.665 3017.945 360.945 ;
        RECT 3018.375 360.665 3018.655 360.945 ;
        RECT 3019.085 360.665 3019.365 360.945 ;
        RECT 3019.795 360.665 3020.075 360.945 ;
        RECT 3025.965 369.895 3026.245 370.175 ;
        RECT 3026.675 369.895 3026.955 370.175 ;
        RECT 3027.385 369.895 3027.665 370.175 ;
        RECT 3028.095 369.895 3028.375 370.175 ;
        RECT 3028.805 369.895 3029.085 370.175 ;
        RECT 3029.515 369.895 3029.795 370.175 ;
        RECT 3030.225 369.895 3030.505 370.175 ;
        RECT 3030.935 369.895 3031.215 370.175 ;
        RECT 3031.645 369.895 3031.925 370.175 ;
        RECT 3032.355 369.895 3032.635 370.175 ;
        RECT 3033.065 369.895 3033.345 370.175 ;
        RECT 3033.775 369.895 3034.055 370.175 ;
        RECT 3034.485 369.895 3034.765 370.175 ;
        RECT 3035.195 369.895 3035.475 370.175 ;
        RECT 3025.965 369.185 3026.245 369.465 ;
        RECT 3026.675 369.185 3026.955 369.465 ;
        RECT 3027.385 369.185 3027.665 369.465 ;
        RECT 3028.095 369.185 3028.375 369.465 ;
        RECT 3028.805 369.185 3029.085 369.465 ;
        RECT 3029.515 369.185 3029.795 369.465 ;
        RECT 3030.225 369.185 3030.505 369.465 ;
        RECT 3030.935 369.185 3031.215 369.465 ;
        RECT 3031.645 369.185 3031.925 369.465 ;
        RECT 3032.355 369.185 3032.635 369.465 ;
        RECT 3033.065 369.185 3033.345 369.465 ;
        RECT 3033.775 369.185 3034.055 369.465 ;
        RECT 3034.485 369.185 3034.765 369.465 ;
        RECT 3035.195 369.185 3035.475 369.465 ;
        RECT 3025.965 368.475 3026.245 368.755 ;
        RECT 3026.675 368.475 3026.955 368.755 ;
        RECT 3027.385 368.475 3027.665 368.755 ;
        RECT 3028.095 368.475 3028.375 368.755 ;
        RECT 3028.805 368.475 3029.085 368.755 ;
        RECT 3029.515 368.475 3029.795 368.755 ;
        RECT 3030.225 368.475 3030.505 368.755 ;
        RECT 3030.935 368.475 3031.215 368.755 ;
        RECT 3031.645 368.475 3031.925 368.755 ;
        RECT 3032.355 368.475 3032.635 368.755 ;
        RECT 3033.065 368.475 3033.345 368.755 ;
        RECT 3033.775 368.475 3034.055 368.755 ;
        RECT 3034.485 368.475 3034.765 368.755 ;
        RECT 3035.195 368.475 3035.475 368.755 ;
        RECT 3025.965 367.765 3026.245 368.045 ;
        RECT 3026.675 367.765 3026.955 368.045 ;
        RECT 3027.385 367.765 3027.665 368.045 ;
        RECT 3028.095 367.765 3028.375 368.045 ;
        RECT 3028.805 367.765 3029.085 368.045 ;
        RECT 3029.515 367.765 3029.795 368.045 ;
        RECT 3030.225 367.765 3030.505 368.045 ;
        RECT 3030.935 367.765 3031.215 368.045 ;
        RECT 3031.645 367.765 3031.925 368.045 ;
        RECT 3032.355 367.765 3032.635 368.045 ;
        RECT 3033.065 367.765 3033.345 368.045 ;
        RECT 3033.775 367.765 3034.055 368.045 ;
        RECT 3034.485 367.765 3034.765 368.045 ;
        RECT 3035.195 367.765 3035.475 368.045 ;
        RECT 3025.965 367.055 3026.245 367.335 ;
        RECT 3026.675 367.055 3026.955 367.335 ;
        RECT 3027.385 367.055 3027.665 367.335 ;
        RECT 3028.095 367.055 3028.375 367.335 ;
        RECT 3028.805 367.055 3029.085 367.335 ;
        RECT 3029.515 367.055 3029.795 367.335 ;
        RECT 3030.225 367.055 3030.505 367.335 ;
        RECT 3030.935 367.055 3031.215 367.335 ;
        RECT 3031.645 367.055 3031.925 367.335 ;
        RECT 3032.355 367.055 3032.635 367.335 ;
        RECT 3033.065 367.055 3033.345 367.335 ;
        RECT 3033.775 367.055 3034.055 367.335 ;
        RECT 3034.485 367.055 3034.765 367.335 ;
        RECT 3035.195 367.055 3035.475 367.335 ;
        RECT 3025.965 366.345 3026.245 366.625 ;
        RECT 3026.675 366.345 3026.955 366.625 ;
        RECT 3027.385 366.345 3027.665 366.625 ;
        RECT 3028.095 366.345 3028.375 366.625 ;
        RECT 3028.805 366.345 3029.085 366.625 ;
        RECT 3029.515 366.345 3029.795 366.625 ;
        RECT 3030.225 366.345 3030.505 366.625 ;
        RECT 3030.935 366.345 3031.215 366.625 ;
        RECT 3031.645 366.345 3031.925 366.625 ;
        RECT 3032.355 366.345 3032.635 366.625 ;
        RECT 3033.065 366.345 3033.345 366.625 ;
        RECT 3033.775 366.345 3034.055 366.625 ;
        RECT 3034.485 366.345 3034.765 366.625 ;
        RECT 3035.195 366.345 3035.475 366.625 ;
        RECT 3025.965 365.635 3026.245 365.915 ;
        RECT 3026.675 365.635 3026.955 365.915 ;
        RECT 3027.385 365.635 3027.665 365.915 ;
        RECT 3028.095 365.635 3028.375 365.915 ;
        RECT 3028.805 365.635 3029.085 365.915 ;
        RECT 3029.515 365.635 3029.795 365.915 ;
        RECT 3030.225 365.635 3030.505 365.915 ;
        RECT 3030.935 365.635 3031.215 365.915 ;
        RECT 3031.645 365.635 3031.925 365.915 ;
        RECT 3032.355 365.635 3032.635 365.915 ;
        RECT 3033.065 365.635 3033.345 365.915 ;
        RECT 3033.775 365.635 3034.055 365.915 ;
        RECT 3034.485 365.635 3034.765 365.915 ;
        RECT 3035.195 365.635 3035.475 365.915 ;
        RECT 3025.965 364.925 3026.245 365.205 ;
        RECT 3026.675 364.925 3026.955 365.205 ;
        RECT 3027.385 364.925 3027.665 365.205 ;
        RECT 3028.095 364.925 3028.375 365.205 ;
        RECT 3028.805 364.925 3029.085 365.205 ;
        RECT 3029.515 364.925 3029.795 365.205 ;
        RECT 3030.225 364.925 3030.505 365.205 ;
        RECT 3030.935 364.925 3031.215 365.205 ;
        RECT 3031.645 364.925 3031.925 365.205 ;
        RECT 3032.355 364.925 3032.635 365.205 ;
        RECT 3033.065 364.925 3033.345 365.205 ;
        RECT 3033.775 364.925 3034.055 365.205 ;
        RECT 3034.485 364.925 3034.765 365.205 ;
        RECT 3035.195 364.925 3035.475 365.205 ;
        RECT 3025.965 364.215 3026.245 364.495 ;
        RECT 3026.675 364.215 3026.955 364.495 ;
        RECT 3027.385 364.215 3027.665 364.495 ;
        RECT 3028.095 364.215 3028.375 364.495 ;
        RECT 3028.805 364.215 3029.085 364.495 ;
        RECT 3029.515 364.215 3029.795 364.495 ;
        RECT 3030.225 364.215 3030.505 364.495 ;
        RECT 3030.935 364.215 3031.215 364.495 ;
        RECT 3031.645 364.215 3031.925 364.495 ;
        RECT 3032.355 364.215 3032.635 364.495 ;
        RECT 3033.065 364.215 3033.345 364.495 ;
        RECT 3033.775 364.215 3034.055 364.495 ;
        RECT 3034.485 364.215 3034.765 364.495 ;
        RECT 3035.195 364.215 3035.475 364.495 ;
        RECT 3025.965 363.505 3026.245 363.785 ;
        RECT 3026.675 363.505 3026.955 363.785 ;
        RECT 3027.385 363.505 3027.665 363.785 ;
        RECT 3028.095 363.505 3028.375 363.785 ;
        RECT 3028.805 363.505 3029.085 363.785 ;
        RECT 3029.515 363.505 3029.795 363.785 ;
        RECT 3030.225 363.505 3030.505 363.785 ;
        RECT 3030.935 363.505 3031.215 363.785 ;
        RECT 3031.645 363.505 3031.925 363.785 ;
        RECT 3032.355 363.505 3032.635 363.785 ;
        RECT 3033.065 363.505 3033.345 363.785 ;
        RECT 3033.775 363.505 3034.055 363.785 ;
        RECT 3034.485 363.505 3034.765 363.785 ;
        RECT 3035.195 363.505 3035.475 363.785 ;
        RECT 3025.965 362.795 3026.245 363.075 ;
        RECT 3026.675 362.795 3026.955 363.075 ;
        RECT 3027.385 362.795 3027.665 363.075 ;
        RECT 3028.095 362.795 3028.375 363.075 ;
        RECT 3028.805 362.795 3029.085 363.075 ;
        RECT 3029.515 362.795 3029.795 363.075 ;
        RECT 3030.225 362.795 3030.505 363.075 ;
        RECT 3030.935 362.795 3031.215 363.075 ;
        RECT 3031.645 362.795 3031.925 363.075 ;
        RECT 3032.355 362.795 3032.635 363.075 ;
        RECT 3033.065 362.795 3033.345 363.075 ;
        RECT 3033.775 362.795 3034.055 363.075 ;
        RECT 3034.485 362.795 3034.765 363.075 ;
        RECT 3035.195 362.795 3035.475 363.075 ;
        RECT 3025.965 362.085 3026.245 362.365 ;
        RECT 3026.675 362.085 3026.955 362.365 ;
        RECT 3027.385 362.085 3027.665 362.365 ;
        RECT 3028.095 362.085 3028.375 362.365 ;
        RECT 3028.805 362.085 3029.085 362.365 ;
        RECT 3029.515 362.085 3029.795 362.365 ;
        RECT 3030.225 362.085 3030.505 362.365 ;
        RECT 3030.935 362.085 3031.215 362.365 ;
        RECT 3031.645 362.085 3031.925 362.365 ;
        RECT 3032.355 362.085 3032.635 362.365 ;
        RECT 3033.065 362.085 3033.345 362.365 ;
        RECT 3033.775 362.085 3034.055 362.365 ;
        RECT 3034.485 362.085 3034.765 362.365 ;
        RECT 3035.195 362.085 3035.475 362.365 ;
        RECT 3025.965 361.375 3026.245 361.655 ;
        RECT 3026.675 361.375 3026.955 361.655 ;
        RECT 3027.385 361.375 3027.665 361.655 ;
        RECT 3028.095 361.375 3028.375 361.655 ;
        RECT 3028.805 361.375 3029.085 361.655 ;
        RECT 3029.515 361.375 3029.795 361.655 ;
        RECT 3030.225 361.375 3030.505 361.655 ;
        RECT 3030.935 361.375 3031.215 361.655 ;
        RECT 3031.645 361.375 3031.925 361.655 ;
        RECT 3032.355 361.375 3032.635 361.655 ;
        RECT 3033.065 361.375 3033.345 361.655 ;
        RECT 3033.775 361.375 3034.055 361.655 ;
        RECT 3034.485 361.375 3034.765 361.655 ;
        RECT 3035.195 361.375 3035.475 361.655 ;
        RECT 3025.965 360.665 3026.245 360.945 ;
        RECT 3026.675 360.665 3026.955 360.945 ;
        RECT 3027.385 360.665 3027.665 360.945 ;
        RECT 3028.095 360.665 3028.375 360.945 ;
        RECT 3028.805 360.665 3029.085 360.945 ;
        RECT 3029.515 360.665 3029.795 360.945 ;
        RECT 3030.225 360.665 3030.505 360.945 ;
        RECT 3030.935 360.665 3031.215 360.945 ;
        RECT 3031.645 360.665 3031.925 360.945 ;
        RECT 3032.355 360.665 3032.635 360.945 ;
        RECT 3033.065 360.665 3033.345 360.945 ;
        RECT 3033.775 360.665 3034.055 360.945 ;
        RECT 3034.485 360.665 3034.765 360.945 ;
        RECT 3035.195 360.665 3035.475 360.945 ;
        RECT 3039.495 369.895 3039.775 370.175 ;
        RECT 3040.205 369.895 3040.485 370.175 ;
        RECT 3040.915 369.895 3041.195 370.175 ;
        RECT 3041.625 369.895 3041.905 370.175 ;
        RECT 3042.335 369.895 3042.615 370.175 ;
        RECT 3043.045 369.895 3043.325 370.175 ;
        RECT 3043.755 369.895 3044.035 370.175 ;
        RECT 3044.465 369.895 3044.745 370.175 ;
        RECT 3045.175 369.895 3045.455 370.175 ;
        RECT 3045.885 369.895 3046.165 370.175 ;
        RECT 3046.595 369.895 3046.875 370.175 ;
        RECT 3047.305 369.895 3047.585 370.175 ;
        RECT 3048.015 369.895 3048.295 370.175 ;
        RECT 3048.725 369.895 3049.005 370.175 ;
        RECT 3039.495 369.185 3039.775 369.465 ;
        RECT 3040.205 369.185 3040.485 369.465 ;
        RECT 3040.915 369.185 3041.195 369.465 ;
        RECT 3041.625 369.185 3041.905 369.465 ;
        RECT 3042.335 369.185 3042.615 369.465 ;
        RECT 3043.045 369.185 3043.325 369.465 ;
        RECT 3043.755 369.185 3044.035 369.465 ;
        RECT 3044.465 369.185 3044.745 369.465 ;
        RECT 3045.175 369.185 3045.455 369.465 ;
        RECT 3045.885 369.185 3046.165 369.465 ;
        RECT 3046.595 369.185 3046.875 369.465 ;
        RECT 3047.305 369.185 3047.585 369.465 ;
        RECT 3048.015 369.185 3048.295 369.465 ;
        RECT 3048.725 369.185 3049.005 369.465 ;
        RECT 3039.495 368.475 3039.775 368.755 ;
        RECT 3040.205 368.475 3040.485 368.755 ;
        RECT 3040.915 368.475 3041.195 368.755 ;
        RECT 3041.625 368.475 3041.905 368.755 ;
        RECT 3042.335 368.475 3042.615 368.755 ;
        RECT 3043.045 368.475 3043.325 368.755 ;
        RECT 3043.755 368.475 3044.035 368.755 ;
        RECT 3044.465 368.475 3044.745 368.755 ;
        RECT 3045.175 368.475 3045.455 368.755 ;
        RECT 3045.885 368.475 3046.165 368.755 ;
        RECT 3046.595 368.475 3046.875 368.755 ;
        RECT 3047.305 368.475 3047.585 368.755 ;
        RECT 3048.015 368.475 3048.295 368.755 ;
        RECT 3048.725 368.475 3049.005 368.755 ;
        RECT 3039.495 367.765 3039.775 368.045 ;
        RECT 3040.205 367.765 3040.485 368.045 ;
        RECT 3040.915 367.765 3041.195 368.045 ;
        RECT 3041.625 367.765 3041.905 368.045 ;
        RECT 3042.335 367.765 3042.615 368.045 ;
        RECT 3043.045 367.765 3043.325 368.045 ;
        RECT 3043.755 367.765 3044.035 368.045 ;
        RECT 3044.465 367.765 3044.745 368.045 ;
        RECT 3045.175 367.765 3045.455 368.045 ;
        RECT 3045.885 367.765 3046.165 368.045 ;
        RECT 3046.595 367.765 3046.875 368.045 ;
        RECT 3047.305 367.765 3047.585 368.045 ;
        RECT 3048.015 367.765 3048.295 368.045 ;
        RECT 3048.725 367.765 3049.005 368.045 ;
        RECT 3039.495 367.055 3039.775 367.335 ;
        RECT 3040.205 367.055 3040.485 367.335 ;
        RECT 3040.915 367.055 3041.195 367.335 ;
        RECT 3041.625 367.055 3041.905 367.335 ;
        RECT 3042.335 367.055 3042.615 367.335 ;
        RECT 3043.045 367.055 3043.325 367.335 ;
        RECT 3043.755 367.055 3044.035 367.335 ;
        RECT 3044.465 367.055 3044.745 367.335 ;
        RECT 3045.175 367.055 3045.455 367.335 ;
        RECT 3045.885 367.055 3046.165 367.335 ;
        RECT 3046.595 367.055 3046.875 367.335 ;
        RECT 3047.305 367.055 3047.585 367.335 ;
        RECT 3048.015 367.055 3048.295 367.335 ;
        RECT 3048.725 367.055 3049.005 367.335 ;
        RECT 3039.495 366.345 3039.775 366.625 ;
        RECT 3040.205 366.345 3040.485 366.625 ;
        RECT 3040.915 366.345 3041.195 366.625 ;
        RECT 3041.625 366.345 3041.905 366.625 ;
        RECT 3042.335 366.345 3042.615 366.625 ;
        RECT 3043.045 366.345 3043.325 366.625 ;
        RECT 3043.755 366.345 3044.035 366.625 ;
        RECT 3044.465 366.345 3044.745 366.625 ;
        RECT 3045.175 366.345 3045.455 366.625 ;
        RECT 3045.885 366.345 3046.165 366.625 ;
        RECT 3046.595 366.345 3046.875 366.625 ;
        RECT 3047.305 366.345 3047.585 366.625 ;
        RECT 3048.015 366.345 3048.295 366.625 ;
        RECT 3048.725 366.345 3049.005 366.625 ;
        RECT 3039.495 365.635 3039.775 365.915 ;
        RECT 3040.205 365.635 3040.485 365.915 ;
        RECT 3040.915 365.635 3041.195 365.915 ;
        RECT 3041.625 365.635 3041.905 365.915 ;
        RECT 3042.335 365.635 3042.615 365.915 ;
        RECT 3043.045 365.635 3043.325 365.915 ;
        RECT 3043.755 365.635 3044.035 365.915 ;
        RECT 3044.465 365.635 3044.745 365.915 ;
        RECT 3045.175 365.635 3045.455 365.915 ;
        RECT 3045.885 365.635 3046.165 365.915 ;
        RECT 3046.595 365.635 3046.875 365.915 ;
        RECT 3047.305 365.635 3047.585 365.915 ;
        RECT 3048.015 365.635 3048.295 365.915 ;
        RECT 3048.725 365.635 3049.005 365.915 ;
        RECT 3039.495 364.925 3039.775 365.205 ;
        RECT 3040.205 364.925 3040.485 365.205 ;
        RECT 3040.915 364.925 3041.195 365.205 ;
        RECT 3041.625 364.925 3041.905 365.205 ;
        RECT 3042.335 364.925 3042.615 365.205 ;
        RECT 3043.045 364.925 3043.325 365.205 ;
        RECT 3043.755 364.925 3044.035 365.205 ;
        RECT 3044.465 364.925 3044.745 365.205 ;
        RECT 3045.175 364.925 3045.455 365.205 ;
        RECT 3045.885 364.925 3046.165 365.205 ;
        RECT 3046.595 364.925 3046.875 365.205 ;
        RECT 3047.305 364.925 3047.585 365.205 ;
        RECT 3048.015 364.925 3048.295 365.205 ;
        RECT 3048.725 364.925 3049.005 365.205 ;
        RECT 3039.495 364.215 3039.775 364.495 ;
        RECT 3040.205 364.215 3040.485 364.495 ;
        RECT 3040.915 364.215 3041.195 364.495 ;
        RECT 3041.625 364.215 3041.905 364.495 ;
        RECT 3042.335 364.215 3042.615 364.495 ;
        RECT 3043.045 364.215 3043.325 364.495 ;
        RECT 3043.755 364.215 3044.035 364.495 ;
        RECT 3044.465 364.215 3044.745 364.495 ;
        RECT 3045.175 364.215 3045.455 364.495 ;
        RECT 3045.885 364.215 3046.165 364.495 ;
        RECT 3046.595 364.215 3046.875 364.495 ;
        RECT 3047.305 364.215 3047.585 364.495 ;
        RECT 3048.015 364.215 3048.295 364.495 ;
        RECT 3048.725 364.215 3049.005 364.495 ;
        RECT 3039.495 363.505 3039.775 363.785 ;
        RECT 3040.205 363.505 3040.485 363.785 ;
        RECT 3040.915 363.505 3041.195 363.785 ;
        RECT 3041.625 363.505 3041.905 363.785 ;
        RECT 3042.335 363.505 3042.615 363.785 ;
        RECT 3043.045 363.505 3043.325 363.785 ;
        RECT 3043.755 363.505 3044.035 363.785 ;
        RECT 3044.465 363.505 3044.745 363.785 ;
        RECT 3045.175 363.505 3045.455 363.785 ;
        RECT 3045.885 363.505 3046.165 363.785 ;
        RECT 3046.595 363.505 3046.875 363.785 ;
        RECT 3047.305 363.505 3047.585 363.785 ;
        RECT 3048.015 363.505 3048.295 363.785 ;
        RECT 3048.725 363.505 3049.005 363.785 ;
        RECT 3039.495 362.795 3039.775 363.075 ;
        RECT 3040.205 362.795 3040.485 363.075 ;
        RECT 3040.915 362.795 3041.195 363.075 ;
        RECT 3041.625 362.795 3041.905 363.075 ;
        RECT 3042.335 362.795 3042.615 363.075 ;
        RECT 3043.045 362.795 3043.325 363.075 ;
        RECT 3043.755 362.795 3044.035 363.075 ;
        RECT 3044.465 362.795 3044.745 363.075 ;
        RECT 3045.175 362.795 3045.455 363.075 ;
        RECT 3045.885 362.795 3046.165 363.075 ;
        RECT 3046.595 362.795 3046.875 363.075 ;
        RECT 3047.305 362.795 3047.585 363.075 ;
        RECT 3048.015 362.795 3048.295 363.075 ;
        RECT 3048.725 362.795 3049.005 363.075 ;
        RECT 3039.495 362.085 3039.775 362.365 ;
        RECT 3040.205 362.085 3040.485 362.365 ;
        RECT 3040.915 362.085 3041.195 362.365 ;
        RECT 3041.625 362.085 3041.905 362.365 ;
        RECT 3042.335 362.085 3042.615 362.365 ;
        RECT 3043.045 362.085 3043.325 362.365 ;
        RECT 3043.755 362.085 3044.035 362.365 ;
        RECT 3044.465 362.085 3044.745 362.365 ;
        RECT 3045.175 362.085 3045.455 362.365 ;
        RECT 3045.885 362.085 3046.165 362.365 ;
        RECT 3046.595 362.085 3046.875 362.365 ;
        RECT 3047.305 362.085 3047.585 362.365 ;
        RECT 3048.015 362.085 3048.295 362.365 ;
        RECT 3048.725 362.085 3049.005 362.365 ;
        RECT 3039.495 361.375 3039.775 361.655 ;
        RECT 3040.205 361.375 3040.485 361.655 ;
        RECT 3040.915 361.375 3041.195 361.655 ;
        RECT 3041.625 361.375 3041.905 361.655 ;
        RECT 3042.335 361.375 3042.615 361.655 ;
        RECT 3043.045 361.375 3043.325 361.655 ;
        RECT 3043.755 361.375 3044.035 361.655 ;
        RECT 3044.465 361.375 3044.745 361.655 ;
        RECT 3045.175 361.375 3045.455 361.655 ;
        RECT 3045.885 361.375 3046.165 361.655 ;
        RECT 3046.595 361.375 3046.875 361.655 ;
        RECT 3047.305 361.375 3047.585 361.655 ;
        RECT 3048.015 361.375 3048.295 361.655 ;
        RECT 3048.725 361.375 3049.005 361.655 ;
        RECT 3039.495 360.665 3039.775 360.945 ;
        RECT 3040.205 360.665 3040.485 360.945 ;
        RECT 3040.915 360.665 3041.195 360.945 ;
        RECT 3041.625 360.665 3041.905 360.945 ;
        RECT 3042.335 360.665 3042.615 360.945 ;
        RECT 3043.045 360.665 3043.325 360.945 ;
        RECT 3043.755 360.665 3044.035 360.945 ;
        RECT 3044.465 360.665 3044.745 360.945 ;
        RECT 3045.175 360.665 3045.455 360.945 ;
        RECT 3045.885 360.665 3046.165 360.945 ;
        RECT 3046.595 360.665 3046.875 360.945 ;
        RECT 3047.305 360.665 3047.585 360.945 ;
        RECT 3048.015 360.665 3048.295 360.945 ;
        RECT 3048.725 360.665 3049.005 360.945 ;
        RECT 3051.345 369.895 3051.625 370.175 ;
        RECT 3052.055 369.895 3052.335 370.175 ;
        RECT 3052.765 369.895 3053.045 370.175 ;
        RECT 3053.475 369.895 3053.755 370.175 ;
        RECT 3054.185 369.895 3054.465 370.175 ;
        RECT 3054.895 369.895 3055.175 370.175 ;
        RECT 3055.605 369.895 3055.885 370.175 ;
        RECT 3056.315 369.895 3056.595 370.175 ;
        RECT 3057.025 369.895 3057.305 370.175 ;
        RECT 3057.735 369.895 3058.015 370.175 ;
        RECT 3058.445 369.895 3058.725 370.175 ;
        RECT 3059.155 369.895 3059.435 370.175 ;
        RECT 3059.865 369.895 3060.145 370.175 ;
        RECT 3060.575 369.895 3060.855 370.175 ;
        RECT 3051.345 369.185 3051.625 369.465 ;
        RECT 3052.055 369.185 3052.335 369.465 ;
        RECT 3052.765 369.185 3053.045 369.465 ;
        RECT 3053.475 369.185 3053.755 369.465 ;
        RECT 3054.185 369.185 3054.465 369.465 ;
        RECT 3054.895 369.185 3055.175 369.465 ;
        RECT 3055.605 369.185 3055.885 369.465 ;
        RECT 3056.315 369.185 3056.595 369.465 ;
        RECT 3057.025 369.185 3057.305 369.465 ;
        RECT 3057.735 369.185 3058.015 369.465 ;
        RECT 3058.445 369.185 3058.725 369.465 ;
        RECT 3059.155 369.185 3059.435 369.465 ;
        RECT 3059.865 369.185 3060.145 369.465 ;
        RECT 3060.575 369.185 3060.855 369.465 ;
        RECT 3051.345 368.475 3051.625 368.755 ;
        RECT 3052.055 368.475 3052.335 368.755 ;
        RECT 3052.765 368.475 3053.045 368.755 ;
        RECT 3053.475 368.475 3053.755 368.755 ;
        RECT 3054.185 368.475 3054.465 368.755 ;
        RECT 3054.895 368.475 3055.175 368.755 ;
        RECT 3055.605 368.475 3055.885 368.755 ;
        RECT 3056.315 368.475 3056.595 368.755 ;
        RECT 3057.025 368.475 3057.305 368.755 ;
        RECT 3057.735 368.475 3058.015 368.755 ;
        RECT 3058.445 368.475 3058.725 368.755 ;
        RECT 3059.155 368.475 3059.435 368.755 ;
        RECT 3059.865 368.475 3060.145 368.755 ;
        RECT 3060.575 368.475 3060.855 368.755 ;
        RECT 3051.345 367.765 3051.625 368.045 ;
        RECT 3052.055 367.765 3052.335 368.045 ;
        RECT 3052.765 367.765 3053.045 368.045 ;
        RECT 3053.475 367.765 3053.755 368.045 ;
        RECT 3054.185 367.765 3054.465 368.045 ;
        RECT 3054.895 367.765 3055.175 368.045 ;
        RECT 3055.605 367.765 3055.885 368.045 ;
        RECT 3056.315 367.765 3056.595 368.045 ;
        RECT 3057.025 367.765 3057.305 368.045 ;
        RECT 3057.735 367.765 3058.015 368.045 ;
        RECT 3058.445 367.765 3058.725 368.045 ;
        RECT 3059.155 367.765 3059.435 368.045 ;
        RECT 3059.865 367.765 3060.145 368.045 ;
        RECT 3060.575 367.765 3060.855 368.045 ;
        RECT 3051.345 367.055 3051.625 367.335 ;
        RECT 3052.055 367.055 3052.335 367.335 ;
        RECT 3052.765 367.055 3053.045 367.335 ;
        RECT 3053.475 367.055 3053.755 367.335 ;
        RECT 3054.185 367.055 3054.465 367.335 ;
        RECT 3054.895 367.055 3055.175 367.335 ;
        RECT 3055.605 367.055 3055.885 367.335 ;
        RECT 3056.315 367.055 3056.595 367.335 ;
        RECT 3057.025 367.055 3057.305 367.335 ;
        RECT 3057.735 367.055 3058.015 367.335 ;
        RECT 3058.445 367.055 3058.725 367.335 ;
        RECT 3059.155 367.055 3059.435 367.335 ;
        RECT 3059.865 367.055 3060.145 367.335 ;
        RECT 3060.575 367.055 3060.855 367.335 ;
        RECT 3051.345 366.345 3051.625 366.625 ;
        RECT 3052.055 366.345 3052.335 366.625 ;
        RECT 3052.765 366.345 3053.045 366.625 ;
        RECT 3053.475 366.345 3053.755 366.625 ;
        RECT 3054.185 366.345 3054.465 366.625 ;
        RECT 3054.895 366.345 3055.175 366.625 ;
        RECT 3055.605 366.345 3055.885 366.625 ;
        RECT 3056.315 366.345 3056.595 366.625 ;
        RECT 3057.025 366.345 3057.305 366.625 ;
        RECT 3057.735 366.345 3058.015 366.625 ;
        RECT 3058.445 366.345 3058.725 366.625 ;
        RECT 3059.155 366.345 3059.435 366.625 ;
        RECT 3059.865 366.345 3060.145 366.625 ;
        RECT 3060.575 366.345 3060.855 366.625 ;
        RECT 3051.345 365.635 3051.625 365.915 ;
        RECT 3052.055 365.635 3052.335 365.915 ;
        RECT 3052.765 365.635 3053.045 365.915 ;
        RECT 3053.475 365.635 3053.755 365.915 ;
        RECT 3054.185 365.635 3054.465 365.915 ;
        RECT 3054.895 365.635 3055.175 365.915 ;
        RECT 3055.605 365.635 3055.885 365.915 ;
        RECT 3056.315 365.635 3056.595 365.915 ;
        RECT 3057.025 365.635 3057.305 365.915 ;
        RECT 3057.735 365.635 3058.015 365.915 ;
        RECT 3058.445 365.635 3058.725 365.915 ;
        RECT 3059.155 365.635 3059.435 365.915 ;
        RECT 3059.865 365.635 3060.145 365.915 ;
        RECT 3060.575 365.635 3060.855 365.915 ;
        RECT 3051.345 364.925 3051.625 365.205 ;
        RECT 3052.055 364.925 3052.335 365.205 ;
        RECT 3052.765 364.925 3053.045 365.205 ;
        RECT 3053.475 364.925 3053.755 365.205 ;
        RECT 3054.185 364.925 3054.465 365.205 ;
        RECT 3054.895 364.925 3055.175 365.205 ;
        RECT 3055.605 364.925 3055.885 365.205 ;
        RECT 3056.315 364.925 3056.595 365.205 ;
        RECT 3057.025 364.925 3057.305 365.205 ;
        RECT 3057.735 364.925 3058.015 365.205 ;
        RECT 3058.445 364.925 3058.725 365.205 ;
        RECT 3059.155 364.925 3059.435 365.205 ;
        RECT 3059.865 364.925 3060.145 365.205 ;
        RECT 3060.575 364.925 3060.855 365.205 ;
        RECT 3051.345 364.215 3051.625 364.495 ;
        RECT 3052.055 364.215 3052.335 364.495 ;
        RECT 3052.765 364.215 3053.045 364.495 ;
        RECT 3053.475 364.215 3053.755 364.495 ;
        RECT 3054.185 364.215 3054.465 364.495 ;
        RECT 3054.895 364.215 3055.175 364.495 ;
        RECT 3055.605 364.215 3055.885 364.495 ;
        RECT 3056.315 364.215 3056.595 364.495 ;
        RECT 3057.025 364.215 3057.305 364.495 ;
        RECT 3057.735 364.215 3058.015 364.495 ;
        RECT 3058.445 364.215 3058.725 364.495 ;
        RECT 3059.155 364.215 3059.435 364.495 ;
        RECT 3059.865 364.215 3060.145 364.495 ;
        RECT 3060.575 364.215 3060.855 364.495 ;
        RECT 3051.345 363.505 3051.625 363.785 ;
        RECT 3052.055 363.505 3052.335 363.785 ;
        RECT 3052.765 363.505 3053.045 363.785 ;
        RECT 3053.475 363.505 3053.755 363.785 ;
        RECT 3054.185 363.505 3054.465 363.785 ;
        RECT 3054.895 363.505 3055.175 363.785 ;
        RECT 3055.605 363.505 3055.885 363.785 ;
        RECT 3056.315 363.505 3056.595 363.785 ;
        RECT 3057.025 363.505 3057.305 363.785 ;
        RECT 3057.735 363.505 3058.015 363.785 ;
        RECT 3058.445 363.505 3058.725 363.785 ;
        RECT 3059.155 363.505 3059.435 363.785 ;
        RECT 3059.865 363.505 3060.145 363.785 ;
        RECT 3060.575 363.505 3060.855 363.785 ;
        RECT 3051.345 362.795 3051.625 363.075 ;
        RECT 3052.055 362.795 3052.335 363.075 ;
        RECT 3052.765 362.795 3053.045 363.075 ;
        RECT 3053.475 362.795 3053.755 363.075 ;
        RECT 3054.185 362.795 3054.465 363.075 ;
        RECT 3054.895 362.795 3055.175 363.075 ;
        RECT 3055.605 362.795 3055.885 363.075 ;
        RECT 3056.315 362.795 3056.595 363.075 ;
        RECT 3057.025 362.795 3057.305 363.075 ;
        RECT 3057.735 362.795 3058.015 363.075 ;
        RECT 3058.445 362.795 3058.725 363.075 ;
        RECT 3059.155 362.795 3059.435 363.075 ;
        RECT 3059.865 362.795 3060.145 363.075 ;
        RECT 3060.575 362.795 3060.855 363.075 ;
        RECT 3051.345 362.085 3051.625 362.365 ;
        RECT 3052.055 362.085 3052.335 362.365 ;
        RECT 3052.765 362.085 3053.045 362.365 ;
        RECT 3053.475 362.085 3053.755 362.365 ;
        RECT 3054.185 362.085 3054.465 362.365 ;
        RECT 3054.895 362.085 3055.175 362.365 ;
        RECT 3055.605 362.085 3055.885 362.365 ;
        RECT 3056.315 362.085 3056.595 362.365 ;
        RECT 3057.025 362.085 3057.305 362.365 ;
        RECT 3057.735 362.085 3058.015 362.365 ;
        RECT 3058.445 362.085 3058.725 362.365 ;
        RECT 3059.155 362.085 3059.435 362.365 ;
        RECT 3059.865 362.085 3060.145 362.365 ;
        RECT 3060.575 362.085 3060.855 362.365 ;
        RECT 3051.345 361.375 3051.625 361.655 ;
        RECT 3052.055 361.375 3052.335 361.655 ;
        RECT 3052.765 361.375 3053.045 361.655 ;
        RECT 3053.475 361.375 3053.755 361.655 ;
        RECT 3054.185 361.375 3054.465 361.655 ;
        RECT 3054.895 361.375 3055.175 361.655 ;
        RECT 3055.605 361.375 3055.885 361.655 ;
        RECT 3056.315 361.375 3056.595 361.655 ;
        RECT 3057.025 361.375 3057.305 361.655 ;
        RECT 3057.735 361.375 3058.015 361.655 ;
        RECT 3058.445 361.375 3058.725 361.655 ;
        RECT 3059.155 361.375 3059.435 361.655 ;
        RECT 3059.865 361.375 3060.145 361.655 ;
        RECT 3060.575 361.375 3060.855 361.655 ;
        RECT 3051.345 360.665 3051.625 360.945 ;
        RECT 3052.055 360.665 3052.335 360.945 ;
        RECT 3052.765 360.665 3053.045 360.945 ;
        RECT 3053.475 360.665 3053.755 360.945 ;
        RECT 3054.185 360.665 3054.465 360.945 ;
        RECT 3054.895 360.665 3055.175 360.945 ;
        RECT 3055.605 360.665 3055.885 360.945 ;
        RECT 3056.315 360.665 3056.595 360.945 ;
        RECT 3057.025 360.665 3057.305 360.945 ;
        RECT 3057.735 360.665 3058.015 360.945 ;
        RECT 3058.445 360.665 3058.725 360.945 ;
        RECT 3059.155 360.665 3059.435 360.945 ;
        RECT 3059.865 360.665 3060.145 360.945 ;
        RECT 3060.575 360.665 3060.855 360.945 ;
        RECT 3064.495 369.895 3064.775 370.175 ;
        RECT 3065.205 369.895 3065.485 370.175 ;
        RECT 3065.915 369.895 3066.195 370.175 ;
        RECT 3066.625 369.895 3066.905 370.175 ;
        RECT 3067.335 369.895 3067.615 370.175 ;
        RECT 3068.045 369.895 3068.325 370.175 ;
        RECT 3068.755 369.895 3069.035 370.175 ;
        RECT 3069.465 369.895 3069.745 370.175 ;
        RECT 3070.175 369.895 3070.455 370.175 ;
        RECT 3070.885 369.895 3071.165 370.175 ;
        RECT 3071.595 369.895 3071.875 370.175 ;
        RECT 3072.305 369.895 3072.585 370.175 ;
        RECT 3073.015 369.895 3073.295 370.175 ;
        RECT 3064.495 369.185 3064.775 369.465 ;
        RECT 3065.205 369.185 3065.485 369.465 ;
        RECT 3065.915 369.185 3066.195 369.465 ;
        RECT 3066.625 369.185 3066.905 369.465 ;
        RECT 3067.335 369.185 3067.615 369.465 ;
        RECT 3068.045 369.185 3068.325 369.465 ;
        RECT 3068.755 369.185 3069.035 369.465 ;
        RECT 3069.465 369.185 3069.745 369.465 ;
        RECT 3070.175 369.185 3070.455 369.465 ;
        RECT 3070.885 369.185 3071.165 369.465 ;
        RECT 3071.595 369.185 3071.875 369.465 ;
        RECT 3072.305 369.185 3072.585 369.465 ;
        RECT 3073.015 369.185 3073.295 369.465 ;
        RECT 3064.495 368.475 3064.775 368.755 ;
        RECT 3065.205 368.475 3065.485 368.755 ;
        RECT 3065.915 368.475 3066.195 368.755 ;
        RECT 3066.625 368.475 3066.905 368.755 ;
        RECT 3067.335 368.475 3067.615 368.755 ;
        RECT 3068.045 368.475 3068.325 368.755 ;
        RECT 3068.755 368.475 3069.035 368.755 ;
        RECT 3069.465 368.475 3069.745 368.755 ;
        RECT 3070.175 368.475 3070.455 368.755 ;
        RECT 3070.885 368.475 3071.165 368.755 ;
        RECT 3071.595 368.475 3071.875 368.755 ;
        RECT 3072.305 368.475 3072.585 368.755 ;
        RECT 3073.015 368.475 3073.295 368.755 ;
        RECT 3064.495 367.765 3064.775 368.045 ;
        RECT 3065.205 367.765 3065.485 368.045 ;
        RECT 3065.915 367.765 3066.195 368.045 ;
        RECT 3066.625 367.765 3066.905 368.045 ;
        RECT 3067.335 367.765 3067.615 368.045 ;
        RECT 3068.045 367.765 3068.325 368.045 ;
        RECT 3068.755 367.765 3069.035 368.045 ;
        RECT 3069.465 367.765 3069.745 368.045 ;
        RECT 3070.175 367.765 3070.455 368.045 ;
        RECT 3070.885 367.765 3071.165 368.045 ;
        RECT 3071.595 367.765 3071.875 368.045 ;
        RECT 3072.305 367.765 3072.585 368.045 ;
        RECT 3073.015 367.765 3073.295 368.045 ;
        RECT 3064.495 367.055 3064.775 367.335 ;
        RECT 3065.205 367.055 3065.485 367.335 ;
        RECT 3065.915 367.055 3066.195 367.335 ;
        RECT 3066.625 367.055 3066.905 367.335 ;
        RECT 3067.335 367.055 3067.615 367.335 ;
        RECT 3068.045 367.055 3068.325 367.335 ;
        RECT 3068.755 367.055 3069.035 367.335 ;
        RECT 3069.465 367.055 3069.745 367.335 ;
        RECT 3070.175 367.055 3070.455 367.335 ;
        RECT 3070.885 367.055 3071.165 367.335 ;
        RECT 3071.595 367.055 3071.875 367.335 ;
        RECT 3072.305 367.055 3072.585 367.335 ;
        RECT 3073.015 367.055 3073.295 367.335 ;
        RECT 3064.495 366.345 3064.775 366.625 ;
        RECT 3065.205 366.345 3065.485 366.625 ;
        RECT 3065.915 366.345 3066.195 366.625 ;
        RECT 3066.625 366.345 3066.905 366.625 ;
        RECT 3067.335 366.345 3067.615 366.625 ;
        RECT 3068.045 366.345 3068.325 366.625 ;
        RECT 3068.755 366.345 3069.035 366.625 ;
        RECT 3069.465 366.345 3069.745 366.625 ;
        RECT 3070.175 366.345 3070.455 366.625 ;
        RECT 3070.885 366.345 3071.165 366.625 ;
        RECT 3071.595 366.345 3071.875 366.625 ;
        RECT 3072.305 366.345 3072.585 366.625 ;
        RECT 3073.015 366.345 3073.295 366.625 ;
        RECT 3064.495 365.635 3064.775 365.915 ;
        RECT 3065.205 365.635 3065.485 365.915 ;
        RECT 3065.915 365.635 3066.195 365.915 ;
        RECT 3066.625 365.635 3066.905 365.915 ;
        RECT 3067.335 365.635 3067.615 365.915 ;
        RECT 3068.045 365.635 3068.325 365.915 ;
        RECT 3068.755 365.635 3069.035 365.915 ;
        RECT 3069.465 365.635 3069.745 365.915 ;
        RECT 3070.175 365.635 3070.455 365.915 ;
        RECT 3070.885 365.635 3071.165 365.915 ;
        RECT 3071.595 365.635 3071.875 365.915 ;
        RECT 3072.305 365.635 3072.585 365.915 ;
        RECT 3073.015 365.635 3073.295 365.915 ;
        RECT 3064.495 364.925 3064.775 365.205 ;
        RECT 3065.205 364.925 3065.485 365.205 ;
        RECT 3065.915 364.925 3066.195 365.205 ;
        RECT 3066.625 364.925 3066.905 365.205 ;
        RECT 3067.335 364.925 3067.615 365.205 ;
        RECT 3068.045 364.925 3068.325 365.205 ;
        RECT 3068.755 364.925 3069.035 365.205 ;
        RECT 3069.465 364.925 3069.745 365.205 ;
        RECT 3070.175 364.925 3070.455 365.205 ;
        RECT 3070.885 364.925 3071.165 365.205 ;
        RECT 3071.595 364.925 3071.875 365.205 ;
        RECT 3072.305 364.925 3072.585 365.205 ;
        RECT 3073.015 364.925 3073.295 365.205 ;
        RECT 3064.495 364.215 3064.775 364.495 ;
        RECT 3065.205 364.215 3065.485 364.495 ;
        RECT 3065.915 364.215 3066.195 364.495 ;
        RECT 3066.625 364.215 3066.905 364.495 ;
        RECT 3067.335 364.215 3067.615 364.495 ;
        RECT 3068.045 364.215 3068.325 364.495 ;
        RECT 3068.755 364.215 3069.035 364.495 ;
        RECT 3069.465 364.215 3069.745 364.495 ;
        RECT 3070.175 364.215 3070.455 364.495 ;
        RECT 3070.885 364.215 3071.165 364.495 ;
        RECT 3071.595 364.215 3071.875 364.495 ;
        RECT 3072.305 364.215 3072.585 364.495 ;
        RECT 3073.015 364.215 3073.295 364.495 ;
        RECT 3064.495 363.505 3064.775 363.785 ;
        RECT 3065.205 363.505 3065.485 363.785 ;
        RECT 3065.915 363.505 3066.195 363.785 ;
        RECT 3066.625 363.505 3066.905 363.785 ;
        RECT 3067.335 363.505 3067.615 363.785 ;
        RECT 3068.045 363.505 3068.325 363.785 ;
        RECT 3068.755 363.505 3069.035 363.785 ;
        RECT 3069.465 363.505 3069.745 363.785 ;
        RECT 3070.175 363.505 3070.455 363.785 ;
        RECT 3070.885 363.505 3071.165 363.785 ;
        RECT 3071.595 363.505 3071.875 363.785 ;
        RECT 3072.305 363.505 3072.585 363.785 ;
        RECT 3073.015 363.505 3073.295 363.785 ;
        RECT 3064.495 362.795 3064.775 363.075 ;
        RECT 3065.205 362.795 3065.485 363.075 ;
        RECT 3065.915 362.795 3066.195 363.075 ;
        RECT 3066.625 362.795 3066.905 363.075 ;
        RECT 3067.335 362.795 3067.615 363.075 ;
        RECT 3068.045 362.795 3068.325 363.075 ;
        RECT 3068.755 362.795 3069.035 363.075 ;
        RECT 3069.465 362.795 3069.745 363.075 ;
        RECT 3070.175 362.795 3070.455 363.075 ;
        RECT 3070.885 362.795 3071.165 363.075 ;
        RECT 3071.595 362.795 3071.875 363.075 ;
        RECT 3072.305 362.795 3072.585 363.075 ;
        RECT 3073.015 362.795 3073.295 363.075 ;
        RECT 3064.495 362.085 3064.775 362.365 ;
        RECT 3065.205 362.085 3065.485 362.365 ;
        RECT 3065.915 362.085 3066.195 362.365 ;
        RECT 3066.625 362.085 3066.905 362.365 ;
        RECT 3067.335 362.085 3067.615 362.365 ;
        RECT 3068.045 362.085 3068.325 362.365 ;
        RECT 3068.755 362.085 3069.035 362.365 ;
        RECT 3069.465 362.085 3069.745 362.365 ;
        RECT 3070.175 362.085 3070.455 362.365 ;
        RECT 3070.885 362.085 3071.165 362.365 ;
        RECT 3071.595 362.085 3071.875 362.365 ;
        RECT 3072.305 362.085 3072.585 362.365 ;
        RECT 3073.015 362.085 3073.295 362.365 ;
        RECT 3064.495 361.375 3064.775 361.655 ;
        RECT 3065.205 361.375 3065.485 361.655 ;
        RECT 3065.915 361.375 3066.195 361.655 ;
        RECT 3066.625 361.375 3066.905 361.655 ;
        RECT 3067.335 361.375 3067.615 361.655 ;
        RECT 3068.045 361.375 3068.325 361.655 ;
        RECT 3068.755 361.375 3069.035 361.655 ;
        RECT 3069.465 361.375 3069.745 361.655 ;
        RECT 3070.175 361.375 3070.455 361.655 ;
        RECT 3070.885 361.375 3071.165 361.655 ;
        RECT 3071.595 361.375 3071.875 361.655 ;
        RECT 3072.305 361.375 3072.585 361.655 ;
        RECT 3073.015 361.375 3073.295 361.655 ;
        RECT 3064.495 360.665 3064.775 360.945 ;
        RECT 3065.205 360.665 3065.485 360.945 ;
        RECT 3065.915 360.665 3066.195 360.945 ;
        RECT 3066.625 360.665 3066.905 360.945 ;
        RECT 3067.335 360.665 3067.615 360.945 ;
        RECT 3068.045 360.665 3068.325 360.945 ;
        RECT 3068.755 360.665 3069.035 360.945 ;
        RECT 3069.465 360.665 3069.745 360.945 ;
        RECT 3070.175 360.665 3070.455 360.945 ;
        RECT 3070.885 360.665 3071.165 360.945 ;
        RECT 3071.595 360.665 3071.875 360.945 ;
        RECT 3072.305 360.665 3072.585 360.945 ;
        RECT 3073.015 360.665 3073.295 360.945 ;
      LAYER Metal4 ;
        RECT 1896.360 4698.600 1900.080 4708.600 ;
        RECT 1908.760 4698.600 1919.010 4708.600 ;
        RECT 1920.610 4698.600 1930.860 4708.600 ;
        RECT 1934.140 4698.600 1944.390 4708.600 ;
        RECT 1945.990 4698.600 1956.240 4708.600 ;
        RECT 1959.140 4698.600 1968.640 4708.600 ;
        RECT 2996.360 4698.600 3005.860 4708.600 ;
        RECT 3008.760 4698.600 3019.010 4708.600 ;
        RECT 3025.100 4698.600 3030.860 4708.600 ;
        RECT 3034.140 4698.600 3044.390 4708.600 ;
        RECT 3045.990 4698.600 3056.240 4708.600 ;
        RECT 3059.140 4698.600 3068.640 4708.600 ;
        RECT 369.330 4392.970 369.610 4393.250 ;
        RECT 370.040 4392.970 370.320 4393.250 ;
        RECT 370.750 4392.970 371.030 4393.250 ;
        RECT 371.460 4392.970 371.740 4393.250 ;
        RECT 372.170 4392.970 372.450 4393.250 ;
        RECT 372.880 4392.970 373.160 4393.250 ;
        RECT 373.590 4392.970 373.870 4393.250 ;
        RECT 374.300 4392.970 374.580 4393.250 ;
        RECT 375.010 4392.970 375.290 4393.250 ;
        RECT 375.720 4392.970 376.000 4393.250 ;
        RECT 376.430 4392.970 376.710 4393.250 ;
        RECT 377.140 4392.970 377.420 4393.250 ;
        RECT 377.850 4392.970 378.130 4393.250 ;
        RECT 378.560 4392.970 378.840 4393.250 ;
        RECT 369.330 4392.260 369.610 4392.540 ;
        RECT 370.040 4392.260 370.320 4392.540 ;
        RECT 370.750 4392.260 371.030 4392.540 ;
        RECT 371.460 4392.260 371.740 4392.540 ;
        RECT 372.170 4392.260 372.450 4392.540 ;
        RECT 372.880 4392.260 373.160 4392.540 ;
        RECT 373.590 4392.260 373.870 4392.540 ;
        RECT 374.300 4392.260 374.580 4392.540 ;
        RECT 375.010 4392.260 375.290 4392.540 ;
        RECT 375.720 4392.260 376.000 4392.540 ;
        RECT 376.430 4392.260 376.710 4392.540 ;
        RECT 377.140 4392.260 377.420 4392.540 ;
        RECT 377.850 4392.260 378.130 4392.540 ;
        RECT 378.560 4392.260 378.840 4392.540 ;
        RECT 369.330 4391.550 369.610 4391.830 ;
        RECT 370.040 4391.550 370.320 4391.830 ;
        RECT 370.750 4391.550 371.030 4391.830 ;
        RECT 371.460 4391.550 371.740 4391.830 ;
        RECT 372.170 4391.550 372.450 4391.830 ;
        RECT 372.880 4391.550 373.160 4391.830 ;
        RECT 373.590 4391.550 373.870 4391.830 ;
        RECT 374.300 4391.550 374.580 4391.830 ;
        RECT 375.010 4391.550 375.290 4391.830 ;
        RECT 375.720 4391.550 376.000 4391.830 ;
        RECT 376.430 4391.550 376.710 4391.830 ;
        RECT 377.140 4391.550 377.420 4391.830 ;
        RECT 377.850 4391.550 378.130 4391.830 ;
        RECT 378.560 4391.550 378.840 4391.830 ;
        RECT 369.330 4390.840 369.610 4391.120 ;
        RECT 370.040 4390.840 370.320 4391.120 ;
        RECT 370.750 4390.840 371.030 4391.120 ;
        RECT 371.460 4390.840 371.740 4391.120 ;
        RECT 372.170 4390.840 372.450 4391.120 ;
        RECT 372.880 4390.840 373.160 4391.120 ;
        RECT 373.590 4390.840 373.870 4391.120 ;
        RECT 374.300 4390.840 374.580 4391.120 ;
        RECT 375.010 4390.840 375.290 4391.120 ;
        RECT 375.720 4390.840 376.000 4391.120 ;
        RECT 376.430 4390.840 376.710 4391.120 ;
        RECT 377.140 4390.840 377.420 4391.120 ;
        RECT 377.850 4390.840 378.130 4391.120 ;
        RECT 378.560 4390.840 378.840 4391.120 ;
        RECT 369.330 4390.130 369.610 4390.410 ;
        RECT 370.040 4390.130 370.320 4390.410 ;
        RECT 370.750 4390.130 371.030 4390.410 ;
        RECT 371.460 4390.130 371.740 4390.410 ;
        RECT 372.170 4390.130 372.450 4390.410 ;
        RECT 372.880 4390.130 373.160 4390.410 ;
        RECT 373.590 4390.130 373.870 4390.410 ;
        RECT 374.300 4390.130 374.580 4390.410 ;
        RECT 375.010 4390.130 375.290 4390.410 ;
        RECT 375.720 4390.130 376.000 4390.410 ;
        RECT 376.430 4390.130 376.710 4390.410 ;
        RECT 377.140 4390.130 377.420 4390.410 ;
        RECT 377.850 4390.130 378.130 4390.410 ;
        RECT 378.560 4390.130 378.840 4390.410 ;
        RECT 369.330 4389.420 369.610 4389.700 ;
        RECT 370.040 4389.420 370.320 4389.700 ;
        RECT 370.750 4389.420 371.030 4389.700 ;
        RECT 371.460 4389.420 371.740 4389.700 ;
        RECT 372.170 4389.420 372.450 4389.700 ;
        RECT 372.880 4389.420 373.160 4389.700 ;
        RECT 373.590 4389.420 373.870 4389.700 ;
        RECT 374.300 4389.420 374.580 4389.700 ;
        RECT 375.010 4389.420 375.290 4389.700 ;
        RECT 375.720 4389.420 376.000 4389.700 ;
        RECT 376.430 4389.420 376.710 4389.700 ;
        RECT 377.140 4389.420 377.420 4389.700 ;
        RECT 377.850 4389.420 378.130 4389.700 ;
        RECT 378.560 4389.420 378.840 4389.700 ;
        RECT 369.330 4388.710 369.610 4388.990 ;
        RECT 370.040 4388.710 370.320 4388.990 ;
        RECT 370.750 4388.710 371.030 4388.990 ;
        RECT 371.460 4388.710 371.740 4388.990 ;
        RECT 372.170 4388.710 372.450 4388.990 ;
        RECT 372.880 4388.710 373.160 4388.990 ;
        RECT 373.590 4388.710 373.870 4388.990 ;
        RECT 374.300 4388.710 374.580 4388.990 ;
        RECT 375.010 4388.710 375.290 4388.990 ;
        RECT 375.720 4388.710 376.000 4388.990 ;
        RECT 376.430 4388.710 376.710 4388.990 ;
        RECT 377.140 4388.710 377.420 4388.990 ;
        RECT 377.850 4388.710 378.130 4388.990 ;
        RECT 378.560 4388.710 378.840 4388.990 ;
        RECT 369.330 4388.000 369.610 4388.280 ;
        RECT 370.040 4388.000 370.320 4388.280 ;
        RECT 370.750 4388.000 371.030 4388.280 ;
        RECT 371.460 4388.000 371.740 4388.280 ;
        RECT 372.170 4388.000 372.450 4388.280 ;
        RECT 372.880 4388.000 373.160 4388.280 ;
        RECT 373.590 4388.000 373.870 4388.280 ;
        RECT 374.300 4388.000 374.580 4388.280 ;
        RECT 375.010 4388.000 375.290 4388.280 ;
        RECT 375.720 4388.000 376.000 4388.280 ;
        RECT 376.430 4388.000 376.710 4388.280 ;
        RECT 377.140 4388.000 377.420 4388.280 ;
        RECT 377.850 4388.000 378.130 4388.280 ;
        RECT 378.560 4388.000 378.840 4388.280 ;
        RECT 3500.200 4388.050 3500.480 4388.330 ;
        RECT 3500.910 4388.050 3501.190 4388.330 ;
        RECT 3501.620 4388.050 3501.900 4388.330 ;
        RECT 3502.330 4388.050 3502.610 4388.330 ;
        RECT 3503.040 4388.050 3503.320 4388.330 ;
        RECT 3503.750 4388.050 3504.030 4388.330 ;
        RECT 3504.460 4388.050 3504.740 4388.330 ;
        RECT 3505.170 4388.050 3505.450 4388.330 ;
        RECT 3505.880 4388.050 3506.160 4388.330 ;
        RECT 3506.590 4388.050 3506.870 4388.330 ;
        RECT 3507.300 4388.050 3507.580 4388.330 ;
        RECT 3508.010 4388.050 3508.290 4388.330 ;
        RECT 3508.720 4388.050 3509.000 4388.330 ;
        RECT 3509.430 4388.050 3509.710 4388.330 ;
        RECT 369.330 4387.290 369.610 4387.570 ;
        RECT 370.040 4387.290 370.320 4387.570 ;
        RECT 370.750 4387.290 371.030 4387.570 ;
        RECT 371.460 4387.290 371.740 4387.570 ;
        RECT 372.170 4387.290 372.450 4387.570 ;
        RECT 372.880 4387.290 373.160 4387.570 ;
        RECT 373.590 4387.290 373.870 4387.570 ;
        RECT 374.300 4387.290 374.580 4387.570 ;
        RECT 375.010 4387.290 375.290 4387.570 ;
        RECT 375.720 4387.290 376.000 4387.570 ;
        RECT 376.430 4387.290 376.710 4387.570 ;
        RECT 377.140 4387.290 377.420 4387.570 ;
        RECT 377.850 4387.290 378.130 4387.570 ;
        RECT 378.560 4387.290 378.840 4387.570 ;
        RECT 3500.200 4387.340 3500.480 4387.620 ;
        RECT 3500.910 4387.340 3501.190 4387.620 ;
        RECT 3501.620 4387.340 3501.900 4387.620 ;
        RECT 3502.330 4387.340 3502.610 4387.620 ;
        RECT 3503.040 4387.340 3503.320 4387.620 ;
        RECT 3503.750 4387.340 3504.030 4387.620 ;
        RECT 3504.460 4387.340 3504.740 4387.620 ;
        RECT 3505.170 4387.340 3505.450 4387.620 ;
        RECT 3505.880 4387.340 3506.160 4387.620 ;
        RECT 3506.590 4387.340 3506.870 4387.620 ;
        RECT 3507.300 4387.340 3507.580 4387.620 ;
        RECT 3508.010 4387.340 3508.290 4387.620 ;
        RECT 3508.720 4387.340 3509.000 4387.620 ;
        RECT 3509.430 4387.340 3509.710 4387.620 ;
        RECT 369.330 4386.580 369.610 4386.860 ;
        RECT 370.040 4386.580 370.320 4386.860 ;
        RECT 370.750 4386.580 371.030 4386.860 ;
        RECT 371.460 4386.580 371.740 4386.860 ;
        RECT 372.170 4386.580 372.450 4386.860 ;
        RECT 372.880 4386.580 373.160 4386.860 ;
        RECT 373.590 4386.580 373.870 4386.860 ;
        RECT 374.300 4386.580 374.580 4386.860 ;
        RECT 375.010 4386.580 375.290 4386.860 ;
        RECT 375.720 4386.580 376.000 4386.860 ;
        RECT 376.430 4386.580 376.710 4386.860 ;
        RECT 377.140 4386.580 377.420 4386.860 ;
        RECT 377.850 4386.580 378.130 4386.860 ;
        RECT 378.560 4386.580 378.840 4386.860 ;
        RECT 3500.200 4386.630 3500.480 4386.910 ;
        RECT 3500.910 4386.630 3501.190 4386.910 ;
        RECT 3501.620 4386.630 3501.900 4386.910 ;
        RECT 3502.330 4386.630 3502.610 4386.910 ;
        RECT 3503.040 4386.630 3503.320 4386.910 ;
        RECT 3503.750 4386.630 3504.030 4386.910 ;
        RECT 3504.460 4386.630 3504.740 4386.910 ;
        RECT 3505.170 4386.630 3505.450 4386.910 ;
        RECT 3505.880 4386.630 3506.160 4386.910 ;
        RECT 3506.590 4386.630 3506.870 4386.910 ;
        RECT 3507.300 4386.630 3507.580 4386.910 ;
        RECT 3508.010 4386.630 3508.290 4386.910 ;
        RECT 3508.720 4386.630 3509.000 4386.910 ;
        RECT 3509.430 4386.630 3509.710 4386.910 ;
        RECT 369.330 4385.870 369.610 4386.150 ;
        RECT 370.040 4385.870 370.320 4386.150 ;
        RECT 370.750 4385.870 371.030 4386.150 ;
        RECT 371.460 4385.870 371.740 4386.150 ;
        RECT 372.170 4385.870 372.450 4386.150 ;
        RECT 372.880 4385.870 373.160 4386.150 ;
        RECT 373.590 4385.870 373.870 4386.150 ;
        RECT 374.300 4385.870 374.580 4386.150 ;
        RECT 375.010 4385.870 375.290 4386.150 ;
        RECT 375.720 4385.870 376.000 4386.150 ;
        RECT 376.430 4385.870 376.710 4386.150 ;
        RECT 377.140 4385.870 377.420 4386.150 ;
        RECT 377.850 4385.870 378.130 4386.150 ;
        RECT 378.560 4385.870 378.840 4386.150 ;
        RECT 3500.200 4385.920 3500.480 4386.200 ;
        RECT 3500.910 4385.920 3501.190 4386.200 ;
        RECT 3501.620 4385.920 3501.900 4386.200 ;
        RECT 3502.330 4385.920 3502.610 4386.200 ;
        RECT 3503.040 4385.920 3503.320 4386.200 ;
        RECT 3503.750 4385.920 3504.030 4386.200 ;
        RECT 3504.460 4385.920 3504.740 4386.200 ;
        RECT 3505.170 4385.920 3505.450 4386.200 ;
        RECT 3505.880 4385.920 3506.160 4386.200 ;
        RECT 3506.590 4385.920 3506.870 4386.200 ;
        RECT 3507.300 4385.920 3507.580 4386.200 ;
        RECT 3508.010 4385.920 3508.290 4386.200 ;
        RECT 3508.720 4385.920 3509.000 4386.200 ;
        RECT 3509.430 4385.920 3509.710 4386.200 ;
        RECT 369.330 4385.160 369.610 4385.440 ;
        RECT 370.040 4385.160 370.320 4385.440 ;
        RECT 370.750 4385.160 371.030 4385.440 ;
        RECT 371.460 4385.160 371.740 4385.440 ;
        RECT 372.170 4385.160 372.450 4385.440 ;
        RECT 372.880 4385.160 373.160 4385.440 ;
        RECT 373.590 4385.160 373.870 4385.440 ;
        RECT 374.300 4385.160 374.580 4385.440 ;
        RECT 375.010 4385.160 375.290 4385.440 ;
        RECT 375.720 4385.160 376.000 4385.440 ;
        RECT 376.430 4385.160 376.710 4385.440 ;
        RECT 377.140 4385.160 377.420 4385.440 ;
        RECT 377.850 4385.160 378.130 4385.440 ;
        RECT 378.560 4385.160 378.840 4385.440 ;
        RECT 3500.200 4385.210 3500.480 4385.490 ;
        RECT 3500.910 4385.210 3501.190 4385.490 ;
        RECT 3501.620 4385.210 3501.900 4385.490 ;
        RECT 3502.330 4385.210 3502.610 4385.490 ;
        RECT 3503.040 4385.210 3503.320 4385.490 ;
        RECT 3503.750 4385.210 3504.030 4385.490 ;
        RECT 3504.460 4385.210 3504.740 4385.490 ;
        RECT 3505.170 4385.210 3505.450 4385.490 ;
        RECT 3505.880 4385.210 3506.160 4385.490 ;
        RECT 3506.590 4385.210 3506.870 4385.490 ;
        RECT 3507.300 4385.210 3507.580 4385.490 ;
        RECT 3508.010 4385.210 3508.290 4385.490 ;
        RECT 3508.720 4385.210 3509.000 4385.490 ;
        RECT 3509.430 4385.210 3509.710 4385.490 ;
        RECT 369.330 4384.450 369.610 4384.730 ;
        RECT 370.040 4384.450 370.320 4384.730 ;
        RECT 370.750 4384.450 371.030 4384.730 ;
        RECT 371.460 4384.450 371.740 4384.730 ;
        RECT 372.170 4384.450 372.450 4384.730 ;
        RECT 372.880 4384.450 373.160 4384.730 ;
        RECT 373.590 4384.450 373.870 4384.730 ;
        RECT 374.300 4384.450 374.580 4384.730 ;
        RECT 375.010 4384.450 375.290 4384.730 ;
        RECT 375.720 4384.450 376.000 4384.730 ;
        RECT 376.430 4384.450 376.710 4384.730 ;
        RECT 377.140 4384.450 377.420 4384.730 ;
        RECT 377.850 4384.450 378.130 4384.730 ;
        RECT 378.560 4384.450 378.840 4384.730 ;
        RECT 3500.200 4384.500 3500.480 4384.780 ;
        RECT 3500.910 4384.500 3501.190 4384.780 ;
        RECT 3501.620 4384.500 3501.900 4384.780 ;
        RECT 3502.330 4384.500 3502.610 4384.780 ;
        RECT 3503.040 4384.500 3503.320 4384.780 ;
        RECT 3503.750 4384.500 3504.030 4384.780 ;
        RECT 3504.460 4384.500 3504.740 4384.780 ;
        RECT 3505.170 4384.500 3505.450 4384.780 ;
        RECT 3505.880 4384.500 3506.160 4384.780 ;
        RECT 3506.590 4384.500 3506.870 4384.780 ;
        RECT 3507.300 4384.500 3507.580 4384.780 ;
        RECT 3508.010 4384.500 3508.290 4384.780 ;
        RECT 3508.720 4384.500 3509.000 4384.780 ;
        RECT 3509.430 4384.500 3509.710 4384.780 ;
        RECT 3500.200 4383.790 3500.480 4384.070 ;
        RECT 3500.910 4383.790 3501.190 4384.070 ;
        RECT 3501.620 4383.790 3501.900 4384.070 ;
        RECT 3502.330 4383.790 3502.610 4384.070 ;
        RECT 3503.040 4383.790 3503.320 4384.070 ;
        RECT 3503.750 4383.790 3504.030 4384.070 ;
        RECT 3504.460 4383.790 3504.740 4384.070 ;
        RECT 3505.170 4383.790 3505.450 4384.070 ;
        RECT 3505.880 4383.790 3506.160 4384.070 ;
        RECT 3506.590 4383.790 3506.870 4384.070 ;
        RECT 3507.300 4383.790 3507.580 4384.070 ;
        RECT 3508.010 4383.790 3508.290 4384.070 ;
        RECT 3508.720 4383.790 3509.000 4384.070 ;
        RECT 3509.430 4383.790 3509.710 4384.070 ;
        RECT 3500.200 4383.080 3500.480 4383.360 ;
        RECT 3500.910 4383.080 3501.190 4383.360 ;
        RECT 3501.620 4383.080 3501.900 4383.360 ;
        RECT 3502.330 4383.080 3502.610 4383.360 ;
        RECT 3503.040 4383.080 3503.320 4383.360 ;
        RECT 3503.750 4383.080 3504.030 4383.360 ;
        RECT 3504.460 4383.080 3504.740 4383.360 ;
        RECT 3505.170 4383.080 3505.450 4383.360 ;
        RECT 3505.880 4383.080 3506.160 4383.360 ;
        RECT 3506.590 4383.080 3506.870 4383.360 ;
        RECT 3507.300 4383.080 3507.580 4383.360 ;
        RECT 3508.010 4383.080 3508.290 4383.360 ;
        RECT 3508.720 4383.080 3509.000 4383.360 ;
        RECT 3509.430 4383.080 3509.710 4383.360 ;
        RECT 3500.200 4382.370 3500.480 4382.650 ;
        RECT 3500.910 4382.370 3501.190 4382.650 ;
        RECT 3501.620 4382.370 3501.900 4382.650 ;
        RECT 3502.330 4382.370 3502.610 4382.650 ;
        RECT 3503.040 4382.370 3503.320 4382.650 ;
        RECT 3503.750 4382.370 3504.030 4382.650 ;
        RECT 3504.460 4382.370 3504.740 4382.650 ;
        RECT 3505.170 4382.370 3505.450 4382.650 ;
        RECT 3505.880 4382.370 3506.160 4382.650 ;
        RECT 3506.590 4382.370 3506.870 4382.650 ;
        RECT 3507.300 4382.370 3507.580 4382.650 ;
        RECT 3508.010 4382.370 3508.290 4382.650 ;
        RECT 3508.720 4382.370 3509.000 4382.650 ;
        RECT 3509.430 4382.370 3509.710 4382.650 ;
        RECT 3500.200 4381.660 3500.480 4381.940 ;
        RECT 3500.910 4381.660 3501.190 4381.940 ;
        RECT 3501.620 4381.660 3501.900 4381.940 ;
        RECT 3502.330 4381.660 3502.610 4381.940 ;
        RECT 3503.040 4381.660 3503.320 4381.940 ;
        RECT 3503.750 4381.660 3504.030 4381.940 ;
        RECT 3504.460 4381.660 3504.740 4381.940 ;
        RECT 3505.170 4381.660 3505.450 4381.940 ;
        RECT 3505.880 4381.660 3506.160 4381.940 ;
        RECT 3506.590 4381.660 3506.870 4381.940 ;
        RECT 3507.300 4381.660 3507.580 4381.940 ;
        RECT 3508.010 4381.660 3508.290 4381.940 ;
        RECT 3508.720 4381.660 3509.000 4381.940 ;
        RECT 3509.430 4381.660 3509.710 4381.940 ;
        RECT 3500.200 4380.950 3500.480 4381.230 ;
        RECT 3500.910 4380.950 3501.190 4381.230 ;
        RECT 3501.620 4380.950 3501.900 4381.230 ;
        RECT 3502.330 4380.950 3502.610 4381.230 ;
        RECT 3503.040 4380.950 3503.320 4381.230 ;
        RECT 3503.750 4380.950 3504.030 4381.230 ;
        RECT 3504.460 4380.950 3504.740 4381.230 ;
        RECT 3505.170 4380.950 3505.450 4381.230 ;
        RECT 3505.880 4380.950 3506.160 4381.230 ;
        RECT 3506.590 4380.950 3506.870 4381.230 ;
        RECT 3507.300 4380.950 3507.580 4381.230 ;
        RECT 3508.010 4380.950 3508.290 4381.230 ;
        RECT 3508.720 4380.950 3509.000 4381.230 ;
        RECT 3509.430 4380.950 3509.710 4381.230 ;
        RECT 369.275 4380.565 369.555 4380.845 ;
        RECT 369.985 4380.565 370.265 4380.845 ;
        RECT 370.695 4380.565 370.975 4380.845 ;
        RECT 371.405 4380.565 371.685 4380.845 ;
        RECT 372.115 4380.565 372.395 4380.845 ;
        RECT 372.825 4380.565 373.105 4380.845 ;
        RECT 373.535 4380.565 373.815 4380.845 ;
        RECT 374.245 4380.565 374.525 4380.845 ;
        RECT 374.955 4380.565 375.235 4380.845 ;
        RECT 375.665 4380.565 375.945 4380.845 ;
        RECT 376.375 4380.565 376.655 4380.845 ;
        RECT 377.085 4380.565 377.365 4380.845 ;
        RECT 377.795 4380.565 378.075 4380.845 ;
        RECT 378.505 4380.565 378.785 4380.845 ;
        RECT 3500.200 4380.240 3500.480 4380.520 ;
        RECT 3500.910 4380.240 3501.190 4380.520 ;
        RECT 3501.620 4380.240 3501.900 4380.520 ;
        RECT 3502.330 4380.240 3502.610 4380.520 ;
        RECT 3503.040 4380.240 3503.320 4380.520 ;
        RECT 3503.750 4380.240 3504.030 4380.520 ;
        RECT 3504.460 4380.240 3504.740 4380.520 ;
        RECT 3505.170 4380.240 3505.450 4380.520 ;
        RECT 3505.880 4380.240 3506.160 4380.520 ;
        RECT 3506.590 4380.240 3506.870 4380.520 ;
        RECT 3507.300 4380.240 3507.580 4380.520 ;
        RECT 3508.010 4380.240 3508.290 4380.520 ;
        RECT 3508.720 4380.240 3509.000 4380.520 ;
        RECT 3509.430 4380.240 3509.710 4380.520 ;
        RECT 369.275 4379.855 369.555 4380.135 ;
        RECT 369.985 4379.855 370.265 4380.135 ;
        RECT 370.695 4379.855 370.975 4380.135 ;
        RECT 371.405 4379.855 371.685 4380.135 ;
        RECT 372.115 4379.855 372.395 4380.135 ;
        RECT 372.825 4379.855 373.105 4380.135 ;
        RECT 373.535 4379.855 373.815 4380.135 ;
        RECT 374.245 4379.855 374.525 4380.135 ;
        RECT 374.955 4379.855 375.235 4380.135 ;
        RECT 375.665 4379.855 375.945 4380.135 ;
        RECT 376.375 4379.855 376.655 4380.135 ;
        RECT 377.085 4379.855 377.365 4380.135 ;
        RECT 377.795 4379.855 378.075 4380.135 ;
        RECT 378.505 4379.855 378.785 4380.135 ;
        RECT 3500.200 4379.530 3500.480 4379.810 ;
        RECT 3500.910 4379.530 3501.190 4379.810 ;
        RECT 3501.620 4379.530 3501.900 4379.810 ;
        RECT 3502.330 4379.530 3502.610 4379.810 ;
        RECT 3503.040 4379.530 3503.320 4379.810 ;
        RECT 3503.750 4379.530 3504.030 4379.810 ;
        RECT 3504.460 4379.530 3504.740 4379.810 ;
        RECT 3505.170 4379.530 3505.450 4379.810 ;
        RECT 3505.880 4379.530 3506.160 4379.810 ;
        RECT 3506.590 4379.530 3506.870 4379.810 ;
        RECT 3507.300 4379.530 3507.580 4379.810 ;
        RECT 3508.010 4379.530 3508.290 4379.810 ;
        RECT 3508.720 4379.530 3509.000 4379.810 ;
        RECT 3509.430 4379.530 3509.710 4379.810 ;
        RECT 369.275 4379.145 369.555 4379.425 ;
        RECT 369.985 4379.145 370.265 4379.425 ;
        RECT 370.695 4379.145 370.975 4379.425 ;
        RECT 371.405 4379.145 371.685 4379.425 ;
        RECT 372.115 4379.145 372.395 4379.425 ;
        RECT 372.825 4379.145 373.105 4379.425 ;
        RECT 373.535 4379.145 373.815 4379.425 ;
        RECT 374.245 4379.145 374.525 4379.425 ;
        RECT 374.955 4379.145 375.235 4379.425 ;
        RECT 375.665 4379.145 375.945 4379.425 ;
        RECT 376.375 4379.145 376.655 4379.425 ;
        RECT 377.085 4379.145 377.365 4379.425 ;
        RECT 377.795 4379.145 378.075 4379.425 ;
        RECT 378.505 4379.145 378.785 4379.425 ;
        RECT 369.275 4378.435 369.555 4378.715 ;
        RECT 369.985 4378.435 370.265 4378.715 ;
        RECT 370.695 4378.435 370.975 4378.715 ;
        RECT 371.405 4378.435 371.685 4378.715 ;
        RECT 372.115 4378.435 372.395 4378.715 ;
        RECT 372.825 4378.435 373.105 4378.715 ;
        RECT 373.535 4378.435 373.815 4378.715 ;
        RECT 374.245 4378.435 374.525 4378.715 ;
        RECT 374.955 4378.435 375.235 4378.715 ;
        RECT 375.665 4378.435 375.945 4378.715 ;
        RECT 376.375 4378.435 376.655 4378.715 ;
        RECT 377.085 4378.435 377.365 4378.715 ;
        RECT 377.795 4378.435 378.075 4378.715 ;
        RECT 378.505 4378.435 378.785 4378.715 ;
        RECT 369.275 4377.725 369.555 4378.005 ;
        RECT 369.985 4377.725 370.265 4378.005 ;
        RECT 370.695 4377.725 370.975 4378.005 ;
        RECT 371.405 4377.725 371.685 4378.005 ;
        RECT 372.115 4377.725 372.395 4378.005 ;
        RECT 372.825 4377.725 373.105 4378.005 ;
        RECT 373.535 4377.725 373.815 4378.005 ;
        RECT 374.245 4377.725 374.525 4378.005 ;
        RECT 374.955 4377.725 375.235 4378.005 ;
        RECT 375.665 4377.725 375.945 4378.005 ;
        RECT 376.375 4377.725 376.655 4378.005 ;
        RECT 377.085 4377.725 377.365 4378.005 ;
        RECT 377.795 4377.725 378.075 4378.005 ;
        RECT 378.505 4377.725 378.785 4378.005 ;
        RECT 369.275 4377.015 369.555 4377.295 ;
        RECT 369.985 4377.015 370.265 4377.295 ;
        RECT 370.695 4377.015 370.975 4377.295 ;
        RECT 371.405 4377.015 371.685 4377.295 ;
        RECT 372.115 4377.015 372.395 4377.295 ;
        RECT 372.825 4377.015 373.105 4377.295 ;
        RECT 373.535 4377.015 373.815 4377.295 ;
        RECT 374.245 4377.015 374.525 4377.295 ;
        RECT 374.955 4377.015 375.235 4377.295 ;
        RECT 375.665 4377.015 375.945 4377.295 ;
        RECT 376.375 4377.015 376.655 4377.295 ;
        RECT 377.085 4377.015 377.365 4377.295 ;
        RECT 377.795 4377.015 378.075 4377.295 ;
        RECT 378.505 4377.015 378.785 4377.295 ;
        RECT 369.275 4376.305 369.555 4376.585 ;
        RECT 369.985 4376.305 370.265 4376.585 ;
        RECT 370.695 4376.305 370.975 4376.585 ;
        RECT 371.405 4376.305 371.685 4376.585 ;
        RECT 372.115 4376.305 372.395 4376.585 ;
        RECT 372.825 4376.305 373.105 4376.585 ;
        RECT 373.535 4376.305 373.815 4376.585 ;
        RECT 374.245 4376.305 374.525 4376.585 ;
        RECT 374.955 4376.305 375.235 4376.585 ;
        RECT 375.665 4376.305 375.945 4376.585 ;
        RECT 376.375 4376.305 376.655 4376.585 ;
        RECT 377.085 4376.305 377.365 4376.585 ;
        RECT 377.795 4376.305 378.075 4376.585 ;
        RECT 378.505 4376.305 378.785 4376.585 ;
        RECT 369.275 4375.595 369.555 4375.875 ;
        RECT 369.985 4375.595 370.265 4375.875 ;
        RECT 370.695 4375.595 370.975 4375.875 ;
        RECT 371.405 4375.595 371.685 4375.875 ;
        RECT 372.115 4375.595 372.395 4375.875 ;
        RECT 372.825 4375.595 373.105 4375.875 ;
        RECT 373.535 4375.595 373.815 4375.875 ;
        RECT 374.245 4375.595 374.525 4375.875 ;
        RECT 374.955 4375.595 375.235 4375.875 ;
        RECT 375.665 4375.595 375.945 4375.875 ;
        RECT 376.375 4375.595 376.655 4375.875 ;
        RECT 377.085 4375.595 377.365 4375.875 ;
        RECT 377.795 4375.595 378.075 4375.875 ;
        RECT 378.505 4375.595 378.785 4375.875 ;
        RECT 3500.255 4375.615 3500.535 4375.895 ;
        RECT 3500.965 4375.615 3501.245 4375.895 ;
        RECT 3501.675 4375.615 3501.955 4375.895 ;
        RECT 3502.385 4375.615 3502.665 4375.895 ;
        RECT 3503.095 4375.615 3503.375 4375.895 ;
        RECT 3503.805 4375.615 3504.085 4375.895 ;
        RECT 3504.515 4375.615 3504.795 4375.895 ;
        RECT 3505.225 4375.615 3505.505 4375.895 ;
        RECT 3505.935 4375.615 3506.215 4375.895 ;
        RECT 3506.645 4375.615 3506.925 4375.895 ;
        RECT 3507.355 4375.615 3507.635 4375.895 ;
        RECT 3508.065 4375.615 3508.345 4375.895 ;
        RECT 3508.775 4375.615 3509.055 4375.895 ;
        RECT 3509.485 4375.615 3509.765 4375.895 ;
        RECT 369.275 4374.885 369.555 4375.165 ;
        RECT 369.985 4374.885 370.265 4375.165 ;
        RECT 370.695 4374.885 370.975 4375.165 ;
        RECT 371.405 4374.885 371.685 4375.165 ;
        RECT 372.115 4374.885 372.395 4375.165 ;
        RECT 372.825 4374.885 373.105 4375.165 ;
        RECT 373.535 4374.885 373.815 4375.165 ;
        RECT 374.245 4374.885 374.525 4375.165 ;
        RECT 374.955 4374.885 375.235 4375.165 ;
        RECT 375.665 4374.885 375.945 4375.165 ;
        RECT 376.375 4374.885 376.655 4375.165 ;
        RECT 377.085 4374.885 377.365 4375.165 ;
        RECT 377.795 4374.885 378.075 4375.165 ;
        RECT 378.505 4374.885 378.785 4375.165 ;
        RECT 3500.255 4374.905 3500.535 4375.185 ;
        RECT 3500.965 4374.905 3501.245 4375.185 ;
        RECT 3501.675 4374.905 3501.955 4375.185 ;
        RECT 3502.385 4374.905 3502.665 4375.185 ;
        RECT 3503.095 4374.905 3503.375 4375.185 ;
        RECT 3503.805 4374.905 3504.085 4375.185 ;
        RECT 3504.515 4374.905 3504.795 4375.185 ;
        RECT 3505.225 4374.905 3505.505 4375.185 ;
        RECT 3505.935 4374.905 3506.215 4375.185 ;
        RECT 3506.645 4374.905 3506.925 4375.185 ;
        RECT 3507.355 4374.905 3507.635 4375.185 ;
        RECT 3508.065 4374.905 3508.345 4375.185 ;
        RECT 3508.775 4374.905 3509.055 4375.185 ;
        RECT 3509.485 4374.905 3509.765 4375.185 ;
        RECT 369.275 4374.175 369.555 4374.455 ;
        RECT 369.985 4374.175 370.265 4374.455 ;
        RECT 370.695 4374.175 370.975 4374.455 ;
        RECT 371.405 4374.175 371.685 4374.455 ;
        RECT 372.115 4374.175 372.395 4374.455 ;
        RECT 372.825 4374.175 373.105 4374.455 ;
        RECT 373.535 4374.175 373.815 4374.455 ;
        RECT 374.245 4374.175 374.525 4374.455 ;
        RECT 374.955 4374.175 375.235 4374.455 ;
        RECT 375.665 4374.175 375.945 4374.455 ;
        RECT 376.375 4374.175 376.655 4374.455 ;
        RECT 377.085 4374.175 377.365 4374.455 ;
        RECT 377.795 4374.175 378.075 4374.455 ;
        RECT 378.505 4374.175 378.785 4374.455 ;
        RECT 3500.255 4374.195 3500.535 4374.475 ;
        RECT 3500.965 4374.195 3501.245 4374.475 ;
        RECT 3501.675 4374.195 3501.955 4374.475 ;
        RECT 3502.385 4374.195 3502.665 4374.475 ;
        RECT 3503.095 4374.195 3503.375 4374.475 ;
        RECT 3503.805 4374.195 3504.085 4374.475 ;
        RECT 3504.515 4374.195 3504.795 4374.475 ;
        RECT 3505.225 4374.195 3505.505 4374.475 ;
        RECT 3505.935 4374.195 3506.215 4374.475 ;
        RECT 3506.645 4374.195 3506.925 4374.475 ;
        RECT 3507.355 4374.195 3507.635 4374.475 ;
        RECT 3508.065 4374.195 3508.345 4374.475 ;
        RECT 3508.775 4374.195 3509.055 4374.475 ;
        RECT 3509.485 4374.195 3509.765 4374.475 ;
        RECT 369.275 4373.465 369.555 4373.745 ;
        RECT 369.985 4373.465 370.265 4373.745 ;
        RECT 370.695 4373.465 370.975 4373.745 ;
        RECT 371.405 4373.465 371.685 4373.745 ;
        RECT 372.115 4373.465 372.395 4373.745 ;
        RECT 372.825 4373.465 373.105 4373.745 ;
        RECT 373.535 4373.465 373.815 4373.745 ;
        RECT 374.245 4373.465 374.525 4373.745 ;
        RECT 374.955 4373.465 375.235 4373.745 ;
        RECT 375.665 4373.465 375.945 4373.745 ;
        RECT 376.375 4373.465 376.655 4373.745 ;
        RECT 377.085 4373.465 377.365 4373.745 ;
        RECT 377.795 4373.465 378.075 4373.745 ;
        RECT 378.505 4373.465 378.785 4373.745 ;
        RECT 3500.255 4373.485 3500.535 4373.765 ;
        RECT 3500.965 4373.485 3501.245 4373.765 ;
        RECT 3501.675 4373.485 3501.955 4373.765 ;
        RECT 3502.385 4373.485 3502.665 4373.765 ;
        RECT 3503.095 4373.485 3503.375 4373.765 ;
        RECT 3503.805 4373.485 3504.085 4373.765 ;
        RECT 3504.515 4373.485 3504.795 4373.765 ;
        RECT 3505.225 4373.485 3505.505 4373.765 ;
        RECT 3505.935 4373.485 3506.215 4373.765 ;
        RECT 3506.645 4373.485 3506.925 4373.765 ;
        RECT 3507.355 4373.485 3507.635 4373.765 ;
        RECT 3508.065 4373.485 3508.345 4373.765 ;
        RECT 3508.775 4373.485 3509.055 4373.765 ;
        RECT 3509.485 4373.485 3509.765 4373.765 ;
        RECT 369.275 4372.755 369.555 4373.035 ;
        RECT 369.985 4372.755 370.265 4373.035 ;
        RECT 370.695 4372.755 370.975 4373.035 ;
        RECT 371.405 4372.755 371.685 4373.035 ;
        RECT 372.115 4372.755 372.395 4373.035 ;
        RECT 372.825 4372.755 373.105 4373.035 ;
        RECT 373.535 4372.755 373.815 4373.035 ;
        RECT 374.245 4372.755 374.525 4373.035 ;
        RECT 374.955 4372.755 375.235 4373.035 ;
        RECT 375.665 4372.755 375.945 4373.035 ;
        RECT 376.375 4372.755 376.655 4373.035 ;
        RECT 377.085 4372.755 377.365 4373.035 ;
        RECT 377.795 4372.755 378.075 4373.035 ;
        RECT 378.505 4372.755 378.785 4373.035 ;
        RECT 3500.255 4372.775 3500.535 4373.055 ;
        RECT 3500.965 4372.775 3501.245 4373.055 ;
        RECT 3501.675 4372.775 3501.955 4373.055 ;
        RECT 3502.385 4372.775 3502.665 4373.055 ;
        RECT 3503.095 4372.775 3503.375 4373.055 ;
        RECT 3503.805 4372.775 3504.085 4373.055 ;
        RECT 3504.515 4372.775 3504.795 4373.055 ;
        RECT 3505.225 4372.775 3505.505 4373.055 ;
        RECT 3505.935 4372.775 3506.215 4373.055 ;
        RECT 3506.645 4372.775 3506.925 4373.055 ;
        RECT 3507.355 4372.775 3507.635 4373.055 ;
        RECT 3508.065 4372.775 3508.345 4373.055 ;
        RECT 3508.775 4372.775 3509.055 4373.055 ;
        RECT 3509.485 4372.775 3509.765 4373.055 ;
        RECT 369.275 4372.045 369.555 4372.325 ;
        RECT 369.985 4372.045 370.265 4372.325 ;
        RECT 370.695 4372.045 370.975 4372.325 ;
        RECT 371.405 4372.045 371.685 4372.325 ;
        RECT 372.115 4372.045 372.395 4372.325 ;
        RECT 372.825 4372.045 373.105 4372.325 ;
        RECT 373.535 4372.045 373.815 4372.325 ;
        RECT 374.245 4372.045 374.525 4372.325 ;
        RECT 374.955 4372.045 375.235 4372.325 ;
        RECT 375.665 4372.045 375.945 4372.325 ;
        RECT 376.375 4372.045 376.655 4372.325 ;
        RECT 377.085 4372.045 377.365 4372.325 ;
        RECT 377.795 4372.045 378.075 4372.325 ;
        RECT 378.505 4372.045 378.785 4372.325 ;
        RECT 3500.255 4372.065 3500.535 4372.345 ;
        RECT 3500.965 4372.065 3501.245 4372.345 ;
        RECT 3501.675 4372.065 3501.955 4372.345 ;
        RECT 3502.385 4372.065 3502.665 4372.345 ;
        RECT 3503.095 4372.065 3503.375 4372.345 ;
        RECT 3503.805 4372.065 3504.085 4372.345 ;
        RECT 3504.515 4372.065 3504.795 4372.345 ;
        RECT 3505.225 4372.065 3505.505 4372.345 ;
        RECT 3505.935 4372.065 3506.215 4372.345 ;
        RECT 3506.645 4372.065 3506.925 4372.345 ;
        RECT 3507.355 4372.065 3507.635 4372.345 ;
        RECT 3508.065 4372.065 3508.345 4372.345 ;
        RECT 3508.775 4372.065 3509.055 4372.345 ;
        RECT 3509.485 4372.065 3509.765 4372.345 ;
        RECT 369.275 4371.335 369.555 4371.615 ;
        RECT 369.985 4371.335 370.265 4371.615 ;
        RECT 370.695 4371.335 370.975 4371.615 ;
        RECT 371.405 4371.335 371.685 4371.615 ;
        RECT 372.115 4371.335 372.395 4371.615 ;
        RECT 372.825 4371.335 373.105 4371.615 ;
        RECT 373.535 4371.335 373.815 4371.615 ;
        RECT 374.245 4371.335 374.525 4371.615 ;
        RECT 374.955 4371.335 375.235 4371.615 ;
        RECT 375.665 4371.335 375.945 4371.615 ;
        RECT 376.375 4371.335 376.655 4371.615 ;
        RECT 377.085 4371.335 377.365 4371.615 ;
        RECT 377.795 4371.335 378.075 4371.615 ;
        RECT 378.505 4371.335 378.785 4371.615 ;
        RECT 3500.255 4371.355 3500.535 4371.635 ;
        RECT 3500.965 4371.355 3501.245 4371.635 ;
        RECT 3501.675 4371.355 3501.955 4371.635 ;
        RECT 3502.385 4371.355 3502.665 4371.635 ;
        RECT 3503.095 4371.355 3503.375 4371.635 ;
        RECT 3503.805 4371.355 3504.085 4371.635 ;
        RECT 3504.515 4371.355 3504.795 4371.635 ;
        RECT 3505.225 4371.355 3505.505 4371.635 ;
        RECT 3505.935 4371.355 3506.215 4371.635 ;
        RECT 3506.645 4371.355 3506.925 4371.635 ;
        RECT 3507.355 4371.355 3507.635 4371.635 ;
        RECT 3508.065 4371.355 3508.345 4371.635 ;
        RECT 3508.775 4371.355 3509.055 4371.635 ;
        RECT 3509.485 4371.355 3509.765 4371.635 ;
        RECT 3500.255 4370.645 3500.535 4370.925 ;
        RECT 3500.965 4370.645 3501.245 4370.925 ;
        RECT 3501.675 4370.645 3501.955 4370.925 ;
        RECT 3502.385 4370.645 3502.665 4370.925 ;
        RECT 3503.095 4370.645 3503.375 4370.925 ;
        RECT 3503.805 4370.645 3504.085 4370.925 ;
        RECT 3504.515 4370.645 3504.795 4370.925 ;
        RECT 3505.225 4370.645 3505.505 4370.925 ;
        RECT 3505.935 4370.645 3506.215 4370.925 ;
        RECT 3506.645 4370.645 3506.925 4370.925 ;
        RECT 3507.355 4370.645 3507.635 4370.925 ;
        RECT 3508.065 4370.645 3508.345 4370.925 ;
        RECT 3508.775 4370.645 3509.055 4370.925 ;
        RECT 3509.485 4370.645 3509.765 4370.925 ;
        RECT 3500.255 4369.935 3500.535 4370.215 ;
        RECT 3500.965 4369.935 3501.245 4370.215 ;
        RECT 3501.675 4369.935 3501.955 4370.215 ;
        RECT 3502.385 4369.935 3502.665 4370.215 ;
        RECT 3503.095 4369.935 3503.375 4370.215 ;
        RECT 3503.805 4369.935 3504.085 4370.215 ;
        RECT 3504.515 4369.935 3504.795 4370.215 ;
        RECT 3505.225 4369.935 3505.505 4370.215 ;
        RECT 3505.935 4369.935 3506.215 4370.215 ;
        RECT 3506.645 4369.935 3506.925 4370.215 ;
        RECT 3507.355 4369.935 3507.635 4370.215 ;
        RECT 3508.065 4369.935 3508.345 4370.215 ;
        RECT 3508.775 4369.935 3509.055 4370.215 ;
        RECT 3509.485 4369.935 3509.765 4370.215 ;
        RECT 3500.255 4369.225 3500.535 4369.505 ;
        RECT 3500.965 4369.225 3501.245 4369.505 ;
        RECT 3501.675 4369.225 3501.955 4369.505 ;
        RECT 3502.385 4369.225 3502.665 4369.505 ;
        RECT 3503.095 4369.225 3503.375 4369.505 ;
        RECT 3503.805 4369.225 3504.085 4369.505 ;
        RECT 3504.515 4369.225 3504.795 4369.505 ;
        RECT 3505.225 4369.225 3505.505 4369.505 ;
        RECT 3505.935 4369.225 3506.215 4369.505 ;
        RECT 3506.645 4369.225 3506.925 4369.505 ;
        RECT 3507.355 4369.225 3507.635 4369.505 ;
        RECT 3508.065 4369.225 3508.345 4369.505 ;
        RECT 3508.775 4369.225 3509.055 4369.505 ;
        RECT 3509.485 4369.225 3509.765 4369.505 ;
        RECT 369.275 4368.715 369.555 4368.995 ;
        RECT 369.985 4368.715 370.265 4368.995 ;
        RECT 370.695 4368.715 370.975 4368.995 ;
        RECT 371.405 4368.715 371.685 4368.995 ;
        RECT 372.115 4368.715 372.395 4368.995 ;
        RECT 372.825 4368.715 373.105 4368.995 ;
        RECT 373.535 4368.715 373.815 4368.995 ;
        RECT 374.245 4368.715 374.525 4368.995 ;
        RECT 374.955 4368.715 375.235 4368.995 ;
        RECT 375.665 4368.715 375.945 4368.995 ;
        RECT 376.375 4368.715 376.655 4368.995 ;
        RECT 377.085 4368.715 377.365 4368.995 ;
        RECT 377.795 4368.715 378.075 4368.995 ;
        RECT 378.505 4368.715 378.785 4368.995 ;
        RECT 3500.255 4368.515 3500.535 4368.795 ;
        RECT 3500.965 4368.515 3501.245 4368.795 ;
        RECT 3501.675 4368.515 3501.955 4368.795 ;
        RECT 3502.385 4368.515 3502.665 4368.795 ;
        RECT 3503.095 4368.515 3503.375 4368.795 ;
        RECT 3503.805 4368.515 3504.085 4368.795 ;
        RECT 3504.515 4368.515 3504.795 4368.795 ;
        RECT 3505.225 4368.515 3505.505 4368.795 ;
        RECT 3505.935 4368.515 3506.215 4368.795 ;
        RECT 3506.645 4368.515 3506.925 4368.795 ;
        RECT 3507.355 4368.515 3507.635 4368.795 ;
        RECT 3508.065 4368.515 3508.345 4368.795 ;
        RECT 3508.775 4368.515 3509.055 4368.795 ;
        RECT 3509.485 4368.515 3509.765 4368.795 ;
        RECT 369.275 4368.005 369.555 4368.285 ;
        RECT 369.985 4368.005 370.265 4368.285 ;
        RECT 370.695 4368.005 370.975 4368.285 ;
        RECT 371.405 4368.005 371.685 4368.285 ;
        RECT 372.115 4368.005 372.395 4368.285 ;
        RECT 372.825 4368.005 373.105 4368.285 ;
        RECT 373.535 4368.005 373.815 4368.285 ;
        RECT 374.245 4368.005 374.525 4368.285 ;
        RECT 374.955 4368.005 375.235 4368.285 ;
        RECT 375.665 4368.005 375.945 4368.285 ;
        RECT 376.375 4368.005 376.655 4368.285 ;
        RECT 377.085 4368.005 377.365 4368.285 ;
        RECT 377.795 4368.005 378.075 4368.285 ;
        RECT 378.505 4368.005 378.785 4368.285 ;
        RECT 3500.255 4367.805 3500.535 4368.085 ;
        RECT 3500.965 4367.805 3501.245 4368.085 ;
        RECT 3501.675 4367.805 3501.955 4368.085 ;
        RECT 3502.385 4367.805 3502.665 4368.085 ;
        RECT 3503.095 4367.805 3503.375 4368.085 ;
        RECT 3503.805 4367.805 3504.085 4368.085 ;
        RECT 3504.515 4367.805 3504.795 4368.085 ;
        RECT 3505.225 4367.805 3505.505 4368.085 ;
        RECT 3505.935 4367.805 3506.215 4368.085 ;
        RECT 3506.645 4367.805 3506.925 4368.085 ;
        RECT 3507.355 4367.805 3507.635 4368.085 ;
        RECT 3508.065 4367.805 3508.345 4368.085 ;
        RECT 3508.775 4367.805 3509.055 4368.085 ;
        RECT 3509.485 4367.805 3509.765 4368.085 ;
        RECT 369.275 4367.295 369.555 4367.575 ;
        RECT 369.985 4367.295 370.265 4367.575 ;
        RECT 370.695 4367.295 370.975 4367.575 ;
        RECT 371.405 4367.295 371.685 4367.575 ;
        RECT 372.115 4367.295 372.395 4367.575 ;
        RECT 372.825 4367.295 373.105 4367.575 ;
        RECT 373.535 4367.295 373.815 4367.575 ;
        RECT 374.245 4367.295 374.525 4367.575 ;
        RECT 374.955 4367.295 375.235 4367.575 ;
        RECT 375.665 4367.295 375.945 4367.575 ;
        RECT 376.375 4367.295 376.655 4367.575 ;
        RECT 377.085 4367.295 377.365 4367.575 ;
        RECT 377.795 4367.295 378.075 4367.575 ;
        RECT 378.505 4367.295 378.785 4367.575 ;
        RECT 3500.255 4367.095 3500.535 4367.375 ;
        RECT 3500.965 4367.095 3501.245 4367.375 ;
        RECT 3501.675 4367.095 3501.955 4367.375 ;
        RECT 3502.385 4367.095 3502.665 4367.375 ;
        RECT 3503.095 4367.095 3503.375 4367.375 ;
        RECT 3503.805 4367.095 3504.085 4367.375 ;
        RECT 3504.515 4367.095 3504.795 4367.375 ;
        RECT 3505.225 4367.095 3505.505 4367.375 ;
        RECT 3505.935 4367.095 3506.215 4367.375 ;
        RECT 3506.645 4367.095 3506.925 4367.375 ;
        RECT 3507.355 4367.095 3507.635 4367.375 ;
        RECT 3508.065 4367.095 3508.345 4367.375 ;
        RECT 3508.775 4367.095 3509.055 4367.375 ;
        RECT 3509.485 4367.095 3509.765 4367.375 ;
        RECT 369.275 4366.585 369.555 4366.865 ;
        RECT 369.985 4366.585 370.265 4366.865 ;
        RECT 370.695 4366.585 370.975 4366.865 ;
        RECT 371.405 4366.585 371.685 4366.865 ;
        RECT 372.115 4366.585 372.395 4366.865 ;
        RECT 372.825 4366.585 373.105 4366.865 ;
        RECT 373.535 4366.585 373.815 4366.865 ;
        RECT 374.245 4366.585 374.525 4366.865 ;
        RECT 374.955 4366.585 375.235 4366.865 ;
        RECT 375.665 4366.585 375.945 4366.865 ;
        RECT 376.375 4366.585 376.655 4366.865 ;
        RECT 377.085 4366.585 377.365 4366.865 ;
        RECT 377.795 4366.585 378.075 4366.865 ;
        RECT 378.505 4366.585 378.785 4366.865 ;
        RECT 3500.255 4366.385 3500.535 4366.665 ;
        RECT 3500.965 4366.385 3501.245 4366.665 ;
        RECT 3501.675 4366.385 3501.955 4366.665 ;
        RECT 3502.385 4366.385 3502.665 4366.665 ;
        RECT 3503.095 4366.385 3503.375 4366.665 ;
        RECT 3503.805 4366.385 3504.085 4366.665 ;
        RECT 3504.515 4366.385 3504.795 4366.665 ;
        RECT 3505.225 4366.385 3505.505 4366.665 ;
        RECT 3505.935 4366.385 3506.215 4366.665 ;
        RECT 3506.645 4366.385 3506.925 4366.665 ;
        RECT 3507.355 4366.385 3507.635 4366.665 ;
        RECT 3508.065 4366.385 3508.345 4366.665 ;
        RECT 3508.775 4366.385 3509.055 4366.665 ;
        RECT 3509.485 4366.385 3509.765 4366.665 ;
        RECT 369.275 4365.875 369.555 4366.155 ;
        RECT 369.985 4365.875 370.265 4366.155 ;
        RECT 370.695 4365.875 370.975 4366.155 ;
        RECT 371.405 4365.875 371.685 4366.155 ;
        RECT 372.115 4365.875 372.395 4366.155 ;
        RECT 372.825 4365.875 373.105 4366.155 ;
        RECT 373.535 4365.875 373.815 4366.155 ;
        RECT 374.245 4365.875 374.525 4366.155 ;
        RECT 374.955 4365.875 375.235 4366.155 ;
        RECT 375.665 4365.875 375.945 4366.155 ;
        RECT 376.375 4365.875 376.655 4366.155 ;
        RECT 377.085 4365.875 377.365 4366.155 ;
        RECT 377.795 4365.875 378.075 4366.155 ;
        RECT 378.505 4365.875 378.785 4366.155 ;
        RECT 369.275 4365.165 369.555 4365.445 ;
        RECT 369.985 4365.165 370.265 4365.445 ;
        RECT 370.695 4365.165 370.975 4365.445 ;
        RECT 371.405 4365.165 371.685 4365.445 ;
        RECT 372.115 4365.165 372.395 4365.445 ;
        RECT 372.825 4365.165 373.105 4365.445 ;
        RECT 373.535 4365.165 373.815 4365.445 ;
        RECT 374.245 4365.165 374.525 4365.445 ;
        RECT 374.955 4365.165 375.235 4365.445 ;
        RECT 375.665 4365.165 375.945 4365.445 ;
        RECT 376.375 4365.165 376.655 4365.445 ;
        RECT 377.085 4365.165 377.365 4365.445 ;
        RECT 377.795 4365.165 378.075 4365.445 ;
        RECT 378.505 4365.165 378.785 4365.445 ;
        RECT 369.275 4364.455 369.555 4364.735 ;
        RECT 369.985 4364.455 370.265 4364.735 ;
        RECT 370.695 4364.455 370.975 4364.735 ;
        RECT 371.405 4364.455 371.685 4364.735 ;
        RECT 372.115 4364.455 372.395 4364.735 ;
        RECT 372.825 4364.455 373.105 4364.735 ;
        RECT 373.535 4364.455 373.815 4364.735 ;
        RECT 374.245 4364.455 374.525 4364.735 ;
        RECT 374.955 4364.455 375.235 4364.735 ;
        RECT 375.665 4364.455 375.945 4364.735 ;
        RECT 376.375 4364.455 376.655 4364.735 ;
        RECT 377.085 4364.455 377.365 4364.735 ;
        RECT 377.795 4364.455 378.075 4364.735 ;
        RECT 378.505 4364.455 378.785 4364.735 ;
        RECT 369.275 4363.745 369.555 4364.025 ;
        RECT 369.985 4363.745 370.265 4364.025 ;
        RECT 370.695 4363.745 370.975 4364.025 ;
        RECT 371.405 4363.745 371.685 4364.025 ;
        RECT 372.115 4363.745 372.395 4364.025 ;
        RECT 372.825 4363.745 373.105 4364.025 ;
        RECT 373.535 4363.745 373.815 4364.025 ;
        RECT 374.245 4363.745 374.525 4364.025 ;
        RECT 374.955 4363.745 375.235 4364.025 ;
        RECT 375.665 4363.745 375.945 4364.025 ;
        RECT 376.375 4363.745 376.655 4364.025 ;
        RECT 377.085 4363.745 377.365 4364.025 ;
        RECT 377.795 4363.745 378.075 4364.025 ;
        RECT 378.505 4363.745 378.785 4364.025 ;
        RECT 3500.255 4363.765 3500.535 4364.045 ;
        RECT 3500.965 4363.765 3501.245 4364.045 ;
        RECT 3501.675 4363.765 3501.955 4364.045 ;
        RECT 3502.385 4363.765 3502.665 4364.045 ;
        RECT 3503.095 4363.765 3503.375 4364.045 ;
        RECT 3503.805 4363.765 3504.085 4364.045 ;
        RECT 3504.515 4363.765 3504.795 4364.045 ;
        RECT 3505.225 4363.765 3505.505 4364.045 ;
        RECT 3505.935 4363.765 3506.215 4364.045 ;
        RECT 3506.645 4363.765 3506.925 4364.045 ;
        RECT 3507.355 4363.765 3507.635 4364.045 ;
        RECT 3508.065 4363.765 3508.345 4364.045 ;
        RECT 3508.775 4363.765 3509.055 4364.045 ;
        RECT 3509.485 4363.765 3509.765 4364.045 ;
        RECT 369.275 4363.035 369.555 4363.315 ;
        RECT 369.985 4363.035 370.265 4363.315 ;
        RECT 370.695 4363.035 370.975 4363.315 ;
        RECT 371.405 4363.035 371.685 4363.315 ;
        RECT 372.115 4363.035 372.395 4363.315 ;
        RECT 372.825 4363.035 373.105 4363.315 ;
        RECT 373.535 4363.035 373.815 4363.315 ;
        RECT 374.245 4363.035 374.525 4363.315 ;
        RECT 374.955 4363.035 375.235 4363.315 ;
        RECT 375.665 4363.035 375.945 4363.315 ;
        RECT 376.375 4363.035 376.655 4363.315 ;
        RECT 377.085 4363.035 377.365 4363.315 ;
        RECT 377.795 4363.035 378.075 4363.315 ;
        RECT 378.505 4363.035 378.785 4363.315 ;
        RECT 3500.255 4363.055 3500.535 4363.335 ;
        RECT 3500.965 4363.055 3501.245 4363.335 ;
        RECT 3501.675 4363.055 3501.955 4363.335 ;
        RECT 3502.385 4363.055 3502.665 4363.335 ;
        RECT 3503.095 4363.055 3503.375 4363.335 ;
        RECT 3503.805 4363.055 3504.085 4363.335 ;
        RECT 3504.515 4363.055 3504.795 4363.335 ;
        RECT 3505.225 4363.055 3505.505 4363.335 ;
        RECT 3505.935 4363.055 3506.215 4363.335 ;
        RECT 3506.645 4363.055 3506.925 4363.335 ;
        RECT 3507.355 4363.055 3507.635 4363.335 ;
        RECT 3508.065 4363.055 3508.345 4363.335 ;
        RECT 3508.775 4363.055 3509.055 4363.335 ;
        RECT 3509.485 4363.055 3509.765 4363.335 ;
        RECT 369.275 4362.325 369.555 4362.605 ;
        RECT 369.985 4362.325 370.265 4362.605 ;
        RECT 370.695 4362.325 370.975 4362.605 ;
        RECT 371.405 4362.325 371.685 4362.605 ;
        RECT 372.115 4362.325 372.395 4362.605 ;
        RECT 372.825 4362.325 373.105 4362.605 ;
        RECT 373.535 4362.325 373.815 4362.605 ;
        RECT 374.245 4362.325 374.525 4362.605 ;
        RECT 374.955 4362.325 375.235 4362.605 ;
        RECT 375.665 4362.325 375.945 4362.605 ;
        RECT 376.375 4362.325 376.655 4362.605 ;
        RECT 377.085 4362.325 377.365 4362.605 ;
        RECT 377.795 4362.325 378.075 4362.605 ;
        RECT 378.505 4362.325 378.785 4362.605 ;
        RECT 3500.255 4362.345 3500.535 4362.625 ;
        RECT 3500.965 4362.345 3501.245 4362.625 ;
        RECT 3501.675 4362.345 3501.955 4362.625 ;
        RECT 3502.385 4362.345 3502.665 4362.625 ;
        RECT 3503.095 4362.345 3503.375 4362.625 ;
        RECT 3503.805 4362.345 3504.085 4362.625 ;
        RECT 3504.515 4362.345 3504.795 4362.625 ;
        RECT 3505.225 4362.345 3505.505 4362.625 ;
        RECT 3505.935 4362.345 3506.215 4362.625 ;
        RECT 3506.645 4362.345 3506.925 4362.625 ;
        RECT 3507.355 4362.345 3507.635 4362.625 ;
        RECT 3508.065 4362.345 3508.345 4362.625 ;
        RECT 3508.775 4362.345 3509.055 4362.625 ;
        RECT 3509.485 4362.345 3509.765 4362.625 ;
        RECT 369.275 4361.615 369.555 4361.895 ;
        RECT 369.985 4361.615 370.265 4361.895 ;
        RECT 370.695 4361.615 370.975 4361.895 ;
        RECT 371.405 4361.615 371.685 4361.895 ;
        RECT 372.115 4361.615 372.395 4361.895 ;
        RECT 372.825 4361.615 373.105 4361.895 ;
        RECT 373.535 4361.615 373.815 4361.895 ;
        RECT 374.245 4361.615 374.525 4361.895 ;
        RECT 374.955 4361.615 375.235 4361.895 ;
        RECT 375.665 4361.615 375.945 4361.895 ;
        RECT 376.375 4361.615 376.655 4361.895 ;
        RECT 377.085 4361.615 377.365 4361.895 ;
        RECT 377.795 4361.615 378.075 4361.895 ;
        RECT 378.505 4361.615 378.785 4361.895 ;
        RECT 3500.255 4361.635 3500.535 4361.915 ;
        RECT 3500.965 4361.635 3501.245 4361.915 ;
        RECT 3501.675 4361.635 3501.955 4361.915 ;
        RECT 3502.385 4361.635 3502.665 4361.915 ;
        RECT 3503.095 4361.635 3503.375 4361.915 ;
        RECT 3503.805 4361.635 3504.085 4361.915 ;
        RECT 3504.515 4361.635 3504.795 4361.915 ;
        RECT 3505.225 4361.635 3505.505 4361.915 ;
        RECT 3505.935 4361.635 3506.215 4361.915 ;
        RECT 3506.645 4361.635 3506.925 4361.915 ;
        RECT 3507.355 4361.635 3507.635 4361.915 ;
        RECT 3508.065 4361.635 3508.345 4361.915 ;
        RECT 3508.775 4361.635 3509.055 4361.915 ;
        RECT 3509.485 4361.635 3509.765 4361.915 ;
        RECT 369.275 4360.905 369.555 4361.185 ;
        RECT 369.985 4360.905 370.265 4361.185 ;
        RECT 370.695 4360.905 370.975 4361.185 ;
        RECT 371.405 4360.905 371.685 4361.185 ;
        RECT 372.115 4360.905 372.395 4361.185 ;
        RECT 372.825 4360.905 373.105 4361.185 ;
        RECT 373.535 4360.905 373.815 4361.185 ;
        RECT 374.245 4360.905 374.525 4361.185 ;
        RECT 374.955 4360.905 375.235 4361.185 ;
        RECT 375.665 4360.905 375.945 4361.185 ;
        RECT 376.375 4360.905 376.655 4361.185 ;
        RECT 377.085 4360.905 377.365 4361.185 ;
        RECT 377.795 4360.905 378.075 4361.185 ;
        RECT 378.505 4360.905 378.785 4361.185 ;
        RECT 3500.255 4360.925 3500.535 4361.205 ;
        RECT 3500.965 4360.925 3501.245 4361.205 ;
        RECT 3501.675 4360.925 3501.955 4361.205 ;
        RECT 3502.385 4360.925 3502.665 4361.205 ;
        RECT 3503.095 4360.925 3503.375 4361.205 ;
        RECT 3503.805 4360.925 3504.085 4361.205 ;
        RECT 3504.515 4360.925 3504.795 4361.205 ;
        RECT 3505.225 4360.925 3505.505 4361.205 ;
        RECT 3505.935 4360.925 3506.215 4361.205 ;
        RECT 3506.645 4360.925 3506.925 4361.205 ;
        RECT 3507.355 4360.925 3507.635 4361.205 ;
        RECT 3508.065 4360.925 3508.345 4361.205 ;
        RECT 3508.775 4360.925 3509.055 4361.205 ;
        RECT 3509.485 4360.925 3509.765 4361.205 ;
        RECT 369.275 4360.195 369.555 4360.475 ;
        RECT 369.985 4360.195 370.265 4360.475 ;
        RECT 370.695 4360.195 370.975 4360.475 ;
        RECT 371.405 4360.195 371.685 4360.475 ;
        RECT 372.115 4360.195 372.395 4360.475 ;
        RECT 372.825 4360.195 373.105 4360.475 ;
        RECT 373.535 4360.195 373.815 4360.475 ;
        RECT 374.245 4360.195 374.525 4360.475 ;
        RECT 374.955 4360.195 375.235 4360.475 ;
        RECT 375.665 4360.195 375.945 4360.475 ;
        RECT 376.375 4360.195 376.655 4360.475 ;
        RECT 377.085 4360.195 377.365 4360.475 ;
        RECT 377.795 4360.195 378.075 4360.475 ;
        RECT 378.505 4360.195 378.785 4360.475 ;
        RECT 3500.255 4360.215 3500.535 4360.495 ;
        RECT 3500.965 4360.215 3501.245 4360.495 ;
        RECT 3501.675 4360.215 3501.955 4360.495 ;
        RECT 3502.385 4360.215 3502.665 4360.495 ;
        RECT 3503.095 4360.215 3503.375 4360.495 ;
        RECT 3503.805 4360.215 3504.085 4360.495 ;
        RECT 3504.515 4360.215 3504.795 4360.495 ;
        RECT 3505.225 4360.215 3505.505 4360.495 ;
        RECT 3505.935 4360.215 3506.215 4360.495 ;
        RECT 3506.645 4360.215 3506.925 4360.495 ;
        RECT 3507.355 4360.215 3507.635 4360.495 ;
        RECT 3508.065 4360.215 3508.345 4360.495 ;
        RECT 3508.775 4360.215 3509.055 4360.495 ;
        RECT 3509.485 4360.215 3509.765 4360.495 ;
        RECT 369.275 4359.485 369.555 4359.765 ;
        RECT 369.985 4359.485 370.265 4359.765 ;
        RECT 370.695 4359.485 370.975 4359.765 ;
        RECT 371.405 4359.485 371.685 4359.765 ;
        RECT 372.115 4359.485 372.395 4359.765 ;
        RECT 372.825 4359.485 373.105 4359.765 ;
        RECT 373.535 4359.485 373.815 4359.765 ;
        RECT 374.245 4359.485 374.525 4359.765 ;
        RECT 374.955 4359.485 375.235 4359.765 ;
        RECT 375.665 4359.485 375.945 4359.765 ;
        RECT 376.375 4359.485 376.655 4359.765 ;
        RECT 377.085 4359.485 377.365 4359.765 ;
        RECT 377.795 4359.485 378.075 4359.765 ;
        RECT 378.505 4359.485 378.785 4359.765 ;
        RECT 3500.255 4359.505 3500.535 4359.785 ;
        RECT 3500.965 4359.505 3501.245 4359.785 ;
        RECT 3501.675 4359.505 3501.955 4359.785 ;
        RECT 3502.385 4359.505 3502.665 4359.785 ;
        RECT 3503.095 4359.505 3503.375 4359.785 ;
        RECT 3503.805 4359.505 3504.085 4359.785 ;
        RECT 3504.515 4359.505 3504.795 4359.785 ;
        RECT 3505.225 4359.505 3505.505 4359.785 ;
        RECT 3505.935 4359.505 3506.215 4359.785 ;
        RECT 3506.645 4359.505 3506.925 4359.785 ;
        RECT 3507.355 4359.505 3507.635 4359.785 ;
        RECT 3508.065 4359.505 3508.345 4359.785 ;
        RECT 3508.775 4359.505 3509.055 4359.785 ;
        RECT 3509.485 4359.505 3509.765 4359.785 ;
        RECT 3500.255 4358.795 3500.535 4359.075 ;
        RECT 3500.965 4358.795 3501.245 4359.075 ;
        RECT 3501.675 4358.795 3501.955 4359.075 ;
        RECT 3502.385 4358.795 3502.665 4359.075 ;
        RECT 3503.095 4358.795 3503.375 4359.075 ;
        RECT 3503.805 4358.795 3504.085 4359.075 ;
        RECT 3504.515 4358.795 3504.795 4359.075 ;
        RECT 3505.225 4358.795 3505.505 4359.075 ;
        RECT 3505.935 4358.795 3506.215 4359.075 ;
        RECT 3506.645 4358.795 3506.925 4359.075 ;
        RECT 3507.355 4358.795 3507.635 4359.075 ;
        RECT 3508.065 4358.795 3508.345 4359.075 ;
        RECT 3508.775 4358.795 3509.055 4359.075 ;
        RECT 3509.485 4358.795 3509.765 4359.075 ;
        RECT 3500.255 4358.085 3500.535 4358.365 ;
        RECT 3500.965 4358.085 3501.245 4358.365 ;
        RECT 3501.675 4358.085 3501.955 4358.365 ;
        RECT 3502.385 4358.085 3502.665 4358.365 ;
        RECT 3503.095 4358.085 3503.375 4358.365 ;
        RECT 3503.805 4358.085 3504.085 4358.365 ;
        RECT 3504.515 4358.085 3504.795 4358.365 ;
        RECT 3505.225 4358.085 3505.505 4358.365 ;
        RECT 3505.935 4358.085 3506.215 4358.365 ;
        RECT 3506.645 4358.085 3506.925 4358.365 ;
        RECT 3507.355 4358.085 3507.635 4358.365 ;
        RECT 3508.065 4358.085 3508.345 4358.365 ;
        RECT 3508.775 4358.085 3509.055 4358.365 ;
        RECT 3509.485 4358.085 3509.765 4358.365 ;
        RECT 3500.255 4357.375 3500.535 4357.655 ;
        RECT 3500.965 4357.375 3501.245 4357.655 ;
        RECT 3501.675 4357.375 3501.955 4357.655 ;
        RECT 3502.385 4357.375 3502.665 4357.655 ;
        RECT 3503.095 4357.375 3503.375 4357.655 ;
        RECT 3503.805 4357.375 3504.085 4357.655 ;
        RECT 3504.515 4357.375 3504.795 4357.655 ;
        RECT 3505.225 4357.375 3505.505 4357.655 ;
        RECT 3505.935 4357.375 3506.215 4357.655 ;
        RECT 3506.645 4357.375 3506.925 4357.655 ;
        RECT 3507.355 4357.375 3507.635 4357.655 ;
        RECT 3508.065 4357.375 3508.345 4357.655 ;
        RECT 3508.775 4357.375 3509.055 4357.655 ;
        RECT 3509.485 4357.375 3509.765 4357.655 ;
        RECT 3500.255 4356.665 3500.535 4356.945 ;
        RECT 3500.965 4356.665 3501.245 4356.945 ;
        RECT 3501.675 4356.665 3501.955 4356.945 ;
        RECT 3502.385 4356.665 3502.665 4356.945 ;
        RECT 3503.095 4356.665 3503.375 4356.945 ;
        RECT 3503.805 4356.665 3504.085 4356.945 ;
        RECT 3504.515 4356.665 3504.795 4356.945 ;
        RECT 3505.225 4356.665 3505.505 4356.945 ;
        RECT 3505.935 4356.665 3506.215 4356.945 ;
        RECT 3506.645 4356.665 3506.925 4356.945 ;
        RECT 3507.355 4356.665 3507.635 4356.945 ;
        RECT 3508.065 4356.665 3508.345 4356.945 ;
        RECT 3508.775 4356.665 3509.055 4356.945 ;
        RECT 3509.485 4356.665 3509.765 4356.945 ;
        RECT 3500.255 4355.955 3500.535 4356.235 ;
        RECT 3500.965 4355.955 3501.245 4356.235 ;
        RECT 3501.675 4355.955 3501.955 4356.235 ;
        RECT 3502.385 4355.955 3502.665 4356.235 ;
        RECT 3503.095 4355.955 3503.375 4356.235 ;
        RECT 3503.805 4355.955 3504.085 4356.235 ;
        RECT 3504.515 4355.955 3504.795 4356.235 ;
        RECT 3505.225 4355.955 3505.505 4356.235 ;
        RECT 3505.935 4355.955 3506.215 4356.235 ;
        RECT 3506.645 4355.955 3506.925 4356.235 ;
        RECT 3507.355 4355.955 3507.635 4356.235 ;
        RECT 3508.065 4355.955 3508.345 4356.235 ;
        RECT 3508.775 4355.955 3509.055 4356.235 ;
        RECT 3509.485 4355.955 3509.765 4356.235 ;
        RECT 369.275 4355.185 369.555 4355.465 ;
        RECT 369.985 4355.185 370.265 4355.465 ;
        RECT 370.695 4355.185 370.975 4355.465 ;
        RECT 371.405 4355.185 371.685 4355.465 ;
        RECT 372.115 4355.185 372.395 4355.465 ;
        RECT 372.825 4355.185 373.105 4355.465 ;
        RECT 373.535 4355.185 373.815 4355.465 ;
        RECT 374.245 4355.185 374.525 4355.465 ;
        RECT 374.955 4355.185 375.235 4355.465 ;
        RECT 375.665 4355.185 375.945 4355.465 ;
        RECT 376.375 4355.185 376.655 4355.465 ;
        RECT 377.085 4355.185 377.365 4355.465 ;
        RECT 377.795 4355.185 378.075 4355.465 ;
        RECT 378.505 4355.185 378.785 4355.465 ;
        RECT 3500.255 4355.245 3500.535 4355.525 ;
        RECT 3500.965 4355.245 3501.245 4355.525 ;
        RECT 3501.675 4355.245 3501.955 4355.525 ;
        RECT 3502.385 4355.245 3502.665 4355.525 ;
        RECT 3503.095 4355.245 3503.375 4355.525 ;
        RECT 3503.805 4355.245 3504.085 4355.525 ;
        RECT 3504.515 4355.245 3504.795 4355.525 ;
        RECT 3505.225 4355.245 3505.505 4355.525 ;
        RECT 3505.935 4355.245 3506.215 4355.525 ;
        RECT 3506.645 4355.245 3506.925 4355.525 ;
        RECT 3507.355 4355.245 3507.635 4355.525 ;
        RECT 3508.065 4355.245 3508.345 4355.525 ;
        RECT 3508.775 4355.245 3509.055 4355.525 ;
        RECT 3509.485 4355.245 3509.765 4355.525 ;
        RECT 369.275 4354.475 369.555 4354.755 ;
        RECT 369.985 4354.475 370.265 4354.755 ;
        RECT 370.695 4354.475 370.975 4354.755 ;
        RECT 371.405 4354.475 371.685 4354.755 ;
        RECT 372.115 4354.475 372.395 4354.755 ;
        RECT 372.825 4354.475 373.105 4354.755 ;
        RECT 373.535 4354.475 373.815 4354.755 ;
        RECT 374.245 4354.475 374.525 4354.755 ;
        RECT 374.955 4354.475 375.235 4354.755 ;
        RECT 375.665 4354.475 375.945 4354.755 ;
        RECT 376.375 4354.475 376.655 4354.755 ;
        RECT 377.085 4354.475 377.365 4354.755 ;
        RECT 377.795 4354.475 378.075 4354.755 ;
        RECT 378.505 4354.475 378.785 4354.755 ;
        RECT 3500.255 4354.535 3500.535 4354.815 ;
        RECT 3500.965 4354.535 3501.245 4354.815 ;
        RECT 3501.675 4354.535 3501.955 4354.815 ;
        RECT 3502.385 4354.535 3502.665 4354.815 ;
        RECT 3503.095 4354.535 3503.375 4354.815 ;
        RECT 3503.805 4354.535 3504.085 4354.815 ;
        RECT 3504.515 4354.535 3504.795 4354.815 ;
        RECT 3505.225 4354.535 3505.505 4354.815 ;
        RECT 3505.935 4354.535 3506.215 4354.815 ;
        RECT 3506.645 4354.535 3506.925 4354.815 ;
        RECT 3507.355 4354.535 3507.635 4354.815 ;
        RECT 3508.065 4354.535 3508.345 4354.815 ;
        RECT 3508.775 4354.535 3509.055 4354.815 ;
        RECT 3509.485 4354.535 3509.765 4354.815 ;
        RECT 369.275 4353.765 369.555 4354.045 ;
        RECT 369.985 4353.765 370.265 4354.045 ;
        RECT 370.695 4353.765 370.975 4354.045 ;
        RECT 371.405 4353.765 371.685 4354.045 ;
        RECT 372.115 4353.765 372.395 4354.045 ;
        RECT 372.825 4353.765 373.105 4354.045 ;
        RECT 373.535 4353.765 373.815 4354.045 ;
        RECT 374.245 4353.765 374.525 4354.045 ;
        RECT 374.955 4353.765 375.235 4354.045 ;
        RECT 375.665 4353.765 375.945 4354.045 ;
        RECT 376.375 4353.765 376.655 4354.045 ;
        RECT 377.085 4353.765 377.365 4354.045 ;
        RECT 377.795 4353.765 378.075 4354.045 ;
        RECT 378.505 4353.765 378.785 4354.045 ;
        RECT 369.275 4353.055 369.555 4353.335 ;
        RECT 369.985 4353.055 370.265 4353.335 ;
        RECT 370.695 4353.055 370.975 4353.335 ;
        RECT 371.405 4353.055 371.685 4353.335 ;
        RECT 372.115 4353.055 372.395 4353.335 ;
        RECT 372.825 4353.055 373.105 4353.335 ;
        RECT 373.535 4353.055 373.815 4353.335 ;
        RECT 374.245 4353.055 374.525 4353.335 ;
        RECT 374.955 4353.055 375.235 4353.335 ;
        RECT 375.665 4353.055 375.945 4353.335 ;
        RECT 376.375 4353.055 376.655 4353.335 ;
        RECT 377.085 4353.055 377.365 4353.335 ;
        RECT 377.795 4353.055 378.075 4353.335 ;
        RECT 378.505 4353.055 378.785 4353.335 ;
        RECT 369.275 4352.345 369.555 4352.625 ;
        RECT 369.985 4352.345 370.265 4352.625 ;
        RECT 370.695 4352.345 370.975 4352.625 ;
        RECT 371.405 4352.345 371.685 4352.625 ;
        RECT 372.115 4352.345 372.395 4352.625 ;
        RECT 372.825 4352.345 373.105 4352.625 ;
        RECT 373.535 4352.345 373.815 4352.625 ;
        RECT 374.245 4352.345 374.525 4352.625 ;
        RECT 374.955 4352.345 375.235 4352.625 ;
        RECT 375.665 4352.345 375.945 4352.625 ;
        RECT 376.375 4352.345 376.655 4352.625 ;
        RECT 377.085 4352.345 377.365 4352.625 ;
        RECT 377.795 4352.345 378.075 4352.625 ;
        RECT 378.505 4352.345 378.785 4352.625 ;
        RECT 369.275 4351.635 369.555 4351.915 ;
        RECT 369.985 4351.635 370.265 4351.915 ;
        RECT 370.695 4351.635 370.975 4351.915 ;
        RECT 371.405 4351.635 371.685 4351.915 ;
        RECT 372.115 4351.635 372.395 4351.915 ;
        RECT 372.825 4351.635 373.105 4351.915 ;
        RECT 373.535 4351.635 373.815 4351.915 ;
        RECT 374.245 4351.635 374.525 4351.915 ;
        RECT 374.955 4351.635 375.235 4351.915 ;
        RECT 375.665 4351.635 375.945 4351.915 ;
        RECT 376.375 4351.635 376.655 4351.915 ;
        RECT 377.085 4351.635 377.365 4351.915 ;
        RECT 377.795 4351.635 378.075 4351.915 ;
        RECT 378.505 4351.635 378.785 4351.915 ;
        RECT 369.275 4350.925 369.555 4351.205 ;
        RECT 369.985 4350.925 370.265 4351.205 ;
        RECT 370.695 4350.925 370.975 4351.205 ;
        RECT 371.405 4350.925 371.685 4351.205 ;
        RECT 372.115 4350.925 372.395 4351.205 ;
        RECT 372.825 4350.925 373.105 4351.205 ;
        RECT 373.535 4350.925 373.815 4351.205 ;
        RECT 374.245 4350.925 374.525 4351.205 ;
        RECT 374.955 4350.925 375.235 4351.205 ;
        RECT 375.665 4350.925 375.945 4351.205 ;
        RECT 376.375 4350.925 376.655 4351.205 ;
        RECT 377.085 4350.925 377.365 4351.205 ;
        RECT 377.795 4350.925 378.075 4351.205 ;
        RECT 378.505 4350.925 378.785 4351.205 ;
        RECT 369.275 4350.215 369.555 4350.495 ;
        RECT 369.985 4350.215 370.265 4350.495 ;
        RECT 370.695 4350.215 370.975 4350.495 ;
        RECT 371.405 4350.215 371.685 4350.495 ;
        RECT 372.115 4350.215 372.395 4350.495 ;
        RECT 372.825 4350.215 373.105 4350.495 ;
        RECT 373.535 4350.215 373.815 4350.495 ;
        RECT 374.245 4350.215 374.525 4350.495 ;
        RECT 374.955 4350.215 375.235 4350.495 ;
        RECT 375.665 4350.215 375.945 4350.495 ;
        RECT 376.375 4350.215 376.655 4350.495 ;
        RECT 377.085 4350.215 377.365 4350.495 ;
        RECT 377.795 4350.215 378.075 4350.495 ;
        RECT 378.505 4350.215 378.785 4350.495 ;
        RECT 3500.255 4350.235 3500.535 4350.515 ;
        RECT 3500.965 4350.235 3501.245 4350.515 ;
        RECT 3501.675 4350.235 3501.955 4350.515 ;
        RECT 3502.385 4350.235 3502.665 4350.515 ;
        RECT 3503.095 4350.235 3503.375 4350.515 ;
        RECT 3503.805 4350.235 3504.085 4350.515 ;
        RECT 3504.515 4350.235 3504.795 4350.515 ;
        RECT 3505.225 4350.235 3505.505 4350.515 ;
        RECT 3505.935 4350.235 3506.215 4350.515 ;
        RECT 3506.645 4350.235 3506.925 4350.515 ;
        RECT 3507.355 4350.235 3507.635 4350.515 ;
        RECT 3508.065 4350.235 3508.345 4350.515 ;
        RECT 3508.775 4350.235 3509.055 4350.515 ;
        RECT 3509.485 4350.235 3509.765 4350.515 ;
        RECT 369.275 4349.505 369.555 4349.785 ;
        RECT 369.985 4349.505 370.265 4349.785 ;
        RECT 370.695 4349.505 370.975 4349.785 ;
        RECT 371.405 4349.505 371.685 4349.785 ;
        RECT 372.115 4349.505 372.395 4349.785 ;
        RECT 372.825 4349.505 373.105 4349.785 ;
        RECT 373.535 4349.505 373.815 4349.785 ;
        RECT 374.245 4349.505 374.525 4349.785 ;
        RECT 374.955 4349.505 375.235 4349.785 ;
        RECT 375.665 4349.505 375.945 4349.785 ;
        RECT 376.375 4349.505 376.655 4349.785 ;
        RECT 377.085 4349.505 377.365 4349.785 ;
        RECT 377.795 4349.505 378.075 4349.785 ;
        RECT 378.505 4349.505 378.785 4349.785 ;
        RECT 3500.255 4349.525 3500.535 4349.805 ;
        RECT 3500.965 4349.525 3501.245 4349.805 ;
        RECT 3501.675 4349.525 3501.955 4349.805 ;
        RECT 3502.385 4349.525 3502.665 4349.805 ;
        RECT 3503.095 4349.525 3503.375 4349.805 ;
        RECT 3503.805 4349.525 3504.085 4349.805 ;
        RECT 3504.515 4349.525 3504.795 4349.805 ;
        RECT 3505.225 4349.525 3505.505 4349.805 ;
        RECT 3505.935 4349.525 3506.215 4349.805 ;
        RECT 3506.645 4349.525 3506.925 4349.805 ;
        RECT 3507.355 4349.525 3507.635 4349.805 ;
        RECT 3508.065 4349.525 3508.345 4349.805 ;
        RECT 3508.775 4349.525 3509.055 4349.805 ;
        RECT 3509.485 4349.525 3509.765 4349.805 ;
        RECT 369.275 4348.795 369.555 4349.075 ;
        RECT 369.985 4348.795 370.265 4349.075 ;
        RECT 370.695 4348.795 370.975 4349.075 ;
        RECT 371.405 4348.795 371.685 4349.075 ;
        RECT 372.115 4348.795 372.395 4349.075 ;
        RECT 372.825 4348.795 373.105 4349.075 ;
        RECT 373.535 4348.795 373.815 4349.075 ;
        RECT 374.245 4348.795 374.525 4349.075 ;
        RECT 374.955 4348.795 375.235 4349.075 ;
        RECT 375.665 4348.795 375.945 4349.075 ;
        RECT 376.375 4348.795 376.655 4349.075 ;
        RECT 377.085 4348.795 377.365 4349.075 ;
        RECT 377.795 4348.795 378.075 4349.075 ;
        RECT 378.505 4348.795 378.785 4349.075 ;
        RECT 3500.255 4348.815 3500.535 4349.095 ;
        RECT 3500.965 4348.815 3501.245 4349.095 ;
        RECT 3501.675 4348.815 3501.955 4349.095 ;
        RECT 3502.385 4348.815 3502.665 4349.095 ;
        RECT 3503.095 4348.815 3503.375 4349.095 ;
        RECT 3503.805 4348.815 3504.085 4349.095 ;
        RECT 3504.515 4348.815 3504.795 4349.095 ;
        RECT 3505.225 4348.815 3505.505 4349.095 ;
        RECT 3505.935 4348.815 3506.215 4349.095 ;
        RECT 3506.645 4348.815 3506.925 4349.095 ;
        RECT 3507.355 4348.815 3507.635 4349.095 ;
        RECT 3508.065 4348.815 3508.345 4349.095 ;
        RECT 3508.775 4348.815 3509.055 4349.095 ;
        RECT 3509.485 4348.815 3509.765 4349.095 ;
        RECT 369.275 4348.085 369.555 4348.365 ;
        RECT 369.985 4348.085 370.265 4348.365 ;
        RECT 370.695 4348.085 370.975 4348.365 ;
        RECT 371.405 4348.085 371.685 4348.365 ;
        RECT 372.115 4348.085 372.395 4348.365 ;
        RECT 372.825 4348.085 373.105 4348.365 ;
        RECT 373.535 4348.085 373.815 4348.365 ;
        RECT 374.245 4348.085 374.525 4348.365 ;
        RECT 374.955 4348.085 375.235 4348.365 ;
        RECT 375.665 4348.085 375.945 4348.365 ;
        RECT 376.375 4348.085 376.655 4348.365 ;
        RECT 377.085 4348.085 377.365 4348.365 ;
        RECT 377.795 4348.085 378.075 4348.365 ;
        RECT 378.505 4348.085 378.785 4348.365 ;
        RECT 3500.255 4348.105 3500.535 4348.385 ;
        RECT 3500.965 4348.105 3501.245 4348.385 ;
        RECT 3501.675 4348.105 3501.955 4348.385 ;
        RECT 3502.385 4348.105 3502.665 4348.385 ;
        RECT 3503.095 4348.105 3503.375 4348.385 ;
        RECT 3503.805 4348.105 3504.085 4348.385 ;
        RECT 3504.515 4348.105 3504.795 4348.385 ;
        RECT 3505.225 4348.105 3505.505 4348.385 ;
        RECT 3505.935 4348.105 3506.215 4348.385 ;
        RECT 3506.645 4348.105 3506.925 4348.385 ;
        RECT 3507.355 4348.105 3507.635 4348.385 ;
        RECT 3508.065 4348.105 3508.345 4348.385 ;
        RECT 3508.775 4348.105 3509.055 4348.385 ;
        RECT 3509.485 4348.105 3509.765 4348.385 ;
        RECT 369.275 4347.375 369.555 4347.655 ;
        RECT 369.985 4347.375 370.265 4347.655 ;
        RECT 370.695 4347.375 370.975 4347.655 ;
        RECT 371.405 4347.375 371.685 4347.655 ;
        RECT 372.115 4347.375 372.395 4347.655 ;
        RECT 372.825 4347.375 373.105 4347.655 ;
        RECT 373.535 4347.375 373.815 4347.655 ;
        RECT 374.245 4347.375 374.525 4347.655 ;
        RECT 374.955 4347.375 375.235 4347.655 ;
        RECT 375.665 4347.375 375.945 4347.655 ;
        RECT 376.375 4347.375 376.655 4347.655 ;
        RECT 377.085 4347.375 377.365 4347.655 ;
        RECT 377.795 4347.375 378.075 4347.655 ;
        RECT 378.505 4347.375 378.785 4347.655 ;
        RECT 3500.255 4347.395 3500.535 4347.675 ;
        RECT 3500.965 4347.395 3501.245 4347.675 ;
        RECT 3501.675 4347.395 3501.955 4347.675 ;
        RECT 3502.385 4347.395 3502.665 4347.675 ;
        RECT 3503.095 4347.395 3503.375 4347.675 ;
        RECT 3503.805 4347.395 3504.085 4347.675 ;
        RECT 3504.515 4347.395 3504.795 4347.675 ;
        RECT 3505.225 4347.395 3505.505 4347.675 ;
        RECT 3505.935 4347.395 3506.215 4347.675 ;
        RECT 3506.645 4347.395 3506.925 4347.675 ;
        RECT 3507.355 4347.395 3507.635 4347.675 ;
        RECT 3508.065 4347.395 3508.345 4347.675 ;
        RECT 3508.775 4347.395 3509.055 4347.675 ;
        RECT 3509.485 4347.395 3509.765 4347.675 ;
        RECT 369.275 4346.665 369.555 4346.945 ;
        RECT 369.985 4346.665 370.265 4346.945 ;
        RECT 370.695 4346.665 370.975 4346.945 ;
        RECT 371.405 4346.665 371.685 4346.945 ;
        RECT 372.115 4346.665 372.395 4346.945 ;
        RECT 372.825 4346.665 373.105 4346.945 ;
        RECT 373.535 4346.665 373.815 4346.945 ;
        RECT 374.245 4346.665 374.525 4346.945 ;
        RECT 374.955 4346.665 375.235 4346.945 ;
        RECT 375.665 4346.665 375.945 4346.945 ;
        RECT 376.375 4346.665 376.655 4346.945 ;
        RECT 377.085 4346.665 377.365 4346.945 ;
        RECT 377.795 4346.665 378.075 4346.945 ;
        RECT 378.505 4346.665 378.785 4346.945 ;
        RECT 3500.255 4346.685 3500.535 4346.965 ;
        RECT 3500.965 4346.685 3501.245 4346.965 ;
        RECT 3501.675 4346.685 3501.955 4346.965 ;
        RECT 3502.385 4346.685 3502.665 4346.965 ;
        RECT 3503.095 4346.685 3503.375 4346.965 ;
        RECT 3503.805 4346.685 3504.085 4346.965 ;
        RECT 3504.515 4346.685 3504.795 4346.965 ;
        RECT 3505.225 4346.685 3505.505 4346.965 ;
        RECT 3505.935 4346.685 3506.215 4346.965 ;
        RECT 3506.645 4346.685 3506.925 4346.965 ;
        RECT 3507.355 4346.685 3507.635 4346.965 ;
        RECT 3508.065 4346.685 3508.345 4346.965 ;
        RECT 3508.775 4346.685 3509.055 4346.965 ;
        RECT 3509.485 4346.685 3509.765 4346.965 ;
        RECT 369.275 4345.955 369.555 4346.235 ;
        RECT 369.985 4345.955 370.265 4346.235 ;
        RECT 370.695 4345.955 370.975 4346.235 ;
        RECT 371.405 4345.955 371.685 4346.235 ;
        RECT 372.115 4345.955 372.395 4346.235 ;
        RECT 372.825 4345.955 373.105 4346.235 ;
        RECT 373.535 4345.955 373.815 4346.235 ;
        RECT 374.245 4345.955 374.525 4346.235 ;
        RECT 374.955 4345.955 375.235 4346.235 ;
        RECT 375.665 4345.955 375.945 4346.235 ;
        RECT 376.375 4345.955 376.655 4346.235 ;
        RECT 377.085 4345.955 377.365 4346.235 ;
        RECT 377.795 4345.955 378.075 4346.235 ;
        RECT 378.505 4345.955 378.785 4346.235 ;
        RECT 3500.255 4345.975 3500.535 4346.255 ;
        RECT 3500.965 4345.975 3501.245 4346.255 ;
        RECT 3501.675 4345.975 3501.955 4346.255 ;
        RECT 3502.385 4345.975 3502.665 4346.255 ;
        RECT 3503.095 4345.975 3503.375 4346.255 ;
        RECT 3503.805 4345.975 3504.085 4346.255 ;
        RECT 3504.515 4345.975 3504.795 4346.255 ;
        RECT 3505.225 4345.975 3505.505 4346.255 ;
        RECT 3505.935 4345.975 3506.215 4346.255 ;
        RECT 3506.645 4345.975 3506.925 4346.255 ;
        RECT 3507.355 4345.975 3507.635 4346.255 ;
        RECT 3508.065 4345.975 3508.345 4346.255 ;
        RECT 3508.775 4345.975 3509.055 4346.255 ;
        RECT 3509.485 4345.975 3509.765 4346.255 ;
        RECT 3500.255 4345.265 3500.535 4345.545 ;
        RECT 3500.965 4345.265 3501.245 4345.545 ;
        RECT 3501.675 4345.265 3501.955 4345.545 ;
        RECT 3502.385 4345.265 3502.665 4345.545 ;
        RECT 3503.095 4345.265 3503.375 4345.545 ;
        RECT 3503.805 4345.265 3504.085 4345.545 ;
        RECT 3504.515 4345.265 3504.795 4345.545 ;
        RECT 3505.225 4345.265 3505.505 4345.545 ;
        RECT 3505.935 4345.265 3506.215 4345.545 ;
        RECT 3506.645 4345.265 3506.925 4345.545 ;
        RECT 3507.355 4345.265 3507.635 4345.545 ;
        RECT 3508.065 4345.265 3508.345 4345.545 ;
        RECT 3508.775 4345.265 3509.055 4345.545 ;
        RECT 3509.485 4345.265 3509.765 4345.545 ;
        RECT 3500.255 4344.555 3500.535 4344.835 ;
        RECT 3500.965 4344.555 3501.245 4344.835 ;
        RECT 3501.675 4344.555 3501.955 4344.835 ;
        RECT 3502.385 4344.555 3502.665 4344.835 ;
        RECT 3503.095 4344.555 3503.375 4344.835 ;
        RECT 3503.805 4344.555 3504.085 4344.835 ;
        RECT 3504.515 4344.555 3504.795 4344.835 ;
        RECT 3505.225 4344.555 3505.505 4344.835 ;
        RECT 3505.935 4344.555 3506.215 4344.835 ;
        RECT 3506.645 4344.555 3506.925 4344.835 ;
        RECT 3507.355 4344.555 3507.635 4344.835 ;
        RECT 3508.065 4344.555 3508.345 4344.835 ;
        RECT 3508.775 4344.555 3509.055 4344.835 ;
        RECT 3509.485 4344.555 3509.765 4344.835 ;
        RECT 3500.255 4343.845 3500.535 4344.125 ;
        RECT 3500.965 4343.845 3501.245 4344.125 ;
        RECT 3501.675 4343.845 3501.955 4344.125 ;
        RECT 3502.385 4343.845 3502.665 4344.125 ;
        RECT 3503.095 4343.845 3503.375 4344.125 ;
        RECT 3503.805 4343.845 3504.085 4344.125 ;
        RECT 3504.515 4343.845 3504.795 4344.125 ;
        RECT 3505.225 4343.845 3505.505 4344.125 ;
        RECT 3505.935 4343.845 3506.215 4344.125 ;
        RECT 3506.645 4343.845 3506.925 4344.125 ;
        RECT 3507.355 4343.845 3507.635 4344.125 ;
        RECT 3508.065 4343.845 3508.345 4344.125 ;
        RECT 3508.775 4343.845 3509.055 4344.125 ;
        RECT 3509.485 4343.845 3509.765 4344.125 ;
        RECT 369.275 4343.335 369.555 4343.615 ;
        RECT 369.985 4343.335 370.265 4343.615 ;
        RECT 370.695 4343.335 370.975 4343.615 ;
        RECT 371.405 4343.335 371.685 4343.615 ;
        RECT 372.115 4343.335 372.395 4343.615 ;
        RECT 372.825 4343.335 373.105 4343.615 ;
        RECT 373.535 4343.335 373.815 4343.615 ;
        RECT 374.245 4343.335 374.525 4343.615 ;
        RECT 374.955 4343.335 375.235 4343.615 ;
        RECT 375.665 4343.335 375.945 4343.615 ;
        RECT 376.375 4343.335 376.655 4343.615 ;
        RECT 377.085 4343.335 377.365 4343.615 ;
        RECT 377.795 4343.335 378.075 4343.615 ;
        RECT 378.505 4343.335 378.785 4343.615 ;
        RECT 3500.255 4343.135 3500.535 4343.415 ;
        RECT 3500.965 4343.135 3501.245 4343.415 ;
        RECT 3501.675 4343.135 3501.955 4343.415 ;
        RECT 3502.385 4343.135 3502.665 4343.415 ;
        RECT 3503.095 4343.135 3503.375 4343.415 ;
        RECT 3503.805 4343.135 3504.085 4343.415 ;
        RECT 3504.515 4343.135 3504.795 4343.415 ;
        RECT 3505.225 4343.135 3505.505 4343.415 ;
        RECT 3505.935 4343.135 3506.215 4343.415 ;
        RECT 3506.645 4343.135 3506.925 4343.415 ;
        RECT 3507.355 4343.135 3507.635 4343.415 ;
        RECT 3508.065 4343.135 3508.345 4343.415 ;
        RECT 3508.775 4343.135 3509.055 4343.415 ;
        RECT 3509.485 4343.135 3509.765 4343.415 ;
        RECT 369.275 4342.625 369.555 4342.905 ;
        RECT 369.985 4342.625 370.265 4342.905 ;
        RECT 370.695 4342.625 370.975 4342.905 ;
        RECT 371.405 4342.625 371.685 4342.905 ;
        RECT 372.115 4342.625 372.395 4342.905 ;
        RECT 372.825 4342.625 373.105 4342.905 ;
        RECT 373.535 4342.625 373.815 4342.905 ;
        RECT 374.245 4342.625 374.525 4342.905 ;
        RECT 374.955 4342.625 375.235 4342.905 ;
        RECT 375.665 4342.625 375.945 4342.905 ;
        RECT 376.375 4342.625 376.655 4342.905 ;
        RECT 377.085 4342.625 377.365 4342.905 ;
        RECT 377.795 4342.625 378.075 4342.905 ;
        RECT 378.505 4342.625 378.785 4342.905 ;
        RECT 3500.255 4342.425 3500.535 4342.705 ;
        RECT 3500.965 4342.425 3501.245 4342.705 ;
        RECT 3501.675 4342.425 3501.955 4342.705 ;
        RECT 3502.385 4342.425 3502.665 4342.705 ;
        RECT 3503.095 4342.425 3503.375 4342.705 ;
        RECT 3503.805 4342.425 3504.085 4342.705 ;
        RECT 3504.515 4342.425 3504.795 4342.705 ;
        RECT 3505.225 4342.425 3505.505 4342.705 ;
        RECT 3505.935 4342.425 3506.215 4342.705 ;
        RECT 3506.645 4342.425 3506.925 4342.705 ;
        RECT 3507.355 4342.425 3507.635 4342.705 ;
        RECT 3508.065 4342.425 3508.345 4342.705 ;
        RECT 3508.775 4342.425 3509.055 4342.705 ;
        RECT 3509.485 4342.425 3509.765 4342.705 ;
        RECT 369.275 4341.915 369.555 4342.195 ;
        RECT 369.985 4341.915 370.265 4342.195 ;
        RECT 370.695 4341.915 370.975 4342.195 ;
        RECT 371.405 4341.915 371.685 4342.195 ;
        RECT 372.115 4341.915 372.395 4342.195 ;
        RECT 372.825 4341.915 373.105 4342.195 ;
        RECT 373.535 4341.915 373.815 4342.195 ;
        RECT 374.245 4341.915 374.525 4342.195 ;
        RECT 374.955 4341.915 375.235 4342.195 ;
        RECT 375.665 4341.915 375.945 4342.195 ;
        RECT 376.375 4341.915 376.655 4342.195 ;
        RECT 377.085 4341.915 377.365 4342.195 ;
        RECT 377.795 4341.915 378.075 4342.195 ;
        RECT 378.505 4341.915 378.785 4342.195 ;
        RECT 3500.255 4341.715 3500.535 4341.995 ;
        RECT 3500.965 4341.715 3501.245 4341.995 ;
        RECT 3501.675 4341.715 3501.955 4341.995 ;
        RECT 3502.385 4341.715 3502.665 4341.995 ;
        RECT 3503.095 4341.715 3503.375 4341.995 ;
        RECT 3503.805 4341.715 3504.085 4341.995 ;
        RECT 3504.515 4341.715 3504.795 4341.995 ;
        RECT 3505.225 4341.715 3505.505 4341.995 ;
        RECT 3505.935 4341.715 3506.215 4341.995 ;
        RECT 3506.645 4341.715 3506.925 4341.995 ;
        RECT 3507.355 4341.715 3507.635 4341.995 ;
        RECT 3508.065 4341.715 3508.345 4341.995 ;
        RECT 3508.775 4341.715 3509.055 4341.995 ;
        RECT 3509.485 4341.715 3509.765 4341.995 ;
        RECT 369.275 4341.205 369.555 4341.485 ;
        RECT 369.985 4341.205 370.265 4341.485 ;
        RECT 370.695 4341.205 370.975 4341.485 ;
        RECT 371.405 4341.205 371.685 4341.485 ;
        RECT 372.115 4341.205 372.395 4341.485 ;
        RECT 372.825 4341.205 373.105 4341.485 ;
        RECT 373.535 4341.205 373.815 4341.485 ;
        RECT 374.245 4341.205 374.525 4341.485 ;
        RECT 374.955 4341.205 375.235 4341.485 ;
        RECT 375.665 4341.205 375.945 4341.485 ;
        RECT 376.375 4341.205 376.655 4341.485 ;
        RECT 377.085 4341.205 377.365 4341.485 ;
        RECT 377.795 4341.205 378.075 4341.485 ;
        RECT 378.505 4341.205 378.785 4341.485 ;
        RECT 3500.255 4341.005 3500.535 4341.285 ;
        RECT 3500.965 4341.005 3501.245 4341.285 ;
        RECT 3501.675 4341.005 3501.955 4341.285 ;
        RECT 3502.385 4341.005 3502.665 4341.285 ;
        RECT 3503.095 4341.005 3503.375 4341.285 ;
        RECT 3503.805 4341.005 3504.085 4341.285 ;
        RECT 3504.515 4341.005 3504.795 4341.285 ;
        RECT 3505.225 4341.005 3505.505 4341.285 ;
        RECT 3505.935 4341.005 3506.215 4341.285 ;
        RECT 3506.645 4341.005 3506.925 4341.285 ;
        RECT 3507.355 4341.005 3507.635 4341.285 ;
        RECT 3508.065 4341.005 3508.345 4341.285 ;
        RECT 3508.775 4341.005 3509.055 4341.285 ;
        RECT 3509.485 4341.005 3509.765 4341.285 ;
        RECT 369.275 4340.495 369.555 4340.775 ;
        RECT 369.985 4340.495 370.265 4340.775 ;
        RECT 370.695 4340.495 370.975 4340.775 ;
        RECT 371.405 4340.495 371.685 4340.775 ;
        RECT 372.115 4340.495 372.395 4340.775 ;
        RECT 372.825 4340.495 373.105 4340.775 ;
        RECT 373.535 4340.495 373.815 4340.775 ;
        RECT 374.245 4340.495 374.525 4340.775 ;
        RECT 374.955 4340.495 375.235 4340.775 ;
        RECT 375.665 4340.495 375.945 4340.775 ;
        RECT 376.375 4340.495 376.655 4340.775 ;
        RECT 377.085 4340.495 377.365 4340.775 ;
        RECT 377.795 4340.495 378.075 4340.775 ;
        RECT 378.505 4340.495 378.785 4340.775 ;
        RECT 369.275 4339.785 369.555 4340.065 ;
        RECT 369.985 4339.785 370.265 4340.065 ;
        RECT 370.695 4339.785 370.975 4340.065 ;
        RECT 371.405 4339.785 371.685 4340.065 ;
        RECT 372.115 4339.785 372.395 4340.065 ;
        RECT 372.825 4339.785 373.105 4340.065 ;
        RECT 373.535 4339.785 373.815 4340.065 ;
        RECT 374.245 4339.785 374.525 4340.065 ;
        RECT 374.955 4339.785 375.235 4340.065 ;
        RECT 375.665 4339.785 375.945 4340.065 ;
        RECT 376.375 4339.785 376.655 4340.065 ;
        RECT 377.085 4339.785 377.365 4340.065 ;
        RECT 377.795 4339.785 378.075 4340.065 ;
        RECT 378.505 4339.785 378.785 4340.065 ;
        RECT 369.275 4339.075 369.555 4339.355 ;
        RECT 369.985 4339.075 370.265 4339.355 ;
        RECT 370.695 4339.075 370.975 4339.355 ;
        RECT 371.405 4339.075 371.685 4339.355 ;
        RECT 372.115 4339.075 372.395 4339.355 ;
        RECT 372.825 4339.075 373.105 4339.355 ;
        RECT 373.535 4339.075 373.815 4339.355 ;
        RECT 374.245 4339.075 374.525 4339.355 ;
        RECT 374.955 4339.075 375.235 4339.355 ;
        RECT 375.665 4339.075 375.945 4339.355 ;
        RECT 376.375 4339.075 376.655 4339.355 ;
        RECT 377.085 4339.075 377.365 4339.355 ;
        RECT 377.795 4339.075 378.075 4339.355 ;
        RECT 378.505 4339.075 378.785 4339.355 ;
        RECT 369.275 4338.365 369.555 4338.645 ;
        RECT 369.985 4338.365 370.265 4338.645 ;
        RECT 370.695 4338.365 370.975 4338.645 ;
        RECT 371.405 4338.365 371.685 4338.645 ;
        RECT 372.115 4338.365 372.395 4338.645 ;
        RECT 372.825 4338.365 373.105 4338.645 ;
        RECT 373.535 4338.365 373.815 4338.645 ;
        RECT 374.245 4338.365 374.525 4338.645 ;
        RECT 374.955 4338.365 375.235 4338.645 ;
        RECT 375.665 4338.365 375.945 4338.645 ;
        RECT 376.375 4338.365 376.655 4338.645 ;
        RECT 377.085 4338.365 377.365 4338.645 ;
        RECT 377.795 4338.365 378.075 4338.645 ;
        RECT 378.505 4338.365 378.785 4338.645 ;
        RECT 3500.255 4338.385 3500.535 4338.665 ;
        RECT 3500.965 4338.385 3501.245 4338.665 ;
        RECT 3501.675 4338.385 3501.955 4338.665 ;
        RECT 3502.385 4338.385 3502.665 4338.665 ;
        RECT 3503.095 4338.385 3503.375 4338.665 ;
        RECT 3503.805 4338.385 3504.085 4338.665 ;
        RECT 3504.515 4338.385 3504.795 4338.665 ;
        RECT 3505.225 4338.385 3505.505 4338.665 ;
        RECT 3505.935 4338.385 3506.215 4338.665 ;
        RECT 3506.645 4338.385 3506.925 4338.665 ;
        RECT 3507.355 4338.385 3507.635 4338.665 ;
        RECT 3508.065 4338.385 3508.345 4338.665 ;
        RECT 3508.775 4338.385 3509.055 4338.665 ;
        RECT 3509.485 4338.385 3509.765 4338.665 ;
        RECT 369.275 4337.655 369.555 4337.935 ;
        RECT 369.985 4337.655 370.265 4337.935 ;
        RECT 370.695 4337.655 370.975 4337.935 ;
        RECT 371.405 4337.655 371.685 4337.935 ;
        RECT 372.115 4337.655 372.395 4337.935 ;
        RECT 372.825 4337.655 373.105 4337.935 ;
        RECT 373.535 4337.655 373.815 4337.935 ;
        RECT 374.245 4337.655 374.525 4337.935 ;
        RECT 374.955 4337.655 375.235 4337.935 ;
        RECT 375.665 4337.655 375.945 4337.935 ;
        RECT 376.375 4337.655 376.655 4337.935 ;
        RECT 377.085 4337.655 377.365 4337.935 ;
        RECT 377.795 4337.655 378.075 4337.935 ;
        RECT 378.505 4337.655 378.785 4337.935 ;
        RECT 3500.255 4337.675 3500.535 4337.955 ;
        RECT 3500.965 4337.675 3501.245 4337.955 ;
        RECT 3501.675 4337.675 3501.955 4337.955 ;
        RECT 3502.385 4337.675 3502.665 4337.955 ;
        RECT 3503.095 4337.675 3503.375 4337.955 ;
        RECT 3503.805 4337.675 3504.085 4337.955 ;
        RECT 3504.515 4337.675 3504.795 4337.955 ;
        RECT 3505.225 4337.675 3505.505 4337.955 ;
        RECT 3505.935 4337.675 3506.215 4337.955 ;
        RECT 3506.645 4337.675 3506.925 4337.955 ;
        RECT 3507.355 4337.675 3507.635 4337.955 ;
        RECT 3508.065 4337.675 3508.345 4337.955 ;
        RECT 3508.775 4337.675 3509.055 4337.955 ;
        RECT 3509.485 4337.675 3509.765 4337.955 ;
        RECT 369.275 4336.945 369.555 4337.225 ;
        RECT 369.985 4336.945 370.265 4337.225 ;
        RECT 370.695 4336.945 370.975 4337.225 ;
        RECT 371.405 4336.945 371.685 4337.225 ;
        RECT 372.115 4336.945 372.395 4337.225 ;
        RECT 372.825 4336.945 373.105 4337.225 ;
        RECT 373.535 4336.945 373.815 4337.225 ;
        RECT 374.245 4336.945 374.525 4337.225 ;
        RECT 374.955 4336.945 375.235 4337.225 ;
        RECT 375.665 4336.945 375.945 4337.225 ;
        RECT 376.375 4336.945 376.655 4337.225 ;
        RECT 377.085 4336.945 377.365 4337.225 ;
        RECT 377.795 4336.945 378.075 4337.225 ;
        RECT 378.505 4336.945 378.785 4337.225 ;
        RECT 3500.255 4336.965 3500.535 4337.245 ;
        RECT 3500.965 4336.965 3501.245 4337.245 ;
        RECT 3501.675 4336.965 3501.955 4337.245 ;
        RECT 3502.385 4336.965 3502.665 4337.245 ;
        RECT 3503.095 4336.965 3503.375 4337.245 ;
        RECT 3503.805 4336.965 3504.085 4337.245 ;
        RECT 3504.515 4336.965 3504.795 4337.245 ;
        RECT 3505.225 4336.965 3505.505 4337.245 ;
        RECT 3505.935 4336.965 3506.215 4337.245 ;
        RECT 3506.645 4336.965 3506.925 4337.245 ;
        RECT 3507.355 4336.965 3507.635 4337.245 ;
        RECT 3508.065 4336.965 3508.345 4337.245 ;
        RECT 3508.775 4336.965 3509.055 4337.245 ;
        RECT 3509.485 4336.965 3509.765 4337.245 ;
        RECT 369.275 4336.235 369.555 4336.515 ;
        RECT 369.985 4336.235 370.265 4336.515 ;
        RECT 370.695 4336.235 370.975 4336.515 ;
        RECT 371.405 4336.235 371.685 4336.515 ;
        RECT 372.115 4336.235 372.395 4336.515 ;
        RECT 372.825 4336.235 373.105 4336.515 ;
        RECT 373.535 4336.235 373.815 4336.515 ;
        RECT 374.245 4336.235 374.525 4336.515 ;
        RECT 374.955 4336.235 375.235 4336.515 ;
        RECT 375.665 4336.235 375.945 4336.515 ;
        RECT 376.375 4336.235 376.655 4336.515 ;
        RECT 377.085 4336.235 377.365 4336.515 ;
        RECT 377.795 4336.235 378.075 4336.515 ;
        RECT 378.505 4336.235 378.785 4336.515 ;
        RECT 3500.255 4336.255 3500.535 4336.535 ;
        RECT 3500.965 4336.255 3501.245 4336.535 ;
        RECT 3501.675 4336.255 3501.955 4336.535 ;
        RECT 3502.385 4336.255 3502.665 4336.535 ;
        RECT 3503.095 4336.255 3503.375 4336.535 ;
        RECT 3503.805 4336.255 3504.085 4336.535 ;
        RECT 3504.515 4336.255 3504.795 4336.535 ;
        RECT 3505.225 4336.255 3505.505 4336.535 ;
        RECT 3505.935 4336.255 3506.215 4336.535 ;
        RECT 3506.645 4336.255 3506.925 4336.535 ;
        RECT 3507.355 4336.255 3507.635 4336.535 ;
        RECT 3508.065 4336.255 3508.345 4336.535 ;
        RECT 3508.775 4336.255 3509.055 4336.535 ;
        RECT 3509.485 4336.255 3509.765 4336.535 ;
        RECT 369.275 4335.525 369.555 4335.805 ;
        RECT 369.985 4335.525 370.265 4335.805 ;
        RECT 370.695 4335.525 370.975 4335.805 ;
        RECT 371.405 4335.525 371.685 4335.805 ;
        RECT 372.115 4335.525 372.395 4335.805 ;
        RECT 372.825 4335.525 373.105 4335.805 ;
        RECT 373.535 4335.525 373.815 4335.805 ;
        RECT 374.245 4335.525 374.525 4335.805 ;
        RECT 374.955 4335.525 375.235 4335.805 ;
        RECT 375.665 4335.525 375.945 4335.805 ;
        RECT 376.375 4335.525 376.655 4335.805 ;
        RECT 377.085 4335.525 377.365 4335.805 ;
        RECT 377.795 4335.525 378.075 4335.805 ;
        RECT 378.505 4335.525 378.785 4335.805 ;
        RECT 3500.255 4335.545 3500.535 4335.825 ;
        RECT 3500.965 4335.545 3501.245 4335.825 ;
        RECT 3501.675 4335.545 3501.955 4335.825 ;
        RECT 3502.385 4335.545 3502.665 4335.825 ;
        RECT 3503.095 4335.545 3503.375 4335.825 ;
        RECT 3503.805 4335.545 3504.085 4335.825 ;
        RECT 3504.515 4335.545 3504.795 4335.825 ;
        RECT 3505.225 4335.545 3505.505 4335.825 ;
        RECT 3505.935 4335.545 3506.215 4335.825 ;
        RECT 3506.645 4335.545 3506.925 4335.825 ;
        RECT 3507.355 4335.545 3507.635 4335.825 ;
        RECT 3508.065 4335.545 3508.345 4335.825 ;
        RECT 3508.775 4335.545 3509.055 4335.825 ;
        RECT 3509.485 4335.545 3509.765 4335.825 ;
        RECT 369.275 4334.815 369.555 4335.095 ;
        RECT 369.985 4334.815 370.265 4335.095 ;
        RECT 370.695 4334.815 370.975 4335.095 ;
        RECT 371.405 4334.815 371.685 4335.095 ;
        RECT 372.115 4334.815 372.395 4335.095 ;
        RECT 372.825 4334.815 373.105 4335.095 ;
        RECT 373.535 4334.815 373.815 4335.095 ;
        RECT 374.245 4334.815 374.525 4335.095 ;
        RECT 374.955 4334.815 375.235 4335.095 ;
        RECT 375.665 4334.815 375.945 4335.095 ;
        RECT 376.375 4334.815 376.655 4335.095 ;
        RECT 377.085 4334.815 377.365 4335.095 ;
        RECT 377.795 4334.815 378.075 4335.095 ;
        RECT 378.505 4334.815 378.785 4335.095 ;
        RECT 3500.255 4334.835 3500.535 4335.115 ;
        RECT 3500.965 4334.835 3501.245 4335.115 ;
        RECT 3501.675 4334.835 3501.955 4335.115 ;
        RECT 3502.385 4334.835 3502.665 4335.115 ;
        RECT 3503.095 4334.835 3503.375 4335.115 ;
        RECT 3503.805 4334.835 3504.085 4335.115 ;
        RECT 3504.515 4334.835 3504.795 4335.115 ;
        RECT 3505.225 4334.835 3505.505 4335.115 ;
        RECT 3505.935 4334.835 3506.215 4335.115 ;
        RECT 3506.645 4334.835 3506.925 4335.115 ;
        RECT 3507.355 4334.835 3507.635 4335.115 ;
        RECT 3508.065 4334.835 3508.345 4335.115 ;
        RECT 3508.775 4334.835 3509.055 4335.115 ;
        RECT 3509.485 4334.835 3509.765 4335.115 ;
        RECT 369.275 4334.105 369.555 4334.385 ;
        RECT 369.985 4334.105 370.265 4334.385 ;
        RECT 370.695 4334.105 370.975 4334.385 ;
        RECT 371.405 4334.105 371.685 4334.385 ;
        RECT 372.115 4334.105 372.395 4334.385 ;
        RECT 372.825 4334.105 373.105 4334.385 ;
        RECT 373.535 4334.105 373.815 4334.385 ;
        RECT 374.245 4334.105 374.525 4334.385 ;
        RECT 374.955 4334.105 375.235 4334.385 ;
        RECT 375.665 4334.105 375.945 4334.385 ;
        RECT 376.375 4334.105 376.655 4334.385 ;
        RECT 377.085 4334.105 377.365 4334.385 ;
        RECT 377.795 4334.105 378.075 4334.385 ;
        RECT 378.505 4334.105 378.785 4334.385 ;
        RECT 3500.255 4334.125 3500.535 4334.405 ;
        RECT 3500.965 4334.125 3501.245 4334.405 ;
        RECT 3501.675 4334.125 3501.955 4334.405 ;
        RECT 3502.385 4334.125 3502.665 4334.405 ;
        RECT 3503.095 4334.125 3503.375 4334.405 ;
        RECT 3503.805 4334.125 3504.085 4334.405 ;
        RECT 3504.515 4334.125 3504.795 4334.405 ;
        RECT 3505.225 4334.125 3505.505 4334.405 ;
        RECT 3505.935 4334.125 3506.215 4334.405 ;
        RECT 3506.645 4334.125 3506.925 4334.405 ;
        RECT 3507.355 4334.125 3507.635 4334.405 ;
        RECT 3508.065 4334.125 3508.345 4334.405 ;
        RECT 3508.775 4334.125 3509.055 4334.405 ;
        RECT 3509.485 4334.125 3509.765 4334.405 ;
        RECT 3500.255 4333.415 3500.535 4333.695 ;
        RECT 3500.965 4333.415 3501.245 4333.695 ;
        RECT 3501.675 4333.415 3501.955 4333.695 ;
        RECT 3502.385 4333.415 3502.665 4333.695 ;
        RECT 3503.095 4333.415 3503.375 4333.695 ;
        RECT 3503.805 4333.415 3504.085 4333.695 ;
        RECT 3504.515 4333.415 3504.795 4333.695 ;
        RECT 3505.225 4333.415 3505.505 4333.695 ;
        RECT 3505.935 4333.415 3506.215 4333.695 ;
        RECT 3506.645 4333.415 3506.925 4333.695 ;
        RECT 3507.355 4333.415 3507.635 4333.695 ;
        RECT 3508.065 4333.415 3508.345 4333.695 ;
        RECT 3508.775 4333.415 3509.055 4333.695 ;
        RECT 3509.485 4333.415 3509.765 4333.695 ;
        RECT 3500.255 4332.705 3500.535 4332.985 ;
        RECT 3500.965 4332.705 3501.245 4332.985 ;
        RECT 3501.675 4332.705 3501.955 4332.985 ;
        RECT 3502.385 4332.705 3502.665 4332.985 ;
        RECT 3503.095 4332.705 3503.375 4332.985 ;
        RECT 3503.805 4332.705 3504.085 4332.985 ;
        RECT 3504.515 4332.705 3504.795 4332.985 ;
        RECT 3505.225 4332.705 3505.505 4332.985 ;
        RECT 3505.935 4332.705 3506.215 4332.985 ;
        RECT 3506.645 4332.705 3506.925 4332.985 ;
        RECT 3507.355 4332.705 3507.635 4332.985 ;
        RECT 3508.065 4332.705 3508.345 4332.985 ;
        RECT 3508.775 4332.705 3509.055 4332.985 ;
        RECT 3509.485 4332.705 3509.765 4332.985 ;
        RECT 3500.255 4331.995 3500.535 4332.275 ;
        RECT 3500.965 4331.995 3501.245 4332.275 ;
        RECT 3501.675 4331.995 3501.955 4332.275 ;
        RECT 3502.385 4331.995 3502.665 4332.275 ;
        RECT 3503.095 4331.995 3503.375 4332.275 ;
        RECT 3503.805 4331.995 3504.085 4332.275 ;
        RECT 3504.515 4331.995 3504.795 4332.275 ;
        RECT 3505.225 4331.995 3505.505 4332.275 ;
        RECT 3505.935 4331.995 3506.215 4332.275 ;
        RECT 3506.645 4331.995 3506.925 4332.275 ;
        RECT 3507.355 4331.995 3507.635 4332.275 ;
        RECT 3508.065 4331.995 3508.345 4332.275 ;
        RECT 3508.775 4331.995 3509.055 4332.275 ;
        RECT 3509.485 4331.995 3509.765 4332.275 ;
        RECT 3500.255 4331.285 3500.535 4331.565 ;
        RECT 3500.965 4331.285 3501.245 4331.565 ;
        RECT 3501.675 4331.285 3501.955 4331.565 ;
        RECT 3502.385 4331.285 3502.665 4331.565 ;
        RECT 3503.095 4331.285 3503.375 4331.565 ;
        RECT 3503.805 4331.285 3504.085 4331.565 ;
        RECT 3504.515 4331.285 3504.795 4331.565 ;
        RECT 3505.225 4331.285 3505.505 4331.565 ;
        RECT 3505.935 4331.285 3506.215 4331.565 ;
        RECT 3506.645 4331.285 3506.925 4331.565 ;
        RECT 3507.355 4331.285 3507.635 4331.565 ;
        RECT 3508.065 4331.285 3508.345 4331.565 ;
        RECT 3508.775 4331.285 3509.055 4331.565 ;
        RECT 3509.485 4331.285 3509.765 4331.565 ;
        RECT 3500.255 4330.575 3500.535 4330.855 ;
        RECT 3500.965 4330.575 3501.245 4330.855 ;
        RECT 3501.675 4330.575 3501.955 4330.855 ;
        RECT 3502.385 4330.575 3502.665 4330.855 ;
        RECT 3503.095 4330.575 3503.375 4330.855 ;
        RECT 3503.805 4330.575 3504.085 4330.855 ;
        RECT 3504.515 4330.575 3504.795 4330.855 ;
        RECT 3505.225 4330.575 3505.505 4330.855 ;
        RECT 3505.935 4330.575 3506.215 4330.855 ;
        RECT 3506.645 4330.575 3506.925 4330.855 ;
        RECT 3507.355 4330.575 3507.635 4330.855 ;
        RECT 3508.065 4330.575 3508.345 4330.855 ;
        RECT 3508.775 4330.575 3509.055 4330.855 ;
        RECT 3509.485 4330.575 3509.765 4330.855 ;
        RECT 369.330 4330.190 369.610 4330.470 ;
        RECT 370.040 4330.190 370.320 4330.470 ;
        RECT 370.750 4330.190 371.030 4330.470 ;
        RECT 371.460 4330.190 371.740 4330.470 ;
        RECT 372.170 4330.190 372.450 4330.470 ;
        RECT 372.880 4330.190 373.160 4330.470 ;
        RECT 373.590 4330.190 373.870 4330.470 ;
        RECT 374.300 4330.190 374.580 4330.470 ;
        RECT 375.010 4330.190 375.290 4330.470 ;
        RECT 375.720 4330.190 376.000 4330.470 ;
        RECT 376.430 4330.190 376.710 4330.470 ;
        RECT 377.140 4330.190 377.420 4330.470 ;
        RECT 377.850 4330.190 378.130 4330.470 ;
        RECT 378.560 4330.190 378.840 4330.470 ;
        RECT 3500.255 4329.865 3500.535 4330.145 ;
        RECT 3500.965 4329.865 3501.245 4330.145 ;
        RECT 3501.675 4329.865 3501.955 4330.145 ;
        RECT 3502.385 4329.865 3502.665 4330.145 ;
        RECT 3503.095 4329.865 3503.375 4330.145 ;
        RECT 3503.805 4329.865 3504.085 4330.145 ;
        RECT 3504.515 4329.865 3504.795 4330.145 ;
        RECT 3505.225 4329.865 3505.505 4330.145 ;
        RECT 3505.935 4329.865 3506.215 4330.145 ;
        RECT 3506.645 4329.865 3506.925 4330.145 ;
        RECT 3507.355 4329.865 3507.635 4330.145 ;
        RECT 3508.065 4329.865 3508.345 4330.145 ;
        RECT 3508.775 4329.865 3509.055 4330.145 ;
        RECT 3509.485 4329.865 3509.765 4330.145 ;
        RECT 369.330 4329.480 369.610 4329.760 ;
        RECT 370.040 4329.480 370.320 4329.760 ;
        RECT 370.750 4329.480 371.030 4329.760 ;
        RECT 371.460 4329.480 371.740 4329.760 ;
        RECT 372.170 4329.480 372.450 4329.760 ;
        RECT 372.880 4329.480 373.160 4329.760 ;
        RECT 373.590 4329.480 373.870 4329.760 ;
        RECT 374.300 4329.480 374.580 4329.760 ;
        RECT 375.010 4329.480 375.290 4329.760 ;
        RECT 375.720 4329.480 376.000 4329.760 ;
        RECT 376.430 4329.480 376.710 4329.760 ;
        RECT 377.140 4329.480 377.420 4329.760 ;
        RECT 377.850 4329.480 378.130 4329.760 ;
        RECT 378.560 4329.480 378.840 4329.760 ;
        RECT 3500.255 4329.155 3500.535 4329.435 ;
        RECT 3500.965 4329.155 3501.245 4329.435 ;
        RECT 3501.675 4329.155 3501.955 4329.435 ;
        RECT 3502.385 4329.155 3502.665 4329.435 ;
        RECT 3503.095 4329.155 3503.375 4329.435 ;
        RECT 3503.805 4329.155 3504.085 4329.435 ;
        RECT 3504.515 4329.155 3504.795 4329.435 ;
        RECT 3505.225 4329.155 3505.505 4329.435 ;
        RECT 3505.935 4329.155 3506.215 4329.435 ;
        RECT 3506.645 4329.155 3506.925 4329.435 ;
        RECT 3507.355 4329.155 3507.635 4329.435 ;
        RECT 3508.065 4329.155 3508.345 4329.435 ;
        RECT 3508.775 4329.155 3509.055 4329.435 ;
        RECT 3509.485 4329.155 3509.765 4329.435 ;
        RECT 369.330 4328.770 369.610 4329.050 ;
        RECT 370.040 4328.770 370.320 4329.050 ;
        RECT 370.750 4328.770 371.030 4329.050 ;
        RECT 371.460 4328.770 371.740 4329.050 ;
        RECT 372.170 4328.770 372.450 4329.050 ;
        RECT 372.880 4328.770 373.160 4329.050 ;
        RECT 373.590 4328.770 373.870 4329.050 ;
        RECT 374.300 4328.770 374.580 4329.050 ;
        RECT 375.010 4328.770 375.290 4329.050 ;
        RECT 375.720 4328.770 376.000 4329.050 ;
        RECT 376.430 4328.770 376.710 4329.050 ;
        RECT 377.140 4328.770 377.420 4329.050 ;
        RECT 377.850 4328.770 378.130 4329.050 ;
        RECT 378.560 4328.770 378.840 4329.050 ;
        RECT 369.330 4328.060 369.610 4328.340 ;
        RECT 370.040 4328.060 370.320 4328.340 ;
        RECT 370.750 4328.060 371.030 4328.340 ;
        RECT 371.460 4328.060 371.740 4328.340 ;
        RECT 372.170 4328.060 372.450 4328.340 ;
        RECT 372.880 4328.060 373.160 4328.340 ;
        RECT 373.590 4328.060 373.870 4328.340 ;
        RECT 374.300 4328.060 374.580 4328.340 ;
        RECT 375.010 4328.060 375.290 4328.340 ;
        RECT 375.720 4328.060 376.000 4328.340 ;
        RECT 376.430 4328.060 376.710 4328.340 ;
        RECT 377.140 4328.060 377.420 4328.340 ;
        RECT 377.850 4328.060 378.130 4328.340 ;
        RECT 378.560 4328.060 378.840 4328.340 ;
        RECT 369.330 4327.350 369.610 4327.630 ;
        RECT 370.040 4327.350 370.320 4327.630 ;
        RECT 370.750 4327.350 371.030 4327.630 ;
        RECT 371.460 4327.350 371.740 4327.630 ;
        RECT 372.170 4327.350 372.450 4327.630 ;
        RECT 372.880 4327.350 373.160 4327.630 ;
        RECT 373.590 4327.350 373.870 4327.630 ;
        RECT 374.300 4327.350 374.580 4327.630 ;
        RECT 375.010 4327.350 375.290 4327.630 ;
        RECT 375.720 4327.350 376.000 4327.630 ;
        RECT 376.430 4327.350 376.710 4327.630 ;
        RECT 377.140 4327.350 377.420 4327.630 ;
        RECT 377.850 4327.350 378.130 4327.630 ;
        RECT 378.560 4327.350 378.840 4327.630 ;
        RECT 369.330 4326.640 369.610 4326.920 ;
        RECT 370.040 4326.640 370.320 4326.920 ;
        RECT 370.750 4326.640 371.030 4326.920 ;
        RECT 371.460 4326.640 371.740 4326.920 ;
        RECT 372.170 4326.640 372.450 4326.920 ;
        RECT 372.880 4326.640 373.160 4326.920 ;
        RECT 373.590 4326.640 373.870 4326.920 ;
        RECT 374.300 4326.640 374.580 4326.920 ;
        RECT 375.010 4326.640 375.290 4326.920 ;
        RECT 375.720 4326.640 376.000 4326.920 ;
        RECT 376.430 4326.640 376.710 4326.920 ;
        RECT 377.140 4326.640 377.420 4326.920 ;
        RECT 377.850 4326.640 378.130 4326.920 ;
        RECT 378.560 4326.640 378.840 4326.920 ;
        RECT 369.330 4325.930 369.610 4326.210 ;
        RECT 370.040 4325.930 370.320 4326.210 ;
        RECT 370.750 4325.930 371.030 4326.210 ;
        RECT 371.460 4325.930 371.740 4326.210 ;
        RECT 372.170 4325.930 372.450 4326.210 ;
        RECT 372.880 4325.930 373.160 4326.210 ;
        RECT 373.590 4325.930 373.870 4326.210 ;
        RECT 374.300 4325.930 374.580 4326.210 ;
        RECT 375.010 4325.930 375.290 4326.210 ;
        RECT 375.720 4325.930 376.000 4326.210 ;
        RECT 376.430 4325.930 376.710 4326.210 ;
        RECT 377.140 4325.930 377.420 4326.210 ;
        RECT 377.850 4325.930 378.130 4326.210 ;
        RECT 378.560 4325.930 378.840 4326.210 ;
        RECT 369.330 4325.220 369.610 4325.500 ;
        RECT 370.040 4325.220 370.320 4325.500 ;
        RECT 370.750 4325.220 371.030 4325.500 ;
        RECT 371.460 4325.220 371.740 4325.500 ;
        RECT 372.170 4325.220 372.450 4325.500 ;
        RECT 372.880 4325.220 373.160 4325.500 ;
        RECT 373.590 4325.220 373.870 4325.500 ;
        RECT 374.300 4325.220 374.580 4325.500 ;
        RECT 375.010 4325.220 375.290 4325.500 ;
        RECT 375.720 4325.220 376.000 4325.500 ;
        RECT 376.430 4325.220 376.710 4325.500 ;
        RECT 377.140 4325.220 377.420 4325.500 ;
        RECT 377.850 4325.220 378.130 4325.500 ;
        RECT 378.560 4325.220 378.840 4325.500 ;
        RECT 3500.200 4325.270 3500.480 4325.550 ;
        RECT 3500.910 4325.270 3501.190 4325.550 ;
        RECT 3501.620 4325.270 3501.900 4325.550 ;
        RECT 3502.330 4325.270 3502.610 4325.550 ;
        RECT 3503.040 4325.270 3503.320 4325.550 ;
        RECT 3503.750 4325.270 3504.030 4325.550 ;
        RECT 3504.460 4325.270 3504.740 4325.550 ;
        RECT 3505.170 4325.270 3505.450 4325.550 ;
        RECT 3505.880 4325.270 3506.160 4325.550 ;
        RECT 3506.590 4325.270 3506.870 4325.550 ;
        RECT 3507.300 4325.270 3507.580 4325.550 ;
        RECT 3508.010 4325.270 3508.290 4325.550 ;
        RECT 3508.720 4325.270 3509.000 4325.550 ;
        RECT 3509.430 4325.270 3509.710 4325.550 ;
        RECT 369.330 4324.510 369.610 4324.790 ;
        RECT 370.040 4324.510 370.320 4324.790 ;
        RECT 370.750 4324.510 371.030 4324.790 ;
        RECT 371.460 4324.510 371.740 4324.790 ;
        RECT 372.170 4324.510 372.450 4324.790 ;
        RECT 372.880 4324.510 373.160 4324.790 ;
        RECT 373.590 4324.510 373.870 4324.790 ;
        RECT 374.300 4324.510 374.580 4324.790 ;
        RECT 375.010 4324.510 375.290 4324.790 ;
        RECT 375.720 4324.510 376.000 4324.790 ;
        RECT 376.430 4324.510 376.710 4324.790 ;
        RECT 377.140 4324.510 377.420 4324.790 ;
        RECT 377.850 4324.510 378.130 4324.790 ;
        RECT 378.560 4324.510 378.840 4324.790 ;
        RECT 3500.200 4324.560 3500.480 4324.840 ;
        RECT 3500.910 4324.560 3501.190 4324.840 ;
        RECT 3501.620 4324.560 3501.900 4324.840 ;
        RECT 3502.330 4324.560 3502.610 4324.840 ;
        RECT 3503.040 4324.560 3503.320 4324.840 ;
        RECT 3503.750 4324.560 3504.030 4324.840 ;
        RECT 3504.460 4324.560 3504.740 4324.840 ;
        RECT 3505.170 4324.560 3505.450 4324.840 ;
        RECT 3505.880 4324.560 3506.160 4324.840 ;
        RECT 3506.590 4324.560 3506.870 4324.840 ;
        RECT 3507.300 4324.560 3507.580 4324.840 ;
        RECT 3508.010 4324.560 3508.290 4324.840 ;
        RECT 3508.720 4324.560 3509.000 4324.840 ;
        RECT 3509.430 4324.560 3509.710 4324.840 ;
        RECT 369.330 4323.800 369.610 4324.080 ;
        RECT 370.040 4323.800 370.320 4324.080 ;
        RECT 370.750 4323.800 371.030 4324.080 ;
        RECT 371.460 4323.800 371.740 4324.080 ;
        RECT 372.170 4323.800 372.450 4324.080 ;
        RECT 372.880 4323.800 373.160 4324.080 ;
        RECT 373.590 4323.800 373.870 4324.080 ;
        RECT 374.300 4323.800 374.580 4324.080 ;
        RECT 375.010 4323.800 375.290 4324.080 ;
        RECT 375.720 4323.800 376.000 4324.080 ;
        RECT 376.430 4323.800 376.710 4324.080 ;
        RECT 377.140 4323.800 377.420 4324.080 ;
        RECT 377.850 4323.800 378.130 4324.080 ;
        RECT 378.560 4323.800 378.840 4324.080 ;
        RECT 3500.200 4323.850 3500.480 4324.130 ;
        RECT 3500.910 4323.850 3501.190 4324.130 ;
        RECT 3501.620 4323.850 3501.900 4324.130 ;
        RECT 3502.330 4323.850 3502.610 4324.130 ;
        RECT 3503.040 4323.850 3503.320 4324.130 ;
        RECT 3503.750 4323.850 3504.030 4324.130 ;
        RECT 3504.460 4323.850 3504.740 4324.130 ;
        RECT 3505.170 4323.850 3505.450 4324.130 ;
        RECT 3505.880 4323.850 3506.160 4324.130 ;
        RECT 3506.590 4323.850 3506.870 4324.130 ;
        RECT 3507.300 4323.850 3507.580 4324.130 ;
        RECT 3508.010 4323.850 3508.290 4324.130 ;
        RECT 3508.720 4323.850 3509.000 4324.130 ;
        RECT 3509.430 4323.850 3509.710 4324.130 ;
        RECT 369.330 4323.090 369.610 4323.370 ;
        RECT 370.040 4323.090 370.320 4323.370 ;
        RECT 370.750 4323.090 371.030 4323.370 ;
        RECT 371.460 4323.090 371.740 4323.370 ;
        RECT 372.170 4323.090 372.450 4323.370 ;
        RECT 372.880 4323.090 373.160 4323.370 ;
        RECT 373.590 4323.090 373.870 4323.370 ;
        RECT 374.300 4323.090 374.580 4323.370 ;
        RECT 375.010 4323.090 375.290 4323.370 ;
        RECT 375.720 4323.090 376.000 4323.370 ;
        RECT 376.430 4323.090 376.710 4323.370 ;
        RECT 377.140 4323.090 377.420 4323.370 ;
        RECT 377.850 4323.090 378.130 4323.370 ;
        RECT 378.560 4323.090 378.840 4323.370 ;
        RECT 3500.200 4323.140 3500.480 4323.420 ;
        RECT 3500.910 4323.140 3501.190 4323.420 ;
        RECT 3501.620 4323.140 3501.900 4323.420 ;
        RECT 3502.330 4323.140 3502.610 4323.420 ;
        RECT 3503.040 4323.140 3503.320 4323.420 ;
        RECT 3503.750 4323.140 3504.030 4323.420 ;
        RECT 3504.460 4323.140 3504.740 4323.420 ;
        RECT 3505.170 4323.140 3505.450 4323.420 ;
        RECT 3505.880 4323.140 3506.160 4323.420 ;
        RECT 3506.590 4323.140 3506.870 4323.420 ;
        RECT 3507.300 4323.140 3507.580 4323.420 ;
        RECT 3508.010 4323.140 3508.290 4323.420 ;
        RECT 3508.720 4323.140 3509.000 4323.420 ;
        RECT 3509.430 4323.140 3509.710 4323.420 ;
        RECT 369.330 4322.380 369.610 4322.660 ;
        RECT 370.040 4322.380 370.320 4322.660 ;
        RECT 370.750 4322.380 371.030 4322.660 ;
        RECT 371.460 4322.380 371.740 4322.660 ;
        RECT 372.170 4322.380 372.450 4322.660 ;
        RECT 372.880 4322.380 373.160 4322.660 ;
        RECT 373.590 4322.380 373.870 4322.660 ;
        RECT 374.300 4322.380 374.580 4322.660 ;
        RECT 375.010 4322.380 375.290 4322.660 ;
        RECT 375.720 4322.380 376.000 4322.660 ;
        RECT 376.430 4322.380 376.710 4322.660 ;
        RECT 377.140 4322.380 377.420 4322.660 ;
        RECT 377.850 4322.380 378.130 4322.660 ;
        RECT 378.560 4322.380 378.840 4322.660 ;
        RECT 3500.200 4322.430 3500.480 4322.710 ;
        RECT 3500.910 4322.430 3501.190 4322.710 ;
        RECT 3501.620 4322.430 3501.900 4322.710 ;
        RECT 3502.330 4322.430 3502.610 4322.710 ;
        RECT 3503.040 4322.430 3503.320 4322.710 ;
        RECT 3503.750 4322.430 3504.030 4322.710 ;
        RECT 3504.460 4322.430 3504.740 4322.710 ;
        RECT 3505.170 4322.430 3505.450 4322.710 ;
        RECT 3505.880 4322.430 3506.160 4322.710 ;
        RECT 3506.590 4322.430 3506.870 4322.710 ;
        RECT 3507.300 4322.430 3507.580 4322.710 ;
        RECT 3508.010 4322.430 3508.290 4322.710 ;
        RECT 3508.720 4322.430 3509.000 4322.710 ;
        RECT 3509.430 4322.430 3509.710 4322.710 ;
        RECT 369.330 4321.670 369.610 4321.950 ;
        RECT 370.040 4321.670 370.320 4321.950 ;
        RECT 370.750 4321.670 371.030 4321.950 ;
        RECT 371.460 4321.670 371.740 4321.950 ;
        RECT 372.170 4321.670 372.450 4321.950 ;
        RECT 372.880 4321.670 373.160 4321.950 ;
        RECT 373.590 4321.670 373.870 4321.950 ;
        RECT 374.300 4321.670 374.580 4321.950 ;
        RECT 375.010 4321.670 375.290 4321.950 ;
        RECT 375.720 4321.670 376.000 4321.950 ;
        RECT 376.430 4321.670 376.710 4321.950 ;
        RECT 377.140 4321.670 377.420 4321.950 ;
        RECT 377.850 4321.670 378.130 4321.950 ;
        RECT 378.560 4321.670 378.840 4321.950 ;
        RECT 3500.200 4321.720 3500.480 4322.000 ;
        RECT 3500.910 4321.720 3501.190 4322.000 ;
        RECT 3501.620 4321.720 3501.900 4322.000 ;
        RECT 3502.330 4321.720 3502.610 4322.000 ;
        RECT 3503.040 4321.720 3503.320 4322.000 ;
        RECT 3503.750 4321.720 3504.030 4322.000 ;
        RECT 3504.460 4321.720 3504.740 4322.000 ;
        RECT 3505.170 4321.720 3505.450 4322.000 ;
        RECT 3505.880 4321.720 3506.160 4322.000 ;
        RECT 3506.590 4321.720 3506.870 4322.000 ;
        RECT 3507.300 4321.720 3507.580 4322.000 ;
        RECT 3508.010 4321.720 3508.290 4322.000 ;
        RECT 3508.720 4321.720 3509.000 4322.000 ;
        RECT 3509.430 4321.720 3509.710 4322.000 ;
        RECT 3500.200 4321.010 3500.480 4321.290 ;
        RECT 3500.910 4321.010 3501.190 4321.290 ;
        RECT 3501.620 4321.010 3501.900 4321.290 ;
        RECT 3502.330 4321.010 3502.610 4321.290 ;
        RECT 3503.040 4321.010 3503.320 4321.290 ;
        RECT 3503.750 4321.010 3504.030 4321.290 ;
        RECT 3504.460 4321.010 3504.740 4321.290 ;
        RECT 3505.170 4321.010 3505.450 4321.290 ;
        RECT 3505.880 4321.010 3506.160 4321.290 ;
        RECT 3506.590 4321.010 3506.870 4321.290 ;
        RECT 3507.300 4321.010 3507.580 4321.290 ;
        RECT 3508.010 4321.010 3508.290 4321.290 ;
        RECT 3508.720 4321.010 3509.000 4321.290 ;
        RECT 3509.430 4321.010 3509.710 4321.290 ;
        RECT 3500.200 4320.300 3500.480 4320.580 ;
        RECT 3500.910 4320.300 3501.190 4320.580 ;
        RECT 3501.620 4320.300 3501.900 4320.580 ;
        RECT 3502.330 4320.300 3502.610 4320.580 ;
        RECT 3503.040 4320.300 3503.320 4320.580 ;
        RECT 3503.750 4320.300 3504.030 4320.580 ;
        RECT 3504.460 4320.300 3504.740 4320.580 ;
        RECT 3505.170 4320.300 3505.450 4320.580 ;
        RECT 3505.880 4320.300 3506.160 4320.580 ;
        RECT 3506.590 4320.300 3506.870 4320.580 ;
        RECT 3507.300 4320.300 3507.580 4320.580 ;
        RECT 3508.010 4320.300 3508.290 4320.580 ;
        RECT 3508.720 4320.300 3509.000 4320.580 ;
        RECT 3509.430 4320.300 3509.710 4320.580 ;
        RECT 3500.200 4319.590 3500.480 4319.870 ;
        RECT 3500.910 4319.590 3501.190 4319.870 ;
        RECT 3501.620 4319.590 3501.900 4319.870 ;
        RECT 3502.330 4319.590 3502.610 4319.870 ;
        RECT 3503.040 4319.590 3503.320 4319.870 ;
        RECT 3503.750 4319.590 3504.030 4319.870 ;
        RECT 3504.460 4319.590 3504.740 4319.870 ;
        RECT 3505.170 4319.590 3505.450 4319.870 ;
        RECT 3505.880 4319.590 3506.160 4319.870 ;
        RECT 3506.590 4319.590 3506.870 4319.870 ;
        RECT 3507.300 4319.590 3507.580 4319.870 ;
        RECT 3508.010 4319.590 3508.290 4319.870 ;
        RECT 3508.720 4319.590 3509.000 4319.870 ;
        RECT 3509.430 4319.590 3509.710 4319.870 ;
        RECT 3500.200 4318.880 3500.480 4319.160 ;
        RECT 3500.910 4318.880 3501.190 4319.160 ;
        RECT 3501.620 4318.880 3501.900 4319.160 ;
        RECT 3502.330 4318.880 3502.610 4319.160 ;
        RECT 3503.040 4318.880 3503.320 4319.160 ;
        RECT 3503.750 4318.880 3504.030 4319.160 ;
        RECT 3504.460 4318.880 3504.740 4319.160 ;
        RECT 3505.170 4318.880 3505.450 4319.160 ;
        RECT 3505.880 4318.880 3506.160 4319.160 ;
        RECT 3506.590 4318.880 3506.870 4319.160 ;
        RECT 3507.300 4318.880 3507.580 4319.160 ;
        RECT 3508.010 4318.880 3508.290 4319.160 ;
        RECT 3508.720 4318.880 3509.000 4319.160 ;
        RECT 3509.430 4318.880 3509.710 4319.160 ;
        RECT 3500.200 4318.170 3500.480 4318.450 ;
        RECT 3500.910 4318.170 3501.190 4318.450 ;
        RECT 3501.620 4318.170 3501.900 4318.450 ;
        RECT 3502.330 4318.170 3502.610 4318.450 ;
        RECT 3503.040 4318.170 3503.320 4318.450 ;
        RECT 3503.750 4318.170 3504.030 4318.450 ;
        RECT 3504.460 4318.170 3504.740 4318.450 ;
        RECT 3505.170 4318.170 3505.450 4318.450 ;
        RECT 3505.880 4318.170 3506.160 4318.450 ;
        RECT 3506.590 4318.170 3506.870 4318.450 ;
        RECT 3507.300 4318.170 3507.580 4318.450 ;
        RECT 3508.010 4318.170 3508.290 4318.450 ;
        RECT 3508.720 4318.170 3509.000 4318.450 ;
        RECT 3509.430 4318.170 3509.710 4318.450 ;
        RECT 3500.200 4317.460 3500.480 4317.740 ;
        RECT 3500.910 4317.460 3501.190 4317.740 ;
        RECT 3501.620 4317.460 3501.900 4317.740 ;
        RECT 3502.330 4317.460 3502.610 4317.740 ;
        RECT 3503.040 4317.460 3503.320 4317.740 ;
        RECT 3503.750 4317.460 3504.030 4317.740 ;
        RECT 3504.460 4317.460 3504.740 4317.740 ;
        RECT 3505.170 4317.460 3505.450 4317.740 ;
        RECT 3505.880 4317.460 3506.160 4317.740 ;
        RECT 3506.590 4317.460 3506.870 4317.740 ;
        RECT 3507.300 4317.460 3507.580 4317.740 ;
        RECT 3508.010 4317.460 3508.290 4317.740 ;
        RECT 3508.720 4317.460 3509.000 4317.740 ;
        RECT 3509.430 4317.460 3509.710 4317.740 ;
        RECT 3500.200 4316.750 3500.480 4317.030 ;
        RECT 3500.910 4316.750 3501.190 4317.030 ;
        RECT 3501.620 4316.750 3501.900 4317.030 ;
        RECT 3502.330 4316.750 3502.610 4317.030 ;
        RECT 3503.040 4316.750 3503.320 4317.030 ;
        RECT 3503.750 4316.750 3504.030 4317.030 ;
        RECT 3504.460 4316.750 3504.740 4317.030 ;
        RECT 3505.170 4316.750 3505.450 4317.030 ;
        RECT 3505.880 4316.750 3506.160 4317.030 ;
        RECT 3506.590 4316.750 3506.870 4317.030 ;
        RECT 3507.300 4316.750 3507.580 4317.030 ;
        RECT 3508.010 4316.750 3508.290 4317.030 ;
        RECT 3508.720 4316.750 3509.000 4317.030 ;
        RECT 3509.430 4316.750 3509.710 4317.030 ;
        RECT 369.330 4187.970 369.610 4188.250 ;
        RECT 370.040 4187.970 370.320 4188.250 ;
        RECT 370.750 4187.970 371.030 4188.250 ;
        RECT 371.460 4187.970 371.740 4188.250 ;
        RECT 372.170 4187.970 372.450 4188.250 ;
        RECT 372.880 4187.970 373.160 4188.250 ;
        RECT 373.590 4187.970 373.870 4188.250 ;
        RECT 374.300 4187.970 374.580 4188.250 ;
        RECT 375.010 4187.970 375.290 4188.250 ;
        RECT 375.720 4187.970 376.000 4188.250 ;
        RECT 376.430 4187.970 376.710 4188.250 ;
        RECT 369.330 4187.260 369.610 4187.540 ;
        RECT 370.040 4187.260 370.320 4187.540 ;
        RECT 370.750 4187.260 371.030 4187.540 ;
        RECT 371.460 4187.260 371.740 4187.540 ;
        RECT 372.170 4187.260 372.450 4187.540 ;
        RECT 372.880 4187.260 373.160 4187.540 ;
        RECT 373.590 4187.260 373.870 4187.540 ;
        RECT 374.300 4187.260 374.580 4187.540 ;
        RECT 375.010 4187.260 375.290 4187.540 ;
        RECT 375.720 4187.260 376.000 4187.540 ;
        RECT 376.430 4187.260 376.710 4187.540 ;
        RECT 369.330 4186.550 369.610 4186.830 ;
        RECT 370.040 4186.550 370.320 4186.830 ;
        RECT 370.750 4186.550 371.030 4186.830 ;
        RECT 371.460 4186.550 371.740 4186.830 ;
        RECT 372.170 4186.550 372.450 4186.830 ;
        RECT 372.880 4186.550 373.160 4186.830 ;
        RECT 373.590 4186.550 373.870 4186.830 ;
        RECT 374.300 4186.550 374.580 4186.830 ;
        RECT 375.010 4186.550 375.290 4186.830 ;
        RECT 375.720 4186.550 376.000 4186.830 ;
        RECT 376.430 4186.550 376.710 4186.830 ;
        RECT 369.330 4185.840 369.610 4186.120 ;
        RECT 370.040 4185.840 370.320 4186.120 ;
        RECT 370.750 4185.840 371.030 4186.120 ;
        RECT 371.460 4185.840 371.740 4186.120 ;
        RECT 372.170 4185.840 372.450 4186.120 ;
        RECT 372.880 4185.840 373.160 4186.120 ;
        RECT 373.590 4185.840 373.870 4186.120 ;
        RECT 374.300 4185.840 374.580 4186.120 ;
        RECT 375.010 4185.840 375.290 4186.120 ;
        RECT 375.720 4185.840 376.000 4186.120 ;
        RECT 376.430 4185.840 376.710 4186.120 ;
        RECT 369.330 4185.130 369.610 4185.410 ;
        RECT 370.040 4185.130 370.320 4185.410 ;
        RECT 370.750 4185.130 371.030 4185.410 ;
        RECT 371.460 4185.130 371.740 4185.410 ;
        RECT 372.170 4185.130 372.450 4185.410 ;
        RECT 372.880 4185.130 373.160 4185.410 ;
        RECT 373.590 4185.130 373.870 4185.410 ;
        RECT 374.300 4185.130 374.580 4185.410 ;
        RECT 375.010 4185.130 375.290 4185.410 ;
        RECT 375.720 4185.130 376.000 4185.410 ;
        RECT 376.430 4185.130 376.710 4185.410 ;
        RECT 369.330 4184.420 369.610 4184.700 ;
        RECT 370.040 4184.420 370.320 4184.700 ;
        RECT 370.750 4184.420 371.030 4184.700 ;
        RECT 371.460 4184.420 371.740 4184.700 ;
        RECT 372.170 4184.420 372.450 4184.700 ;
        RECT 372.880 4184.420 373.160 4184.700 ;
        RECT 373.590 4184.420 373.870 4184.700 ;
        RECT 374.300 4184.420 374.580 4184.700 ;
        RECT 375.010 4184.420 375.290 4184.700 ;
        RECT 375.720 4184.420 376.000 4184.700 ;
        RECT 376.430 4184.420 376.710 4184.700 ;
        RECT 369.330 4183.710 369.610 4183.990 ;
        RECT 370.040 4183.710 370.320 4183.990 ;
        RECT 370.750 4183.710 371.030 4183.990 ;
        RECT 371.460 4183.710 371.740 4183.990 ;
        RECT 372.170 4183.710 372.450 4183.990 ;
        RECT 372.880 4183.710 373.160 4183.990 ;
        RECT 373.590 4183.710 373.870 4183.990 ;
        RECT 374.300 4183.710 374.580 4183.990 ;
        RECT 375.010 4183.710 375.290 4183.990 ;
        RECT 375.720 4183.710 376.000 4183.990 ;
        RECT 376.430 4183.710 376.710 4183.990 ;
        RECT 369.330 4183.000 369.610 4183.280 ;
        RECT 370.040 4183.000 370.320 4183.280 ;
        RECT 370.750 4183.000 371.030 4183.280 ;
        RECT 371.460 4183.000 371.740 4183.280 ;
        RECT 372.170 4183.000 372.450 4183.280 ;
        RECT 372.880 4183.000 373.160 4183.280 ;
        RECT 373.590 4183.000 373.870 4183.280 ;
        RECT 374.300 4183.000 374.580 4183.280 ;
        RECT 375.010 4183.000 375.290 4183.280 ;
        RECT 375.720 4183.000 376.000 4183.280 ;
        RECT 376.430 4183.000 376.710 4183.280 ;
        RECT 369.330 4182.290 369.610 4182.570 ;
        RECT 370.040 4182.290 370.320 4182.570 ;
        RECT 370.750 4182.290 371.030 4182.570 ;
        RECT 371.460 4182.290 371.740 4182.570 ;
        RECT 372.170 4182.290 372.450 4182.570 ;
        RECT 372.880 4182.290 373.160 4182.570 ;
        RECT 373.590 4182.290 373.870 4182.570 ;
        RECT 374.300 4182.290 374.580 4182.570 ;
        RECT 375.010 4182.290 375.290 4182.570 ;
        RECT 375.720 4182.290 376.000 4182.570 ;
        RECT 376.430 4182.290 376.710 4182.570 ;
        RECT 369.330 4181.580 369.610 4181.860 ;
        RECT 370.040 4181.580 370.320 4181.860 ;
        RECT 370.750 4181.580 371.030 4181.860 ;
        RECT 371.460 4181.580 371.740 4181.860 ;
        RECT 372.170 4181.580 372.450 4181.860 ;
        RECT 372.880 4181.580 373.160 4181.860 ;
        RECT 373.590 4181.580 373.870 4181.860 ;
        RECT 374.300 4181.580 374.580 4181.860 ;
        RECT 375.010 4181.580 375.290 4181.860 ;
        RECT 375.720 4181.580 376.000 4181.860 ;
        RECT 376.430 4181.580 376.710 4181.860 ;
        RECT 369.330 4180.870 369.610 4181.150 ;
        RECT 370.040 4180.870 370.320 4181.150 ;
        RECT 370.750 4180.870 371.030 4181.150 ;
        RECT 371.460 4180.870 371.740 4181.150 ;
        RECT 372.170 4180.870 372.450 4181.150 ;
        RECT 372.880 4180.870 373.160 4181.150 ;
        RECT 373.590 4180.870 373.870 4181.150 ;
        RECT 374.300 4180.870 374.580 4181.150 ;
        RECT 375.010 4180.870 375.290 4181.150 ;
        RECT 375.720 4180.870 376.000 4181.150 ;
        RECT 376.430 4180.870 376.710 4181.150 ;
        RECT 369.330 4180.160 369.610 4180.440 ;
        RECT 370.040 4180.160 370.320 4180.440 ;
        RECT 370.750 4180.160 371.030 4180.440 ;
        RECT 371.460 4180.160 371.740 4180.440 ;
        RECT 372.170 4180.160 372.450 4180.440 ;
        RECT 372.880 4180.160 373.160 4180.440 ;
        RECT 373.590 4180.160 373.870 4180.440 ;
        RECT 374.300 4180.160 374.580 4180.440 ;
        RECT 375.010 4180.160 375.290 4180.440 ;
        RECT 375.720 4180.160 376.000 4180.440 ;
        RECT 376.430 4180.160 376.710 4180.440 ;
        RECT 369.330 4179.450 369.610 4179.730 ;
        RECT 370.040 4179.450 370.320 4179.730 ;
        RECT 370.750 4179.450 371.030 4179.730 ;
        RECT 371.460 4179.450 371.740 4179.730 ;
        RECT 372.170 4179.450 372.450 4179.730 ;
        RECT 372.880 4179.450 373.160 4179.730 ;
        RECT 373.590 4179.450 373.870 4179.730 ;
        RECT 374.300 4179.450 374.580 4179.730 ;
        RECT 375.010 4179.450 375.290 4179.730 ;
        RECT 375.720 4179.450 376.000 4179.730 ;
        RECT 376.430 4179.450 376.710 4179.730 ;
        RECT 369.275 4175.565 369.555 4175.845 ;
        RECT 369.985 4175.565 370.265 4175.845 ;
        RECT 370.695 4175.565 370.975 4175.845 ;
        RECT 371.405 4175.565 371.685 4175.845 ;
        RECT 372.115 4175.565 372.395 4175.845 ;
        RECT 372.825 4175.565 373.105 4175.845 ;
        RECT 373.535 4175.565 373.815 4175.845 ;
        RECT 374.245 4175.565 374.525 4175.845 ;
        RECT 374.955 4175.565 375.235 4175.845 ;
        RECT 375.665 4175.565 375.945 4175.845 ;
        RECT 376.375 4175.565 376.655 4175.845 ;
        RECT 369.275 4174.855 369.555 4175.135 ;
        RECT 369.985 4174.855 370.265 4175.135 ;
        RECT 370.695 4174.855 370.975 4175.135 ;
        RECT 371.405 4174.855 371.685 4175.135 ;
        RECT 372.115 4174.855 372.395 4175.135 ;
        RECT 372.825 4174.855 373.105 4175.135 ;
        RECT 373.535 4174.855 373.815 4175.135 ;
        RECT 374.245 4174.855 374.525 4175.135 ;
        RECT 374.955 4174.855 375.235 4175.135 ;
        RECT 375.665 4174.855 375.945 4175.135 ;
        RECT 376.375 4174.855 376.655 4175.135 ;
        RECT 369.275 4174.145 369.555 4174.425 ;
        RECT 369.985 4174.145 370.265 4174.425 ;
        RECT 370.695 4174.145 370.975 4174.425 ;
        RECT 371.405 4174.145 371.685 4174.425 ;
        RECT 372.115 4174.145 372.395 4174.425 ;
        RECT 372.825 4174.145 373.105 4174.425 ;
        RECT 373.535 4174.145 373.815 4174.425 ;
        RECT 374.245 4174.145 374.525 4174.425 ;
        RECT 374.955 4174.145 375.235 4174.425 ;
        RECT 375.665 4174.145 375.945 4174.425 ;
        RECT 376.375 4174.145 376.655 4174.425 ;
        RECT 369.275 4173.435 369.555 4173.715 ;
        RECT 369.985 4173.435 370.265 4173.715 ;
        RECT 370.695 4173.435 370.975 4173.715 ;
        RECT 371.405 4173.435 371.685 4173.715 ;
        RECT 372.115 4173.435 372.395 4173.715 ;
        RECT 372.825 4173.435 373.105 4173.715 ;
        RECT 373.535 4173.435 373.815 4173.715 ;
        RECT 374.245 4173.435 374.525 4173.715 ;
        RECT 374.955 4173.435 375.235 4173.715 ;
        RECT 375.665 4173.435 375.945 4173.715 ;
        RECT 376.375 4173.435 376.655 4173.715 ;
        RECT 369.275 4172.725 369.555 4173.005 ;
        RECT 369.985 4172.725 370.265 4173.005 ;
        RECT 370.695 4172.725 370.975 4173.005 ;
        RECT 371.405 4172.725 371.685 4173.005 ;
        RECT 372.115 4172.725 372.395 4173.005 ;
        RECT 372.825 4172.725 373.105 4173.005 ;
        RECT 373.535 4172.725 373.815 4173.005 ;
        RECT 374.245 4172.725 374.525 4173.005 ;
        RECT 374.955 4172.725 375.235 4173.005 ;
        RECT 375.665 4172.725 375.945 4173.005 ;
        RECT 376.375 4172.725 376.655 4173.005 ;
        RECT 369.275 4172.015 369.555 4172.295 ;
        RECT 369.985 4172.015 370.265 4172.295 ;
        RECT 370.695 4172.015 370.975 4172.295 ;
        RECT 371.405 4172.015 371.685 4172.295 ;
        RECT 372.115 4172.015 372.395 4172.295 ;
        RECT 372.825 4172.015 373.105 4172.295 ;
        RECT 373.535 4172.015 373.815 4172.295 ;
        RECT 374.245 4172.015 374.525 4172.295 ;
        RECT 374.955 4172.015 375.235 4172.295 ;
        RECT 375.665 4172.015 375.945 4172.295 ;
        RECT 376.375 4172.015 376.655 4172.295 ;
        RECT 369.275 4171.305 369.555 4171.585 ;
        RECT 369.985 4171.305 370.265 4171.585 ;
        RECT 370.695 4171.305 370.975 4171.585 ;
        RECT 371.405 4171.305 371.685 4171.585 ;
        RECT 372.115 4171.305 372.395 4171.585 ;
        RECT 372.825 4171.305 373.105 4171.585 ;
        RECT 373.535 4171.305 373.815 4171.585 ;
        RECT 374.245 4171.305 374.525 4171.585 ;
        RECT 374.955 4171.305 375.235 4171.585 ;
        RECT 375.665 4171.305 375.945 4171.585 ;
        RECT 376.375 4171.305 376.655 4171.585 ;
        RECT 369.275 4170.595 369.555 4170.875 ;
        RECT 369.985 4170.595 370.265 4170.875 ;
        RECT 370.695 4170.595 370.975 4170.875 ;
        RECT 371.405 4170.595 371.685 4170.875 ;
        RECT 372.115 4170.595 372.395 4170.875 ;
        RECT 372.825 4170.595 373.105 4170.875 ;
        RECT 373.535 4170.595 373.815 4170.875 ;
        RECT 374.245 4170.595 374.525 4170.875 ;
        RECT 374.955 4170.595 375.235 4170.875 ;
        RECT 375.665 4170.595 375.945 4170.875 ;
        RECT 376.375 4170.595 376.655 4170.875 ;
        RECT 369.275 4169.885 369.555 4170.165 ;
        RECT 369.985 4169.885 370.265 4170.165 ;
        RECT 370.695 4169.885 370.975 4170.165 ;
        RECT 371.405 4169.885 371.685 4170.165 ;
        RECT 372.115 4169.885 372.395 4170.165 ;
        RECT 372.825 4169.885 373.105 4170.165 ;
        RECT 373.535 4169.885 373.815 4170.165 ;
        RECT 374.245 4169.885 374.525 4170.165 ;
        RECT 374.955 4169.885 375.235 4170.165 ;
        RECT 375.665 4169.885 375.945 4170.165 ;
        RECT 376.375 4169.885 376.655 4170.165 ;
        RECT 369.275 4169.175 369.555 4169.455 ;
        RECT 369.985 4169.175 370.265 4169.455 ;
        RECT 370.695 4169.175 370.975 4169.455 ;
        RECT 371.405 4169.175 371.685 4169.455 ;
        RECT 372.115 4169.175 372.395 4169.455 ;
        RECT 372.825 4169.175 373.105 4169.455 ;
        RECT 373.535 4169.175 373.815 4169.455 ;
        RECT 374.245 4169.175 374.525 4169.455 ;
        RECT 374.955 4169.175 375.235 4169.455 ;
        RECT 375.665 4169.175 375.945 4169.455 ;
        RECT 376.375 4169.175 376.655 4169.455 ;
        RECT 369.275 4168.465 369.555 4168.745 ;
        RECT 369.985 4168.465 370.265 4168.745 ;
        RECT 370.695 4168.465 370.975 4168.745 ;
        RECT 371.405 4168.465 371.685 4168.745 ;
        RECT 372.115 4168.465 372.395 4168.745 ;
        RECT 372.825 4168.465 373.105 4168.745 ;
        RECT 373.535 4168.465 373.815 4168.745 ;
        RECT 374.245 4168.465 374.525 4168.745 ;
        RECT 374.955 4168.465 375.235 4168.745 ;
        RECT 375.665 4168.465 375.945 4168.745 ;
        RECT 376.375 4168.465 376.655 4168.745 ;
        RECT 369.275 4167.755 369.555 4168.035 ;
        RECT 369.985 4167.755 370.265 4168.035 ;
        RECT 370.695 4167.755 370.975 4168.035 ;
        RECT 371.405 4167.755 371.685 4168.035 ;
        RECT 372.115 4167.755 372.395 4168.035 ;
        RECT 372.825 4167.755 373.105 4168.035 ;
        RECT 373.535 4167.755 373.815 4168.035 ;
        RECT 374.245 4167.755 374.525 4168.035 ;
        RECT 374.955 4167.755 375.235 4168.035 ;
        RECT 375.665 4167.755 375.945 4168.035 ;
        RECT 376.375 4167.755 376.655 4168.035 ;
        RECT 369.275 4167.045 369.555 4167.325 ;
        RECT 369.985 4167.045 370.265 4167.325 ;
        RECT 370.695 4167.045 370.975 4167.325 ;
        RECT 371.405 4167.045 371.685 4167.325 ;
        RECT 372.115 4167.045 372.395 4167.325 ;
        RECT 372.825 4167.045 373.105 4167.325 ;
        RECT 373.535 4167.045 373.815 4167.325 ;
        RECT 374.245 4167.045 374.525 4167.325 ;
        RECT 374.955 4167.045 375.235 4167.325 ;
        RECT 375.665 4167.045 375.945 4167.325 ;
        RECT 376.375 4167.045 376.655 4167.325 ;
        RECT 369.275 4166.335 369.555 4166.615 ;
        RECT 369.985 4166.335 370.265 4166.615 ;
        RECT 370.695 4166.335 370.975 4166.615 ;
        RECT 371.405 4166.335 371.685 4166.615 ;
        RECT 372.115 4166.335 372.395 4166.615 ;
        RECT 372.825 4166.335 373.105 4166.615 ;
        RECT 373.535 4166.335 373.815 4166.615 ;
        RECT 374.245 4166.335 374.525 4166.615 ;
        RECT 374.955 4166.335 375.235 4166.615 ;
        RECT 375.665 4166.335 375.945 4166.615 ;
        RECT 376.375 4166.335 376.655 4166.615 ;
        RECT 369.275 4163.715 369.555 4163.995 ;
        RECT 369.985 4163.715 370.265 4163.995 ;
        RECT 370.695 4163.715 370.975 4163.995 ;
        RECT 371.405 4163.715 371.685 4163.995 ;
        RECT 372.115 4163.715 372.395 4163.995 ;
        RECT 372.825 4163.715 373.105 4163.995 ;
        RECT 373.535 4163.715 373.815 4163.995 ;
        RECT 374.245 4163.715 374.525 4163.995 ;
        RECT 374.955 4163.715 375.235 4163.995 ;
        RECT 375.665 4163.715 375.945 4163.995 ;
        RECT 376.375 4163.715 376.655 4163.995 ;
        RECT 369.275 4163.005 369.555 4163.285 ;
        RECT 369.985 4163.005 370.265 4163.285 ;
        RECT 370.695 4163.005 370.975 4163.285 ;
        RECT 371.405 4163.005 371.685 4163.285 ;
        RECT 372.115 4163.005 372.395 4163.285 ;
        RECT 372.825 4163.005 373.105 4163.285 ;
        RECT 373.535 4163.005 373.815 4163.285 ;
        RECT 374.245 4163.005 374.525 4163.285 ;
        RECT 374.955 4163.005 375.235 4163.285 ;
        RECT 375.665 4163.005 375.945 4163.285 ;
        RECT 376.375 4163.005 376.655 4163.285 ;
        RECT 369.275 4162.295 369.555 4162.575 ;
        RECT 369.985 4162.295 370.265 4162.575 ;
        RECT 370.695 4162.295 370.975 4162.575 ;
        RECT 371.405 4162.295 371.685 4162.575 ;
        RECT 372.115 4162.295 372.395 4162.575 ;
        RECT 372.825 4162.295 373.105 4162.575 ;
        RECT 373.535 4162.295 373.815 4162.575 ;
        RECT 374.245 4162.295 374.525 4162.575 ;
        RECT 374.955 4162.295 375.235 4162.575 ;
        RECT 375.665 4162.295 375.945 4162.575 ;
        RECT 376.375 4162.295 376.655 4162.575 ;
        RECT 369.275 4161.585 369.555 4161.865 ;
        RECT 369.985 4161.585 370.265 4161.865 ;
        RECT 370.695 4161.585 370.975 4161.865 ;
        RECT 371.405 4161.585 371.685 4161.865 ;
        RECT 372.115 4161.585 372.395 4161.865 ;
        RECT 372.825 4161.585 373.105 4161.865 ;
        RECT 373.535 4161.585 373.815 4161.865 ;
        RECT 374.245 4161.585 374.525 4161.865 ;
        RECT 374.955 4161.585 375.235 4161.865 ;
        RECT 375.665 4161.585 375.945 4161.865 ;
        RECT 376.375 4161.585 376.655 4161.865 ;
        RECT 369.275 4160.875 369.555 4161.155 ;
        RECT 369.985 4160.875 370.265 4161.155 ;
        RECT 370.695 4160.875 370.975 4161.155 ;
        RECT 371.405 4160.875 371.685 4161.155 ;
        RECT 372.115 4160.875 372.395 4161.155 ;
        RECT 372.825 4160.875 373.105 4161.155 ;
        RECT 373.535 4160.875 373.815 4161.155 ;
        RECT 374.245 4160.875 374.525 4161.155 ;
        RECT 374.955 4160.875 375.235 4161.155 ;
        RECT 375.665 4160.875 375.945 4161.155 ;
        RECT 376.375 4160.875 376.655 4161.155 ;
        RECT 369.275 4160.165 369.555 4160.445 ;
        RECT 369.985 4160.165 370.265 4160.445 ;
        RECT 370.695 4160.165 370.975 4160.445 ;
        RECT 371.405 4160.165 371.685 4160.445 ;
        RECT 372.115 4160.165 372.395 4160.445 ;
        RECT 372.825 4160.165 373.105 4160.445 ;
        RECT 373.535 4160.165 373.815 4160.445 ;
        RECT 374.245 4160.165 374.525 4160.445 ;
        RECT 374.955 4160.165 375.235 4160.445 ;
        RECT 375.665 4160.165 375.945 4160.445 ;
        RECT 376.375 4160.165 376.655 4160.445 ;
        RECT 369.275 4159.455 369.555 4159.735 ;
        RECT 369.985 4159.455 370.265 4159.735 ;
        RECT 370.695 4159.455 370.975 4159.735 ;
        RECT 371.405 4159.455 371.685 4159.735 ;
        RECT 372.115 4159.455 372.395 4159.735 ;
        RECT 372.825 4159.455 373.105 4159.735 ;
        RECT 373.535 4159.455 373.815 4159.735 ;
        RECT 374.245 4159.455 374.525 4159.735 ;
        RECT 374.955 4159.455 375.235 4159.735 ;
        RECT 375.665 4159.455 375.945 4159.735 ;
        RECT 376.375 4159.455 376.655 4159.735 ;
        RECT 369.275 4158.745 369.555 4159.025 ;
        RECT 369.985 4158.745 370.265 4159.025 ;
        RECT 370.695 4158.745 370.975 4159.025 ;
        RECT 371.405 4158.745 371.685 4159.025 ;
        RECT 372.115 4158.745 372.395 4159.025 ;
        RECT 372.825 4158.745 373.105 4159.025 ;
        RECT 373.535 4158.745 373.815 4159.025 ;
        RECT 374.245 4158.745 374.525 4159.025 ;
        RECT 374.955 4158.745 375.235 4159.025 ;
        RECT 375.665 4158.745 375.945 4159.025 ;
        RECT 376.375 4158.745 376.655 4159.025 ;
        RECT 369.275 4158.035 369.555 4158.315 ;
        RECT 369.985 4158.035 370.265 4158.315 ;
        RECT 370.695 4158.035 370.975 4158.315 ;
        RECT 371.405 4158.035 371.685 4158.315 ;
        RECT 372.115 4158.035 372.395 4158.315 ;
        RECT 372.825 4158.035 373.105 4158.315 ;
        RECT 373.535 4158.035 373.815 4158.315 ;
        RECT 374.245 4158.035 374.525 4158.315 ;
        RECT 374.955 4158.035 375.235 4158.315 ;
        RECT 375.665 4158.035 375.945 4158.315 ;
        RECT 376.375 4158.035 376.655 4158.315 ;
        RECT 369.275 4157.325 369.555 4157.605 ;
        RECT 369.985 4157.325 370.265 4157.605 ;
        RECT 370.695 4157.325 370.975 4157.605 ;
        RECT 371.405 4157.325 371.685 4157.605 ;
        RECT 372.115 4157.325 372.395 4157.605 ;
        RECT 372.825 4157.325 373.105 4157.605 ;
        RECT 373.535 4157.325 373.815 4157.605 ;
        RECT 374.245 4157.325 374.525 4157.605 ;
        RECT 374.955 4157.325 375.235 4157.605 ;
        RECT 375.665 4157.325 375.945 4157.605 ;
        RECT 376.375 4157.325 376.655 4157.605 ;
        RECT 369.275 4156.615 369.555 4156.895 ;
        RECT 369.985 4156.615 370.265 4156.895 ;
        RECT 370.695 4156.615 370.975 4156.895 ;
        RECT 371.405 4156.615 371.685 4156.895 ;
        RECT 372.115 4156.615 372.395 4156.895 ;
        RECT 372.825 4156.615 373.105 4156.895 ;
        RECT 373.535 4156.615 373.815 4156.895 ;
        RECT 374.245 4156.615 374.525 4156.895 ;
        RECT 374.955 4156.615 375.235 4156.895 ;
        RECT 375.665 4156.615 375.945 4156.895 ;
        RECT 376.375 4156.615 376.655 4156.895 ;
        RECT 369.275 4155.905 369.555 4156.185 ;
        RECT 369.985 4155.905 370.265 4156.185 ;
        RECT 370.695 4155.905 370.975 4156.185 ;
        RECT 371.405 4155.905 371.685 4156.185 ;
        RECT 372.115 4155.905 372.395 4156.185 ;
        RECT 372.825 4155.905 373.105 4156.185 ;
        RECT 373.535 4155.905 373.815 4156.185 ;
        RECT 374.245 4155.905 374.525 4156.185 ;
        RECT 374.955 4155.905 375.235 4156.185 ;
        RECT 375.665 4155.905 375.945 4156.185 ;
        RECT 376.375 4155.905 376.655 4156.185 ;
        RECT 369.275 4155.195 369.555 4155.475 ;
        RECT 369.985 4155.195 370.265 4155.475 ;
        RECT 370.695 4155.195 370.975 4155.475 ;
        RECT 371.405 4155.195 371.685 4155.475 ;
        RECT 372.115 4155.195 372.395 4155.475 ;
        RECT 372.825 4155.195 373.105 4155.475 ;
        RECT 373.535 4155.195 373.815 4155.475 ;
        RECT 374.245 4155.195 374.525 4155.475 ;
        RECT 374.955 4155.195 375.235 4155.475 ;
        RECT 375.665 4155.195 375.945 4155.475 ;
        RECT 376.375 4155.195 376.655 4155.475 ;
        RECT 369.275 4154.485 369.555 4154.765 ;
        RECT 369.985 4154.485 370.265 4154.765 ;
        RECT 370.695 4154.485 370.975 4154.765 ;
        RECT 371.405 4154.485 371.685 4154.765 ;
        RECT 372.115 4154.485 372.395 4154.765 ;
        RECT 372.825 4154.485 373.105 4154.765 ;
        RECT 373.535 4154.485 373.815 4154.765 ;
        RECT 374.245 4154.485 374.525 4154.765 ;
        RECT 374.955 4154.485 375.235 4154.765 ;
        RECT 375.665 4154.485 375.945 4154.765 ;
        RECT 376.375 4154.485 376.655 4154.765 ;
        RECT 369.275 4150.185 369.555 4150.465 ;
        RECT 369.985 4150.185 370.265 4150.465 ;
        RECT 370.695 4150.185 370.975 4150.465 ;
        RECT 371.405 4150.185 371.685 4150.465 ;
        RECT 372.115 4150.185 372.395 4150.465 ;
        RECT 372.825 4150.185 373.105 4150.465 ;
        RECT 373.535 4150.185 373.815 4150.465 ;
        RECT 374.245 4150.185 374.525 4150.465 ;
        RECT 374.955 4150.185 375.235 4150.465 ;
        RECT 375.665 4150.185 375.945 4150.465 ;
        RECT 376.375 4150.185 376.655 4150.465 ;
        RECT 369.275 4149.475 369.555 4149.755 ;
        RECT 369.985 4149.475 370.265 4149.755 ;
        RECT 370.695 4149.475 370.975 4149.755 ;
        RECT 371.405 4149.475 371.685 4149.755 ;
        RECT 372.115 4149.475 372.395 4149.755 ;
        RECT 372.825 4149.475 373.105 4149.755 ;
        RECT 373.535 4149.475 373.815 4149.755 ;
        RECT 374.245 4149.475 374.525 4149.755 ;
        RECT 374.955 4149.475 375.235 4149.755 ;
        RECT 375.665 4149.475 375.945 4149.755 ;
        RECT 376.375 4149.475 376.655 4149.755 ;
        RECT 369.275 4148.765 369.555 4149.045 ;
        RECT 369.985 4148.765 370.265 4149.045 ;
        RECT 370.695 4148.765 370.975 4149.045 ;
        RECT 371.405 4148.765 371.685 4149.045 ;
        RECT 372.115 4148.765 372.395 4149.045 ;
        RECT 372.825 4148.765 373.105 4149.045 ;
        RECT 373.535 4148.765 373.815 4149.045 ;
        RECT 374.245 4148.765 374.525 4149.045 ;
        RECT 374.955 4148.765 375.235 4149.045 ;
        RECT 375.665 4148.765 375.945 4149.045 ;
        RECT 376.375 4148.765 376.655 4149.045 ;
        RECT 369.275 4148.055 369.555 4148.335 ;
        RECT 369.985 4148.055 370.265 4148.335 ;
        RECT 370.695 4148.055 370.975 4148.335 ;
        RECT 371.405 4148.055 371.685 4148.335 ;
        RECT 372.115 4148.055 372.395 4148.335 ;
        RECT 372.825 4148.055 373.105 4148.335 ;
        RECT 373.535 4148.055 373.815 4148.335 ;
        RECT 374.245 4148.055 374.525 4148.335 ;
        RECT 374.955 4148.055 375.235 4148.335 ;
        RECT 375.665 4148.055 375.945 4148.335 ;
        RECT 376.375 4148.055 376.655 4148.335 ;
        RECT 369.275 4147.345 369.555 4147.625 ;
        RECT 369.985 4147.345 370.265 4147.625 ;
        RECT 370.695 4147.345 370.975 4147.625 ;
        RECT 371.405 4147.345 371.685 4147.625 ;
        RECT 372.115 4147.345 372.395 4147.625 ;
        RECT 372.825 4147.345 373.105 4147.625 ;
        RECT 373.535 4147.345 373.815 4147.625 ;
        RECT 374.245 4147.345 374.525 4147.625 ;
        RECT 374.955 4147.345 375.235 4147.625 ;
        RECT 375.665 4147.345 375.945 4147.625 ;
        RECT 376.375 4147.345 376.655 4147.625 ;
        RECT 369.275 4146.635 369.555 4146.915 ;
        RECT 369.985 4146.635 370.265 4146.915 ;
        RECT 370.695 4146.635 370.975 4146.915 ;
        RECT 371.405 4146.635 371.685 4146.915 ;
        RECT 372.115 4146.635 372.395 4146.915 ;
        RECT 372.825 4146.635 373.105 4146.915 ;
        RECT 373.535 4146.635 373.815 4146.915 ;
        RECT 374.245 4146.635 374.525 4146.915 ;
        RECT 374.955 4146.635 375.235 4146.915 ;
        RECT 375.665 4146.635 375.945 4146.915 ;
        RECT 376.375 4146.635 376.655 4146.915 ;
        RECT 369.275 4145.925 369.555 4146.205 ;
        RECT 369.985 4145.925 370.265 4146.205 ;
        RECT 370.695 4145.925 370.975 4146.205 ;
        RECT 371.405 4145.925 371.685 4146.205 ;
        RECT 372.115 4145.925 372.395 4146.205 ;
        RECT 372.825 4145.925 373.105 4146.205 ;
        RECT 373.535 4145.925 373.815 4146.205 ;
        RECT 374.245 4145.925 374.525 4146.205 ;
        RECT 374.955 4145.925 375.235 4146.205 ;
        RECT 375.665 4145.925 375.945 4146.205 ;
        RECT 376.375 4145.925 376.655 4146.205 ;
        RECT 369.275 4145.215 369.555 4145.495 ;
        RECT 369.985 4145.215 370.265 4145.495 ;
        RECT 370.695 4145.215 370.975 4145.495 ;
        RECT 371.405 4145.215 371.685 4145.495 ;
        RECT 372.115 4145.215 372.395 4145.495 ;
        RECT 372.825 4145.215 373.105 4145.495 ;
        RECT 373.535 4145.215 373.815 4145.495 ;
        RECT 374.245 4145.215 374.525 4145.495 ;
        RECT 374.955 4145.215 375.235 4145.495 ;
        RECT 375.665 4145.215 375.945 4145.495 ;
        RECT 376.375 4145.215 376.655 4145.495 ;
        RECT 369.275 4144.505 369.555 4144.785 ;
        RECT 369.985 4144.505 370.265 4144.785 ;
        RECT 370.695 4144.505 370.975 4144.785 ;
        RECT 371.405 4144.505 371.685 4144.785 ;
        RECT 372.115 4144.505 372.395 4144.785 ;
        RECT 372.825 4144.505 373.105 4144.785 ;
        RECT 373.535 4144.505 373.815 4144.785 ;
        RECT 374.245 4144.505 374.525 4144.785 ;
        RECT 374.955 4144.505 375.235 4144.785 ;
        RECT 375.665 4144.505 375.945 4144.785 ;
        RECT 376.375 4144.505 376.655 4144.785 ;
        RECT 369.275 4143.795 369.555 4144.075 ;
        RECT 369.985 4143.795 370.265 4144.075 ;
        RECT 370.695 4143.795 370.975 4144.075 ;
        RECT 371.405 4143.795 371.685 4144.075 ;
        RECT 372.115 4143.795 372.395 4144.075 ;
        RECT 372.825 4143.795 373.105 4144.075 ;
        RECT 373.535 4143.795 373.815 4144.075 ;
        RECT 374.245 4143.795 374.525 4144.075 ;
        RECT 374.955 4143.795 375.235 4144.075 ;
        RECT 375.665 4143.795 375.945 4144.075 ;
        RECT 376.375 4143.795 376.655 4144.075 ;
        RECT 369.275 4143.085 369.555 4143.365 ;
        RECT 369.985 4143.085 370.265 4143.365 ;
        RECT 370.695 4143.085 370.975 4143.365 ;
        RECT 371.405 4143.085 371.685 4143.365 ;
        RECT 372.115 4143.085 372.395 4143.365 ;
        RECT 372.825 4143.085 373.105 4143.365 ;
        RECT 373.535 4143.085 373.815 4143.365 ;
        RECT 374.245 4143.085 374.525 4143.365 ;
        RECT 374.955 4143.085 375.235 4143.365 ;
        RECT 375.665 4143.085 375.945 4143.365 ;
        RECT 376.375 4143.085 376.655 4143.365 ;
        RECT 369.275 4142.375 369.555 4142.655 ;
        RECT 369.985 4142.375 370.265 4142.655 ;
        RECT 370.695 4142.375 370.975 4142.655 ;
        RECT 371.405 4142.375 371.685 4142.655 ;
        RECT 372.115 4142.375 372.395 4142.655 ;
        RECT 372.825 4142.375 373.105 4142.655 ;
        RECT 373.535 4142.375 373.815 4142.655 ;
        RECT 374.245 4142.375 374.525 4142.655 ;
        RECT 374.955 4142.375 375.235 4142.655 ;
        RECT 375.665 4142.375 375.945 4142.655 ;
        RECT 376.375 4142.375 376.655 4142.655 ;
        RECT 369.275 4141.665 369.555 4141.945 ;
        RECT 369.985 4141.665 370.265 4141.945 ;
        RECT 370.695 4141.665 370.975 4141.945 ;
        RECT 371.405 4141.665 371.685 4141.945 ;
        RECT 372.115 4141.665 372.395 4141.945 ;
        RECT 372.825 4141.665 373.105 4141.945 ;
        RECT 373.535 4141.665 373.815 4141.945 ;
        RECT 374.245 4141.665 374.525 4141.945 ;
        RECT 374.955 4141.665 375.235 4141.945 ;
        RECT 375.665 4141.665 375.945 4141.945 ;
        RECT 376.375 4141.665 376.655 4141.945 ;
        RECT 369.275 4140.955 369.555 4141.235 ;
        RECT 369.985 4140.955 370.265 4141.235 ;
        RECT 370.695 4140.955 370.975 4141.235 ;
        RECT 371.405 4140.955 371.685 4141.235 ;
        RECT 372.115 4140.955 372.395 4141.235 ;
        RECT 372.825 4140.955 373.105 4141.235 ;
        RECT 373.535 4140.955 373.815 4141.235 ;
        RECT 374.245 4140.955 374.525 4141.235 ;
        RECT 374.955 4140.955 375.235 4141.235 ;
        RECT 375.665 4140.955 375.945 4141.235 ;
        RECT 376.375 4140.955 376.655 4141.235 ;
        RECT 369.275 4138.335 369.555 4138.615 ;
        RECT 369.985 4138.335 370.265 4138.615 ;
        RECT 370.695 4138.335 370.975 4138.615 ;
        RECT 371.405 4138.335 371.685 4138.615 ;
        RECT 372.115 4138.335 372.395 4138.615 ;
        RECT 372.825 4138.335 373.105 4138.615 ;
        RECT 373.535 4138.335 373.815 4138.615 ;
        RECT 374.245 4138.335 374.525 4138.615 ;
        RECT 374.955 4138.335 375.235 4138.615 ;
        RECT 375.665 4138.335 375.945 4138.615 ;
        RECT 376.375 4138.335 376.655 4138.615 ;
        RECT 369.275 4137.625 369.555 4137.905 ;
        RECT 369.985 4137.625 370.265 4137.905 ;
        RECT 370.695 4137.625 370.975 4137.905 ;
        RECT 371.405 4137.625 371.685 4137.905 ;
        RECT 372.115 4137.625 372.395 4137.905 ;
        RECT 372.825 4137.625 373.105 4137.905 ;
        RECT 373.535 4137.625 373.815 4137.905 ;
        RECT 374.245 4137.625 374.525 4137.905 ;
        RECT 374.955 4137.625 375.235 4137.905 ;
        RECT 375.665 4137.625 375.945 4137.905 ;
        RECT 376.375 4137.625 376.655 4137.905 ;
        RECT 369.275 4136.915 369.555 4137.195 ;
        RECT 369.985 4136.915 370.265 4137.195 ;
        RECT 370.695 4136.915 370.975 4137.195 ;
        RECT 371.405 4136.915 371.685 4137.195 ;
        RECT 372.115 4136.915 372.395 4137.195 ;
        RECT 372.825 4136.915 373.105 4137.195 ;
        RECT 373.535 4136.915 373.815 4137.195 ;
        RECT 374.245 4136.915 374.525 4137.195 ;
        RECT 374.955 4136.915 375.235 4137.195 ;
        RECT 375.665 4136.915 375.945 4137.195 ;
        RECT 376.375 4136.915 376.655 4137.195 ;
        RECT 369.275 4136.205 369.555 4136.485 ;
        RECT 369.985 4136.205 370.265 4136.485 ;
        RECT 370.695 4136.205 370.975 4136.485 ;
        RECT 371.405 4136.205 371.685 4136.485 ;
        RECT 372.115 4136.205 372.395 4136.485 ;
        RECT 372.825 4136.205 373.105 4136.485 ;
        RECT 373.535 4136.205 373.815 4136.485 ;
        RECT 374.245 4136.205 374.525 4136.485 ;
        RECT 374.955 4136.205 375.235 4136.485 ;
        RECT 375.665 4136.205 375.945 4136.485 ;
        RECT 376.375 4136.205 376.655 4136.485 ;
        RECT 369.275 4135.495 369.555 4135.775 ;
        RECT 369.985 4135.495 370.265 4135.775 ;
        RECT 370.695 4135.495 370.975 4135.775 ;
        RECT 371.405 4135.495 371.685 4135.775 ;
        RECT 372.115 4135.495 372.395 4135.775 ;
        RECT 372.825 4135.495 373.105 4135.775 ;
        RECT 373.535 4135.495 373.815 4135.775 ;
        RECT 374.245 4135.495 374.525 4135.775 ;
        RECT 374.955 4135.495 375.235 4135.775 ;
        RECT 375.665 4135.495 375.945 4135.775 ;
        RECT 376.375 4135.495 376.655 4135.775 ;
        RECT 369.275 4134.785 369.555 4135.065 ;
        RECT 369.985 4134.785 370.265 4135.065 ;
        RECT 370.695 4134.785 370.975 4135.065 ;
        RECT 371.405 4134.785 371.685 4135.065 ;
        RECT 372.115 4134.785 372.395 4135.065 ;
        RECT 372.825 4134.785 373.105 4135.065 ;
        RECT 373.535 4134.785 373.815 4135.065 ;
        RECT 374.245 4134.785 374.525 4135.065 ;
        RECT 374.955 4134.785 375.235 4135.065 ;
        RECT 375.665 4134.785 375.945 4135.065 ;
        RECT 376.375 4134.785 376.655 4135.065 ;
        RECT 369.275 4134.075 369.555 4134.355 ;
        RECT 369.985 4134.075 370.265 4134.355 ;
        RECT 370.695 4134.075 370.975 4134.355 ;
        RECT 371.405 4134.075 371.685 4134.355 ;
        RECT 372.115 4134.075 372.395 4134.355 ;
        RECT 372.825 4134.075 373.105 4134.355 ;
        RECT 373.535 4134.075 373.815 4134.355 ;
        RECT 374.245 4134.075 374.525 4134.355 ;
        RECT 374.955 4134.075 375.235 4134.355 ;
        RECT 375.665 4134.075 375.945 4134.355 ;
        RECT 376.375 4134.075 376.655 4134.355 ;
        RECT 369.275 4133.365 369.555 4133.645 ;
        RECT 369.985 4133.365 370.265 4133.645 ;
        RECT 370.695 4133.365 370.975 4133.645 ;
        RECT 371.405 4133.365 371.685 4133.645 ;
        RECT 372.115 4133.365 372.395 4133.645 ;
        RECT 372.825 4133.365 373.105 4133.645 ;
        RECT 373.535 4133.365 373.815 4133.645 ;
        RECT 374.245 4133.365 374.525 4133.645 ;
        RECT 374.955 4133.365 375.235 4133.645 ;
        RECT 375.665 4133.365 375.945 4133.645 ;
        RECT 376.375 4133.365 376.655 4133.645 ;
        RECT 369.275 4132.655 369.555 4132.935 ;
        RECT 369.985 4132.655 370.265 4132.935 ;
        RECT 370.695 4132.655 370.975 4132.935 ;
        RECT 371.405 4132.655 371.685 4132.935 ;
        RECT 372.115 4132.655 372.395 4132.935 ;
        RECT 372.825 4132.655 373.105 4132.935 ;
        RECT 373.535 4132.655 373.815 4132.935 ;
        RECT 374.245 4132.655 374.525 4132.935 ;
        RECT 374.955 4132.655 375.235 4132.935 ;
        RECT 375.665 4132.655 375.945 4132.935 ;
        RECT 376.375 4132.655 376.655 4132.935 ;
        RECT 369.275 4131.945 369.555 4132.225 ;
        RECT 369.985 4131.945 370.265 4132.225 ;
        RECT 370.695 4131.945 370.975 4132.225 ;
        RECT 371.405 4131.945 371.685 4132.225 ;
        RECT 372.115 4131.945 372.395 4132.225 ;
        RECT 372.825 4131.945 373.105 4132.225 ;
        RECT 373.535 4131.945 373.815 4132.225 ;
        RECT 374.245 4131.945 374.525 4132.225 ;
        RECT 374.955 4131.945 375.235 4132.225 ;
        RECT 375.665 4131.945 375.945 4132.225 ;
        RECT 376.375 4131.945 376.655 4132.225 ;
        RECT 369.275 4131.235 369.555 4131.515 ;
        RECT 369.985 4131.235 370.265 4131.515 ;
        RECT 370.695 4131.235 370.975 4131.515 ;
        RECT 371.405 4131.235 371.685 4131.515 ;
        RECT 372.115 4131.235 372.395 4131.515 ;
        RECT 372.825 4131.235 373.105 4131.515 ;
        RECT 373.535 4131.235 373.815 4131.515 ;
        RECT 374.245 4131.235 374.525 4131.515 ;
        RECT 374.955 4131.235 375.235 4131.515 ;
        RECT 375.665 4131.235 375.945 4131.515 ;
        RECT 376.375 4131.235 376.655 4131.515 ;
        RECT 369.275 4130.525 369.555 4130.805 ;
        RECT 369.985 4130.525 370.265 4130.805 ;
        RECT 370.695 4130.525 370.975 4130.805 ;
        RECT 371.405 4130.525 371.685 4130.805 ;
        RECT 372.115 4130.525 372.395 4130.805 ;
        RECT 372.825 4130.525 373.105 4130.805 ;
        RECT 373.535 4130.525 373.815 4130.805 ;
        RECT 374.245 4130.525 374.525 4130.805 ;
        RECT 374.955 4130.525 375.235 4130.805 ;
        RECT 375.665 4130.525 375.945 4130.805 ;
        RECT 376.375 4130.525 376.655 4130.805 ;
        RECT 369.275 4129.815 369.555 4130.095 ;
        RECT 369.985 4129.815 370.265 4130.095 ;
        RECT 370.695 4129.815 370.975 4130.095 ;
        RECT 371.405 4129.815 371.685 4130.095 ;
        RECT 372.115 4129.815 372.395 4130.095 ;
        RECT 372.825 4129.815 373.105 4130.095 ;
        RECT 373.535 4129.815 373.815 4130.095 ;
        RECT 374.245 4129.815 374.525 4130.095 ;
        RECT 374.955 4129.815 375.235 4130.095 ;
        RECT 375.665 4129.815 375.945 4130.095 ;
        RECT 376.375 4129.815 376.655 4130.095 ;
        RECT 369.275 4129.105 369.555 4129.385 ;
        RECT 369.985 4129.105 370.265 4129.385 ;
        RECT 370.695 4129.105 370.975 4129.385 ;
        RECT 371.405 4129.105 371.685 4129.385 ;
        RECT 372.115 4129.105 372.395 4129.385 ;
        RECT 372.825 4129.105 373.105 4129.385 ;
        RECT 373.535 4129.105 373.815 4129.385 ;
        RECT 374.245 4129.105 374.525 4129.385 ;
        RECT 374.955 4129.105 375.235 4129.385 ;
        RECT 375.665 4129.105 375.945 4129.385 ;
        RECT 376.375 4129.105 376.655 4129.385 ;
        RECT 369.330 4125.190 369.610 4125.470 ;
        RECT 370.040 4125.190 370.320 4125.470 ;
        RECT 370.750 4125.190 371.030 4125.470 ;
        RECT 371.460 4125.190 371.740 4125.470 ;
        RECT 372.170 4125.190 372.450 4125.470 ;
        RECT 372.880 4125.190 373.160 4125.470 ;
        RECT 373.590 4125.190 373.870 4125.470 ;
        RECT 374.300 4125.190 374.580 4125.470 ;
        RECT 375.010 4125.190 375.290 4125.470 ;
        RECT 375.720 4125.190 376.000 4125.470 ;
        RECT 376.430 4125.190 376.710 4125.470 ;
        RECT 369.330 4124.480 369.610 4124.760 ;
        RECT 370.040 4124.480 370.320 4124.760 ;
        RECT 370.750 4124.480 371.030 4124.760 ;
        RECT 371.460 4124.480 371.740 4124.760 ;
        RECT 372.170 4124.480 372.450 4124.760 ;
        RECT 372.880 4124.480 373.160 4124.760 ;
        RECT 373.590 4124.480 373.870 4124.760 ;
        RECT 374.300 4124.480 374.580 4124.760 ;
        RECT 375.010 4124.480 375.290 4124.760 ;
        RECT 375.720 4124.480 376.000 4124.760 ;
        RECT 376.430 4124.480 376.710 4124.760 ;
        RECT 369.330 4123.770 369.610 4124.050 ;
        RECT 370.040 4123.770 370.320 4124.050 ;
        RECT 370.750 4123.770 371.030 4124.050 ;
        RECT 371.460 4123.770 371.740 4124.050 ;
        RECT 372.170 4123.770 372.450 4124.050 ;
        RECT 372.880 4123.770 373.160 4124.050 ;
        RECT 373.590 4123.770 373.870 4124.050 ;
        RECT 374.300 4123.770 374.580 4124.050 ;
        RECT 375.010 4123.770 375.290 4124.050 ;
        RECT 375.720 4123.770 376.000 4124.050 ;
        RECT 376.430 4123.770 376.710 4124.050 ;
        RECT 369.330 4123.060 369.610 4123.340 ;
        RECT 370.040 4123.060 370.320 4123.340 ;
        RECT 370.750 4123.060 371.030 4123.340 ;
        RECT 371.460 4123.060 371.740 4123.340 ;
        RECT 372.170 4123.060 372.450 4123.340 ;
        RECT 372.880 4123.060 373.160 4123.340 ;
        RECT 373.590 4123.060 373.870 4123.340 ;
        RECT 374.300 4123.060 374.580 4123.340 ;
        RECT 375.010 4123.060 375.290 4123.340 ;
        RECT 375.720 4123.060 376.000 4123.340 ;
        RECT 376.430 4123.060 376.710 4123.340 ;
        RECT 369.330 4122.350 369.610 4122.630 ;
        RECT 370.040 4122.350 370.320 4122.630 ;
        RECT 370.750 4122.350 371.030 4122.630 ;
        RECT 371.460 4122.350 371.740 4122.630 ;
        RECT 372.170 4122.350 372.450 4122.630 ;
        RECT 372.880 4122.350 373.160 4122.630 ;
        RECT 373.590 4122.350 373.870 4122.630 ;
        RECT 374.300 4122.350 374.580 4122.630 ;
        RECT 375.010 4122.350 375.290 4122.630 ;
        RECT 375.720 4122.350 376.000 4122.630 ;
        RECT 376.430 4122.350 376.710 4122.630 ;
        RECT 369.330 4121.640 369.610 4121.920 ;
        RECT 370.040 4121.640 370.320 4121.920 ;
        RECT 370.750 4121.640 371.030 4121.920 ;
        RECT 371.460 4121.640 371.740 4121.920 ;
        RECT 372.170 4121.640 372.450 4121.920 ;
        RECT 372.880 4121.640 373.160 4121.920 ;
        RECT 373.590 4121.640 373.870 4121.920 ;
        RECT 374.300 4121.640 374.580 4121.920 ;
        RECT 375.010 4121.640 375.290 4121.920 ;
        RECT 375.720 4121.640 376.000 4121.920 ;
        RECT 376.430 4121.640 376.710 4121.920 ;
        RECT 369.330 4120.930 369.610 4121.210 ;
        RECT 370.040 4120.930 370.320 4121.210 ;
        RECT 370.750 4120.930 371.030 4121.210 ;
        RECT 371.460 4120.930 371.740 4121.210 ;
        RECT 372.170 4120.930 372.450 4121.210 ;
        RECT 372.880 4120.930 373.160 4121.210 ;
        RECT 373.590 4120.930 373.870 4121.210 ;
        RECT 374.300 4120.930 374.580 4121.210 ;
        RECT 375.010 4120.930 375.290 4121.210 ;
        RECT 375.720 4120.930 376.000 4121.210 ;
        RECT 376.430 4120.930 376.710 4121.210 ;
        RECT 369.330 4120.220 369.610 4120.500 ;
        RECT 370.040 4120.220 370.320 4120.500 ;
        RECT 370.750 4120.220 371.030 4120.500 ;
        RECT 371.460 4120.220 371.740 4120.500 ;
        RECT 372.170 4120.220 372.450 4120.500 ;
        RECT 372.880 4120.220 373.160 4120.500 ;
        RECT 373.590 4120.220 373.870 4120.500 ;
        RECT 374.300 4120.220 374.580 4120.500 ;
        RECT 375.010 4120.220 375.290 4120.500 ;
        RECT 375.720 4120.220 376.000 4120.500 ;
        RECT 376.430 4120.220 376.710 4120.500 ;
        RECT 369.330 4119.510 369.610 4119.790 ;
        RECT 370.040 4119.510 370.320 4119.790 ;
        RECT 370.750 4119.510 371.030 4119.790 ;
        RECT 371.460 4119.510 371.740 4119.790 ;
        RECT 372.170 4119.510 372.450 4119.790 ;
        RECT 372.880 4119.510 373.160 4119.790 ;
        RECT 373.590 4119.510 373.870 4119.790 ;
        RECT 374.300 4119.510 374.580 4119.790 ;
        RECT 375.010 4119.510 375.290 4119.790 ;
        RECT 375.720 4119.510 376.000 4119.790 ;
        RECT 376.430 4119.510 376.710 4119.790 ;
        RECT 369.330 4118.800 369.610 4119.080 ;
        RECT 370.040 4118.800 370.320 4119.080 ;
        RECT 370.750 4118.800 371.030 4119.080 ;
        RECT 371.460 4118.800 371.740 4119.080 ;
        RECT 372.170 4118.800 372.450 4119.080 ;
        RECT 372.880 4118.800 373.160 4119.080 ;
        RECT 373.590 4118.800 373.870 4119.080 ;
        RECT 374.300 4118.800 374.580 4119.080 ;
        RECT 375.010 4118.800 375.290 4119.080 ;
        RECT 375.720 4118.800 376.000 4119.080 ;
        RECT 376.430 4118.800 376.710 4119.080 ;
        RECT 369.330 4118.090 369.610 4118.370 ;
        RECT 370.040 4118.090 370.320 4118.370 ;
        RECT 370.750 4118.090 371.030 4118.370 ;
        RECT 371.460 4118.090 371.740 4118.370 ;
        RECT 372.170 4118.090 372.450 4118.370 ;
        RECT 372.880 4118.090 373.160 4118.370 ;
        RECT 373.590 4118.090 373.870 4118.370 ;
        RECT 374.300 4118.090 374.580 4118.370 ;
        RECT 375.010 4118.090 375.290 4118.370 ;
        RECT 375.720 4118.090 376.000 4118.370 ;
        RECT 376.430 4118.090 376.710 4118.370 ;
        RECT 369.330 4117.380 369.610 4117.660 ;
        RECT 370.040 4117.380 370.320 4117.660 ;
        RECT 370.750 4117.380 371.030 4117.660 ;
        RECT 371.460 4117.380 371.740 4117.660 ;
        RECT 372.170 4117.380 372.450 4117.660 ;
        RECT 372.880 4117.380 373.160 4117.660 ;
        RECT 373.590 4117.380 373.870 4117.660 ;
        RECT 374.300 4117.380 374.580 4117.660 ;
        RECT 375.010 4117.380 375.290 4117.660 ;
        RECT 375.720 4117.380 376.000 4117.660 ;
        RECT 376.430 4117.380 376.710 4117.660 ;
        RECT 369.330 4116.670 369.610 4116.950 ;
        RECT 370.040 4116.670 370.320 4116.950 ;
        RECT 370.750 4116.670 371.030 4116.950 ;
        RECT 371.460 4116.670 371.740 4116.950 ;
        RECT 372.170 4116.670 372.450 4116.950 ;
        RECT 372.880 4116.670 373.160 4116.950 ;
        RECT 373.590 4116.670 373.870 4116.950 ;
        RECT 374.300 4116.670 374.580 4116.950 ;
        RECT 375.010 4116.670 375.290 4116.950 ;
        RECT 375.720 4116.670 376.000 4116.950 ;
        RECT 376.430 4116.670 376.710 4116.950 ;
        RECT 357.330 3982.970 357.610 3983.250 ;
        RECT 358.040 3982.970 358.320 3983.250 ;
        RECT 358.750 3982.970 359.030 3983.250 ;
        RECT 359.460 3982.970 359.740 3983.250 ;
        RECT 360.170 3982.970 360.450 3983.250 ;
        RECT 360.880 3982.970 361.160 3983.250 ;
        RECT 361.590 3982.970 361.870 3983.250 ;
        RECT 362.300 3982.970 362.580 3983.250 ;
        RECT 363.010 3982.970 363.290 3983.250 ;
        RECT 363.720 3982.970 364.000 3983.250 ;
        RECT 364.430 3982.970 364.710 3983.250 ;
        RECT 365.140 3982.970 365.420 3983.250 ;
        RECT 365.850 3982.970 366.130 3983.250 ;
        RECT 366.560 3982.970 366.840 3983.250 ;
        RECT 357.330 3982.260 357.610 3982.540 ;
        RECT 358.040 3982.260 358.320 3982.540 ;
        RECT 358.750 3982.260 359.030 3982.540 ;
        RECT 359.460 3982.260 359.740 3982.540 ;
        RECT 360.170 3982.260 360.450 3982.540 ;
        RECT 360.880 3982.260 361.160 3982.540 ;
        RECT 361.590 3982.260 361.870 3982.540 ;
        RECT 362.300 3982.260 362.580 3982.540 ;
        RECT 363.010 3982.260 363.290 3982.540 ;
        RECT 363.720 3982.260 364.000 3982.540 ;
        RECT 364.430 3982.260 364.710 3982.540 ;
        RECT 365.140 3982.260 365.420 3982.540 ;
        RECT 365.850 3982.260 366.130 3982.540 ;
        RECT 366.560 3982.260 366.840 3982.540 ;
        RECT 357.330 3981.550 357.610 3981.830 ;
        RECT 358.040 3981.550 358.320 3981.830 ;
        RECT 358.750 3981.550 359.030 3981.830 ;
        RECT 359.460 3981.550 359.740 3981.830 ;
        RECT 360.170 3981.550 360.450 3981.830 ;
        RECT 360.880 3981.550 361.160 3981.830 ;
        RECT 361.590 3981.550 361.870 3981.830 ;
        RECT 362.300 3981.550 362.580 3981.830 ;
        RECT 363.010 3981.550 363.290 3981.830 ;
        RECT 363.720 3981.550 364.000 3981.830 ;
        RECT 364.430 3981.550 364.710 3981.830 ;
        RECT 365.140 3981.550 365.420 3981.830 ;
        RECT 365.850 3981.550 366.130 3981.830 ;
        RECT 366.560 3981.550 366.840 3981.830 ;
        RECT 357.330 3980.840 357.610 3981.120 ;
        RECT 358.040 3980.840 358.320 3981.120 ;
        RECT 358.750 3980.840 359.030 3981.120 ;
        RECT 359.460 3980.840 359.740 3981.120 ;
        RECT 360.170 3980.840 360.450 3981.120 ;
        RECT 360.880 3980.840 361.160 3981.120 ;
        RECT 361.590 3980.840 361.870 3981.120 ;
        RECT 362.300 3980.840 362.580 3981.120 ;
        RECT 363.010 3980.840 363.290 3981.120 ;
        RECT 363.720 3980.840 364.000 3981.120 ;
        RECT 364.430 3980.840 364.710 3981.120 ;
        RECT 365.140 3980.840 365.420 3981.120 ;
        RECT 365.850 3980.840 366.130 3981.120 ;
        RECT 366.560 3980.840 366.840 3981.120 ;
        RECT 357.330 3980.130 357.610 3980.410 ;
        RECT 358.040 3980.130 358.320 3980.410 ;
        RECT 358.750 3980.130 359.030 3980.410 ;
        RECT 359.460 3980.130 359.740 3980.410 ;
        RECT 360.170 3980.130 360.450 3980.410 ;
        RECT 360.880 3980.130 361.160 3980.410 ;
        RECT 361.590 3980.130 361.870 3980.410 ;
        RECT 362.300 3980.130 362.580 3980.410 ;
        RECT 363.010 3980.130 363.290 3980.410 ;
        RECT 363.720 3980.130 364.000 3980.410 ;
        RECT 364.430 3980.130 364.710 3980.410 ;
        RECT 365.140 3980.130 365.420 3980.410 ;
        RECT 365.850 3980.130 366.130 3980.410 ;
        RECT 366.560 3980.130 366.840 3980.410 ;
        RECT 357.330 3979.420 357.610 3979.700 ;
        RECT 358.040 3979.420 358.320 3979.700 ;
        RECT 358.750 3979.420 359.030 3979.700 ;
        RECT 359.460 3979.420 359.740 3979.700 ;
        RECT 360.170 3979.420 360.450 3979.700 ;
        RECT 360.880 3979.420 361.160 3979.700 ;
        RECT 361.590 3979.420 361.870 3979.700 ;
        RECT 362.300 3979.420 362.580 3979.700 ;
        RECT 363.010 3979.420 363.290 3979.700 ;
        RECT 363.720 3979.420 364.000 3979.700 ;
        RECT 364.430 3979.420 364.710 3979.700 ;
        RECT 365.140 3979.420 365.420 3979.700 ;
        RECT 365.850 3979.420 366.130 3979.700 ;
        RECT 366.560 3979.420 366.840 3979.700 ;
        RECT 357.330 3978.710 357.610 3978.990 ;
        RECT 358.040 3978.710 358.320 3978.990 ;
        RECT 358.750 3978.710 359.030 3978.990 ;
        RECT 359.460 3978.710 359.740 3978.990 ;
        RECT 360.170 3978.710 360.450 3978.990 ;
        RECT 360.880 3978.710 361.160 3978.990 ;
        RECT 361.590 3978.710 361.870 3978.990 ;
        RECT 362.300 3978.710 362.580 3978.990 ;
        RECT 363.010 3978.710 363.290 3978.990 ;
        RECT 363.720 3978.710 364.000 3978.990 ;
        RECT 364.430 3978.710 364.710 3978.990 ;
        RECT 365.140 3978.710 365.420 3978.990 ;
        RECT 365.850 3978.710 366.130 3978.990 ;
        RECT 366.560 3978.710 366.840 3978.990 ;
        RECT 357.330 3978.000 357.610 3978.280 ;
        RECT 358.040 3978.000 358.320 3978.280 ;
        RECT 358.750 3978.000 359.030 3978.280 ;
        RECT 359.460 3978.000 359.740 3978.280 ;
        RECT 360.170 3978.000 360.450 3978.280 ;
        RECT 360.880 3978.000 361.160 3978.280 ;
        RECT 361.590 3978.000 361.870 3978.280 ;
        RECT 362.300 3978.000 362.580 3978.280 ;
        RECT 363.010 3978.000 363.290 3978.280 ;
        RECT 363.720 3978.000 364.000 3978.280 ;
        RECT 364.430 3978.000 364.710 3978.280 ;
        RECT 365.140 3978.000 365.420 3978.280 ;
        RECT 365.850 3978.000 366.130 3978.280 ;
        RECT 366.560 3978.000 366.840 3978.280 ;
        RECT 357.330 3977.290 357.610 3977.570 ;
        RECT 358.040 3977.290 358.320 3977.570 ;
        RECT 358.750 3977.290 359.030 3977.570 ;
        RECT 359.460 3977.290 359.740 3977.570 ;
        RECT 360.170 3977.290 360.450 3977.570 ;
        RECT 360.880 3977.290 361.160 3977.570 ;
        RECT 361.590 3977.290 361.870 3977.570 ;
        RECT 362.300 3977.290 362.580 3977.570 ;
        RECT 363.010 3977.290 363.290 3977.570 ;
        RECT 363.720 3977.290 364.000 3977.570 ;
        RECT 364.430 3977.290 364.710 3977.570 ;
        RECT 365.140 3977.290 365.420 3977.570 ;
        RECT 365.850 3977.290 366.130 3977.570 ;
        RECT 366.560 3977.290 366.840 3977.570 ;
        RECT 357.330 3976.580 357.610 3976.860 ;
        RECT 358.040 3976.580 358.320 3976.860 ;
        RECT 358.750 3976.580 359.030 3976.860 ;
        RECT 359.460 3976.580 359.740 3976.860 ;
        RECT 360.170 3976.580 360.450 3976.860 ;
        RECT 360.880 3976.580 361.160 3976.860 ;
        RECT 361.590 3976.580 361.870 3976.860 ;
        RECT 362.300 3976.580 362.580 3976.860 ;
        RECT 363.010 3976.580 363.290 3976.860 ;
        RECT 363.720 3976.580 364.000 3976.860 ;
        RECT 364.430 3976.580 364.710 3976.860 ;
        RECT 365.140 3976.580 365.420 3976.860 ;
        RECT 365.850 3976.580 366.130 3976.860 ;
        RECT 366.560 3976.580 366.840 3976.860 ;
        RECT 357.330 3975.870 357.610 3976.150 ;
        RECT 358.040 3975.870 358.320 3976.150 ;
        RECT 358.750 3975.870 359.030 3976.150 ;
        RECT 359.460 3975.870 359.740 3976.150 ;
        RECT 360.170 3975.870 360.450 3976.150 ;
        RECT 360.880 3975.870 361.160 3976.150 ;
        RECT 361.590 3975.870 361.870 3976.150 ;
        RECT 362.300 3975.870 362.580 3976.150 ;
        RECT 363.010 3975.870 363.290 3976.150 ;
        RECT 363.720 3975.870 364.000 3976.150 ;
        RECT 364.430 3975.870 364.710 3976.150 ;
        RECT 365.140 3975.870 365.420 3976.150 ;
        RECT 365.850 3975.870 366.130 3976.150 ;
        RECT 366.560 3975.870 366.840 3976.150 ;
        RECT 357.330 3975.160 357.610 3975.440 ;
        RECT 358.040 3975.160 358.320 3975.440 ;
        RECT 358.750 3975.160 359.030 3975.440 ;
        RECT 359.460 3975.160 359.740 3975.440 ;
        RECT 360.170 3975.160 360.450 3975.440 ;
        RECT 360.880 3975.160 361.160 3975.440 ;
        RECT 361.590 3975.160 361.870 3975.440 ;
        RECT 362.300 3975.160 362.580 3975.440 ;
        RECT 363.010 3975.160 363.290 3975.440 ;
        RECT 363.720 3975.160 364.000 3975.440 ;
        RECT 364.430 3975.160 364.710 3975.440 ;
        RECT 365.140 3975.160 365.420 3975.440 ;
        RECT 365.850 3975.160 366.130 3975.440 ;
        RECT 366.560 3975.160 366.840 3975.440 ;
        RECT 357.330 3974.450 357.610 3974.730 ;
        RECT 358.040 3974.450 358.320 3974.730 ;
        RECT 358.750 3974.450 359.030 3974.730 ;
        RECT 359.460 3974.450 359.740 3974.730 ;
        RECT 360.170 3974.450 360.450 3974.730 ;
        RECT 360.880 3974.450 361.160 3974.730 ;
        RECT 361.590 3974.450 361.870 3974.730 ;
        RECT 362.300 3974.450 362.580 3974.730 ;
        RECT 363.010 3974.450 363.290 3974.730 ;
        RECT 363.720 3974.450 364.000 3974.730 ;
        RECT 364.430 3974.450 364.710 3974.730 ;
        RECT 365.140 3974.450 365.420 3974.730 ;
        RECT 365.850 3974.450 366.130 3974.730 ;
        RECT 366.560 3974.450 366.840 3974.730 ;
        RECT 357.275 3970.565 357.555 3970.845 ;
        RECT 357.985 3970.565 358.265 3970.845 ;
        RECT 358.695 3970.565 358.975 3970.845 ;
        RECT 359.405 3970.565 359.685 3970.845 ;
        RECT 360.115 3970.565 360.395 3970.845 ;
        RECT 360.825 3970.565 361.105 3970.845 ;
        RECT 361.535 3970.565 361.815 3970.845 ;
        RECT 362.245 3970.565 362.525 3970.845 ;
        RECT 362.955 3970.565 363.235 3970.845 ;
        RECT 363.665 3970.565 363.945 3970.845 ;
        RECT 364.375 3970.565 364.655 3970.845 ;
        RECT 365.085 3970.565 365.365 3970.845 ;
        RECT 365.795 3970.565 366.075 3970.845 ;
        RECT 366.505 3970.565 366.785 3970.845 ;
        RECT 357.275 3969.855 357.555 3970.135 ;
        RECT 357.985 3969.855 358.265 3970.135 ;
        RECT 358.695 3969.855 358.975 3970.135 ;
        RECT 359.405 3969.855 359.685 3970.135 ;
        RECT 360.115 3969.855 360.395 3970.135 ;
        RECT 360.825 3969.855 361.105 3970.135 ;
        RECT 361.535 3969.855 361.815 3970.135 ;
        RECT 362.245 3969.855 362.525 3970.135 ;
        RECT 362.955 3969.855 363.235 3970.135 ;
        RECT 363.665 3969.855 363.945 3970.135 ;
        RECT 364.375 3969.855 364.655 3970.135 ;
        RECT 365.085 3969.855 365.365 3970.135 ;
        RECT 365.795 3969.855 366.075 3970.135 ;
        RECT 366.505 3969.855 366.785 3970.135 ;
        RECT 357.275 3969.145 357.555 3969.425 ;
        RECT 357.985 3969.145 358.265 3969.425 ;
        RECT 358.695 3969.145 358.975 3969.425 ;
        RECT 359.405 3969.145 359.685 3969.425 ;
        RECT 360.115 3969.145 360.395 3969.425 ;
        RECT 360.825 3969.145 361.105 3969.425 ;
        RECT 361.535 3969.145 361.815 3969.425 ;
        RECT 362.245 3969.145 362.525 3969.425 ;
        RECT 362.955 3969.145 363.235 3969.425 ;
        RECT 363.665 3969.145 363.945 3969.425 ;
        RECT 364.375 3969.145 364.655 3969.425 ;
        RECT 365.085 3969.145 365.365 3969.425 ;
        RECT 365.795 3969.145 366.075 3969.425 ;
        RECT 366.505 3969.145 366.785 3969.425 ;
        RECT 357.275 3968.435 357.555 3968.715 ;
        RECT 357.985 3968.435 358.265 3968.715 ;
        RECT 358.695 3968.435 358.975 3968.715 ;
        RECT 359.405 3968.435 359.685 3968.715 ;
        RECT 360.115 3968.435 360.395 3968.715 ;
        RECT 360.825 3968.435 361.105 3968.715 ;
        RECT 361.535 3968.435 361.815 3968.715 ;
        RECT 362.245 3968.435 362.525 3968.715 ;
        RECT 362.955 3968.435 363.235 3968.715 ;
        RECT 363.665 3968.435 363.945 3968.715 ;
        RECT 364.375 3968.435 364.655 3968.715 ;
        RECT 365.085 3968.435 365.365 3968.715 ;
        RECT 365.795 3968.435 366.075 3968.715 ;
        RECT 366.505 3968.435 366.785 3968.715 ;
        RECT 357.275 3967.725 357.555 3968.005 ;
        RECT 357.985 3967.725 358.265 3968.005 ;
        RECT 358.695 3967.725 358.975 3968.005 ;
        RECT 359.405 3967.725 359.685 3968.005 ;
        RECT 360.115 3967.725 360.395 3968.005 ;
        RECT 360.825 3967.725 361.105 3968.005 ;
        RECT 361.535 3967.725 361.815 3968.005 ;
        RECT 362.245 3967.725 362.525 3968.005 ;
        RECT 362.955 3967.725 363.235 3968.005 ;
        RECT 363.665 3967.725 363.945 3968.005 ;
        RECT 364.375 3967.725 364.655 3968.005 ;
        RECT 365.085 3967.725 365.365 3968.005 ;
        RECT 365.795 3967.725 366.075 3968.005 ;
        RECT 366.505 3967.725 366.785 3968.005 ;
        RECT 357.275 3967.015 357.555 3967.295 ;
        RECT 357.985 3967.015 358.265 3967.295 ;
        RECT 358.695 3967.015 358.975 3967.295 ;
        RECT 359.405 3967.015 359.685 3967.295 ;
        RECT 360.115 3967.015 360.395 3967.295 ;
        RECT 360.825 3967.015 361.105 3967.295 ;
        RECT 361.535 3967.015 361.815 3967.295 ;
        RECT 362.245 3967.015 362.525 3967.295 ;
        RECT 362.955 3967.015 363.235 3967.295 ;
        RECT 363.665 3967.015 363.945 3967.295 ;
        RECT 364.375 3967.015 364.655 3967.295 ;
        RECT 365.085 3967.015 365.365 3967.295 ;
        RECT 365.795 3967.015 366.075 3967.295 ;
        RECT 366.505 3967.015 366.785 3967.295 ;
        RECT 357.275 3966.305 357.555 3966.585 ;
        RECT 357.985 3966.305 358.265 3966.585 ;
        RECT 358.695 3966.305 358.975 3966.585 ;
        RECT 359.405 3966.305 359.685 3966.585 ;
        RECT 360.115 3966.305 360.395 3966.585 ;
        RECT 360.825 3966.305 361.105 3966.585 ;
        RECT 361.535 3966.305 361.815 3966.585 ;
        RECT 362.245 3966.305 362.525 3966.585 ;
        RECT 362.955 3966.305 363.235 3966.585 ;
        RECT 363.665 3966.305 363.945 3966.585 ;
        RECT 364.375 3966.305 364.655 3966.585 ;
        RECT 365.085 3966.305 365.365 3966.585 ;
        RECT 365.795 3966.305 366.075 3966.585 ;
        RECT 366.505 3966.305 366.785 3966.585 ;
        RECT 357.275 3965.595 357.555 3965.875 ;
        RECT 357.985 3965.595 358.265 3965.875 ;
        RECT 358.695 3965.595 358.975 3965.875 ;
        RECT 359.405 3965.595 359.685 3965.875 ;
        RECT 360.115 3965.595 360.395 3965.875 ;
        RECT 360.825 3965.595 361.105 3965.875 ;
        RECT 361.535 3965.595 361.815 3965.875 ;
        RECT 362.245 3965.595 362.525 3965.875 ;
        RECT 362.955 3965.595 363.235 3965.875 ;
        RECT 363.665 3965.595 363.945 3965.875 ;
        RECT 364.375 3965.595 364.655 3965.875 ;
        RECT 365.085 3965.595 365.365 3965.875 ;
        RECT 365.795 3965.595 366.075 3965.875 ;
        RECT 366.505 3965.595 366.785 3965.875 ;
        RECT 357.275 3964.885 357.555 3965.165 ;
        RECT 357.985 3964.885 358.265 3965.165 ;
        RECT 358.695 3964.885 358.975 3965.165 ;
        RECT 359.405 3964.885 359.685 3965.165 ;
        RECT 360.115 3964.885 360.395 3965.165 ;
        RECT 360.825 3964.885 361.105 3965.165 ;
        RECT 361.535 3964.885 361.815 3965.165 ;
        RECT 362.245 3964.885 362.525 3965.165 ;
        RECT 362.955 3964.885 363.235 3965.165 ;
        RECT 363.665 3964.885 363.945 3965.165 ;
        RECT 364.375 3964.885 364.655 3965.165 ;
        RECT 365.085 3964.885 365.365 3965.165 ;
        RECT 365.795 3964.885 366.075 3965.165 ;
        RECT 366.505 3964.885 366.785 3965.165 ;
        RECT 357.275 3964.175 357.555 3964.455 ;
        RECT 357.985 3964.175 358.265 3964.455 ;
        RECT 358.695 3964.175 358.975 3964.455 ;
        RECT 359.405 3964.175 359.685 3964.455 ;
        RECT 360.115 3964.175 360.395 3964.455 ;
        RECT 360.825 3964.175 361.105 3964.455 ;
        RECT 361.535 3964.175 361.815 3964.455 ;
        RECT 362.245 3964.175 362.525 3964.455 ;
        RECT 362.955 3964.175 363.235 3964.455 ;
        RECT 363.665 3964.175 363.945 3964.455 ;
        RECT 364.375 3964.175 364.655 3964.455 ;
        RECT 365.085 3964.175 365.365 3964.455 ;
        RECT 365.795 3964.175 366.075 3964.455 ;
        RECT 366.505 3964.175 366.785 3964.455 ;
        RECT 357.275 3963.465 357.555 3963.745 ;
        RECT 357.985 3963.465 358.265 3963.745 ;
        RECT 358.695 3963.465 358.975 3963.745 ;
        RECT 359.405 3963.465 359.685 3963.745 ;
        RECT 360.115 3963.465 360.395 3963.745 ;
        RECT 360.825 3963.465 361.105 3963.745 ;
        RECT 361.535 3963.465 361.815 3963.745 ;
        RECT 362.245 3963.465 362.525 3963.745 ;
        RECT 362.955 3963.465 363.235 3963.745 ;
        RECT 363.665 3963.465 363.945 3963.745 ;
        RECT 364.375 3963.465 364.655 3963.745 ;
        RECT 365.085 3963.465 365.365 3963.745 ;
        RECT 365.795 3963.465 366.075 3963.745 ;
        RECT 366.505 3963.465 366.785 3963.745 ;
        RECT 357.275 3962.755 357.555 3963.035 ;
        RECT 357.985 3962.755 358.265 3963.035 ;
        RECT 358.695 3962.755 358.975 3963.035 ;
        RECT 359.405 3962.755 359.685 3963.035 ;
        RECT 360.115 3962.755 360.395 3963.035 ;
        RECT 360.825 3962.755 361.105 3963.035 ;
        RECT 361.535 3962.755 361.815 3963.035 ;
        RECT 362.245 3962.755 362.525 3963.035 ;
        RECT 362.955 3962.755 363.235 3963.035 ;
        RECT 363.665 3962.755 363.945 3963.035 ;
        RECT 364.375 3962.755 364.655 3963.035 ;
        RECT 365.085 3962.755 365.365 3963.035 ;
        RECT 365.795 3962.755 366.075 3963.035 ;
        RECT 366.505 3962.755 366.785 3963.035 ;
        RECT 357.275 3962.045 357.555 3962.325 ;
        RECT 357.985 3962.045 358.265 3962.325 ;
        RECT 358.695 3962.045 358.975 3962.325 ;
        RECT 359.405 3962.045 359.685 3962.325 ;
        RECT 360.115 3962.045 360.395 3962.325 ;
        RECT 360.825 3962.045 361.105 3962.325 ;
        RECT 361.535 3962.045 361.815 3962.325 ;
        RECT 362.245 3962.045 362.525 3962.325 ;
        RECT 362.955 3962.045 363.235 3962.325 ;
        RECT 363.665 3962.045 363.945 3962.325 ;
        RECT 364.375 3962.045 364.655 3962.325 ;
        RECT 365.085 3962.045 365.365 3962.325 ;
        RECT 365.795 3962.045 366.075 3962.325 ;
        RECT 366.505 3962.045 366.785 3962.325 ;
        RECT 357.275 3961.335 357.555 3961.615 ;
        RECT 357.985 3961.335 358.265 3961.615 ;
        RECT 358.695 3961.335 358.975 3961.615 ;
        RECT 359.405 3961.335 359.685 3961.615 ;
        RECT 360.115 3961.335 360.395 3961.615 ;
        RECT 360.825 3961.335 361.105 3961.615 ;
        RECT 361.535 3961.335 361.815 3961.615 ;
        RECT 362.245 3961.335 362.525 3961.615 ;
        RECT 362.955 3961.335 363.235 3961.615 ;
        RECT 363.665 3961.335 363.945 3961.615 ;
        RECT 364.375 3961.335 364.655 3961.615 ;
        RECT 365.085 3961.335 365.365 3961.615 ;
        RECT 365.795 3961.335 366.075 3961.615 ;
        RECT 366.505 3961.335 366.785 3961.615 ;
        RECT 357.275 3958.715 357.555 3958.995 ;
        RECT 357.985 3958.715 358.265 3958.995 ;
        RECT 358.695 3958.715 358.975 3958.995 ;
        RECT 359.405 3958.715 359.685 3958.995 ;
        RECT 360.115 3958.715 360.395 3958.995 ;
        RECT 360.825 3958.715 361.105 3958.995 ;
        RECT 361.535 3958.715 361.815 3958.995 ;
        RECT 362.245 3958.715 362.525 3958.995 ;
        RECT 362.955 3958.715 363.235 3958.995 ;
        RECT 363.665 3958.715 363.945 3958.995 ;
        RECT 364.375 3958.715 364.655 3958.995 ;
        RECT 365.085 3958.715 365.365 3958.995 ;
        RECT 365.795 3958.715 366.075 3958.995 ;
        RECT 366.505 3958.715 366.785 3958.995 ;
        RECT 357.275 3958.005 357.555 3958.285 ;
        RECT 357.985 3958.005 358.265 3958.285 ;
        RECT 358.695 3958.005 358.975 3958.285 ;
        RECT 359.405 3958.005 359.685 3958.285 ;
        RECT 360.115 3958.005 360.395 3958.285 ;
        RECT 360.825 3958.005 361.105 3958.285 ;
        RECT 361.535 3958.005 361.815 3958.285 ;
        RECT 362.245 3958.005 362.525 3958.285 ;
        RECT 362.955 3958.005 363.235 3958.285 ;
        RECT 363.665 3958.005 363.945 3958.285 ;
        RECT 364.375 3958.005 364.655 3958.285 ;
        RECT 365.085 3958.005 365.365 3958.285 ;
        RECT 365.795 3958.005 366.075 3958.285 ;
        RECT 366.505 3958.005 366.785 3958.285 ;
        RECT 3500.200 3958.050 3500.480 3958.330 ;
        RECT 3500.910 3958.050 3501.190 3958.330 ;
        RECT 3501.620 3958.050 3501.900 3958.330 ;
        RECT 3502.330 3958.050 3502.610 3958.330 ;
        RECT 3503.040 3958.050 3503.320 3958.330 ;
        RECT 3503.750 3958.050 3504.030 3958.330 ;
        RECT 3504.460 3958.050 3504.740 3958.330 ;
        RECT 3505.170 3958.050 3505.450 3958.330 ;
        RECT 3505.880 3958.050 3506.160 3958.330 ;
        RECT 3506.590 3958.050 3506.870 3958.330 ;
        RECT 3507.300 3958.050 3507.580 3958.330 ;
        RECT 3508.010 3958.050 3508.290 3958.330 ;
        RECT 3508.720 3958.050 3509.000 3958.330 ;
        RECT 3509.430 3958.050 3509.710 3958.330 ;
        RECT 357.275 3957.295 357.555 3957.575 ;
        RECT 357.985 3957.295 358.265 3957.575 ;
        RECT 358.695 3957.295 358.975 3957.575 ;
        RECT 359.405 3957.295 359.685 3957.575 ;
        RECT 360.115 3957.295 360.395 3957.575 ;
        RECT 360.825 3957.295 361.105 3957.575 ;
        RECT 361.535 3957.295 361.815 3957.575 ;
        RECT 362.245 3957.295 362.525 3957.575 ;
        RECT 362.955 3957.295 363.235 3957.575 ;
        RECT 363.665 3957.295 363.945 3957.575 ;
        RECT 364.375 3957.295 364.655 3957.575 ;
        RECT 365.085 3957.295 365.365 3957.575 ;
        RECT 365.795 3957.295 366.075 3957.575 ;
        RECT 366.505 3957.295 366.785 3957.575 ;
        RECT 3500.200 3957.340 3500.480 3957.620 ;
        RECT 3500.910 3957.340 3501.190 3957.620 ;
        RECT 3501.620 3957.340 3501.900 3957.620 ;
        RECT 3502.330 3957.340 3502.610 3957.620 ;
        RECT 3503.040 3957.340 3503.320 3957.620 ;
        RECT 3503.750 3957.340 3504.030 3957.620 ;
        RECT 3504.460 3957.340 3504.740 3957.620 ;
        RECT 3505.170 3957.340 3505.450 3957.620 ;
        RECT 3505.880 3957.340 3506.160 3957.620 ;
        RECT 3506.590 3957.340 3506.870 3957.620 ;
        RECT 3507.300 3957.340 3507.580 3957.620 ;
        RECT 3508.010 3957.340 3508.290 3957.620 ;
        RECT 3508.720 3957.340 3509.000 3957.620 ;
        RECT 3509.430 3957.340 3509.710 3957.620 ;
        RECT 357.275 3956.585 357.555 3956.865 ;
        RECT 357.985 3956.585 358.265 3956.865 ;
        RECT 358.695 3956.585 358.975 3956.865 ;
        RECT 359.405 3956.585 359.685 3956.865 ;
        RECT 360.115 3956.585 360.395 3956.865 ;
        RECT 360.825 3956.585 361.105 3956.865 ;
        RECT 361.535 3956.585 361.815 3956.865 ;
        RECT 362.245 3956.585 362.525 3956.865 ;
        RECT 362.955 3956.585 363.235 3956.865 ;
        RECT 363.665 3956.585 363.945 3956.865 ;
        RECT 364.375 3956.585 364.655 3956.865 ;
        RECT 365.085 3956.585 365.365 3956.865 ;
        RECT 365.795 3956.585 366.075 3956.865 ;
        RECT 366.505 3956.585 366.785 3956.865 ;
        RECT 3500.200 3956.630 3500.480 3956.910 ;
        RECT 3500.910 3956.630 3501.190 3956.910 ;
        RECT 3501.620 3956.630 3501.900 3956.910 ;
        RECT 3502.330 3956.630 3502.610 3956.910 ;
        RECT 3503.040 3956.630 3503.320 3956.910 ;
        RECT 3503.750 3956.630 3504.030 3956.910 ;
        RECT 3504.460 3956.630 3504.740 3956.910 ;
        RECT 3505.170 3956.630 3505.450 3956.910 ;
        RECT 3505.880 3956.630 3506.160 3956.910 ;
        RECT 3506.590 3956.630 3506.870 3956.910 ;
        RECT 3507.300 3956.630 3507.580 3956.910 ;
        RECT 3508.010 3956.630 3508.290 3956.910 ;
        RECT 3508.720 3956.630 3509.000 3956.910 ;
        RECT 3509.430 3956.630 3509.710 3956.910 ;
        RECT 357.275 3955.875 357.555 3956.155 ;
        RECT 357.985 3955.875 358.265 3956.155 ;
        RECT 358.695 3955.875 358.975 3956.155 ;
        RECT 359.405 3955.875 359.685 3956.155 ;
        RECT 360.115 3955.875 360.395 3956.155 ;
        RECT 360.825 3955.875 361.105 3956.155 ;
        RECT 361.535 3955.875 361.815 3956.155 ;
        RECT 362.245 3955.875 362.525 3956.155 ;
        RECT 362.955 3955.875 363.235 3956.155 ;
        RECT 363.665 3955.875 363.945 3956.155 ;
        RECT 364.375 3955.875 364.655 3956.155 ;
        RECT 365.085 3955.875 365.365 3956.155 ;
        RECT 365.795 3955.875 366.075 3956.155 ;
        RECT 366.505 3955.875 366.785 3956.155 ;
        RECT 3500.200 3955.920 3500.480 3956.200 ;
        RECT 3500.910 3955.920 3501.190 3956.200 ;
        RECT 3501.620 3955.920 3501.900 3956.200 ;
        RECT 3502.330 3955.920 3502.610 3956.200 ;
        RECT 3503.040 3955.920 3503.320 3956.200 ;
        RECT 3503.750 3955.920 3504.030 3956.200 ;
        RECT 3504.460 3955.920 3504.740 3956.200 ;
        RECT 3505.170 3955.920 3505.450 3956.200 ;
        RECT 3505.880 3955.920 3506.160 3956.200 ;
        RECT 3506.590 3955.920 3506.870 3956.200 ;
        RECT 3507.300 3955.920 3507.580 3956.200 ;
        RECT 3508.010 3955.920 3508.290 3956.200 ;
        RECT 3508.720 3955.920 3509.000 3956.200 ;
        RECT 3509.430 3955.920 3509.710 3956.200 ;
        RECT 357.275 3955.165 357.555 3955.445 ;
        RECT 357.985 3955.165 358.265 3955.445 ;
        RECT 358.695 3955.165 358.975 3955.445 ;
        RECT 359.405 3955.165 359.685 3955.445 ;
        RECT 360.115 3955.165 360.395 3955.445 ;
        RECT 360.825 3955.165 361.105 3955.445 ;
        RECT 361.535 3955.165 361.815 3955.445 ;
        RECT 362.245 3955.165 362.525 3955.445 ;
        RECT 362.955 3955.165 363.235 3955.445 ;
        RECT 363.665 3955.165 363.945 3955.445 ;
        RECT 364.375 3955.165 364.655 3955.445 ;
        RECT 365.085 3955.165 365.365 3955.445 ;
        RECT 365.795 3955.165 366.075 3955.445 ;
        RECT 366.505 3955.165 366.785 3955.445 ;
        RECT 3500.200 3955.210 3500.480 3955.490 ;
        RECT 3500.910 3955.210 3501.190 3955.490 ;
        RECT 3501.620 3955.210 3501.900 3955.490 ;
        RECT 3502.330 3955.210 3502.610 3955.490 ;
        RECT 3503.040 3955.210 3503.320 3955.490 ;
        RECT 3503.750 3955.210 3504.030 3955.490 ;
        RECT 3504.460 3955.210 3504.740 3955.490 ;
        RECT 3505.170 3955.210 3505.450 3955.490 ;
        RECT 3505.880 3955.210 3506.160 3955.490 ;
        RECT 3506.590 3955.210 3506.870 3955.490 ;
        RECT 3507.300 3955.210 3507.580 3955.490 ;
        RECT 3508.010 3955.210 3508.290 3955.490 ;
        RECT 3508.720 3955.210 3509.000 3955.490 ;
        RECT 3509.430 3955.210 3509.710 3955.490 ;
        RECT 357.275 3954.455 357.555 3954.735 ;
        RECT 357.985 3954.455 358.265 3954.735 ;
        RECT 358.695 3954.455 358.975 3954.735 ;
        RECT 359.405 3954.455 359.685 3954.735 ;
        RECT 360.115 3954.455 360.395 3954.735 ;
        RECT 360.825 3954.455 361.105 3954.735 ;
        RECT 361.535 3954.455 361.815 3954.735 ;
        RECT 362.245 3954.455 362.525 3954.735 ;
        RECT 362.955 3954.455 363.235 3954.735 ;
        RECT 363.665 3954.455 363.945 3954.735 ;
        RECT 364.375 3954.455 364.655 3954.735 ;
        RECT 365.085 3954.455 365.365 3954.735 ;
        RECT 365.795 3954.455 366.075 3954.735 ;
        RECT 366.505 3954.455 366.785 3954.735 ;
        RECT 3500.200 3954.500 3500.480 3954.780 ;
        RECT 3500.910 3954.500 3501.190 3954.780 ;
        RECT 3501.620 3954.500 3501.900 3954.780 ;
        RECT 3502.330 3954.500 3502.610 3954.780 ;
        RECT 3503.040 3954.500 3503.320 3954.780 ;
        RECT 3503.750 3954.500 3504.030 3954.780 ;
        RECT 3504.460 3954.500 3504.740 3954.780 ;
        RECT 3505.170 3954.500 3505.450 3954.780 ;
        RECT 3505.880 3954.500 3506.160 3954.780 ;
        RECT 3506.590 3954.500 3506.870 3954.780 ;
        RECT 3507.300 3954.500 3507.580 3954.780 ;
        RECT 3508.010 3954.500 3508.290 3954.780 ;
        RECT 3508.720 3954.500 3509.000 3954.780 ;
        RECT 3509.430 3954.500 3509.710 3954.780 ;
        RECT 357.275 3953.745 357.555 3954.025 ;
        RECT 357.985 3953.745 358.265 3954.025 ;
        RECT 358.695 3953.745 358.975 3954.025 ;
        RECT 359.405 3953.745 359.685 3954.025 ;
        RECT 360.115 3953.745 360.395 3954.025 ;
        RECT 360.825 3953.745 361.105 3954.025 ;
        RECT 361.535 3953.745 361.815 3954.025 ;
        RECT 362.245 3953.745 362.525 3954.025 ;
        RECT 362.955 3953.745 363.235 3954.025 ;
        RECT 363.665 3953.745 363.945 3954.025 ;
        RECT 364.375 3953.745 364.655 3954.025 ;
        RECT 365.085 3953.745 365.365 3954.025 ;
        RECT 365.795 3953.745 366.075 3954.025 ;
        RECT 366.505 3953.745 366.785 3954.025 ;
        RECT 3500.200 3953.790 3500.480 3954.070 ;
        RECT 3500.910 3953.790 3501.190 3954.070 ;
        RECT 3501.620 3953.790 3501.900 3954.070 ;
        RECT 3502.330 3953.790 3502.610 3954.070 ;
        RECT 3503.040 3953.790 3503.320 3954.070 ;
        RECT 3503.750 3953.790 3504.030 3954.070 ;
        RECT 3504.460 3953.790 3504.740 3954.070 ;
        RECT 3505.170 3953.790 3505.450 3954.070 ;
        RECT 3505.880 3953.790 3506.160 3954.070 ;
        RECT 3506.590 3953.790 3506.870 3954.070 ;
        RECT 3507.300 3953.790 3507.580 3954.070 ;
        RECT 3508.010 3953.790 3508.290 3954.070 ;
        RECT 3508.720 3953.790 3509.000 3954.070 ;
        RECT 3509.430 3953.790 3509.710 3954.070 ;
        RECT 357.275 3953.035 357.555 3953.315 ;
        RECT 357.985 3953.035 358.265 3953.315 ;
        RECT 358.695 3953.035 358.975 3953.315 ;
        RECT 359.405 3953.035 359.685 3953.315 ;
        RECT 360.115 3953.035 360.395 3953.315 ;
        RECT 360.825 3953.035 361.105 3953.315 ;
        RECT 361.535 3953.035 361.815 3953.315 ;
        RECT 362.245 3953.035 362.525 3953.315 ;
        RECT 362.955 3953.035 363.235 3953.315 ;
        RECT 363.665 3953.035 363.945 3953.315 ;
        RECT 364.375 3953.035 364.655 3953.315 ;
        RECT 365.085 3953.035 365.365 3953.315 ;
        RECT 365.795 3953.035 366.075 3953.315 ;
        RECT 366.505 3953.035 366.785 3953.315 ;
        RECT 3500.200 3953.080 3500.480 3953.360 ;
        RECT 3500.910 3953.080 3501.190 3953.360 ;
        RECT 3501.620 3953.080 3501.900 3953.360 ;
        RECT 3502.330 3953.080 3502.610 3953.360 ;
        RECT 3503.040 3953.080 3503.320 3953.360 ;
        RECT 3503.750 3953.080 3504.030 3953.360 ;
        RECT 3504.460 3953.080 3504.740 3953.360 ;
        RECT 3505.170 3953.080 3505.450 3953.360 ;
        RECT 3505.880 3953.080 3506.160 3953.360 ;
        RECT 3506.590 3953.080 3506.870 3953.360 ;
        RECT 3507.300 3953.080 3507.580 3953.360 ;
        RECT 3508.010 3953.080 3508.290 3953.360 ;
        RECT 3508.720 3953.080 3509.000 3953.360 ;
        RECT 3509.430 3953.080 3509.710 3953.360 ;
        RECT 357.275 3952.325 357.555 3952.605 ;
        RECT 357.985 3952.325 358.265 3952.605 ;
        RECT 358.695 3952.325 358.975 3952.605 ;
        RECT 359.405 3952.325 359.685 3952.605 ;
        RECT 360.115 3952.325 360.395 3952.605 ;
        RECT 360.825 3952.325 361.105 3952.605 ;
        RECT 361.535 3952.325 361.815 3952.605 ;
        RECT 362.245 3952.325 362.525 3952.605 ;
        RECT 362.955 3952.325 363.235 3952.605 ;
        RECT 363.665 3952.325 363.945 3952.605 ;
        RECT 364.375 3952.325 364.655 3952.605 ;
        RECT 365.085 3952.325 365.365 3952.605 ;
        RECT 365.795 3952.325 366.075 3952.605 ;
        RECT 366.505 3952.325 366.785 3952.605 ;
        RECT 3500.200 3952.370 3500.480 3952.650 ;
        RECT 3500.910 3952.370 3501.190 3952.650 ;
        RECT 3501.620 3952.370 3501.900 3952.650 ;
        RECT 3502.330 3952.370 3502.610 3952.650 ;
        RECT 3503.040 3952.370 3503.320 3952.650 ;
        RECT 3503.750 3952.370 3504.030 3952.650 ;
        RECT 3504.460 3952.370 3504.740 3952.650 ;
        RECT 3505.170 3952.370 3505.450 3952.650 ;
        RECT 3505.880 3952.370 3506.160 3952.650 ;
        RECT 3506.590 3952.370 3506.870 3952.650 ;
        RECT 3507.300 3952.370 3507.580 3952.650 ;
        RECT 3508.010 3952.370 3508.290 3952.650 ;
        RECT 3508.720 3952.370 3509.000 3952.650 ;
        RECT 3509.430 3952.370 3509.710 3952.650 ;
        RECT 357.275 3951.615 357.555 3951.895 ;
        RECT 357.985 3951.615 358.265 3951.895 ;
        RECT 358.695 3951.615 358.975 3951.895 ;
        RECT 359.405 3951.615 359.685 3951.895 ;
        RECT 360.115 3951.615 360.395 3951.895 ;
        RECT 360.825 3951.615 361.105 3951.895 ;
        RECT 361.535 3951.615 361.815 3951.895 ;
        RECT 362.245 3951.615 362.525 3951.895 ;
        RECT 362.955 3951.615 363.235 3951.895 ;
        RECT 363.665 3951.615 363.945 3951.895 ;
        RECT 364.375 3951.615 364.655 3951.895 ;
        RECT 365.085 3951.615 365.365 3951.895 ;
        RECT 365.795 3951.615 366.075 3951.895 ;
        RECT 366.505 3951.615 366.785 3951.895 ;
        RECT 3500.200 3951.660 3500.480 3951.940 ;
        RECT 3500.910 3951.660 3501.190 3951.940 ;
        RECT 3501.620 3951.660 3501.900 3951.940 ;
        RECT 3502.330 3951.660 3502.610 3951.940 ;
        RECT 3503.040 3951.660 3503.320 3951.940 ;
        RECT 3503.750 3951.660 3504.030 3951.940 ;
        RECT 3504.460 3951.660 3504.740 3951.940 ;
        RECT 3505.170 3951.660 3505.450 3951.940 ;
        RECT 3505.880 3951.660 3506.160 3951.940 ;
        RECT 3506.590 3951.660 3506.870 3951.940 ;
        RECT 3507.300 3951.660 3507.580 3951.940 ;
        RECT 3508.010 3951.660 3508.290 3951.940 ;
        RECT 3508.720 3951.660 3509.000 3951.940 ;
        RECT 3509.430 3951.660 3509.710 3951.940 ;
        RECT 357.275 3950.905 357.555 3951.185 ;
        RECT 357.985 3950.905 358.265 3951.185 ;
        RECT 358.695 3950.905 358.975 3951.185 ;
        RECT 359.405 3950.905 359.685 3951.185 ;
        RECT 360.115 3950.905 360.395 3951.185 ;
        RECT 360.825 3950.905 361.105 3951.185 ;
        RECT 361.535 3950.905 361.815 3951.185 ;
        RECT 362.245 3950.905 362.525 3951.185 ;
        RECT 362.955 3950.905 363.235 3951.185 ;
        RECT 363.665 3950.905 363.945 3951.185 ;
        RECT 364.375 3950.905 364.655 3951.185 ;
        RECT 365.085 3950.905 365.365 3951.185 ;
        RECT 365.795 3950.905 366.075 3951.185 ;
        RECT 366.505 3950.905 366.785 3951.185 ;
        RECT 3500.200 3950.950 3500.480 3951.230 ;
        RECT 3500.910 3950.950 3501.190 3951.230 ;
        RECT 3501.620 3950.950 3501.900 3951.230 ;
        RECT 3502.330 3950.950 3502.610 3951.230 ;
        RECT 3503.040 3950.950 3503.320 3951.230 ;
        RECT 3503.750 3950.950 3504.030 3951.230 ;
        RECT 3504.460 3950.950 3504.740 3951.230 ;
        RECT 3505.170 3950.950 3505.450 3951.230 ;
        RECT 3505.880 3950.950 3506.160 3951.230 ;
        RECT 3506.590 3950.950 3506.870 3951.230 ;
        RECT 3507.300 3950.950 3507.580 3951.230 ;
        RECT 3508.010 3950.950 3508.290 3951.230 ;
        RECT 3508.720 3950.950 3509.000 3951.230 ;
        RECT 3509.430 3950.950 3509.710 3951.230 ;
        RECT 357.275 3950.195 357.555 3950.475 ;
        RECT 357.985 3950.195 358.265 3950.475 ;
        RECT 358.695 3950.195 358.975 3950.475 ;
        RECT 359.405 3950.195 359.685 3950.475 ;
        RECT 360.115 3950.195 360.395 3950.475 ;
        RECT 360.825 3950.195 361.105 3950.475 ;
        RECT 361.535 3950.195 361.815 3950.475 ;
        RECT 362.245 3950.195 362.525 3950.475 ;
        RECT 362.955 3950.195 363.235 3950.475 ;
        RECT 363.665 3950.195 363.945 3950.475 ;
        RECT 364.375 3950.195 364.655 3950.475 ;
        RECT 365.085 3950.195 365.365 3950.475 ;
        RECT 365.795 3950.195 366.075 3950.475 ;
        RECT 366.505 3950.195 366.785 3950.475 ;
        RECT 3500.200 3950.240 3500.480 3950.520 ;
        RECT 3500.910 3950.240 3501.190 3950.520 ;
        RECT 3501.620 3950.240 3501.900 3950.520 ;
        RECT 3502.330 3950.240 3502.610 3950.520 ;
        RECT 3503.040 3950.240 3503.320 3950.520 ;
        RECT 3503.750 3950.240 3504.030 3950.520 ;
        RECT 3504.460 3950.240 3504.740 3950.520 ;
        RECT 3505.170 3950.240 3505.450 3950.520 ;
        RECT 3505.880 3950.240 3506.160 3950.520 ;
        RECT 3506.590 3950.240 3506.870 3950.520 ;
        RECT 3507.300 3950.240 3507.580 3950.520 ;
        RECT 3508.010 3950.240 3508.290 3950.520 ;
        RECT 3508.720 3950.240 3509.000 3950.520 ;
        RECT 3509.430 3950.240 3509.710 3950.520 ;
        RECT 357.275 3949.485 357.555 3949.765 ;
        RECT 357.985 3949.485 358.265 3949.765 ;
        RECT 358.695 3949.485 358.975 3949.765 ;
        RECT 359.405 3949.485 359.685 3949.765 ;
        RECT 360.115 3949.485 360.395 3949.765 ;
        RECT 360.825 3949.485 361.105 3949.765 ;
        RECT 361.535 3949.485 361.815 3949.765 ;
        RECT 362.245 3949.485 362.525 3949.765 ;
        RECT 362.955 3949.485 363.235 3949.765 ;
        RECT 363.665 3949.485 363.945 3949.765 ;
        RECT 364.375 3949.485 364.655 3949.765 ;
        RECT 365.085 3949.485 365.365 3949.765 ;
        RECT 365.795 3949.485 366.075 3949.765 ;
        RECT 366.505 3949.485 366.785 3949.765 ;
        RECT 3500.200 3949.530 3500.480 3949.810 ;
        RECT 3500.910 3949.530 3501.190 3949.810 ;
        RECT 3501.620 3949.530 3501.900 3949.810 ;
        RECT 3502.330 3949.530 3502.610 3949.810 ;
        RECT 3503.040 3949.530 3503.320 3949.810 ;
        RECT 3503.750 3949.530 3504.030 3949.810 ;
        RECT 3504.460 3949.530 3504.740 3949.810 ;
        RECT 3505.170 3949.530 3505.450 3949.810 ;
        RECT 3505.880 3949.530 3506.160 3949.810 ;
        RECT 3506.590 3949.530 3506.870 3949.810 ;
        RECT 3507.300 3949.530 3507.580 3949.810 ;
        RECT 3508.010 3949.530 3508.290 3949.810 ;
        RECT 3508.720 3949.530 3509.000 3949.810 ;
        RECT 3509.430 3949.530 3509.710 3949.810 ;
        RECT 3500.255 3945.615 3500.535 3945.895 ;
        RECT 3500.965 3945.615 3501.245 3945.895 ;
        RECT 3501.675 3945.615 3501.955 3945.895 ;
        RECT 3502.385 3945.615 3502.665 3945.895 ;
        RECT 3503.095 3945.615 3503.375 3945.895 ;
        RECT 3503.805 3945.615 3504.085 3945.895 ;
        RECT 3504.515 3945.615 3504.795 3945.895 ;
        RECT 3505.225 3945.615 3505.505 3945.895 ;
        RECT 3505.935 3945.615 3506.215 3945.895 ;
        RECT 3506.645 3945.615 3506.925 3945.895 ;
        RECT 3507.355 3945.615 3507.635 3945.895 ;
        RECT 3508.065 3945.615 3508.345 3945.895 ;
        RECT 3508.775 3945.615 3509.055 3945.895 ;
        RECT 3509.485 3945.615 3509.765 3945.895 ;
        RECT 357.275 3945.185 357.555 3945.465 ;
        RECT 357.985 3945.185 358.265 3945.465 ;
        RECT 358.695 3945.185 358.975 3945.465 ;
        RECT 359.405 3945.185 359.685 3945.465 ;
        RECT 360.115 3945.185 360.395 3945.465 ;
        RECT 360.825 3945.185 361.105 3945.465 ;
        RECT 361.535 3945.185 361.815 3945.465 ;
        RECT 362.245 3945.185 362.525 3945.465 ;
        RECT 362.955 3945.185 363.235 3945.465 ;
        RECT 363.665 3945.185 363.945 3945.465 ;
        RECT 364.375 3945.185 364.655 3945.465 ;
        RECT 365.085 3945.185 365.365 3945.465 ;
        RECT 365.795 3945.185 366.075 3945.465 ;
        RECT 366.505 3945.185 366.785 3945.465 ;
        RECT 3500.255 3944.905 3500.535 3945.185 ;
        RECT 3500.965 3944.905 3501.245 3945.185 ;
        RECT 3501.675 3944.905 3501.955 3945.185 ;
        RECT 3502.385 3944.905 3502.665 3945.185 ;
        RECT 3503.095 3944.905 3503.375 3945.185 ;
        RECT 3503.805 3944.905 3504.085 3945.185 ;
        RECT 3504.515 3944.905 3504.795 3945.185 ;
        RECT 3505.225 3944.905 3505.505 3945.185 ;
        RECT 3505.935 3944.905 3506.215 3945.185 ;
        RECT 3506.645 3944.905 3506.925 3945.185 ;
        RECT 3507.355 3944.905 3507.635 3945.185 ;
        RECT 3508.065 3944.905 3508.345 3945.185 ;
        RECT 3508.775 3944.905 3509.055 3945.185 ;
        RECT 3509.485 3944.905 3509.765 3945.185 ;
        RECT 357.275 3944.475 357.555 3944.755 ;
        RECT 357.985 3944.475 358.265 3944.755 ;
        RECT 358.695 3944.475 358.975 3944.755 ;
        RECT 359.405 3944.475 359.685 3944.755 ;
        RECT 360.115 3944.475 360.395 3944.755 ;
        RECT 360.825 3944.475 361.105 3944.755 ;
        RECT 361.535 3944.475 361.815 3944.755 ;
        RECT 362.245 3944.475 362.525 3944.755 ;
        RECT 362.955 3944.475 363.235 3944.755 ;
        RECT 363.665 3944.475 363.945 3944.755 ;
        RECT 364.375 3944.475 364.655 3944.755 ;
        RECT 365.085 3944.475 365.365 3944.755 ;
        RECT 365.795 3944.475 366.075 3944.755 ;
        RECT 366.505 3944.475 366.785 3944.755 ;
        RECT 3500.255 3944.195 3500.535 3944.475 ;
        RECT 3500.965 3944.195 3501.245 3944.475 ;
        RECT 3501.675 3944.195 3501.955 3944.475 ;
        RECT 3502.385 3944.195 3502.665 3944.475 ;
        RECT 3503.095 3944.195 3503.375 3944.475 ;
        RECT 3503.805 3944.195 3504.085 3944.475 ;
        RECT 3504.515 3944.195 3504.795 3944.475 ;
        RECT 3505.225 3944.195 3505.505 3944.475 ;
        RECT 3505.935 3944.195 3506.215 3944.475 ;
        RECT 3506.645 3944.195 3506.925 3944.475 ;
        RECT 3507.355 3944.195 3507.635 3944.475 ;
        RECT 3508.065 3944.195 3508.345 3944.475 ;
        RECT 3508.775 3944.195 3509.055 3944.475 ;
        RECT 3509.485 3944.195 3509.765 3944.475 ;
        RECT 357.275 3943.765 357.555 3944.045 ;
        RECT 357.985 3943.765 358.265 3944.045 ;
        RECT 358.695 3943.765 358.975 3944.045 ;
        RECT 359.405 3943.765 359.685 3944.045 ;
        RECT 360.115 3943.765 360.395 3944.045 ;
        RECT 360.825 3943.765 361.105 3944.045 ;
        RECT 361.535 3943.765 361.815 3944.045 ;
        RECT 362.245 3943.765 362.525 3944.045 ;
        RECT 362.955 3943.765 363.235 3944.045 ;
        RECT 363.665 3943.765 363.945 3944.045 ;
        RECT 364.375 3943.765 364.655 3944.045 ;
        RECT 365.085 3943.765 365.365 3944.045 ;
        RECT 365.795 3943.765 366.075 3944.045 ;
        RECT 366.505 3943.765 366.785 3944.045 ;
        RECT 3500.255 3943.485 3500.535 3943.765 ;
        RECT 3500.965 3943.485 3501.245 3943.765 ;
        RECT 3501.675 3943.485 3501.955 3943.765 ;
        RECT 3502.385 3943.485 3502.665 3943.765 ;
        RECT 3503.095 3943.485 3503.375 3943.765 ;
        RECT 3503.805 3943.485 3504.085 3943.765 ;
        RECT 3504.515 3943.485 3504.795 3943.765 ;
        RECT 3505.225 3943.485 3505.505 3943.765 ;
        RECT 3505.935 3943.485 3506.215 3943.765 ;
        RECT 3506.645 3943.485 3506.925 3943.765 ;
        RECT 3507.355 3943.485 3507.635 3943.765 ;
        RECT 3508.065 3943.485 3508.345 3943.765 ;
        RECT 3508.775 3943.485 3509.055 3943.765 ;
        RECT 3509.485 3943.485 3509.765 3943.765 ;
        RECT 357.275 3943.055 357.555 3943.335 ;
        RECT 357.985 3943.055 358.265 3943.335 ;
        RECT 358.695 3943.055 358.975 3943.335 ;
        RECT 359.405 3943.055 359.685 3943.335 ;
        RECT 360.115 3943.055 360.395 3943.335 ;
        RECT 360.825 3943.055 361.105 3943.335 ;
        RECT 361.535 3943.055 361.815 3943.335 ;
        RECT 362.245 3943.055 362.525 3943.335 ;
        RECT 362.955 3943.055 363.235 3943.335 ;
        RECT 363.665 3943.055 363.945 3943.335 ;
        RECT 364.375 3943.055 364.655 3943.335 ;
        RECT 365.085 3943.055 365.365 3943.335 ;
        RECT 365.795 3943.055 366.075 3943.335 ;
        RECT 366.505 3943.055 366.785 3943.335 ;
        RECT 3500.255 3942.775 3500.535 3943.055 ;
        RECT 3500.965 3942.775 3501.245 3943.055 ;
        RECT 3501.675 3942.775 3501.955 3943.055 ;
        RECT 3502.385 3942.775 3502.665 3943.055 ;
        RECT 3503.095 3942.775 3503.375 3943.055 ;
        RECT 3503.805 3942.775 3504.085 3943.055 ;
        RECT 3504.515 3942.775 3504.795 3943.055 ;
        RECT 3505.225 3942.775 3505.505 3943.055 ;
        RECT 3505.935 3942.775 3506.215 3943.055 ;
        RECT 3506.645 3942.775 3506.925 3943.055 ;
        RECT 3507.355 3942.775 3507.635 3943.055 ;
        RECT 3508.065 3942.775 3508.345 3943.055 ;
        RECT 3508.775 3942.775 3509.055 3943.055 ;
        RECT 3509.485 3942.775 3509.765 3943.055 ;
        RECT 357.275 3942.345 357.555 3942.625 ;
        RECT 357.985 3942.345 358.265 3942.625 ;
        RECT 358.695 3942.345 358.975 3942.625 ;
        RECT 359.405 3942.345 359.685 3942.625 ;
        RECT 360.115 3942.345 360.395 3942.625 ;
        RECT 360.825 3942.345 361.105 3942.625 ;
        RECT 361.535 3942.345 361.815 3942.625 ;
        RECT 362.245 3942.345 362.525 3942.625 ;
        RECT 362.955 3942.345 363.235 3942.625 ;
        RECT 363.665 3942.345 363.945 3942.625 ;
        RECT 364.375 3942.345 364.655 3942.625 ;
        RECT 365.085 3942.345 365.365 3942.625 ;
        RECT 365.795 3942.345 366.075 3942.625 ;
        RECT 366.505 3942.345 366.785 3942.625 ;
        RECT 3500.255 3942.065 3500.535 3942.345 ;
        RECT 3500.965 3942.065 3501.245 3942.345 ;
        RECT 3501.675 3942.065 3501.955 3942.345 ;
        RECT 3502.385 3942.065 3502.665 3942.345 ;
        RECT 3503.095 3942.065 3503.375 3942.345 ;
        RECT 3503.805 3942.065 3504.085 3942.345 ;
        RECT 3504.515 3942.065 3504.795 3942.345 ;
        RECT 3505.225 3942.065 3505.505 3942.345 ;
        RECT 3505.935 3942.065 3506.215 3942.345 ;
        RECT 3506.645 3942.065 3506.925 3942.345 ;
        RECT 3507.355 3942.065 3507.635 3942.345 ;
        RECT 3508.065 3942.065 3508.345 3942.345 ;
        RECT 3508.775 3942.065 3509.055 3942.345 ;
        RECT 3509.485 3942.065 3509.765 3942.345 ;
        RECT 357.275 3941.635 357.555 3941.915 ;
        RECT 357.985 3941.635 358.265 3941.915 ;
        RECT 358.695 3941.635 358.975 3941.915 ;
        RECT 359.405 3941.635 359.685 3941.915 ;
        RECT 360.115 3941.635 360.395 3941.915 ;
        RECT 360.825 3941.635 361.105 3941.915 ;
        RECT 361.535 3941.635 361.815 3941.915 ;
        RECT 362.245 3941.635 362.525 3941.915 ;
        RECT 362.955 3941.635 363.235 3941.915 ;
        RECT 363.665 3941.635 363.945 3941.915 ;
        RECT 364.375 3941.635 364.655 3941.915 ;
        RECT 365.085 3941.635 365.365 3941.915 ;
        RECT 365.795 3941.635 366.075 3941.915 ;
        RECT 366.505 3941.635 366.785 3941.915 ;
        RECT 3500.255 3941.355 3500.535 3941.635 ;
        RECT 3500.965 3941.355 3501.245 3941.635 ;
        RECT 3501.675 3941.355 3501.955 3941.635 ;
        RECT 3502.385 3941.355 3502.665 3941.635 ;
        RECT 3503.095 3941.355 3503.375 3941.635 ;
        RECT 3503.805 3941.355 3504.085 3941.635 ;
        RECT 3504.515 3941.355 3504.795 3941.635 ;
        RECT 3505.225 3941.355 3505.505 3941.635 ;
        RECT 3505.935 3941.355 3506.215 3941.635 ;
        RECT 3506.645 3941.355 3506.925 3941.635 ;
        RECT 3507.355 3941.355 3507.635 3941.635 ;
        RECT 3508.065 3941.355 3508.345 3941.635 ;
        RECT 3508.775 3941.355 3509.055 3941.635 ;
        RECT 3509.485 3941.355 3509.765 3941.635 ;
        RECT 357.275 3940.925 357.555 3941.205 ;
        RECT 357.985 3940.925 358.265 3941.205 ;
        RECT 358.695 3940.925 358.975 3941.205 ;
        RECT 359.405 3940.925 359.685 3941.205 ;
        RECT 360.115 3940.925 360.395 3941.205 ;
        RECT 360.825 3940.925 361.105 3941.205 ;
        RECT 361.535 3940.925 361.815 3941.205 ;
        RECT 362.245 3940.925 362.525 3941.205 ;
        RECT 362.955 3940.925 363.235 3941.205 ;
        RECT 363.665 3940.925 363.945 3941.205 ;
        RECT 364.375 3940.925 364.655 3941.205 ;
        RECT 365.085 3940.925 365.365 3941.205 ;
        RECT 365.795 3940.925 366.075 3941.205 ;
        RECT 366.505 3940.925 366.785 3941.205 ;
        RECT 3500.255 3940.645 3500.535 3940.925 ;
        RECT 3500.965 3940.645 3501.245 3940.925 ;
        RECT 3501.675 3940.645 3501.955 3940.925 ;
        RECT 3502.385 3940.645 3502.665 3940.925 ;
        RECT 3503.095 3940.645 3503.375 3940.925 ;
        RECT 3503.805 3940.645 3504.085 3940.925 ;
        RECT 3504.515 3940.645 3504.795 3940.925 ;
        RECT 3505.225 3940.645 3505.505 3940.925 ;
        RECT 3505.935 3940.645 3506.215 3940.925 ;
        RECT 3506.645 3940.645 3506.925 3940.925 ;
        RECT 3507.355 3940.645 3507.635 3940.925 ;
        RECT 3508.065 3940.645 3508.345 3940.925 ;
        RECT 3508.775 3940.645 3509.055 3940.925 ;
        RECT 3509.485 3940.645 3509.765 3940.925 ;
        RECT 357.275 3940.215 357.555 3940.495 ;
        RECT 357.985 3940.215 358.265 3940.495 ;
        RECT 358.695 3940.215 358.975 3940.495 ;
        RECT 359.405 3940.215 359.685 3940.495 ;
        RECT 360.115 3940.215 360.395 3940.495 ;
        RECT 360.825 3940.215 361.105 3940.495 ;
        RECT 361.535 3940.215 361.815 3940.495 ;
        RECT 362.245 3940.215 362.525 3940.495 ;
        RECT 362.955 3940.215 363.235 3940.495 ;
        RECT 363.665 3940.215 363.945 3940.495 ;
        RECT 364.375 3940.215 364.655 3940.495 ;
        RECT 365.085 3940.215 365.365 3940.495 ;
        RECT 365.795 3940.215 366.075 3940.495 ;
        RECT 366.505 3940.215 366.785 3940.495 ;
        RECT 3500.255 3939.935 3500.535 3940.215 ;
        RECT 3500.965 3939.935 3501.245 3940.215 ;
        RECT 3501.675 3939.935 3501.955 3940.215 ;
        RECT 3502.385 3939.935 3502.665 3940.215 ;
        RECT 3503.095 3939.935 3503.375 3940.215 ;
        RECT 3503.805 3939.935 3504.085 3940.215 ;
        RECT 3504.515 3939.935 3504.795 3940.215 ;
        RECT 3505.225 3939.935 3505.505 3940.215 ;
        RECT 3505.935 3939.935 3506.215 3940.215 ;
        RECT 3506.645 3939.935 3506.925 3940.215 ;
        RECT 3507.355 3939.935 3507.635 3940.215 ;
        RECT 3508.065 3939.935 3508.345 3940.215 ;
        RECT 3508.775 3939.935 3509.055 3940.215 ;
        RECT 3509.485 3939.935 3509.765 3940.215 ;
        RECT 357.275 3939.505 357.555 3939.785 ;
        RECT 357.985 3939.505 358.265 3939.785 ;
        RECT 358.695 3939.505 358.975 3939.785 ;
        RECT 359.405 3939.505 359.685 3939.785 ;
        RECT 360.115 3939.505 360.395 3939.785 ;
        RECT 360.825 3939.505 361.105 3939.785 ;
        RECT 361.535 3939.505 361.815 3939.785 ;
        RECT 362.245 3939.505 362.525 3939.785 ;
        RECT 362.955 3939.505 363.235 3939.785 ;
        RECT 363.665 3939.505 363.945 3939.785 ;
        RECT 364.375 3939.505 364.655 3939.785 ;
        RECT 365.085 3939.505 365.365 3939.785 ;
        RECT 365.795 3939.505 366.075 3939.785 ;
        RECT 366.505 3939.505 366.785 3939.785 ;
        RECT 3500.255 3939.225 3500.535 3939.505 ;
        RECT 3500.965 3939.225 3501.245 3939.505 ;
        RECT 3501.675 3939.225 3501.955 3939.505 ;
        RECT 3502.385 3939.225 3502.665 3939.505 ;
        RECT 3503.095 3939.225 3503.375 3939.505 ;
        RECT 3503.805 3939.225 3504.085 3939.505 ;
        RECT 3504.515 3939.225 3504.795 3939.505 ;
        RECT 3505.225 3939.225 3505.505 3939.505 ;
        RECT 3505.935 3939.225 3506.215 3939.505 ;
        RECT 3506.645 3939.225 3506.925 3939.505 ;
        RECT 3507.355 3939.225 3507.635 3939.505 ;
        RECT 3508.065 3939.225 3508.345 3939.505 ;
        RECT 3508.775 3939.225 3509.055 3939.505 ;
        RECT 3509.485 3939.225 3509.765 3939.505 ;
        RECT 357.275 3938.795 357.555 3939.075 ;
        RECT 357.985 3938.795 358.265 3939.075 ;
        RECT 358.695 3938.795 358.975 3939.075 ;
        RECT 359.405 3938.795 359.685 3939.075 ;
        RECT 360.115 3938.795 360.395 3939.075 ;
        RECT 360.825 3938.795 361.105 3939.075 ;
        RECT 361.535 3938.795 361.815 3939.075 ;
        RECT 362.245 3938.795 362.525 3939.075 ;
        RECT 362.955 3938.795 363.235 3939.075 ;
        RECT 363.665 3938.795 363.945 3939.075 ;
        RECT 364.375 3938.795 364.655 3939.075 ;
        RECT 365.085 3938.795 365.365 3939.075 ;
        RECT 365.795 3938.795 366.075 3939.075 ;
        RECT 366.505 3938.795 366.785 3939.075 ;
        RECT 3500.255 3938.515 3500.535 3938.795 ;
        RECT 3500.965 3938.515 3501.245 3938.795 ;
        RECT 3501.675 3938.515 3501.955 3938.795 ;
        RECT 3502.385 3938.515 3502.665 3938.795 ;
        RECT 3503.095 3938.515 3503.375 3938.795 ;
        RECT 3503.805 3938.515 3504.085 3938.795 ;
        RECT 3504.515 3938.515 3504.795 3938.795 ;
        RECT 3505.225 3938.515 3505.505 3938.795 ;
        RECT 3505.935 3938.515 3506.215 3938.795 ;
        RECT 3506.645 3938.515 3506.925 3938.795 ;
        RECT 3507.355 3938.515 3507.635 3938.795 ;
        RECT 3508.065 3938.515 3508.345 3938.795 ;
        RECT 3508.775 3938.515 3509.055 3938.795 ;
        RECT 3509.485 3938.515 3509.765 3938.795 ;
        RECT 357.275 3938.085 357.555 3938.365 ;
        RECT 357.985 3938.085 358.265 3938.365 ;
        RECT 358.695 3938.085 358.975 3938.365 ;
        RECT 359.405 3938.085 359.685 3938.365 ;
        RECT 360.115 3938.085 360.395 3938.365 ;
        RECT 360.825 3938.085 361.105 3938.365 ;
        RECT 361.535 3938.085 361.815 3938.365 ;
        RECT 362.245 3938.085 362.525 3938.365 ;
        RECT 362.955 3938.085 363.235 3938.365 ;
        RECT 363.665 3938.085 363.945 3938.365 ;
        RECT 364.375 3938.085 364.655 3938.365 ;
        RECT 365.085 3938.085 365.365 3938.365 ;
        RECT 365.795 3938.085 366.075 3938.365 ;
        RECT 366.505 3938.085 366.785 3938.365 ;
        RECT 3500.255 3937.805 3500.535 3938.085 ;
        RECT 3500.965 3937.805 3501.245 3938.085 ;
        RECT 3501.675 3937.805 3501.955 3938.085 ;
        RECT 3502.385 3937.805 3502.665 3938.085 ;
        RECT 3503.095 3937.805 3503.375 3938.085 ;
        RECT 3503.805 3937.805 3504.085 3938.085 ;
        RECT 3504.515 3937.805 3504.795 3938.085 ;
        RECT 3505.225 3937.805 3505.505 3938.085 ;
        RECT 3505.935 3937.805 3506.215 3938.085 ;
        RECT 3506.645 3937.805 3506.925 3938.085 ;
        RECT 3507.355 3937.805 3507.635 3938.085 ;
        RECT 3508.065 3937.805 3508.345 3938.085 ;
        RECT 3508.775 3937.805 3509.055 3938.085 ;
        RECT 3509.485 3937.805 3509.765 3938.085 ;
        RECT 357.275 3937.375 357.555 3937.655 ;
        RECT 357.985 3937.375 358.265 3937.655 ;
        RECT 358.695 3937.375 358.975 3937.655 ;
        RECT 359.405 3937.375 359.685 3937.655 ;
        RECT 360.115 3937.375 360.395 3937.655 ;
        RECT 360.825 3937.375 361.105 3937.655 ;
        RECT 361.535 3937.375 361.815 3937.655 ;
        RECT 362.245 3937.375 362.525 3937.655 ;
        RECT 362.955 3937.375 363.235 3937.655 ;
        RECT 363.665 3937.375 363.945 3937.655 ;
        RECT 364.375 3937.375 364.655 3937.655 ;
        RECT 365.085 3937.375 365.365 3937.655 ;
        RECT 365.795 3937.375 366.075 3937.655 ;
        RECT 366.505 3937.375 366.785 3937.655 ;
        RECT 3500.255 3937.095 3500.535 3937.375 ;
        RECT 3500.965 3937.095 3501.245 3937.375 ;
        RECT 3501.675 3937.095 3501.955 3937.375 ;
        RECT 3502.385 3937.095 3502.665 3937.375 ;
        RECT 3503.095 3937.095 3503.375 3937.375 ;
        RECT 3503.805 3937.095 3504.085 3937.375 ;
        RECT 3504.515 3937.095 3504.795 3937.375 ;
        RECT 3505.225 3937.095 3505.505 3937.375 ;
        RECT 3505.935 3937.095 3506.215 3937.375 ;
        RECT 3506.645 3937.095 3506.925 3937.375 ;
        RECT 3507.355 3937.095 3507.635 3937.375 ;
        RECT 3508.065 3937.095 3508.345 3937.375 ;
        RECT 3508.775 3937.095 3509.055 3937.375 ;
        RECT 3509.485 3937.095 3509.765 3937.375 ;
        RECT 357.275 3936.665 357.555 3936.945 ;
        RECT 357.985 3936.665 358.265 3936.945 ;
        RECT 358.695 3936.665 358.975 3936.945 ;
        RECT 359.405 3936.665 359.685 3936.945 ;
        RECT 360.115 3936.665 360.395 3936.945 ;
        RECT 360.825 3936.665 361.105 3936.945 ;
        RECT 361.535 3936.665 361.815 3936.945 ;
        RECT 362.245 3936.665 362.525 3936.945 ;
        RECT 362.955 3936.665 363.235 3936.945 ;
        RECT 363.665 3936.665 363.945 3936.945 ;
        RECT 364.375 3936.665 364.655 3936.945 ;
        RECT 365.085 3936.665 365.365 3936.945 ;
        RECT 365.795 3936.665 366.075 3936.945 ;
        RECT 366.505 3936.665 366.785 3936.945 ;
        RECT 3500.255 3936.385 3500.535 3936.665 ;
        RECT 3500.965 3936.385 3501.245 3936.665 ;
        RECT 3501.675 3936.385 3501.955 3936.665 ;
        RECT 3502.385 3936.385 3502.665 3936.665 ;
        RECT 3503.095 3936.385 3503.375 3936.665 ;
        RECT 3503.805 3936.385 3504.085 3936.665 ;
        RECT 3504.515 3936.385 3504.795 3936.665 ;
        RECT 3505.225 3936.385 3505.505 3936.665 ;
        RECT 3505.935 3936.385 3506.215 3936.665 ;
        RECT 3506.645 3936.385 3506.925 3936.665 ;
        RECT 3507.355 3936.385 3507.635 3936.665 ;
        RECT 3508.065 3936.385 3508.345 3936.665 ;
        RECT 3508.775 3936.385 3509.055 3936.665 ;
        RECT 3509.485 3936.385 3509.765 3936.665 ;
        RECT 357.275 3935.955 357.555 3936.235 ;
        RECT 357.985 3935.955 358.265 3936.235 ;
        RECT 358.695 3935.955 358.975 3936.235 ;
        RECT 359.405 3935.955 359.685 3936.235 ;
        RECT 360.115 3935.955 360.395 3936.235 ;
        RECT 360.825 3935.955 361.105 3936.235 ;
        RECT 361.535 3935.955 361.815 3936.235 ;
        RECT 362.245 3935.955 362.525 3936.235 ;
        RECT 362.955 3935.955 363.235 3936.235 ;
        RECT 363.665 3935.955 363.945 3936.235 ;
        RECT 364.375 3935.955 364.655 3936.235 ;
        RECT 365.085 3935.955 365.365 3936.235 ;
        RECT 365.795 3935.955 366.075 3936.235 ;
        RECT 366.505 3935.955 366.785 3936.235 ;
        RECT 3500.255 3933.765 3500.535 3934.045 ;
        RECT 3500.965 3933.765 3501.245 3934.045 ;
        RECT 3501.675 3933.765 3501.955 3934.045 ;
        RECT 3502.385 3933.765 3502.665 3934.045 ;
        RECT 3503.095 3933.765 3503.375 3934.045 ;
        RECT 3503.805 3933.765 3504.085 3934.045 ;
        RECT 3504.515 3933.765 3504.795 3934.045 ;
        RECT 3505.225 3933.765 3505.505 3934.045 ;
        RECT 3505.935 3933.765 3506.215 3934.045 ;
        RECT 3506.645 3933.765 3506.925 3934.045 ;
        RECT 3507.355 3933.765 3507.635 3934.045 ;
        RECT 3508.065 3933.765 3508.345 3934.045 ;
        RECT 3508.775 3933.765 3509.055 3934.045 ;
        RECT 3509.485 3933.765 3509.765 3934.045 ;
        RECT 357.275 3933.335 357.555 3933.615 ;
        RECT 357.985 3933.335 358.265 3933.615 ;
        RECT 358.695 3933.335 358.975 3933.615 ;
        RECT 359.405 3933.335 359.685 3933.615 ;
        RECT 360.115 3933.335 360.395 3933.615 ;
        RECT 360.825 3933.335 361.105 3933.615 ;
        RECT 361.535 3933.335 361.815 3933.615 ;
        RECT 362.245 3933.335 362.525 3933.615 ;
        RECT 362.955 3933.335 363.235 3933.615 ;
        RECT 363.665 3933.335 363.945 3933.615 ;
        RECT 364.375 3933.335 364.655 3933.615 ;
        RECT 365.085 3933.335 365.365 3933.615 ;
        RECT 365.795 3933.335 366.075 3933.615 ;
        RECT 366.505 3933.335 366.785 3933.615 ;
        RECT 3500.255 3933.055 3500.535 3933.335 ;
        RECT 3500.965 3933.055 3501.245 3933.335 ;
        RECT 3501.675 3933.055 3501.955 3933.335 ;
        RECT 3502.385 3933.055 3502.665 3933.335 ;
        RECT 3503.095 3933.055 3503.375 3933.335 ;
        RECT 3503.805 3933.055 3504.085 3933.335 ;
        RECT 3504.515 3933.055 3504.795 3933.335 ;
        RECT 3505.225 3933.055 3505.505 3933.335 ;
        RECT 3505.935 3933.055 3506.215 3933.335 ;
        RECT 3506.645 3933.055 3506.925 3933.335 ;
        RECT 3507.355 3933.055 3507.635 3933.335 ;
        RECT 3508.065 3933.055 3508.345 3933.335 ;
        RECT 3508.775 3933.055 3509.055 3933.335 ;
        RECT 3509.485 3933.055 3509.765 3933.335 ;
        RECT 357.275 3932.625 357.555 3932.905 ;
        RECT 357.985 3932.625 358.265 3932.905 ;
        RECT 358.695 3932.625 358.975 3932.905 ;
        RECT 359.405 3932.625 359.685 3932.905 ;
        RECT 360.115 3932.625 360.395 3932.905 ;
        RECT 360.825 3932.625 361.105 3932.905 ;
        RECT 361.535 3932.625 361.815 3932.905 ;
        RECT 362.245 3932.625 362.525 3932.905 ;
        RECT 362.955 3932.625 363.235 3932.905 ;
        RECT 363.665 3932.625 363.945 3932.905 ;
        RECT 364.375 3932.625 364.655 3932.905 ;
        RECT 365.085 3932.625 365.365 3932.905 ;
        RECT 365.795 3932.625 366.075 3932.905 ;
        RECT 366.505 3932.625 366.785 3932.905 ;
        RECT 3500.255 3932.345 3500.535 3932.625 ;
        RECT 3500.965 3932.345 3501.245 3932.625 ;
        RECT 3501.675 3932.345 3501.955 3932.625 ;
        RECT 3502.385 3932.345 3502.665 3932.625 ;
        RECT 3503.095 3932.345 3503.375 3932.625 ;
        RECT 3503.805 3932.345 3504.085 3932.625 ;
        RECT 3504.515 3932.345 3504.795 3932.625 ;
        RECT 3505.225 3932.345 3505.505 3932.625 ;
        RECT 3505.935 3932.345 3506.215 3932.625 ;
        RECT 3506.645 3932.345 3506.925 3932.625 ;
        RECT 3507.355 3932.345 3507.635 3932.625 ;
        RECT 3508.065 3932.345 3508.345 3932.625 ;
        RECT 3508.775 3932.345 3509.055 3932.625 ;
        RECT 3509.485 3932.345 3509.765 3932.625 ;
        RECT 357.275 3931.915 357.555 3932.195 ;
        RECT 357.985 3931.915 358.265 3932.195 ;
        RECT 358.695 3931.915 358.975 3932.195 ;
        RECT 359.405 3931.915 359.685 3932.195 ;
        RECT 360.115 3931.915 360.395 3932.195 ;
        RECT 360.825 3931.915 361.105 3932.195 ;
        RECT 361.535 3931.915 361.815 3932.195 ;
        RECT 362.245 3931.915 362.525 3932.195 ;
        RECT 362.955 3931.915 363.235 3932.195 ;
        RECT 363.665 3931.915 363.945 3932.195 ;
        RECT 364.375 3931.915 364.655 3932.195 ;
        RECT 365.085 3931.915 365.365 3932.195 ;
        RECT 365.795 3931.915 366.075 3932.195 ;
        RECT 366.505 3931.915 366.785 3932.195 ;
        RECT 3500.255 3931.635 3500.535 3931.915 ;
        RECT 3500.965 3931.635 3501.245 3931.915 ;
        RECT 3501.675 3931.635 3501.955 3931.915 ;
        RECT 3502.385 3931.635 3502.665 3931.915 ;
        RECT 3503.095 3931.635 3503.375 3931.915 ;
        RECT 3503.805 3931.635 3504.085 3931.915 ;
        RECT 3504.515 3931.635 3504.795 3931.915 ;
        RECT 3505.225 3931.635 3505.505 3931.915 ;
        RECT 3505.935 3931.635 3506.215 3931.915 ;
        RECT 3506.645 3931.635 3506.925 3931.915 ;
        RECT 3507.355 3931.635 3507.635 3931.915 ;
        RECT 3508.065 3931.635 3508.345 3931.915 ;
        RECT 3508.775 3931.635 3509.055 3931.915 ;
        RECT 3509.485 3931.635 3509.765 3931.915 ;
        RECT 357.275 3931.205 357.555 3931.485 ;
        RECT 357.985 3931.205 358.265 3931.485 ;
        RECT 358.695 3931.205 358.975 3931.485 ;
        RECT 359.405 3931.205 359.685 3931.485 ;
        RECT 360.115 3931.205 360.395 3931.485 ;
        RECT 360.825 3931.205 361.105 3931.485 ;
        RECT 361.535 3931.205 361.815 3931.485 ;
        RECT 362.245 3931.205 362.525 3931.485 ;
        RECT 362.955 3931.205 363.235 3931.485 ;
        RECT 363.665 3931.205 363.945 3931.485 ;
        RECT 364.375 3931.205 364.655 3931.485 ;
        RECT 365.085 3931.205 365.365 3931.485 ;
        RECT 365.795 3931.205 366.075 3931.485 ;
        RECT 366.505 3931.205 366.785 3931.485 ;
        RECT 3500.255 3930.925 3500.535 3931.205 ;
        RECT 3500.965 3930.925 3501.245 3931.205 ;
        RECT 3501.675 3930.925 3501.955 3931.205 ;
        RECT 3502.385 3930.925 3502.665 3931.205 ;
        RECT 3503.095 3930.925 3503.375 3931.205 ;
        RECT 3503.805 3930.925 3504.085 3931.205 ;
        RECT 3504.515 3930.925 3504.795 3931.205 ;
        RECT 3505.225 3930.925 3505.505 3931.205 ;
        RECT 3505.935 3930.925 3506.215 3931.205 ;
        RECT 3506.645 3930.925 3506.925 3931.205 ;
        RECT 3507.355 3930.925 3507.635 3931.205 ;
        RECT 3508.065 3930.925 3508.345 3931.205 ;
        RECT 3508.775 3930.925 3509.055 3931.205 ;
        RECT 3509.485 3930.925 3509.765 3931.205 ;
        RECT 357.275 3930.495 357.555 3930.775 ;
        RECT 357.985 3930.495 358.265 3930.775 ;
        RECT 358.695 3930.495 358.975 3930.775 ;
        RECT 359.405 3930.495 359.685 3930.775 ;
        RECT 360.115 3930.495 360.395 3930.775 ;
        RECT 360.825 3930.495 361.105 3930.775 ;
        RECT 361.535 3930.495 361.815 3930.775 ;
        RECT 362.245 3930.495 362.525 3930.775 ;
        RECT 362.955 3930.495 363.235 3930.775 ;
        RECT 363.665 3930.495 363.945 3930.775 ;
        RECT 364.375 3930.495 364.655 3930.775 ;
        RECT 365.085 3930.495 365.365 3930.775 ;
        RECT 365.795 3930.495 366.075 3930.775 ;
        RECT 366.505 3930.495 366.785 3930.775 ;
        RECT 3500.255 3930.215 3500.535 3930.495 ;
        RECT 3500.965 3930.215 3501.245 3930.495 ;
        RECT 3501.675 3930.215 3501.955 3930.495 ;
        RECT 3502.385 3930.215 3502.665 3930.495 ;
        RECT 3503.095 3930.215 3503.375 3930.495 ;
        RECT 3503.805 3930.215 3504.085 3930.495 ;
        RECT 3504.515 3930.215 3504.795 3930.495 ;
        RECT 3505.225 3930.215 3505.505 3930.495 ;
        RECT 3505.935 3930.215 3506.215 3930.495 ;
        RECT 3506.645 3930.215 3506.925 3930.495 ;
        RECT 3507.355 3930.215 3507.635 3930.495 ;
        RECT 3508.065 3930.215 3508.345 3930.495 ;
        RECT 3508.775 3930.215 3509.055 3930.495 ;
        RECT 3509.485 3930.215 3509.765 3930.495 ;
        RECT 357.275 3929.785 357.555 3930.065 ;
        RECT 357.985 3929.785 358.265 3930.065 ;
        RECT 358.695 3929.785 358.975 3930.065 ;
        RECT 359.405 3929.785 359.685 3930.065 ;
        RECT 360.115 3929.785 360.395 3930.065 ;
        RECT 360.825 3929.785 361.105 3930.065 ;
        RECT 361.535 3929.785 361.815 3930.065 ;
        RECT 362.245 3929.785 362.525 3930.065 ;
        RECT 362.955 3929.785 363.235 3930.065 ;
        RECT 363.665 3929.785 363.945 3930.065 ;
        RECT 364.375 3929.785 364.655 3930.065 ;
        RECT 365.085 3929.785 365.365 3930.065 ;
        RECT 365.795 3929.785 366.075 3930.065 ;
        RECT 366.505 3929.785 366.785 3930.065 ;
        RECT 3500.255 3929.505 3500.535 3929.785 ;
        RECT 3500.965 3929.505 3501.245 3929.785 ;
        RECT 3501.675 3929.505 3501.955 3929.785 ;
        RECT 3502.385 3929.505 3502.665 3929.785 ;
        RECT 3503.095 3929.505 3503.375 3929.785 ;
        RECT 3503.805 3929.505 3504.085 3929.785 ;
        RECT 3504.515 3929.505 3504.795 3929.785 ;
        RECT 3505.225 3929.505 3505.505 3929.785 ;
        RECT 3505.935 3929.505 3506.215 3929.785 ;
        RECT 3506.645 3929.505 3506.925 3929.785 ;
        RECT 3507.355 3929.505 3507.635 3929.785 ;
        RECT 3508.065 3929.505 3508.345 3929.785 ;
        RECT 3508.775 3929.505 3509.055 3929.785 ;
        RECT 3509.485 3929.505 3509.765 3929.785 ;
        RECT 357.275 3929.075 357.555 3929.355 ;
        RECT 357.985 3929.075 358.265 3929.355 ;
        RECT 358.695 3929.075 358.975 3929.355 ;
        RECT 359.405 3929.075 359.685 3929.355 ;
        RECT 360.115 3929.075 360.395 3929.355 ;
        RECT 360.825 3929.075 361.105 3929.355 ;
        RECT 361.535 3929.075 361.815 3929.355 ;
        RECT 362.245 3929.075 362.525 3929.355 ;
        RECT 362.955 3929.075 363.235 3929.355 ;
        RECT 363.665 3929.075 363.945 3929.355 ;
        RECT 364.375 3929.075 364.655 3929.355 ;
        RECT 365.085 3929.075 365.365 3929.355 ;
        RECT 365.795 3929.075 366.075 3929.355 ;
        RECT 366.505 3929.075 366.785 3929.355 ;
        RECT 3500.255 3928.795 3500.535 3929.075 ;
        RECT 3500.965 3928.795 3501.245 3929.075 ;
        RECT 3501.675 3928.795 3501.955 3929.075 ;
        RECT 3502.385 3928.795 3502.665 3929.075 ;
        RECT 3503.095 3928.795 3503.375 3929.075 ;
        RECT 3503.805 3928.795 3504.085 3929.075 ;
        RECT 3504.515 3928.795 3504.795 3929.075 ;
        RECT 3505.225 3928.795 3505.505 3929.075 ;
        RECT 3505.935 3928.795 3506.215 3929.075 ;
        RECT 3506.645 3928.795 3506.925 3929.075 ;
        RECT 3507.355 3928.795 3507.635 3929.075 ;
        RECT 3508.065 3928.795 3508.345 3929.075 ;
        RECT 3508.775 3928.795 3509.055 3929.075 ;
        RECT 3509.485 3928.795 3509.765 3929.075 ;
        RECT 357.275 3928.365 357.555 3928.645 ;
        RECT 357.985 3928.365 358.265 3928.645 ;
        RECT 358.695 3928.365 358.975 3928.645 ;
        RECT 359.405 3928.365 359.685 3928.645 ;
        RECT 360.115 3928.365 360.395 3928.645 ;
        RECT 360.825 3928.365 361.105 3928.645 ;
        RECT 361.535 3928.365 361.815 3928.645 ;
        RECT 362.245 3928.365 362.525 3928.645 ;
        RECT 362.955 3928.365 363.235 3928.645 ;
        RECT 363.665 3928.365 363.945 3928.645 ;
        RECT 364.375 3928.365 364.655 3928.645 ;
        RECT 365.085 3928.365 365.365 3928.645 ;
        RECT 365.795 3928.365 366.075 3928.645 ;
        RECT 366.505 3928.365 366.785 3928.645 ;
        RECT 3500.255 3928.085 3500.535 3928.365 ;
        RECT 3500.965 3928.085 3501.245 3928.365 ;
        RECT 3501.675 3928.085 3501.955 3928.365 ;
        RECT 3502.385 3928.085 3502.665 3928.365 ;
        RECT 3503.095 3928.085 3503.375 3928.365 ;
        RECT 3503.805 3928.085 3504.085 3928.365 ;
        RECT 3504.515 3928.085 3504.795 3928.365 ;
        RECT 3505.225 3928.085 3505.505 3928.365 ;
        RECT 3505.935 3928.085 3506.215 3928.365 ;
        RECT 3506.645 3928.085 3506.925 3928.365 ;
        RECT 3507.355 3928.085 3507.635 3928.365 ;
        RECT 3508.065 3928.085 3508.345 3928.365 ;
        RECT 3508.775 3928.085 3509.055 3928.365 ;
        RECT 3509.485 3928.085 3509.765 3928.365 ;
        RECT 357.275 3927.655 357.555 3927.935 ;
        RECT 357.985 3927.655 358.265 3927.935 ;
        RECT 358.695 3927.655 358.975 3927.935 ;
        RECT 359.405 3927.655 359.685 3927.935 ;
        RECT 360.115 3927.655 360.395 3927.935 ;
        RECT 360.825 3927.655 361.105 3927.935 ;
        RECT 361.535 3927.655 361.815 3927.935 ;
        RECT 362.245 3927.655 362.525 3927.935 ;
        RECT 362.955 3927.655 363.235 3927.935 ;
        RECT 363.665 3927.655 363.945 3927.935 ;
        RECT 364.375 3927.655 364.655 3927.935 ;
        RECT 365.085 3927.655 365.365 3927.935 ;
        RECT 365.795 3927.655 366.075 3927.935 ;
        RECT 366.505 3927.655 366.785 3927.935 ;
        RECT 3500.255 3927.375 3500.535 3927.655 ;
        RECT 3500.965 3927.375 3501.245 3927.655 ;
        RECT 3501.675 3927.375 3501.955 3927.655 ;
        RECT 3502.385 3927.375 3502.665 3927.655 ;
        RECT 3503.095 3927.375 3503.375 3927.655 ;
        RECT 3503.805 3927.375 3504.085 3927.655 ;
        RECT 3504.515 3927.375 3504.795 3927.655 ;
        RECT 3505.225 3927.375 3505.505 3927.655 ;
        RECT 3505.935 3927.375 3506.215 3927.655 ;
        RECT 3506.645 3927.375 3506.925 3927.655 ;
        RECT 3507.355 3927.375 3507.635 3927.655 ;
        RECT 3508.065 3927.375 3508.345 3927.655 ;
        RECT 3508.775 3927.375 3509.055 3927.655 ;
        RECT 3509.485 3927.375 3509.765 3927.655 ;
        RECT 357.275 3926.945 357.555 3927.225 ;
        RECT 357.985 3926.945 358.265 3927.225 ;
        RECT 358.695 3926.945 358.975 3927.225 ;
        RECT 359.405 3926.945 359.685 3927.225 ;
        RECT 360.115 3926.945 360.395 3927.225 ;
        RECT 360.825 3926.945 361.105 3927.225 ;
        RECT 361.535 3926.945 361.815 3927.225 ;
        RECT 362.245 3926.945 362.525 3927.225 ;
        RECT 362.955 3926.945 363.235 3927.225 ;
        RECT 363.665 3926.945 363.945 3927.225 ;
        RECT 364.375 3926.945 364.655 3927.225 ;
        RECT 365.085 3926.945 365.365 3927.225 ;
        RECT 365.795 3926.945 366.075 3927.225 ;
        RECT 366.505 3926.945 366.785 3927.225 ;
        RECT 3500.255 3926.665 3500.535 3926.945 ;
        RECT 3500.965 3926.665 3501.245 3926.945 ;
        RECT 3501.675 3926.665 3501.955 3926.945 ;
        RECT 3502.385 3926.665 3502.665 3926.945 ;
        RECT 3503.095 3926.665 3503.375 3926.945 ;
        RECT 3503.805 3926.665 3504.085 3926.945 ;
        RECT 3504.515 3926.665 3504.795 3926.945 ;
        RECT 3505.225 3926.665 3505.505 3926.945 ;
        RECT 3505.935 3926.665 3506.215 3926.945 ;
        RECT 3506.645 3926.665 3506.925 3926.945 ;
        RECT 3507.355 3926.665 3507.635 3926.945 ;
        RECT 3508.065 3926.665 3508.345 3926.945 ;
        RECT 3508.775 3926.665 3509.055 3926.945 ;
        RECT 3509.485 3926.665 3509.765 3926.945 ;
        RECT 357.275 3926.235 357.555 3926.515 ;
        RECT 357.985 3926.235 358.265 3926.515 ;
        RECT 358.695 3926.235 358.975 3926.515 ;
        RECT 359.405 3926.235 359.685 3926.515 ;
        RECT 360.115 3926.235 360.395 3926.515 ;
        RECT 360.825 3926.235 361.105 3926.515 ;
        RECT 361.535 3926.235 361.815 3926.515 ;
        RECT 362.245 3926.235 362.525 3926.515 ;
        RECT 362.955 3926.235 363.235 3926.515 ;
        RECT 363.665 3926.235 363.945 3926.515 ;
        RECT 364.375 3926.235 364.655 3926.515 ;
        RECT 365.085 3926.235 365.365 3926.515 ;
        RECT 365.795 3926.235 366.075 3926.515 ;
        RECT 366.505 3926.235 366.785 3926.515 ;
        RECT 3500.255 3925.955 3500.535 3926.235 ;
        RECT 3500.965 3925.955 3501.245 3926.235 ;
        RECT 3501.675 3925.955 3501.955 3926.235 ;
        RECT 3502.385 3925.955 3502.665 3926.235 ;
        RECT 3503.095 3925.955 3503.375 3926.235 ;
        RECT 3503.805 3925.955 3504.085 3926.235 ;
        RECT 3504.515 3925.955 3504.795 3926.235 ;
        RECT 3505.225 3925.955 3505.505 3926.235 ;
        RECT 3505.935 3925.955 3506.215 3926.235 ;
        RECT 3506.645 3925.955 3506.925 3926.235 ;
        RECT 3507.355 3925.955 3507.635 3926.235 ;
        RECT 3508.065 3925.955 3508.345 3926.235 ;
        RECT 3508.775 3925.955 3509.055 3926.235 ;
        RECT 3509.485 3925.955 3509.765 3926.235 ;
        RECT 357.275 3925.525 357.555 3925.805 ;
        RECT 357.985 3925.525 358.265 3925.805 ;
        RECT 358.695 3925.525 358.975 3925.805 ;
        RECT 359.405 3925.525 359.685 3925.805 ;
        RECT 360.115 3925.525 360.395 3925.805 ;
        RECT 360.825 3925.525 361.105 3925.805 ;
        RECT 361.535 3925.525 361.815 3925.805 ;
        RECT 362.245 3925.525 362.525 3925.805 ;
        RECT 362.955 3925.525 363.235 3925.805 ;
        RECT 363.665 3925.525 363.945 3925.805 ;
        RECT 364.375 3925.525 364.655 3925.805 ;
        RECT 365.085 3925.525 365.365 3925.805 ;
        RECT 365.795 3925.525 366.075 3925.805 ;
        RECT 366.505 3925.525 366.785 3925.805 ;
        RECT 3500.255 3925.245 3500.535 3925.525 ;
        RECT 3500.965 3925.245 3501.245 3925.525 ;
        RECT 3501.675 3925.245 3501.955 3925.525 ;
        RECT 3502.385 3925.245 3502.665 3925.525 ;
        RECT 3503.095 3925.245 3503.375 3925.525 ;
        RECT 3503.805 3925.245 3504.085 3925.525 ;
        RECT 3504.515 3925.245 3504.795 3925.525 ;
        RECT 3505.225 3925.245 3505.505 3925.525 ;
        RECT 3505.935 3925.245 3506.215 3925.525 ;
        RECT 3506.645 3925.245 3506.925 3925.525 ;
        RECT 3507.355 3925.245 3507.635 3925.525 ;
        RECT 3508.065 3925.245 3508.345 3925.525 ;
        RECT 3508.775 3925.245 3509.055 3925.525 ;
        RECT 3509.485 3925.245 3509.765 3925.525 ;
        RECT 357.275 3924.815 357.555 3925.095 ;
        RECT 357.985 3924.815 358.265 3925.095 ;
        RECT 358.695 3924.815 358.975 3925.095 ;
        RECT 359.405 3924.815 359.685 3925.095 ;
        RECT 360.115 3924.815 360.395 3925.095 ;
        RECT 360.825 3924.815 361.105 3925.095 ;
        RECT 361.535 3924.815 361.815 3925.095 ;
        RECT 362.245 3924.815 362.525 3925.095 ;
        RECT 362.955 3924.815 363.235 3925.095 ;
        RECT 363.665 3924.815 363.945 3925.095 ;
        RECT 364.375 3924.815 364.655 3925.095 ;
        RECT 365.085 3924.815 365.365 3925.095 ;
        RECT 365.795 3924.815 366.075 3925.095 ;
        RECT 366.505 3924.815 366.785 3925.095 ;
        RECT 3500.255 3924.535 3500.535 3924.815 ;
        RECT 3500.965 3924.535 3501.245 3924.815 ;
        RECT 3501.675 3924.535 3501.955 3924.815 ;
        RECT 3502.385 3924.535 3502.665 3924.815 ;
        RECT 3503.095 3924.535 3503.375 3924.815 ;
        RECT 3503.805 3924.535 3504.085 3924.815 ;
        RECT 3504.515 3924.535 3504.795 3924.815 ;
        RECT 3505.225 3924.535 3505.505 3924.815 ;
        RECT 3505.935 3924.535 3506.215 3924.815 ;
        RECT 3506.645 3924.535 3506.925 3924.815 ;
        RECT 3507.355 3924.535 3507.635 3924.815 ;
        RECT 3508.065 3924.535 3508.345 3924.815 ;
        RECT 3508.775 3924.535 3509.055 3924.815 ;
        RECT 3509.485 3924.535 3509.765 3924.815 ;
        RECT 357.275 3924.105 357.555 3924.385 ;
        RECT 357.985 3924.105 358.265 3924.385 ;
        RECT 358.695 3924.105 358.975 3924.385 ;
        RECT 359.405 3924.105 359.685 3924.385 ;
        RECT 360.115 3924.105 360.395 3924.385 ;
        RECT 360.825 3924.105 361.105 3924.385 ;
        RECT 361.535 3924.105 361.815 3924.385 ;
        RECT 362.245 3924.105 362.525 3924.385 ;
        RECT 362.955 3924.105 363.235 3924.385 ;
        RECT 363.665 3924.105 363.945 3924.385 ;
        RECT 364.375 3924.105 364.655 3924.385 ;
        RECT 365.085 3924.105 365.365 3924.385 ;
        RECT 365.795 3924.105 366.075 3924.385 ;
        RECT 366.505 3924.105 366.785 3924.385 ;
        RECT 357.330 3920.190 357.610 3920.470 ;
        RECT 358.040 3920.190 358.320 3920.470 ;
        RECT 358.750 3920.190 359.030 3920.470 ;
        RECT 359.460 3920.190 359.740 3920.470 ;
        RECT 360.170 3920.190 360.450 3920.470 ;
        RECT 360.880 3920.190 361.160 3920.470 ;
        RECT 361.590 3920.190 361.870 3920.470 ;
        RECT 362.300 3920.190 362.580 3920.470 ;
        RECT 363.010 3920.190 363.290 3920.470 ;
        RECT 363.720 3920.190 364.000 3920.470 ;
        RECT 364.430 3920.190 364.710 3920.470 ;
        RECT 365.140 3920.190 365.420 3920.470 ;
        RECT 365.850 3920.190 366.130 3920.470 ;
        RECT 366.560 3920.190 366.840 3920.470 ;
        RECT 3500.255 3920.235 3500.535 3920.515 ;
        RECT 3500.965 3920.235 3501.245 3920.515 ;
        RECT 3501.675 3920.235 3501.955 3920.515 ;
        RECT 3502.385 3920.235 3502.665 3920.515 ;
        RECT 3503.095 3920.235 3503.375 3920.515 ;
        RECT 3503.805 3920.235 3504.085 3920.515 ;
        RECT 3504.515 3920.235 3504.795 3920.515 ;
        RECT 3505.225 3920.235 3505.505 3920.515 ;
        RECT 3505.935 3920.235 3506.215 3920.515 ;
        RECT 3506.645 3920.235 3506.925 3920.515 ;
        RECT 3507.355 3920.235 3507.635 3920.515 ;
        RECT 3508.065 3920.235 3508.345 3920.515 ;
        RECT 3508.775 3920.235 3509.055 3920.515 ;
        RECT 3509.485 3920.235 3509.765 3920.515 ;
        RECT 357.330 3919.480 357.610 3919.760 ;
        RECT 358.040 3919.480 358.320 3919.760 ;
        RECT 358.750 3919.480 359.030 3919.760 ;
        RECT 359.460 3919.480 359.740 3919.760 ;
        RECT 360.170 3919.480 360.450 3919.760 ;
        RECT 360.880 3919.480 361.160 3919.760 ;
        RECT 361.590 3919.480 361.870 3919.760 ;
        RECT 362.300 3919.480 362.580 3919.760 ;
        RECT 363.010 3919.480 363.290 3919.760 ;
        RECT 363.720 3919.480 364.000 3919.760 ;
        RECT 364.430 3919.480 364.710 3919.760 ;
        RECT 365.140 3919.480 365.420 3919.760 ;
        RECT 365.850 3919.480 366.130 3919.760 ;
        RECT 366.560 3919.480 366.840 3919.760 ;
        RECT 3500.255 3919.525 3500.535 3919.805 ;
        RECT 3500.965 3919.525 3501.245 3919.805 ;
        RECT 3501.675 3919.525 3501.955 3919.805 ;
        RECT 3502.385 3919.525 3502.665 3919.805 ;
        RECT 3503.095 3919.525 3503.375 3919.805 ;
        RECT 3503.805 3919.525 3504.085 3919.805 ;
        RECT 3504.515 3919.525 3504.795 3919.805 ;
        RECT 3505.225 3919.525 3505.505 3919.805 ;
        RECT 3505.935 3919.525 3506.215 3919.805 ;
        RECT 3506.645 3919.525 3506.925 3919.805 ;
        RECT 3507.355 3919.525 3507.635 3919.805 ;
        RECT 3508.065 3919.525 3508.345 3919.805 ;
        RECT 3508.775 3919.525 3509.055 3919.805 ;
        RECT 3509.485 3919.525 3509.765 3919.805 ;
        RECT 357.330 3918.770 357.610 3919.050 ;
        RECT 358.040 3918.770 358.320 3919.050 ;
        RECT 358.750 3918.770 359.030 3919.050 ;
        RECT 359.460 3918.770 359.740 3919.050 ;
        RECT 360.170 3918.770 360.450 3919.050 ;
        RECT 360.880 3918.770 361.160 3919.050 ;
        RECT 361.590 3918.770 361.870 3919.050 ;
        RECT 362.300 3918.770 362.580 3919.050 ;
        RECT 363.010 3918.770 363.290 3919.050 ;
        RECT 363.720 3918.770 364.000 3919.050 ;
        RECT 364.430 3918.770 364.710 3919.050 ;
        RECT 365.140 3918.770 365.420 3919.050 ;
        RECT 365.850 3918.770 366.130 3919.050 ;
        RECT 366.560 3918.770 366.840 3919.050 ;
        RECT 3500.255 3918.815 3500.535 3919.095 ;
        RECT 3500.965 3918.815 3501.245 3919.095 ;
        RECT 3501.675 3918.815 3501.955 3919.095 ;
        RECT 3502.385 3918.815 3502.665 3919.095 ;
        RECT 3503.095 3918.815 3503.375 3919.095 ;
        RECT 3503.805 3918.815 3504.085 3919.095 ;
        RECT 3504.515 3918.815 3504.795 3919.095 ;
        RECT 3505.225 3918.815 3505.505 3919.095 ;
        RECT 3505.935 3918.815 3506.215 3919.095 ;
        RECT 3506.645 3918.815 3506.925 3919.095 ;
        RECT 3507.355 3918.815 3507.635 3919.095 ;
        RECT 3508.065 3918.815 3508.345 3919.095 ;
        RECT 3508.775 3918.815 3509.055 3919.095 ;
        RECT 3509.485 3918.815 3509.765 3919.095 ;
        RECT 357.330 3918.060 357.610 3918.340 ;
        RECT 358.040 3918.060 358.320 3918.340 ;
        RECT 358.750 3918.060 359.030 3918.340 ;
        RECT 359.460 3918.060 359.740 3918.340 ;
        RECT 360.170 3918.060 360.450 3918.340 ;
        RECT 360.880 3918.060 361.160 3918.340 ;
        RECT 361.590 3918.060 361.870 3918.340 ;
        RECT 362.300 3918.060 362.580 3918.340 ;
        RECT 363.010 3918.060 363.290 3918.340 ;
        RECT 363.720 3918.060 364.000 3918.340 ;
        RECT 364.430 3918.060 364.710 3918.340 ;
        RECT 365.140 3918.060 365.420 3918.340 ;
        RECT 365.850 3918.060 366.130 3918.340 ;
        RECT 366.560 3918.060 366.840 3918.340 ;
        RECT 3500.255 3918.105 3500.535 3918.385 ;
        RECT 3500.965 3918.105 3501.245 3918.385 ;
        RECT 3501.675 3918.105 3501.955 3918.385 ;
        RECT 3502.385 3918.105 3502.665 3918.385 ;
        RECT 3503.095 3918.105 3503.375 3918.385 ;
        RECT 3503.805 3918.105 3504.085 3918.385 ;
        RECT 3504.515 3918.105 3504.795 3918.385 ;
        RECT 3505.225 3918.105 3505.505 3918.385 ;
        RECT 3505.935 3918.105 3506.215 3918.385 ;
        RECT 3506.645 3918.105 3506.925 3918.385 ;
        RECT 3507.355 3918.105 3507.635 3918.385 ;
        RECT 3508.065 3918.105 3508.345 3918.385 ;
        RECT 3508.775 3918.105 3509.055 3918.385 ;
        RECT 3509.485 3918.105 3509.765 3918.385 ;
        RECT 357.330 3917.350 357.610 3917.630 ;
        RECT 358.040 3917.350 358.320 3917.630 ;
        RECT 358.750 3917.350 359.030 3917.630 ;
        RECT 359.460 3917.350 359.740 3917.630 ;
        RECT 360.170 3917.350 360.450 3917.630 ;
        RECT 360.880 3917.350 361.160 3917.630 ;
        RECT 361.590 3917.350 361.870 3917.630 ;
        RECT 362.300 3917.350 362.580 3917.630 ;
        RECT 363.010 3917.350 363.290 3917.630 ;
        RECT 363.720 3917.350 364.000 3917.630 ;
        RECT 364.430 3917.350 364.710 3917.630 ;
        RECT 365.140 3917.350 365.420 3917.630 ;
        RECT 365.850 3917.350 366.130 3917.630 ;
        RECT 366.560 3917.350 366.840 3917.630 ;
        RECT 3500.255 3917.395 3500.535 3917.675 ;
        RECT 3500.965 3917.395 3501.245 3917.675 ;
        RECT 3501.675 3917.395 3501.955 3917.675 ;
        RECT 3502.385 3917.395 3502.665 3917.675 ;
        RECT 3503.095 3917.395 3503.375 3917.675 ;
        RECT 3503.805 3917.395 3504.085 3917.675 ;
        RECT 3504.515 3917.395 3504.795 3917.675 ;
        RECT 3505.225 3917.395 3505.505 3917.675 ;
        RECT 3505.935 3917.395 3506.215 3917.675 ;
        RECT 3506.645 3917.395 3506.925 3917.675 ;
        RECT 3507.355 3917.395 3507.635 3917.675 ;
        RECT 3508.065 3917.395 3508.345 3917.675 ;
        RECT 3508.775 3917.395 3509.055 3917.675 ;
        RECT 3509.485 3917.395 3509.765 3917.675 ;
        RECT 357.330 3916.640 357.610 3916.920 ;
        RECT 358.040 3916.640 358.320 3916.920 ;
        RECT 358.750 3916.640 359.030 3916.920 ;
        RECT 359.460 3916.640 359.740 3916.920 ;
        RECT 360.170 3916.640 360.450 3916.920 ;
        RECT 360.880 3916.640 361.160 3916.920 ;
        RECT 361.590 3916.640 361.870 3916.920 ;
        RECT 362.300 3916.640 362.580 3916.920 ;
        RECT 363.010 3916.640 363.290 3916.920 ;
        RECT 363.720 3916.640 364.000 3916.920 ;
        RECT 364.430 3916.640 364.710 3916.920 ;
        RECT 365.140 3916.640 365.420 3916.920 ;
        RECT 365.850 3916.640 366.130 3916.920 ;
        RECT 366.560 3916.640 366.840 3916.920 ;
        RECT 3500.255 3916.685 3500.535 3916.965 ;
        RECT 3500.965 3916.685 3501.245 3916.965 ;
        RECT 3501.675 3916.685 3501.955 3916.965 ;
        RECT 3502.385 3916.685 3502.665 3916.965 ;
        RECT 3503.095 3916.685 3503.375 3916.965 ;
        RECT 3503.805 3916.685 3504.085 3916.965 ;
        RECT 3504.515 3916.685 3504.795 3916.965 ;
        RECT 3505.225 3916.685 3505.505 3916.965 ;
        RECT 3505.935 3916.685 3506.215 3916.965 ;
        RECT 3506.645 3916.685 3506.925 3916.965 ;
        RECT 3507.355 3916.685 3507.635 3916.965 ;
        RECT 3508.065 3916.685 3508.345 3916.965 ;
        RECT 3508.775 3916.685 3509.055 3916.965 ;
        RECT 3509.485 3916.685 3509.765 3916.965 ;
        RECT 357.330 3915.930 357.610 3916.210 ;
        RECT 358.040 3915.930 358.320 3916.210 ;
        RECT 358.750 3915.930 359.030 3916.210 ;
        RECT 359.460 3915.930 359.740 3916.210 ;
        RECT 360.170 3915.930 360.450 3916.210 ;
        RECT 360.880 3915.930 361.160 3916.210 ;
        RECT 361.590 3915.930 361.870 3916.210 ;
        RECT 362.300 3915.930 362.580 3916.210 ;
        RECT 363.010 3915.930 363.290 3916.210 ;
        RECT 363.720 3915.930 364.000 3916.210 ;
        RECT 364.430 3915.930 364.710 3916.210 ;
        RECT 365.140 3915.930 365.420 3916.210 ;
        RECT 365.850 3915.930 366.130 3916.210 ;
        RECT 366.560 3915.930 366.840 3916.210 ;
        RECT 3500.255 3915.975 3500.535 3916.255 ;
        RECT 3500.965 3915.975 3501.245 3916.255 ;
        RECT 3501.675 3915.975 3501.955 3916.255 ;
        RECT 3502.385 3915.975 3502.665 3916.255 ;
        RECT 3503.095 3915.975 3503.375 3916.255 ;
        RECT 3503.805 3915.975 3504.085 3916.255 ;
        RECT 3504.515 3915.975 3504.795 3916.255 ;
        RECT 3505.225 3915.975 3505.505 3916.255 ;
        RECT 3505.935 3915.975 3506.215 3916.255 ;
        RECT 3506.645 3915.975 3506.925 3916.255 ;
        RECT 3507.355 3915.975 3507.635 3916.255 ;
        RECT 3508.065 3915.975 3508.345 3916.255 ;
        RECT 3508.775 3915.975 3509.055 3916.255 ;
        RECT 3509.485 3915.975 3509.765 3916.255 ;
        RECT 357.330 3915.220 357.610 3915.500 ;
        RECT 358.040 3915.220 358.320 3915.500 ;
        RECT 358.750 3915.220 359.030 3915.500 ;
        RECT 359.460 3915.220 359.740 3915.500 ;
        RECT 360.170 3915.220 360.450 3915.500 ;
        RECT 360.880 3915.220 361.160 3915.500 ;
        RECT 361.590 3915.220 361.870 3915.500 ;
        RECT 362.300 3915.220 362.580 3915.500 ;
        RECT 363.010 3915.220 363.290 3915.500 ;
        RECT 363.720 3915.220 364.000 3915.500 ;
        RECT 364.430 3915.220 364.710 3915.500 ;
        RECT 365.140 3915.220 365.420 3915.500 ;
        RECT 365.850 3915.220 366.130 3915.500 ;
        RECT 366.560 3915.220 366.840 3915.500 ;
        RECT 3500.255 3915.265 3500.535 3915.545 ;
        RECT 3500.965 3915.265 3501.245 3915.545 ;
        RECT 3501.675 3915.265 3501.955 3915.545 ;
        RECT 3502.385 3915.265 3502.665 3915.545 ;
        RECT 3503.095 3915.265 3503.375 3915.545 ;
        RECT 3503.805 3915.265 3504.085 3915.545 ;
        RECT 3504.515 3915.265 3504.795 3915.545 ;
        RECT 3505.225 3915.265 3505.505 3915.545 ;
        RECT 3505.935 3915.265 3506.215 3915.545 ;
        RECT 3506.645 3915.265 3506.925 3915.545 ;
        RECT 3507.355 3915.265 3507.635 3915.545 ;
        RECT 3508.065 3915.265 3508.345 3915.545 ;
        RECT 3508.775 3915.265 3509.055 3915.545 ;
        RECT 3509.485 3915.265 3509.765 3915.545 ;
        RECT 357.330 3914.510 357.610 3914.790 ;
        RECT 358.040 3914.510 358.320 3914.790 ;
        RECT 358.750 3914.510 359.030 3914.790 ;
        RECT 359.460 3914.510 359.740 3914.790 ;
        RECT 360.170 3914.510 360.450 3914.790 ;
        RECT 360.880 3914.510 361.160 3914.790 ;
        RECT 361.590 3914.510 361.870 3914.790 ;
        RECT 362.300 3914.510 362.580 3914.790 ;
        RECT 363.010 3914.510 363.290 3914.790 ;
        RECT 363.720 3914.510 364.000 3914.790 ;
        RECT 364.430 3914.510 364.710 3914.790 ;
        RECT 365.140 3914.510 365.420 3914.790 ;
        RECT 365.850 3914.510 366.130 3914.790 ;
        RECT 366.560 3914.510 366.840 3914.790 ;
        RECT 3500.255 3914.555 3500.535 3914.835 ;
        RECT 3500.965 3914.555 3501.245 3914.835 ;
        RECT 3501.675 3914.555 3501.955 3914.835 ;
        RECT 3502.385 3914.555 3502.665 3914.835 ;
        RECT 3503.095 3914.555 3503.375 3914.835 ;
        RECT 3503.805 3914.555 3504.085 3914.835 ;
        RECT 3504.515 3914.555 3504.795 3914.835 ;
        RECT 3505.225 3914.555 3505.505 3914.835 ;
        RECT 3505.935 3914.555 3506.215 3914.835 ;
        RECT 3506.645 3914.555 3506.925 3914.835 ;
        RECT 3507.355 3914.555 3507.635 3914.835 ;
        RECT 3508.065 3914.555 3508.345 3914.835 ;
        RECT 3508.775 3914.555 3509.055 3914.835 ;
        RECT 3509.485 3914.555 3509.765 3914.835 ;
        RECT 357.330 3913.800 357.610 3914.080 ;
        RECT 358.040 3913.800 358.320 3914.080 ;
        RECT 358.750 3913.800 359.030 3914.080 ;
        RECT 359.460 3913.800 359.740 3914.080 ;
        RECT 360.170 3913.800 360.450 3914.080 ;
        RECT 360.880 3913.800 361.160 3914.080 ;
        RECT 361.590 3913.800 361.870 3914.080 ;
        RECT 362.300 3913.800 362.580 3914.080 ;
        RECT 363.010 3913.800 363.290 3914.080 ;
        RECT 363.720 3913.800 364.000 3914.080 ;
        RECT 364.430 3913.800 364.710 3914.080 ;
        RECT 365.140 3913.800 365.420 3914.080 ;
        RECT 365.850 3913.800 366.130 3914.080 ;
        RECT 366.560 3913.800 366.840 3914.080 ;
        RECT 3500.255 3913.845 3500.535 3914.125 ;
        RECT 3500.965 3913.845 3501.245 3914.125 ;
        RECT 3501.675 3913.845 3501.955 3914.125 ;
        RECT 3502.385 3913.845 3502.665 3914.125 ;
        RECT 3503.095 3913.845 3503.375 3914.125 ;
        RECT 3503.805 3913.845 3504.085 3914.125 ;
        RECT 3504.515 3913.845 3504.795 3914.125 ;
        RECT 3505.225 3913.845 3505.505 3914.125 ;
        RECT 3505.935 3913.845 3506.215 3914.125 ;
        RECT 3506.645 3913.845 3506.925 3914.125 ;
        RECT 3507.355 3913.845 3507.635 3914.125 ;
        RECT 3508.065 3913.845 3508.345 3914.125 ;
        RECT 3508.775 3913.845 3509.055 3914.125 ;
        RECT 3509.485 3913.845 3509.765 3914.125 ;
        RECT 357.330 3913.090 357.610 3913.370 ;
        RECT 358.040 3913.090 358.320 3913.370 ;
        RECT 358.750 3913.090 359.030 3913.370 ;
        RECT 359.460 3913.090 359.740 3913.370 ;
        RECT 360.170 3913.090 360.450 3913.370 ;
        RECT 360.880 3913.090 361.160 3913.370 ;
        RECT 361.590 3913.090 361.870 3913.370 ;
        RECT 362.300 3913.090 362.580 3913.370 ;
        RECT 363.010 3913.090 363.290 3913.370 ;
        RECT 363.720 3913.090 364.000 3913.370 ;
        RECT 364.430 3913.090 364.710 3913.370 ;
        RECT 365.140 3913.090 365.420 3913.370 ;
        RECT 365.850 3913.090 366.130 3913.370 ;
        RECT 366.560 3913.090 366.840 3913.370 ;
        RECT 3500.255 3913.135 3500.535 3913.415 ;
        RECT 3500.965 3913.135 3501.245 3913.415 ;
        RECT 3501.675 3913.135 3501.955 3913.415 ;
        RECT 3502.385 3913.135 3502.665 3913.415 ;
        RECT 3503.095 3913.135 3503.375 3913.415 ;
        RECT 3503.805 3913.135 3504.085 3913.415 ;
        RECT 3504.515 3913.135 3504.795 3913.415 ;
        RECT 3505.225 3913.135 3505.505 3913.415 ;
        RECT 3505.935 3913.135 3506.215 3913.415 ;
        RECT 3506.645 3913.135 3506.925 3913.415 ;
        RECT 3507.355 3913.135 3507.635 3913.415 ;
        RECT 3508.065 3913.135 3508.345 3913.415 ;
        RECT 3508.775 3913.135 3509.055 3913.415 ;
        RECT 3509.485 3913.135 3509.765 3913.415 ;
        RECT 357.330 3912.380 357.610 3912.660 ;
        RECT 358.040 3912.380 358.320 3912.660 ;
        RECT 358.750 3912.380 359.030 3912.660 ;
        RECT 359.460 3912.380 359.740 3912.660 ;
        RECT 360.170 3912.380 360.450 3912.660 ;
        RECT 360.880 3912.380 361.160 3912.660 ;
        RECT 361.590 3912.380 361.870 3912.660 ;
        RECT 362.300 3912.380 362.580 3912.660 ;
        RECT 363.010 3912.380 363.290 3912.660 ;
        RECT 363.720 3912.380 364.000 3912.660 ;
        RECT 364.430 3912.380 364.710 3912.660 ;
        RECT 365.140 3912.380 365.420 3912.660 ;
        RECT 365.850 3912.380 366.130 3912.660 ;
        RECT 366.560 3912.380 366.840 3912.660 ;
        RECT 3500.255 3912.425 3500.535 3912.705 ;
        RECT 3500.965 3912.425 3501.245 3912.705 ;
        RECT 3501.675 3912.425 3501.955 3912.705 ;
        RECT 3502.385 3912.425 3502.665 3912.705 ;
        RECT 3503.095 3912.425 3503.375 3912.705 ;
        RECT 3503.805 3912.425 3504.085 3912.705 ;
        RECT 3504.515 3912.425 3504.795 3912.705 ;
        RECT 3505.225 3912.425 3505.505 3912.705 ;
        RECT 3505.935 3912.425 3506.215 3912.705 ;
        RECT 3506.645 3912.425 3506.925 3912.705 ;
        RECT 3507.355 3912.425 3507.635 3912.705 ;
        RECT 3508.065 3912.425 3508.345 3912.705 ;
        RECT 3508.775 3912.425 3509.055 3912.705 ;
        RECT 3509.485 3912.425 3509.765 3912.705 ;
        RECT 357.330 3911.670 357.610 3911.950 ;
        RECT 358.040 3911.670 358.320 3911.950 ;
        RECT 358.750 3911.670 359.030 3911.950 ;
        RECT 359.460 3911.670 359.740 3911.950 ;
        RECT 360.170 3911.670 360.450 3911.950 ;
        RECT 360.880 3911.670 361.160 3911.950 ;
        RECT 361.590 3911.670 361.870 3911.950 ;
        RECT 362.300 3911.670 362.580 3911.950 ;
        RECT 363.010 3911.670 363.290 3911.950 ;
        RECT 363.720 3911.670 364.000 3911.950 ;
        RECT 364.430 3911.670 364.710 3911.950 ;
        RECT 365.140 3911.670 365.420 3911.950 ;
        RECT 365.850 3911.670 366.130 3911.950 ;
        RECT 366.560 3911.670 366.840 3911.950 ;
        RECT 3500.255 3911.715 3500.535 3911.995 ;
        RECT 3500.965 3911.715 3501.245 3911.995 ;
        RECT 3501.675 3911.715 3501.955 3911.995 ;
        RECT 3502.385 3911.715 3502.665 3911.995 ;
        RECT 3503.095 3911.715 3503.375 3911.995 ;
        RECT 3503.805 3911.715 3504.085 3911.995 ;
        RECT 3504.515 3911.715 3504.795 3911.995 ;
        RECT 3505.225 3911.715 3505.505 3911.995 ;
        RECT 3505.935 3911.715 3506.215 3911.995 ;
        RECT 3506.645 3911.715 3506.925 3911.995 ;
        RECT 3507.355 3911.715 3507.635 3911.995 ;
        RECT 3508.065 3911.715 3508.345 3911.995 ;
        RECT 3508.775 3911.715 3509.055 3911.995 ;
        RECT 3509.485 3911.715 3509.765 3911.995 ;
        RECT 3500.255 3911.005 3500.535 3911.285 ;
        RECT 3500.965 3911.005 3501.245 3911.285 ;
        RECT 3501.675 3911.005 3501.955 3911.285 ;
        RECT 3502.385 3911.005 3502.665 3911.285 ;
        RECT 3503.095 3911.005 3503.375 3911.285 ;
        RECT 3503.805 3911.005 3504.085 3911.285 ;
        RECT 3504.515 3911.005 3504.795 3911.285 ;
        RECT 3505.225 3911.005 3505.505 3911.285 ;
        RECT 3505.935 3911.005 3506.215 3911.285 ;
        RECT 3506.645 3911.005 3506.925 3911.285 ;
        RECT 3507.355 3911.005 3507.635 3911.285 ;
        RECT 3508.065 3911.005 3508.345 3911.285 ;
        RECT 3508.775 3911.005 3509.055 3911.285 ;
        RECT 3509.485 3911.005 3509.765 3911.285 ;
        RECT 3500.255 3908.385 3500.535 3908.665 ;
        RECT 3500.965 3908.385 3501.245 3908.665 ;
        RECT 3501.675 3908.385 3501.955 3908.665 ;
        RECT 3502.385 3908.385 3502.665 3908.665 ;
        RECT 3503.095 3908.385 3503.375 3908.665 ;
        RECT 3503.805 3908.385 3504.085 3908.665 ;
        RECT 3504.515 3908.385 3504.795 3908.665 ;
        RECT 3505.225 3908.385 3505.505 3908.665 ;
        RECT 3505.935 3908.385 3506.215 3908.665 ;
        RECT 3506.645 3908.385 3506.925 3908.665 ;
        RECT 3507.355 3908.385 3507.635 3908.665 ;
        RECT 3508.065 3908.385 3508.345 3908.665 ;
        RECT 3508.775 3908.385 3509.055 3908.665 ;
        RECT 3509.485 3908.385 3509.765 3908.665 ;
        RECT 3500.255 3907.675 3500.535 3907.955 ;
        RECT 3500.965 3907.675 3501.245 3907.955 ;
        RECT 3501.675 3907.675 3501.955 3907.955 ;
        RECT 3502.385 3907.675 3502.665 3907.955 ;
        RECT 3503.095 3907.675 3503.375 3907.955 ;
        RECT 3503.805 3907.675 3504.085 3907.955 ;
        RECT 3504.515 3907.675 3504.795 3907.955 ;
        RECT 3505.225 3907.675 3505.505 3907.955 ;
        RECT 3505.935 3907.675 3506.215 3907.955 ;
        RECT 3506.645 3907.675 3506.925 3907.955 ;
        RECT 3507.355 3907.675 3507.635 3907.955 ;
        RECT 3508.065 3907.675 3508.345 3907.955 ;
        RECT 3508.775 3907.675 3509.055 3907.955 ;
        RECT 3509.485 3907.675 3509.765 3907.955 ;
        RECT 3500.255 3906.965 3500.535 3907.245 ;
        RECT 3500.965 3906.965 3501.245 3907.245 ;
        RECT 3501.675 3906.965 3501.955 3907.245 ;
        RECT 3502.385 3906.965 3502.665 3907.245 ;
        RECT 3503.095 3906.965 3503.375 3907.245 ;
        RECT 3503.805 3906.965 3504.085 3907.245 ;
        RECT 3504.515 3906.965 3504.795 3907.245 ;
        RECT 3505.225 3906.965 3505.505 3907.245 ;
        RECT 3505.935 3906.965 3506.215 3907.245 ;
        RECT 3506.645 3906.965 3506.925 3907.245 ;
        RECT 3507.355 3906.965 3507.635 3907.245 ;
        RECT 3508.065 3906.965 3508.345 3907.245 ;
        RECT 3508.775 3906.965 3509.055 3907.245 ;
        RECT 3509.485 3906.965 3509.765 3907.245 ;
        RECT 3500.255 3906.255 3500.535 3906.535 ;
        RECT 3500.965 3906.255 3501.245 3906.535 ;
        RECT 3501.675 3906.255 3501.955 3906.535 ;
        RECT 3502.385 3906.255 3502.665 3906.535 ;
        RECT 3503.095 3906.255 3503.375 3906.535 ;
        RECT 3503.805 3906.255 3504.085 3906.535 ;
        RECT 3504.515 3906.255 3504.795 3906.535 ;
        RECT 3505.225 3906.255 3505.505 3906.535 ;
        RECT 3505.935 3906.255 3506.215 3906.535 ;
        RECT 3506.645 3906.255 3506.925 3906.535 ;
        RECT 3507.355 3906.255 3507.635 3906.535 ;
        RECT 3508.065 3906.255 3508.345 3906.535 ;
        RECT 3508.775 3906.255 3509.055 3906.535 ;
        RECT 3509.485 3906.255 3509.765 3906.535 ;
        RECT 3500.255 3905.545 3500.535 3905.825 ;
        RECT 3500.965 3905.545 3501.245 3905.825 ;
        RECT 3501.675 3905.545 3501.955 3905.825 ;
        RECT 3502.385 3905.545 3502.665 3905.825 ;
        RECT 3503.095 3905.545 3503.375 3905.825 ;
        RECT 3503.805 3905.545 3504.085 3905.825 ;
        RECT 3504.515 3905.545 3504.795 3905.825 ;
        RECT 3505.225 3905.545 3505.505 3905.825 ;
        RECT 3505.935 3905.545 3506.215 3905.825 ;
        RECT 3506.645 3905.545 3506.925 3905.825 ;
        RECT 3507.355 3905.545 3507.635 3905.825 ;
        RECT 3508.065 3905.545 3508.345 3905.825 ;
        RECT 3508.775 3905.545 3509.055 3905.825 ;
        RECT 3509.485 3905.545 3509.765 3905.825 ;
        RECT 3500.255 3904.835 3500.535 3905.115 ;
        RECT 3500.965 3904.835 3501.245 3905.115 ;
        RECT 3501.675 3904.835 3501.955 3905.115 ;
        RECT 3502.385 3904.835 3502.665 3905.115 ;
        RECT 3503.095 3904.835 3503.375 3905.115 ;
        RECT 3503.805 3904.835 3504.085 3905.115 ;
        RECT 3504.515 3904.835 3504.795 3905.115 ;
        RECT 3505.225 3904.835 3505.505 3905.115 ;
        RECT 3505.935 3904.835 3506.215 3905.115 ;
        RECT 3506.645 3904.835 3506.925 3905.115 ;
        RECT 3507.355 3904.835 3507.635 3905.115 ;
        RECT 3508.065 3904.835 3508.345 3905.115 ;
        RECT 3508.775 3904.835 3509.055 3905.115 ;
        RECT 3509.485 3904.835 3509.765 3905.115 ;
        RECT 3500.255 3904.125 3500.535 3904.405 ;
        RECT 3500.965 3904.125 3501.245 3904.405 ;
        RECT 3501.675 3904.125 3501.955 3904.405 ;
        RECT 3502.385 3904.125 3502.665 3904.405 ;
        RECT 3503.095 3904.125 3503.375 3904.405 ;
        RECT 3503.805 3904.125 3504.085 3904.405 ;
        RECT 3504.515 3904.125 3504.795 3904.405 ;
        RECT 3505.225 3904.125 3505.505 3904.405 ;
        RECT 3505.935 3904.125 3506.215 3904.405 ;
        RECT 3506.645 3904.125 3506.925 3904.405 ;
        RECT 3507.355 3904.125 3507.635 3904.405 ;
        RECT 3508.065 3904.125 3508.345 3904.405 ;
        RECT 3508.775 3904.125 3509.055 3904.405 ;
        RECT 3509.485 3904.125 3509.765 3904.405 ;
        RECT 3500.255 3903.415 3500.535 3903.695 ;
        RECT 3500.965 3903.415 3501.245 3903.695 ;
        RECT 3501.675 3903.415 3501.955 3903.695 ;
        RECT 3502.385 3903.415 3502.665 3903.695 ;
        RECT 3503.095 3903.415 3503.375 3903.695 ;
        RECT 3503.805 3903.415 3504.085 3903.695 ;
        RECT 3504.515 3903.415 3504.795 3903.695 ;
        RECT 3505.225 3903.415 3505.505 3903.695 ;
        RECT 3505.935 3903.415 3506.215 3903.695 ;
        RECT 3506.645 3903.415 3506.925 3903.695 ;
        RECT 3507.355 3903.415 3507.635 3903.695 ;
        RECT 3508.065 3903.415 3508.345 3903.695 ;
        RECT 3508.775 3903.415 3509.055 3903.695 ;
        RECT 3509.485 3903.415 3509.765 3903.695 ;
        RECT 3500.255 3902.705 3500.535 3902.985 ;
        RECT 3500.965 3902.705 3501.245 3902.985 ;
        RECT 3501.675 3902.705 3501.955 3902.985 ;
        RECT 3502.385 3902.705 3502.665 3902.985 ;
        RECT 3503.095 3902.705 3503.375 3902.985 ;
        RECT 3503.805 3902.705 3504.085 3902.985 ;
        RECT 3504.515 3902.705 3504.795 3902.985 ;
        RECT 3505.225 3902.705 3505.505 3902.985 ;
        RECT 3505.935 3902.705 3506.215 3902.985 ;
        RECT 3506.645 3902.705 3506.925 3902.985 ;
        RECT 3507.355 3902.705 3507.635 3902.985 ;
        RECT 3508.065 3902.705 3508.345 3902.985 ;
        RECT 3508.775 3902.705 3509.055 3902.985 ;
        RECT 3509.485 3902.705 3509.765 3902.985 ;
        RECT 3500.255 3901.995 3500.535 3902.275 ;
        RECT 3500.965 3901.995 3501.245 3902.275 ;
        RECT 3501.675 3901.995 3501.955 3902.275 ;
        RECT 3502.385 3901.995 3502.665 3902.275 ;
        RECT 3503.095 3901.995 3503.375 3902.275 ;
        RECT 3503.805 3901.995 3504.085 3902.275 ;
        RECT 3504.515 3901.995 3504.795 3902.275 ;
        RECT 3505.225 3901.995 3505.505 3902.275 ;
        RECT 3505.935 3901.995 3506.215 3902.275 ;
        RECT 3506.645 3901.995 3506.925 3902.275 ;
        RECT 3507.355 3901.995 3507.635 3902.275 ;
        RECT 3508.065 3901.995 3508.345 3902.275 ;
        RECT 3508.775 3901.995 3509.055 3902.275 ;
        RECT 3509.485 3901.995 3509.765 3902.275 ;
        RECT 3500.255 3901.285 3500.535 3901.565 ;
        RECT 3500.965 3901.285 3501.245 3901.565 ;
        RECT 3501.675 3901.285 3501.955 3901.565 ;
        RECT 3502.385 3901.285 3502.665 3901.565 ;
        RECT 3503.095 3901.285 3503.375 3901.565 ;
        RECT 3503.805 3901.285 3504.085 3901.565 ;
        RECT 3504.515 3901.285 3504.795 3901.565 ;
        RECT 3505.225 3901.285 3505.505 3901.565 ;
        RECT 3505.935 3901.285 3506.215 3901.565 ;
        RECT 3506.645 3901.285 3506.925 3901.565 ;
        RECT 3507.355 3901.285 3507.635 3901.565 ;
        RECT 3508.065 3901.285 3508.345 3901.565 ;
        RECT 3508.775 3901.285 3509.055 3901.565 ;
        RECT 3509.485 3901.285 3509.765 3901.565 ;
        RECT 3500.255 3900.575 3500.535 3900.855 ;
        RECT 3500.965 3900.575 3501.245 3900.855 ;
        RECT 3501.675 3900.575 3501.955 3900.855 ;
        RECT 3502.385 3900.575 3502.665 3900.855 ;
        RECT 3503.095 3900.575 3503.375 3900.855 ;
        RECT 3503.805 3900.575 3504.085 3900.855 ;
        RECT 3504.515 3900.575 3504.795 3900.855 ;
        RECT 3505.225 3900.575 3505.505 3900.855 ;
        RECT 3505.935 3900.575 3506.215 3900.855 ;
        RECT 3506.645 3900.575 3506.925 3900.855 ;
        RECT 3507.355 3900.575 3507.635 3900.855 ;
        RECT 3508.065 3900.575 3508.345 3900.855 ;
        RECT 3508.775 3900.575 3509.055 3900.855 ;
        RECT 3509.485 3900.575 3509.765 3900.855 ;
        RECT 3500.255 3899.865 3500.535 3900.145 ;
        RECT 3500.965 3899.865 3501.245 3900.145 ;
        RECT 3501.675 3899.865 3501.955 3900.145 ;
        RECT 3502.385 3899.865 3502.665 3900.145 ;
        RECT 3503.095 3899.865 3503.375 3900.145 ;
        RECT 3503.805 3899.865 3504.085 3900.145 ;
        RECT 3504.515 3899.865 3504.795 3900.145 ;
        RECT 3505.225 3899.865 3505.505 3900.145 ;
        RECT 3505.935 3899.865 3506.215 3900.145 ;
        RECT 3506.645 3899.865 3506.925 3900.145 ;
        RECT 3507.355 3899.865 3507.635 3900.145 ;
        RECT 3508.065 3899.865 3508.345 3900.145 ;
        RECT 3508.775 3899.865 3509.055 3900.145 ;
        RECT 3509.485 3899.865 3509.765 3900.145 ;
        RECT 3500.255 3899.155 3500.535 3899.435 ;
        RECT 3500.965 3899.155 3501.245 3899.435 ;
        RECT 3501.675 3899.155 3501.955 3899.435 ;
        RECT 3502.385 3899.155 3502.665 3899.435 ;
        RECT 3503.095 3899.155 3503.375 3899.435 ;
        RECT 3503.805 3899.155 3504.085 3899.435 ;
        RECT 3504.515 3899.155 3504.795 3899.435 ;
        RECT 3505.225 3899.155 3505.505 3899.435 ;
        RECT 3505.935 3899.155 3506.215 3899.435 ;
        RECT 3506.645 3899.155 3506.925 3899.435 ;
        RECT 3507.355 3899.155 3507.635 3899.435 ;
        RECT 3508.065 3899.155 3508.345 3899.435 ;
        RECT 3508.775 3899.155 3509.055 3899.435 ;
        RECT 3509.485 3899.155 3509.765 3899.435 ;
        RECT 3500.200 3895.270 3500.480 3895.550 ;
        RECT 3500.910 3895.270 3501.190 3895.550 ;
        RECT 3501.620 3895.270 3501.900 3895.550 ;
        RECT 3502.330 3895.270 3502.610 3895.550 ;
        RECT 3503.040 3895.270 3503.320 3895.550 ;
        RECT 3503.750 3895.270 3504.030 3895.550 ;
        RECT 3504.460 3895.270 3504.740 3895.550 ;
        RECT 3505.170 3895.270 3505.450 3895.550 ;
        RECT 3505.880 3895.270 3506.160 3895.550 ;
        RECT 3506.590 3895.270 3506.870 3895.550 ;
        RECT 3507.300 3895.270 3507.580 3895.550 ;
        RECT 3508.010 3895.270 3508.290 3895.550 ;
        RECT 3508.720 3895.270 3509.000 3895.550 ;
        RECT 3509.430 3895.270 3509.710 3895.550 ;
        RECT 3500.200 3894.560 3500.480 3894.840 ;
        RECT 3500.910 3894.560 3501.190 3894.840 ;
        RECT 3501.620 3894.560 3501.900 3894.840 ;
        RECT 3502.330 3894.560 3502.610 3894.840 ;
        RECT 3503.040 3894.560 3503.320 3894.840 ;
        RECT 3503.750 3894.560 3504.030 3894.840 ;
        RECT 3504.460 3894.560 3504.740 3894.840 ;
        RECT 3505.170 3894.560 3505.450 3894.840 ;
        RECT 3505.880 3894.560 3506.160 3894.840 ;
        RECT 3506.590 3894.560 3506.870 3894.840 ;
        RECT 3507.300 3894.560 3507.580 3894.840 ;
        RECT 3508.010 3894.560 3508.290 3894.840 ;
        RECT 3508.720 3894.560 3509.000 3894.840 ;
        RECT 3509.430 3894.560 3509.710 3894.840 ;
        RECT 3500.200 3893.850 3500.480 3894.130 ;
        RECT 3500.910 3893.850 3501.190 3894.130 ;
        RECT 3501.620 3893.850 3501.900 3894.130 ;
        RECT 3502.330 3893.850 3502.610 3894.130 ;
        RECT 3503.040 3893.850 3503.320 3894.130 ;
        RECT 3503.750 3893.850 3504.030 3894.130 ;
        RECT 3504.460 3893.850 3504.740 3894.130 ;
        RECT 3505.170 3893.850 3505.450 3894.130 ;
        RECT 3505.880 3893.850 3506.160 3894.130 ;
        RECT 3506.590 3893.850 3506.870 3894.130 ;
        RECT 3507.300 3893.850 3507.580 3894.130 ;
        RECT 3508.010 3893.850 3508.290 3894.130 ;
        RECT 3508.720 3893.850 3509.000 3894.130 ;
        RECT 3509.430 3893.850 3509.710 3894.130 ;
        RECT 3500.200 3893.140 3500.480 3893.420 ;
        RECT 3500.910 3893.140 3501.190 3893.420 ;
        RECT 3501.620 3893.140 3501.900 3893.420 ;
        RECT 3502.330 3893.140 3502.610 3893.420 ;
        RECT 3503.040 3893.140 3503.320 3893.420 ;
        RECT 3503.750 3893.140 3504.030 3893.420 ;
        RECT 3504.460 3893.140 3504.740 3893.420 ;
        RECT 3505.170 3893.140 3505.450 3893.420 ;
        RECT 3505.880 3893.140 3506.160 3893.420 ;
        RECT 3506.590 3893.140 3506.870 3893.420 ;
        RECT 3507.300 3893.140 3507.580 3893.420 ;
        RECT 3508.010 3893.140 3508.290 3893.420 ;
        RECT 3508.720 3893.140 3509.000 3893.420 ;
        RECT 3509.430 3893.140 3509.710 3893.420 ;
        RECT 3500.200 3892.430 3500.480 3892.710 ;
        RECT 3500.910 3892.430 3501.190 3892.710 ;
        RECT 3501.620 3892.430 3501.900 3892.710 ;
        RECT 3502.330 3892.430 3502.610 3892.710 ;
        RECT 3503.040 3892.430 3503.320 3892.710 ;
        RECT 3503.750 3892.430 3504.030 3892.710 ;
        RECT 3504.460 3892.430 3504.740 3892.710 ;
        RECT 3505.170 3892.430 3505.450 3892.710 ;
        RECT 3505.880 3892.430 3506.160 3892.710 ;
        RECT 3506.590 3892.430 3506.870 3892.710 ;
        RECT 3507.300 3892.430 3507.580 3892.710 ;
        RECT 3508.010 3892.430 3508.290 3892.710 ;
        RECT 3508.720 3892.430 3509.000 3892.710 ;
        RECT 3509.430 3892.430 3509.710 3892.710 ;
        RECT 3500.200 3891.720 3500.480 3892.000 ;
        RECT 3500.910 3891.720 3501.190 3892.000 ;
        RECT 3501.620 3891.720 3501.900 3892.000 ;
        RECT 3502.330 3891.720 3502.610 3892.000 ;
        RECT 3503.040 3891.720 3503.320 3892.000 ;
        RECT 3503.750 3891.720 3504.030 3892.000 ;
        RECT 3504.460 3891.720 3504.740 3892.000 ;
        RECT 3505.170 3891.720 3505.450 3892.000 ;
        RECT 3505.880 3891.720 3506.160 3892.000 ;
        RECT 3506.590 3891.720 3506.870 3892.000 ;
        RECT 3507.300 3891.720 3507.580 3892.000 ;
        RECT 3508.010 3891.720 3508.290 3892.000 ;
        RECT 3508.720 3891.720 3509.000 3892.000 ;
        RECT 3509.430 3891.720 3509.710 3892.000 ;
        RECT 3500.200 3891.010 3500.480 3891.290 ;
        RECT 3500.910 3891.010 3501.190 3891.290 ;
        RECT 3501.620 3891.010 3501.900 3891.290 ;
        RECT 3502.330 3891.010 3502.610 3891.290 ;
        RECT 3503.040 3891.010 3503.320 3891.290 ;
        RECT 3503.750 3891.010 3504.030 3891.290 ;
        RECT 3504.460 3891.010 3504.740 3891.290 ;
        RECT 3505.170 3891.010 3505.450 3891.290 ;
        RECT 3505.880 3891.010 3506.160 3891.290 ;
        RECT 3506.590 3891.010 3506.870 3891.290 ;
        RECT 3507.300 3891.010 3507.580 3891.290 ;
        RECT 3508.010 3891.010 3508.290 3891.290 ;
        RECT 3508.720 3891.010 3509.000 3891.290 ;
        RECT 3509.430 3891.010 3509.710 3891.290 ;
        RECT 3500.200 3890.300 3500.480 3890.580 ;
        RECT 3500.910 3890.300 3501.190 3890.580 ;
        RECT 3501.620 3890.300 3501.900 3890.580 ;
        RECT 3502.330 3890.300 3502.610 3890.580 ;
        RECT 3503.040 3890.300 3503.320 3890.580 ;
        RECT 3503.750 3890.300 3504.030 3890.580 ;
        RECT 3504.460 3890.300 3504.740 3890.580 ;
        RECT 3505.170 3890.300 3505.450 3890.580 ;
        RECT 3505.880 3890.300 3506.160 3890.580 ;
        RECT 3506.590 3890.300 3506.870 3890.580 ;
        RECT 3507.300 3890.300 3507.580 3890.580 ;
        RECT 3508.010 3890.300 3508.290 3890.580 ;
        RECT 3508.720 3890.300 3509.000 3890.580 ;
        RECT 3509.430 3890.300 3509.710 3890.580 ;
        RECT 3500.200 3889.590 3500.480 3889.870 ;
        RECT 3500.910 3889.590 3501.190 3889.870 ;
        RECT 3501.620 3889.590 3501.900 3889.870 ;
        RECT 3502.330 3889.590 3502.610 3889.870 ;
        RECT 3503.040 3889.590 3503.320 3889.870 ;
        RECT 3503.750 3889.590 3504.030 3889.870 ;
        RECT 3504.460 3889.590 3504.740 3889.870 ;
        RECT 3505.170 3889.590 3505.450 3889.870 ;
        RECT 3505.880 3889.590 3506.160 3889.870 ;
        RECT 3506.590 3889.590 3506.870 3889.870 ;
        RECT 3507.300 3889.590 3507.580 3889.870 ;
        RECT 3508.010 3889.590 3508.290 3889.870 ;
        RECT 3508.720 3889.590 3509.000 3889.870 ;
        RECT 3509.430 3889.590 3509.710 3889.870 ;
        RECT 3500.200 3888.880 3500.480 3889.160 ;
        RECT 3500.910 3888.880 3501.190 3889.160 ;
        RECT 3501.620 3888.880 3501.900 3889.160 ;
        RECT 3502.330 3888.880 3502.610 3889.160 ;
        RECT 3503.040 3888.880 3503.320 3889.160 ;
        RECT 3503.750 3888.880 3504.030 3889.160 ;
        RECT 3504.460 3888.880 3504.740 3889.160 ;
        RECT 3505.170 3888.880 3505.450 3889.160 ;
        RECT 3505.880 3888.880 3506.160 3889.160 ;
        RECT 3506.590 3888.880 3506.870 3889.160 ;
        RECT 3507.300 3888.880 3507.580 3889.160 ;
        RECT 3508.010 3888.880 3508.290 3889.160 ;
        RECT 3508.720 3888.880 3509.000 3889.160 ;
        RECT 3509.430 3888.880 3509.710 3889.160 ;
        RECT 3500.200 3888.170 3500.480 3888.450 ;
        RECT 3500.910 3888.170 3501.190 3888.450 ;
        RECT 3501.620 3888.170 3501.900 3888.450 ;
        RECT 3502.330 3888.170 3502.610 3888.450 ;
        RECT 3503.040 3888.170 3503.320 3888.450 ;
        RECT 3503.750 3888.170 3504.030 3888.450 ;
        RECT 3504.460 3888.170 3504.740 3888.450 ;
        RECT 3505.170 3888.170 3505.450 3888.450 ;
        RECT 3505.880 3888.170 3506.160 3888.450 ;
        RECT 3506.590 3888.170 3506.870 3888.450 ;
        RECT 3507.300 3888.170 3507.580 3888.450 ;
        RECT 3508.010 3888.170 3508.290 3888.450 ;
        RECT 3508.720 3888.170 3509.000 3888.450 ;
        RECT 3509.430 3888.170 3509.710 3888.450 ;
        RECT 3500.200 3887.460 3500.480 3887.740 ;
        RECT 3500.910 3887.460 3501.190 3887.740 ;
        RECT 3501.620 3887.460 3501.900 3887.740 ;
        RECT 3502.330 3887.460 3502.610 3887.740 ;
        RECT 3503.040 3887.460 3503.320 3887.740 ;
        RECT 3503.750 3887.460 3504.030 3887.740 ;
        RECT 3504.460 3887.460 3504.740 3887.740 ;
        RECT 3505.170 3887.460 3505.450 3887.740 ;
        RECT 3505.880 3887.460 3506.160 3887.740 ;
        RECT 3506.590 3887.460 3506.870 3887.740 ;
        RECT 3507.300 3887.460 3507.580 3887.740 ;
        RECT 3508.010 3887.460 3508.290 3887.740 ;
        RECT 3508.720 3887.460 3509.000 3887.740 ;
        RECT 3509.430 3887.460 3509.710 3887.740 ;
        RECT 3500.200 3886.750 3500.480 3887.030 ;
        RECT 3500.910 3886.750 3501.190 3887.030 ;
        RECT 3501.620 3886.750 3501.900 3887.030 ;
        RECT 3502.330 3886.750 3502.610 3887.030 ;
        RECT 3503.040 3886.750 3503.320 3887.030 ;
        RECT 3503.750 3886.750 3504.030 3887.030 ;
        RECT 3504.460 3886.750 3504.740 3887.030 ;
        RECT 3505.170 3886.750 3505.450 3887.030 ;
        RECT 3505.880 3886.750 3506.160 3887.030 ;
        RECT 3506.590 3886.750 3506.870 3887.030 ;
        RECT 3507.300 3886.750 3507.580 3887.030 ;
        RECT 3508.010 3886.750 3508.290 3887.030 ;
        RECT 3508.720 3886.750 3509.000 3887.030 ;
        RECT 3509.430 3886.750 3509.710 3887.030 ;
        RECT 3500.200 2453.050 3500.480 2453.330 ;
        RECT 3500.910 2453.050 3501.190 2453.330 ;
        RECT 3501.620 2453.050 3501.900 2453.330 ;
        RECT 3502.330 2453.050 3502.610 2453.330 ;
        RECT 3503.040 2453.050 3503.320 2453.330 ;
        RECT 3503.750 2453.050 3504.030 2453.330 ;
        RECT 3504.460 2453.050 3504.740 2453.330 ;
        RECT 3505.170 2453.050 3505.450 2453.330 ;
        RECT 3505.880 2453.050 3506.160 2453.330 ;
        RECT 3506.590 2453.050 3506.870 2453.330 ;
        RECT 3507.300 2453.050 3507.580 2453.330 ;
        RECT 3508.010 2453.050 3508.290 2453.330 ;
        RECT 3508.720 2453.050 3509.000 2453.330 ;
        RECT 3509.430 2453.050 3509.710 2453.330 ;
        RECT 3500.200 2452.340 3500.480 2452.620 ;
        RECT 3500.910 2452.340 3501.190 2452.620 ;
        RECT 3501.620 2452.340 3501.900 2452.620 ;
        RECT 3502.330 2452.340 3502.610 2452.620 ;
        RECT 3503.040 2452.340 3503.320 2452.620 ;
        RECT 3503.750 2452.340 3504.030 2452.620 ;
        RECT 3504.460 2452.340 3504.740 2452.620 ;
        RECT 3505.170 2452.340 3505.450 2452.620 ;
        RECT 3505.880 2452.340 3506.160 2452.620 ;
        RECT 3506.590 2452.340 3506.870 2452.620 ;
        RECT 3507.300 2452.340 3507.580 2452.620 ;
        RECT 3508.010 2452.340 3508.290 2452.620 ;
        RECT 3508.720 2452.340 3509.000 2452.620 ;
        RECT 3509.430 2452.340 3509.710 2452.620 ;
        RECT 3500.200 2451.630 3500.480 2451.910 ;
        RECT 3500.910 2451.630 3501.190 2451.910 ;
        RECT 3501.620 2451.630 3501.900 2451.910 ;
        RECT 3502.330 2451.630 3502.610 2451.910 ;
        RECT 3503.040 2451.630 3503.320 2451.910 ;
        RECT 3503.750 2451.630 3504.030 2451.910 ;
        RECT 3504.460 2451.630 3504.740 2451.910 ;
        RECT 3505.170 2451.630 3505.450 2451.910 ;
        RECT 3505.880 2451.630 3506.160 2451.910 ;
        RECT 3506.590 2451.630 3506.870 2451.910 ;
        RECT 3507.300 2451.630 3507.580 2451.910 ;
        RECT 3508.010 2451.630 3508.290 2451.910 ;
        RECT 3508.720 2451.630 3509.000 2451.910 ;
        RECT 3509.430 2451.630 3509.710 2451.910 ;
        RECT 3500.200 2450.920 3500.480 2451.200 ;
        RECT 3500.910 2450.920 3501.190 2451.200 ;
        RECT 3501.620 2450.920 3501.900 2451.200 ;
        RECT 3502.330 2450.920 3502.610 2451.200 ;
        RECT 3503.040 2450.920 3503.320 2451.200 ;
        RECT 3503.750 2450.920 3504.030 2451.200 ;
        RECT 3504.460 2450.920 3504.740 2451.200 ;
        RECT 3505.170 2450.920 3505.450 2451.200 ;
        RECT 3505.880 2450.920 3506.160 2451.200 ;
        RECT 3506.590 2450.920 3506.870 2451.200 ;
        RECT 3507.300 2450.920 3507.580 2451.200 ;
        RECT 3508.010 2450.920 3508.290 2451.200 ;
        RECT 3508.720 2450.920 3509.000 2451.200 ;
        RECT 3509.430 2450.920 3509.710 2451.200 ;
        RECT 3500.200 2450.210 3500.480 2450.490 ;
        RECT 3500.910 2450.210 3501.190 2450.490 ;
        RECT 3501.620 2450.210 3501.900 2450.490 ;
        RECT 3502.330 2450.210 3502.610 2450.490 ;
        RECT 3503.040 2450.210 3503.320 2450.490 ;
        RECT 3503.750 2450.210 3504.030 2450.490 ;
        RECT 3504.460 2450.210 3504.740 2450.490 ;
        RECT 3505.170 2450.210 3505.450 2450.490 ;
        RECT 3505.880 2450.210 3506.160 2450.490 ;
        RECT 3506.590 2450.210 3506.870 2450.490 ;
        RECT 3507.300 2450.210 3507.580 2450.490 ;
        RECT 3508.010 2450.210 3508.290 2450.490 ;
        RECT 3508.720 2450.210 3509.000 2450.490 ;
        RECT 3509.430 2450.210 3509.710 2450.490 ;
        RECT 3500.200 2449.500 3500.480 2449.780 ;
        RECT 3500.910 2449.500 3501.190 2449.780 ;
        RECT 3501.620 2449.500 3501.900 2449.780 ;
        RECT 3502.330 2449.500 3502.610 2449.780 ;
        RECT 3503.040 2449.500 3503.320 2449.780 ;
        RECT 3503.750 2449.500 3504.030 2449.780 ;
        RECT 3504.460 2449.500 3504.740 2449.780 ;
        RECT 3505.170 2449.500 3505.450 2449.780 ;
        RECT 3505.880 2449.500 3506.160 2449.780 ;
        RECT 3506.590 2449.500 3506.870 2449.780 ;
        RECT 3507.300 2449.500 3507.580 2449.780 ;
        RECT 3508.010 2449.500 3508.290 2449.780 ;
        RECT 3508.720 2449.500 3509.000 2449.780 ;
        RECT 3509.430 2449.500 3509.710 2449.780 ;
        RECT 3500.200 2448.790 3500.480 2449.070 ;
        RECT 3500.910 2448.790 3501.190 2449.070 ;
        RECT 3501.620 2448.790 3501.900 2449.070 ;
        RECT 3502.330 2448.790 3502.610 2449.070 ;
        RECT 3503.040 2448.790 3503.320 2449.070 ;
        RECT 3503.750 2448.790 3504.030 2449.070 ;
        RECT 3504.460 2448.790 3504.740 2449.070 ;
        RECT 3505.170 2448.790 3505.450 2449.070 ;
        RECT 3505.880 2448.790 3506.160 2449.070 ;
        RECT 3506.590 2448.790 3506.870 2449.070 ;
        RECT 3507.300 2448.790 3507.580 2449.070 ;
        RECT 3508.010 2448.790 3508.290 2449.070 ;
        RECT 3508.720 2448.790 3509.000 2449.070 ;
        RECT 3509.430 2448.790 3509.710 2449.070 ;
        RECT 3500.200 2448.080 3500.480 2448.360 ;
        RECT 3500.910 2448.080 3501.190 2448.360 ;
        RECT 3501.620 2448.080 3501.900 2448.360 ;
        RECT 3502.330 2448.080 3502.610 2448.360 ;
        RECT 3503.040 2448.080 3503.320 2448.360 ;
        RECT 3503.750 2448.080 3504.030 2448.360 ;
        RECT 3504.460 2448.080 3504.740 2448.360 ;
        RECT 3505.170 2448.080 3505.450 2448.360 ;
        RECT 3505.880 2448.080 3506.160 2448.360 ;
        RECT 3506.590 2448.080 3506.870 2448.360 ;
        RECT 3507.300 2448.080 3507.580 2448.360 ;
        RECT 3508.010 2448.080 3508.290 2448.360 ;
        RECT 3508.720 2448.080 3509.000 2448.360 ;
        RECT 3509.430 2448.080 3509.710 2448.360 ;
        RECT 3500.200 2447.370 3500.480 2447.650 ;
        RECT 3500.910 2447.370 3501.190 2447.650 ;
        RECT 3501.620 2447.370 3501.900 2447.650 ;
        RECT 3502.330 2447.370 3502.610 2447.650 ;
        RECT 3503.040 2447.370 3503.320 2447.650 ;
        RECT 3503.750 2447.370 3504.030 2447.650 ;
        RECT 3504.460 2447.370 3504.740 2447.650 ;
        RECT 3505.170 2447.370 3505.450 2447.650 ;
        RECT 3505.880 2447.370 3506.160 2447.650 ;
        RECT 3506.590 2447.370 3506.870 2447.650 ;
        RECT 3507.300 2447.370 3507.580 2447.650 ;
        RECT 3508.010 2447.370 3508.290 2447.650 ;
        RECT 3508.720 2447.370 3509.000 2447.650 ;
        RECT 3509.430 2447.370 3509.710 2447.650 ;
        RECT 3500.200 2446.660 3500.480 2446.940 ;
        RECT 3500.910 2446.660 3501.190 2446.940 ;
        RECT 3501.620 2446.660 3501.900 2446.940 ;
        RECT 3502.330 2446.660 3502.610 2446.940 ;
        RECT 3503.040 2446.660 3503.320 2446.940 ;
        RECT 3503.750 2446.660 3504.030 2446.940 ;
        RECT 3504.460 2446.660 3504.740 2446.940 ;
        RECT 3505.170 2446.660 3505.450 2446.940 ;
        RECT 3505.880 2446.660 3506.160 2446.940 ;
        RECT 3506.590 2446.660 3506.870 2446.940 ;
        RECT 3507.300 2446.660 3507.580 2446.940 ;
        RECT 3508.010 2446.660 3508.290 2446.940 ;
        RECT 3508.720 2446.660 3509.000 2446.940 ;
        RECT 3509.430 2446.660 3509.710 2446.940 ;
        RECT 3500.200 2445.950 3500.480 2446.230 ;
        RECT 3500.910 2445.950 3501.190 2446.230 ;
        RECT 3501.620 2445.950 3501.900 2446.230 ;
        RECT 3502.330 2445.950 3502.610 2446.230 ;
        RECT 3503.040 2445.950 3503.320 2446.230 ;
        RECT 3503.750 2445.950 3504.030 2446.230 ;
        RECT 3504.460 2445.950 3504.740 2446.230 ;
        RECT 3505.170 2445.950 3505.450 2446.230 ;
        RECT 3505.880 2445.950 3506.160 2446.230 ;
        RECT 3506.590 2445.950 3506.870 2446.230 ;
        RECT 3507.300 2445.950 3507.580 2446.230 ;
        RECT 3508.010 2445.950 3508.290 2446.230 ;
        RECT 3508.720 2445.950 3509.000 2446.230 ;
        RECT 3509.430 2445.950 3509.710 2446.230 ;
        RECT 3500.200 2445.240 3500.480 2445.520 ;
        RECT 3500.910 2445.240 3501.190 2445.520 ;
        RECT 3501.620 2445.240 3501.900 2445.520 ;
        RECT 3502.330 2445.240 3502.610 2445.520 ;
        RECT 3503.040 2445.240 3503.320 2445.520 ;
        RECT 3503.750 2445.240 3504.030 2445.520 ;
        RECT 3504.460 2445.240 3504.740 2445.520 ;
        RECT 3505.170 2445.240 3505.450 2445.520 ;
        RECT 3505.880 2445.240 3506.160 2445.520 ;
        RECT 3506.590 2445.240 3506.870 2445.520 ;
        RECT 3507.300 2445.240 3507.580 2445.520 ;
        RECT 3508.010 2445.240 3508.290 2445.520 ;
        RECT 3508.720 2445.240 3509.000 2445.520 ;
        RECT 3509.430 2445.240 3509.710 2445.520 ;
        RECT 3500.200 2444.530 3500.480 2444.810 ;
        RECT 3500.910 2444.530 3501.190 2444.810 ;
        RECT 3501.620 2444.530 3501.900 2444.810 ;
        RECT 3502.330 2444.530 3502.610 2444.810 ;
        RECT 3503.040 2444.530 3503.320 2444.810 ;
        RECT 3503.750 2444.530 3504.030 2444.810 ;
        RECT 3504.460 2444.530 3504.740 2444.810 ;
        RECT 3505.170 2444.530 3505.450 2444.810 ;
        RECT 3505.880 2444.530 3506.160 2444.810 ;
        RECT 3506.590 2444.530 3506.870 2444.810 ;
        RECT 3507.300 2444.530 3507.580 2444.810 ;
        RECT 3508.010 2444.530 3508.290 2444.810 ;
        RECT 3508.720 2444.530 3509.000 2444.810 ;
        RECT 3509.430 2444.530 3509.710 2444.810 ;
        RECT 3500.255 2440.615 3500.535 2440.895 ;
        RECT 3500.965 2440.615 3501.245 2440.895 ;
        RECT 3501.675 2440.615 3501.955 2440.895 ;
        RECT 3502.385 2440.615 3502.665 2440.895 ;
        RECT 3503.095 2440.615 3503.375 2440.895 ;
        RECT 3503.805 2440.615 3504.085 2440.895 ;
        RECT 3504.515 2440.615 3504.795 2440.895 ;
        RECT 3505.225 2440.615 3505.505 2440.895 ;
        RECT 3505.935 2440.615 3506.215 2440.895 ;
        RECT 3506.645 2440.615 3506.925 2440.895 ;
        RECT 3507.355 2440.615 3507.635 2440.895 ;
        RECT 3508.065 2440.615 3508.345 2440.895 ;
        RECT 3508.775 2440.615 3509.055 2440.895 ;
        RECT 3509.485 2440.615 3509.765 2440.895 ;
        RECT 3500.255 2439.905 3500.535 2440.185 ;
        RECT 3500.965 2439.905 3501.245 2440.185 ;
        RECT 3501.675 2439.905 3501.955 2440.185 ;
        RECT 3502.385 2439.905 3502.665 2440.185 ;
        RECT 3503.095 2439.905 3503.375 2440.185 ;
        RECT 3503.805 2439.905 3504.085 2440.185 ;
        RECT 3504.515 2439.905 3504.795 2440.185 ;
        RECT 3505.225 2439.905 3505.505 2440.185 ;
        RECT 3505.935 2439.905 3506.215 2440.185 ;
        RECT 3506.645 2439.905 3506.925 2440.185 ;
        RECT 3507.355 2439.905 3507.635 2440.185 ;
        RECT 3508.065 2439.905 3508.345 2440.185 ;
        RECT 3508.775 2439.905 3509.055 2440.185 ;
        RECT 3509.485 2439.905 3509.765 2440.185 ;
        RECT 3500.255 2439.195 3500.535 2439.475 ;
        RECT 3500.965 2439.195 3501.245 2439.475 ;
        RECT 3501.675 2439.195 3501.955 2439.475 ;
        RECT 3502.385 2439.195 3502.665 2439.475 ;
        RECT 3503.095 2439.195 3503.375 2439.475 ;
        RECT 3503.805 2439.195 3504.085 2439.475 ;
        RECT 3504.515 2439.195 3504.795 2439.475 ;
        RECT 3505.225 2439.195 3505.505 2439.475 ;
        RECT 3505.935 2439.195 3506.215 2439.475 ;
        RECT 3506.645 2439.195 3506.925 2439.475 ;
        RECT 3507.355 2439.195 3507.635 2439.475 ;
        RECT 3508.065 2439.195 3508.345 2439.475 ;
        RECT 3508.775 2439.195 3509.055 2439.475 ;
        RECT 3509.485 2439.195 3509.765 2439.475 ;
        RECT 3500.255 2438.485 3500.535 2438.765 ;
        RECT 3500.965 2438.485 3501.245 2438.765 ;
        RECT 3501.675 2438.485 3501.955 2438.765 ;
        RECT 3502.385 2438.485 3502.665 2438.765 ;
        RECT 3503.095 2438.485 3503.375 2438.765 ;
        RECT 3503.805 2438.485 3504.085 2438.765 ;
        RECT 3504.515 2438.485 3504.795 2438.765 ;
        RECT 3505.225 2438.485 3505.505 2438.765 ;
        RECT 3505.935 2438.485 3506.215 2438.765 ;
        RECT 3506.645 2438.485 3506.925 2438.765 ;
        RECT 3507.355 2438.485 3507.635 2438.765 ;
        RECT 3508.065 2438.485 3508.345 2438.765 ;
        RECT 3508.775 2438.485 3509.055 2438.765 ;
        RECT 3509.485 2438.485 3509.765 2438.765 ;
        RECT 3500.255 2437.775 3500.535 2438.055 ;
        RECT 3500.965 2437.775 3501.245 2438.055 ;
        RECT 3501.675 2437.775 3501.955 2438.055 ;
        RECT 3502.385 2437.775 3502.665 2438.055 ;
        RECT 3503.095 2437.775 3503.375 2438.055 ;
        RECT 3503.805 2437.775 3504.085 2438.055 ;
        RECT 3504.515 2437.775 3504.795 2438.055 ;
        RECT 3505.225 2437.775 3505.505 2438.055 ;
        RECT 3505.935 2437.775 3506.215 2438.055 ;
        RECT 3506.645 2437.775 3506.925 2438.055 ;
        RECT 3507.355 2437.775 3507.635 2438.055 ;
        RECT 3508.065 2437.775 3508.345 2438.055 ;
        RECT 3508.775 2437.775 3509.055 2438.055 ;
        RECT 3509.485 2437.775 3509.765 2438.055 ;
        RECT 3500.255 2437.065 3500.535 2437.345 ;
        RECT 3500.965 2437.065 3501.245 2437.345 ;
        RECT 3501.675 2437.065 3501.955 2437.345 ;
        RECT 3502.385 2437.065 3502.665 2437.345 ;
        RECT 3503.095 2437.065 3503.375 2437.345 ;
        RECT 3503.805 2437.065 3504.085 2437.345 ;
        RECT 3504.515 2437.065 3504.795 2437.345 ;
        RECT 3505.225 2437.065 3505.505 2437.345 ;
        RECT 3505.935 2437.065 3506.215 2437.345 ;
        RECT 3506.645 2437.065 3506.925 2437.345 ;
        RECT 3507.355 2437.065 3507.635 2437.345 ;
        RECT 3508.065 2437.065 3508.345 2437.345 ;
        RECT 3508.775 2437.065 3509.055 2437.345 ;
        RECT 3509.485 2437.065 3509.765 2437.345 ;
        RECT 3500.255 2436.355 3500.535 2436.635 ;
        RECT 3500.965 2436.355 3501.245 2436.635 ;
        RECT 3501.675 2436.355 3501.955 2436.635 ;
        RECT 3502.385 2436.355 3502.665 2436.635 ;
        RECT 3503.095 2436.355 3503.375 2436.635 ;
        RECT 3503.805 2436.355 3504.085 2436.635 ;
        RECT 3504.515 2436.355 3504.795 2436.635 ;
        RECT 3505.225 2436.355 3505.505 2436.635 ;
        RECT 3505.935 2436.355 3506.215 2436.635 ;
        RECT 3506.645 2436.355 3506.925 2436.635 ;
        RECT 3507.355 2436.355 3507.635 2436.635 ;
        RECT 3508.065 2436.355 3508.345 2436.635 ;
        RECT 3508.775 2436.355 3509.055 2436.635 ;
        RECT 3509.485 2436.355 3509.765 2436.635 ;
        RECT 3500.255 2435.645 3500.535 2435.925 ;
        RECT 3500.965 2435.645 3501.245 2435.925 ;
        RECT 3501.675 2435.645 3501.955 2435.925 ;
        RECT 3502.385 2435.645 3502.665 2435.925 ;
        RECT 3503.095 2435.645 3503.375 2435.925 ;
        RECT 3503.805 2435.645 3504.085 2435.925 ;
        RECT 3504.515 2435.645 3504.795 2435.925 ;
        RECT 3505.225 2435.645 3505.505 2435.925 ;
        RECT 3505.935 2435.645 3506.215 2435.925 ;
        RECT 3506.645 2435.645 3506.925 2435.925 ;
        RECT 3507.355 2435.645 3507.635 2435.925 ;
        RECT 3508.065 2435.645 3508.345 2435.925 ;
        RECT 3508.775 2435.645 3509.055 2435.925 ;
        RECT 3509.485 2435.645 3509.765 2435.925 ;
        RECT 3500.255 2434.935 3500.535 2435.215 ;
        RECT 3500.965 2434.935 3501.245 2435.215 ;
        RECT 3501.675 2434.935 3501.955 2435.215 ;
        RECT 3502.385 2434.935 3502.665 2435.215 ;
        RECT 3503.095 2434.935 3503.375 2435.215 ;
        RECT 3503.805 2434.935 3504.085 2435.215 ;
        RECT 3504.515 2434.935 3504.795 2435.215 ;
        RECT 3505.225 2434.935 3505.505 2435.215 ;
        RECT 3505.935 2434.935 3506.215 2435.215 ;
        RECT 3506.645 2434.935 3506.925 2435.215 ;
        RECT 3507.355 2434.935 3507.635 2435.215 ;
        RECT 3508.065 2434.935 3508.345 2435.215 ;
        RECT 3508.775 2434.935 3509.055 2435.215 ;
        RECT 3509.485 2434.935 3509.765 2435.215 ;
        RECT 3500.255 2434.225 3500.535 2434.505 ;
        RECT 3500.965 2434.225 3501.245 2434.505 ;
        RECT 3501.675 2434.225 3501.955 2434.505 ;
        RECT 3502.385 2434.225 3502.665 2434.505 ;
        RECT 3503.095 2434.225 3503.375 2434.505 ;
        RECT 3503.805 2434.225 3504.085 2434.505 ;
        RECT 3504.515 2434.225 3504.795 2434.505 ;
        RECT 3505.225 2434.225 3505.505 2434.505 ;
        RECT 3505.935 2434.225 3506.215 2434.505 ;
        RECT 3506.645 2434.225 3506.925 2434.505 ;
        RECT 3507.355 2434.225 3507.635 2434.505 ;
        RECT 3508.065 2434.225 3508.345 2434.505 ;
        RECT 3508.775 2434.225 3509.055 2434.505 ;
        RECT 3509.485 2434.225 3509.765 2434.505 ;
        RECT 3500.255 2433.515 3500.535 2433.795 ;
        RECT 3500.965 2433.515 3501.245 2433.795 ;
        RECT 3501.675 2433.515 3501.955 2433.795 ;
        RECT 3502.385 2433.515 3502.665 2433.795 ;
        RECT 3503.095 2433.515 3503.375 2433.795 ;
        RECT 3503.805 2433.515 3504.085 2433.795 ;
        RECT 3504.515 2433.515 3504.795 2433.795 ;
        RECT 3505.225 2433.515 3505.505 2433.795 ;
        RECT 3505.935 2433.515 3506.215 2433.795 ;
        RECT 3506.645 2433.515 3506.925 2433.795 ;
        RECT 3507.355 2433.515 3507.635 2433.795 ;
        RECT 3508.065 2433.515 3508.345 2433.795 ;
        RECT 3508.775 2433.515 3509.055 2433.795 ;
        RECT 3509.485 2433.515 3509.765 2433.795 ;
        RECT 3500.255 2432.805 3500.535 2433.085 ;
        RECT 3500.965 2432.805 3501.245 2433.085 ;
        RECT 3501.675 2432.805 3501.955 2433.085 ;
        RECT 3502.385 2432.805 3502.665 2433.085 ;
        RECT 3503.095 2432.805 3503.375 2433.085 ;
        RECT 3503.805 2432.805 3504.085 2433.085 ;
        RECT 3504.515 2432.805 3504.795 2433.085 ;
        RECT 3505.225 2432.805 3505.505 2433.085 ;
        RECT 3505.935 2432.805 3506.215 2433.085 ;
        RECT 3506.645 2432.805 3506.925 2433.085 ;
        RECT 3507.355 2432.805 3507.635 2433.085 ;
        RECT 3508.065 2432.805 3508.345 2433.085 ;
        RECT 3508.775 2432.805 3509.055 2433.085 ;
        RECT 3509.485 2432.805 3509.765 2433.085 ;
        RECT 3500.255 2432.095 3500.535 2432.375 ;
        RECT 3500.965 2432.095 3501.245 2432.375 ;
        RECT 3501.675 2432.095 3501.955 2432.375 ;
        RECT 3502.385 2432.095 3502.665 2432.375 ;
        RECT 3503.095 2432.095 3503.375 2432.375 ;
        RECT 3503.805 2432.095 3504.085 2432.375 ;
        RECT 3504.515 2432.095 3504.795 2432.375 ;
        RECT 3505.225 2432.095 3505.505 2432.375 ;
        RECT 3505.935 2432.095 3506.215 2432.375 ;
        RECT 3506.645 2432.095 3506.925 2432.375 ;
        RECT 3507.355 2432.095 3507.635 2432.375 ;
        RECT 3508.065 2432.095 3508.345 2432.375 ;
        RECT 3508.775 2432.095 3509.055 2432.375 ;
        RECT 3509.485 2432.095 3509.765 2432.375 ;
        RECT 3500.255 2431.385 3500.535 2431.665 ;
        RECT 3500.965 2431.385 3501.245 2431.665 ;
        RECT 3501.675 2431.385 3501.955 2431.665 ;
        RECT 3502.385 2431.385 3502.665 2431.665 ;
        RECT 3503.095 2431.385 3503.375 2431.665 ;
        RECT 3503.805 2431.385 3504.085 2431.665 ;
        RECT 3504.515 2431.385 3504.795 2431.665 ;
        RECT 3505.225 2431.385 3505.505 2431.665 ;
        RECT 3505.935 2431.385 3506.215 2431.665 ;
        RECT 3506.645 2431.385 3506.925 2431.665 ;
        RECT 3507.355 2431.385 3507.635 2431.665 ;
        RECT 3508.065 2431.385 3508.345 2431.665 ;
        RECT 3508.775 2431.385 3509.055 2431.665 ;
        RECT 3509.485 2431.385 3509.765 2431.665 ;
        RECT 3500.255 2428.765 3500.535 2429.045 ;
        RECT 3500.965 2428.765 3501.245 2429.045 ;
        RECT 3501.675 2428.765 3501.955 2429.045 ;
        RECT 3502.385 2428.765 3502.665 2429.045 ;
        RECT 3503.095 2428.765 3503.375 2429.045 ;
        RECT 3503.805 2428.765 3504.085 2429.045 ;
        RECT 3504.515 2428.765 3504.795 2429.045 ;
        RECT 3505.225 2428.765 3505.505 2429.045 ;
        RECT 3505.935 2428.765 3506.215 2429.045 ;
        RECT 3506.645 2428.765 3506.925 2429.045 ;
        RECT 3507.355 2428.765 3507.635 2429.045 ;
        RECT 3508.065 2428.765 3508.345 2429.045 ;
        RECT 3508.775 2428.765 3509.055 2429.045 ;
        RECT 3509.485 2428.765 3509.765 2429.045 ;
        RECT 3500.255 2428.055 3500.535 2428.335 ;
        RECT 3500.965 2428.055 3501.245 2428.335 ;
        RECT 3501.675 2428.055 3501.955 2428.335 ;
        RECT 3502.385 2428.055 3502.665 2428.335 ;
        RECT 3503.095 2428.055 3503.375 2428.335 ;
        RECT 3503.805 2428.055 3504.085 2428.335 ;
        RECT 3504.515 2428.055 3504.795 2428.335 ;
        RECT 3505.225 2428.055 3505.505 2428.335 ;
        RECT 3505.935 2428.055 3506.215 2428.335 ;
        RECT 3506.645 2428.055 3506.925 2428.335 ;
        RECT 3507.355 2428.055 3507.635 2428.335 ;
        RECT 3508.065 2428.055 3508.345 2428.335 ;
        RECT 3508.775 2428.055 3509.055 2428.335 ;
        RECT 3509.485 2428.055 3509.765 2428.335 ;
        RECT 3500.255 2427.345 3500.535 2427.625 ;
        RECT 3500.965 2427.345 3501.245 2427.625 ;
        RECT 3501.675 2427.345 3501.955 2427.625 ;
        RECT 3502.385 2427.345 3502.665 2427.625 ;
        RECT 3503.095 2427.345 3503.375 2427.625 ;
        RECT 3503.805 2427.345 3504.085 2427.625 ;
        RECT 3504.515 2427.345 3504.795 2427.625 ;
        RECT 3505.225 2427.345 3505.505 2427.625 ;
        RECT 3505.935 2427.345 3506.215 2427.625 ;
        RECT 3506.645 2427.345 3506.925 2427.625 ;
        RECT 3507.355 2427.345 3507.635 2427.625 ;
        RECT 3508.065 2427.345 3508.345 2427.625 ;
        RECT 3508.775 2427.345 3509.055 2427.625 ;
        RECT 3509.485 2427.345 3509.765 2427.625 ;
        RECT 3500.255 2426.635 3500.535 2426.915 ;
        RECT 3500.965 2426.635 3501.245 2426.915 ;
        RECT 3501.675 2426.635 3501.955 2426.915 ;
        RECT 3502.385 2426.635 3502.665 2426.915 ;
        RECT 3503.095 2426.635 3503.375 2426.915 ;
        RECT 3503.805 2426.635 3504.085 2426.915 ;
        RECT 3504.515 2426.635 3504.795 2426.915 ;
        RECT 3505.225 2426.635 3505.505 2426.915 ;
        RECT 3505.935 2426.635 3506.215 2426.915 ;
        RECT 3506.645 2426.635 3506.925 2426.915 ;
        RECT 3507.355 2426.635 3507.635 2426.915 ;
        RECT 3508.065 2426.635 3508.345 2426.915 ;
        RECT 3508.775 2426.635 3509.055 2426.915 ;
        RECT 3509.485 2426.635 3509.765 2426.915 ;
        RECT 3500.255 2425.925 3500.535 2426.205 ;
        RECT 3500.965 2425.925 3501.245 2426.205 ;
        RECT 3501.675 2425.925 3501.955 2426.205 ;
        RECT 3502.385 2425.925 3502.665 2426.205 ;
        RECT 3503.095 2425.925 3503.375 2426.205 ;
        RECT 3503.805 2425.925 3504.085 2426.205 ;
        RECT 3504.515 2425.925 3504.795 2426.205 ;
        RECT 3505.225 2425.925 3505.505 2426.205 ;
        RECT 3505.935 2425.925 3506.215 2426.205 ;
        RECT 3506.645 2425.925 3506.925 2426.205 ;
        RECT 3507.355 2425.925 3507.635 2426.205 ;
        RECT 3508.065 2425.925 3508.345 2426.205 ;
        RECT 3508.775 2425.925 3509.055 2426.205 ;
        RECT 3509.485 2425.925 3509.765 2426.205 ;
        RECT 3500.255 2425.215 3500.535 2425.495 ;
        RECT 3500.965 2425.215 3501.245 2425.495 ;
        RECT 3501.675 2425.215 3501.955 2425.495 ;
        RECT 3502.385 2425.215 3502.665 2425.495 ;
        RECT 3503.095 2425.215 3503.375 2425.495 ;
        RECT 3503.805 2425.215 3504.085 2425.495 ;
        RECT 3504.515 2425.215 3504.795 2425.495 ;
        RECT 3505.225 2425.215 3505.505 2425.495 ;
        RECT 3505.935 2425.215 3506.215 2425.495 ;
        RECT 3506.645 2425.215 3506.925 2425.495 ;
        RECT 3507.355 2425.215 3507.635 2425.495 ;
        RECT 3508.065 2425.215 3508.345 2425.495 ;
        RECT 3508.775 2425.215 3509.055 2425.495 ;
        RECT 3509.485 2425.215 3509.765 2425.495 ;
        RECT 3500.255 2424.505 3500.535 2424.785 ;
        RECT 3500.965 2424.505 3501.245 2424.785 ;
        RECT 3501.675 2424.505 3501.955 2424.785 ;
        RECT 3502.385 2424.505 3502.665 2424.785 ;
        RECT 3503.095 2424.505 3503.375 2424.785 ;
        RECT 3503.805 2424.505 3504.085 2424.785 ;
        RECT 3504.515 2424.505 3504.795 2424.785 ;
        RECT 3505.225 2424.505 3505.505 2424.785 ;
        RECT 3505.935 2424.505 3506.215 2424.785 ;
        RECT 3506.645 2424.505 3506.925 2424.785 ;
        RECT 3507.355 2424.505 3507.635 2424.785 ;
        RECT 3508.065 2424.505 3508.345 2424.785 ;
        RECT 3508.775 2424.505 3509.055 2424.785 ;
        RECT 3509.485 2424.505 3509.765 2424.785 ;
        RECT 3500.255 2423.795 3500.535 2424.075 ;
        RECT 3500.965 2423.795 3501.245 2424.075 ;
        RECT 3501.675 2423.795 3501.955 2424.075 ;
        RECT 3502.385 2423.795 3502.665 2424.075 ;
        RECT 3503.095 2423.795 3503.375 2424.075 ;
        RECT 3503.805 2423.795 3504.085 2424.075 ;
        RECT 3504.515 2423.795 3504.795 2424.075 ;
        RECT 3505.225 2423.795 3505.505 2424.075 ;
        RECT 3505.935 2423.795 3506.215 2424.075 ;
        RECT 3506.645 2423.795 3506.925 2424.075 ;
        RECT 3507.355 2423.795 3507.635 2424.075 ;
        RECT 3508.065 2423.795 3508.345 2424.075 ;
        RECT 3508.775 2423.795 3509.055 2424.075 ;
        RECT 3509.485 2423.795 3509.765 2424.075 ;
        RECT 3500.255 2423.085 3500.535 2423.365 ;
        RECT 3500.965 2423.085 3501.245 2423.365 ;
        RECT 3501.675 2423.085 3501.955 2423.365 ;
        RECT 3502.385 2423.085 3502.665 2423.365 ;
        RECT 3503.095 2423.085 3503.375 2423.365 ;
        RECT 3503.805 2423.085 3504.085 2423.365 ;
        RECT 3504.515 2423.085 3504.795 2423.365 ;
        RECT 3505.225 2423.085 3505.505 2423.365 ;
        RECT 3505.935 2423.085 3506.215 2423.365 ;
        RECT 3506.645 2423.085 3506.925 2423.365 ;
        RECT 3507.355 2423.085 3507.635 2423.365 ;
        RECT 3508.065 2423.085 3508.345 2423.365 ;
        RECT 3508.775 2423.085 3509.055 2423.365 ;
        RECT 3509.485 2423.085 3509.765 2423.365 ;
        RECT 3500.255 2422.375 3500.535 2422.655 ;
        RECT 3500.965 2422.375 3501.245 2422.655 ;
        RECT 3501.675 2422.375 3501.955 2422.655 ;
        RECT 3502.385 2422.375 3502.665 2422.655 ;
        RECT 3503.095 2422.375 3503.375 2422.655 ;
        RECT 3503.805 2422.375 3504.085 2422.655 ;
        RECT 3504.515 2422.375 3504.795 2422.655 ;
        RECT 3505.225 2422.375 3505.505 2422.655 ;
        RECT 3505.935 2422.375 3506.215 2422.655 ;
        RECT 3506.645 2422.375 3506.925 2422.655 ;
        RECT 3507.355 2422.375 3507.635 2422.655 ;
        RECT 3508.065 2422.375 3508.345 2422.655 ;
        RECT 3508.775 2422.375 3509.055 2422.655 ;
        RECT 3509.485 2422.375 3509.765 2422.655 ;
        RECT 3500.255 2421.665 3500.535 2421.945 ;
        RECT 3500.965 2421.665 3501.245 2421.945 ;
        RECT 3501.675 2421.665 3501.955 2421.945 ;
        RECT 3502.385 2421.665 3502.665 2421.945 ;
        RECT 3503.095 2421.665 3503.375 2421.945 ;
        RECT 3503.805 2421.665 3504.085 2421.945 ;
        RECT 3504.515 2421.665 3504.795 2421.945 ;
        RECT 3505.225 2421.665 3505.505 2421.945 ;
        RECT 3505.935 2421.665 3506.215 2421.945 ;
        RECT 3506.645 2421.665 3506.925 2421.945 ;
        RECT 3507.355 2421.665 3507.635 2421.945 ;
        RECT 3508.065 2421.665 3508.345 2421.945 ;
        RECT 3508.775 2421.665 3509.055 2421.945 ;
        RECT 3509.485 2421.665 3509.765 2421.945 ;
        RECT 3500.255 2420.955 3500.535 2421.235 ;
        RECT 3500.965 2420.955 3501.245 2421.235 ;
        RECT 3501.675 2420.955 3501.955 2421.235 ;
        RECT 3502.385 2420.955 3502.665 2421.235 ;
        RECT 3503.095 2420.955 3503.375 2421.235 ;
        RECT 3503.805 2420.955 3504.085 2421.235 ;
        RECT 3504.515 2420.955 3504.795 2421.235 ;
        RECT 3505.225 2420.955 3505.505 2421.235 ;
        RECT 3505.935 2420.955 3506.215 2421.235 ;
        RECT 3506.645 2420.955 3506.925 2421.235 ;
        RECT 3507.355 2420.955 3507.635 2421.235 ;
        RECT 3508.065 2420.955 3508.345 2421.235 ;
        RECT 3508.775 2420.955 3509.055 2421.235 ;
        RECT 3509.485 2420.955 3509.765 2421.235 ;
        RECT 3500.255 2420.245 3500.535 2420.525 ;
        RECT 3500.965 2420.245 3501.245 2420.525 ;
        RECT 3501.675 2420.245 3501.955 2420.525 ;
        RECT 3502.385 2420.245 3502.665 2420.525 ;
        RECT 3503.095 2420.245 3503.375 2420.525 ;
        RECT 3503.805 2420.245 3504.085 2420.525 ;
        RECT 3504.515 2420.245 3504.795 2420.525 ;
        RECT 3505.225 2420.245 3505.505 2420.525 ;
        RECT 3505.935 2420.245 3506.215 2420.525 ;
        RECT 3506.645 2420.245 3506.925 2420.525 ;
        RECT 3507.355 2420.245 3507.635 2420.525 ;
        RECT 3508.065 2420.245 3508.345 2420.525 ;
        RECT 3508.775 2420.245 3509.055 2420.525 ;
        RECT 3509.485 2420.245 3509.765 2420.525 ;
        RECT 3500.255 2419.535 3500.535 2419.815 ;
        RECT 3500.965 2419.535 3501.245 2419.815 ;
        RECT 3501.675 2419.535 3501.955 2419.815 ;
        RECT 3502.385 2419.535 3502.665 2419.815 ;
        RECT 3503.095 2419.535 3503.375 2419.815 ;
        RECT 3503.805 2419.535 3504.085 2419.815 ;
        RECT 3504.515 2419.535 3504.795 2419.815 ;
        RECT 3505.225 2419.535 3505.505 2419.815 ;
        RECT 3505.935 2419.535 3506.215 2419.815 ;
        RECT 3506.645 2419.535 3506.925 2419.815 ;
        RECT 3507.355 2419.535 3507.635 2419.815 ;
        RECT 3508.065 2419.535 3508.345 2419.815 ;
        RECT 3508.775 2419.535 3509.055 2419.815 ;
        RECT 3509.485 2419.535 3509.765 2419.815 ;
        RECT 3500.255 2415.235 3500.535 2415.515 ;
        RECT 3500.965 2415.235 3501.245 2415.515 ;
        RECT 3501.675 2415.235 3501.955 2415.515 ;
        RECT 3502.385 2415.235 3502.665 2415.515 ;
        RECT 3503.095 2415.235 3503.375 2415.515 ;
        RECT 3503.805 2415.235 3504.085 2415.515 ;
        RECT 3504.515 2415.235 3504.795 2415.515 ;
        RECT 3505.225 2415.235 3505.505 2415.515 ;
        RECT 3505.935 2415.235 3506.215 2415.515 ;
        RECT 3506.645 2415.235 3506.925 2415.515 ;
        RECT 3507.355 2415.235 3507.635 2415.515 ;
        RECT 3508.065 2415.235 3508.345 2415.515 ;
        RECT 3508.775 2415.235 3509.055 2415.515 ;
        RECT 3509.485 2415.235 3509.765 2415.515 ;
        RECT 3500.255 2414.525 3500.535 2414.805 ;
        RECT 3500.965 2414.525 3501.245 2414.805 ;
        RECT 3501.675 2414.525 3501.955 2414.805 ;
        RECT 3502.385 2414.525 3502.665 2414.805 ;
        RECT 3503.095 2414.525 3503.375 2414.805 ;
        RECT 3503.805 2414.525 3504.085 2414.805 ;
        RECT 3504.515 2414.525 3504.795 2414.805 ;
        RECT 3505.225 2414.525 3505.505 2414.805 ;
        RECT 3505.935 2414.525 3506.215 2414.805 ;
        RECT 3506.645 2414.525 3506.925 2414.805 ;
        RECT 3507.355 2414.525 3507.635 2414.805 ;
        RECT 3508.065 2414.525 3508.345 2414.805 ;
        RECT 3508.775 2414.525 3509.055 2414.805 ;
        RECT 3509.485 2414.525 3509.765 2414.805 ;
        RECT 3500.255 2413.815 3500.535 2414.095 ;
        RECT 3500.965 2413.815 3501.245 2414.095 ;
        RECT 3501.675 2413.815 3501.955 2414.095 ;
        RECT 3502.385 2413.815 3502.665 2414.095 ;
        RECT 3503.095 2413.815 3503.375 2414.095 ;
        RECT 3503.805 2413.815 3504.085 2414.095 ;
        RECT 3504.515 2413.815 3504.795 2414.095 ;
        RECT 3505.225 2413.815 3505.505 2414.095 ;
        RECT 3505.935 2413.815 3506.215 2414.095 ;
        RECT 3506.645 2413.815 3506.925 2414.095 ;
        RECT 3507.355 2413.815 3507.635 2414.095 ;
        RECT 3508.065 2413.815 3508.345 2414.095 ;
        RECT 3508.775 2413.815 3509.055 2414.095 ;
        RECT 3509.485 2413.815 3509.765 2414.095 ;
        RECT 3500.255 2413.105 3500.535 2413.385 ;
        RECT 3500.965 2413.105 3501.245 2413.385 ;
        RECT 3501.675 2413.105 3501.955 2413.385 ;
        RECT 3502.385 2413.105 3502.665 2413.385 ;
        RECT 3503.095 2413.105 3503.375 2413.385 ;
        RECT 3503.805 2413.105 3504.085 2413.385 ;
        RECT 3504.515 2413.105 3504.795 2413.385 ;
        RECT 3505.225 2413.105 3505.505 2413.385 ;
        RECT 3505.935 2413.105 3506.215 2413.385 ;
        RECT 3506.645 2413.105 3506.925 2413.385 ;
        RECT 3507.355 2413.105 3507.635 2413.385 ;
        RECT 3508.065 2413.105 3508.345 2413.385 ;
        RECT 3508.775 2413.105 3509.055 2413.385 ;
        RECT 3509.485 2413.105 3509.765 2413.385 ;
        RECT 3500.255 2412.395 3500.535 2412.675 ;
        RECT 3500.965 2412.395 3501.245 2412.675 ;
        RECT 3501.675 2412.395 3501.955 2412.675 ;
        RECT 3502.385 2412.395 3502.665 2412.675 ;
        RECT 3503.095 2412.395 3503.375 2412.675 ;
        RECT 3503.805 2412.395 3504.085 2412.675 ;
        RECT 3504.515 2412.395 3504.795 2412.675 ;
        RECT 3505.225 2412.395 3505.505 2412.675 ;
        RECT 3505.935 2412.395 3506.215 2412.675 ;
        RECT 3506.645 2412.395 3506.925 2412.675 ;
        RECT 3507.355 2412.395 3507.635 2412.675 ;
        RECT 3508.065 2412.395 3508.345 2412.675 ;
        RECT 3508.775 2412.395 3509.055 2412.675 ;
        RECT 3509.485 2412.395 3509.765 2412.675 ;
        RECT 3500.255 2411.685 3500.535 2411.965 ;
        RECT 3500.965 2411.685 3501.245 2411.965 ;
        RECT 3501.675 2411.685 3501.955 2411.965 ;
        RECT 3502.385 2411.685 3502.665 2411.965 ;
        RECT 3503.095 2411.685 3503.375 2411.965 ;
        RECT 3503.805 2411.685 3504.085 2411.965 ;
        RECT 3504.515 2411.685 3504.795 2411.965 ;
        RECT 3505.225 2411.685 3505.505 2411.965 ;
        RECT 3505.935 2411.685 3506.215 2411.965 ;
        RECT 3506.645 2411.685 3506.925 2411.965 ;
        RECT 3507.355 2411.685 3507.635 2411.965 ;
        RECT 3508.065 2411.685 3508.345 2411.965 ;
        RECT 3508.775 2411.685 3509.055 2411.965 ;
        RECT 3509.485 2411.685 3509.765 2411.965 ;
        RECT 3500.255 2410.975 3500.535 2411.255 ;
        RECT 3500.965 2410.975 3501.245 2411.255 ;
        RECT 3501.675 2410.975 3501.955 2411.255 ;
        RECT 3502.385 2410.975 3502.665 2411.255 ;
        RECT 3503.095 2410.975 3503.375 2411.255 ;
        RECT 3503.805 2410.975 3504.085 2411.255 ;
        RECT 3504.515 2410.975 3504.795 2411.255 ;
        RECT 3505.225 2410.975 3505.505 2411.255 ;
        RECT 3505.935 2410.975 3506.215 2411.255 ;
        RECT 3506.645 2410.975 3506.925 2411.255 ;
        RECT 3507.355 2410.975 3507.635 2411.255 ;
        RECT 3508.065 2410.975 3508.345 2411.255 ;
        RECT 3508.775 2410.975 3509.055 2411.255 ;
        RECT 3509.485 2410.975 3509.765 2411.255 ;
        RECT 3500.255 2410.265 3500.535 2410.545 ;
        RECT 3500.965 2410.265 3501.245 2410.545 ;
        RECT 3501.675 2410.265 3501.955 2410.545 ;
        RECT 3502.385 2410.265 3502.665 2410.545 ;
        RECT 3503.095 2410.265 3503.375 2410.545 ;
        RECT 3503.805 2410.265 3504.085 2410.545 ;
        RECT 3504.515 2410.265 3504.795 2410.545 ;
        RECT 3505.225 2410.265 3505.505 2410.545 ;
        RECT 3505.935 2410.265 3506.215 2410.545 ;
        RECT 3506.645 2410.265 3506.925 2410.545 ;
        RECT 3507.355 2410.265 3507.635 2410.545 ;
        RECT 3508.065 2410.265 3508.345 2410.545 ;
        RECT 3508.775 2410.265 3509.055 2410.545 ;
        RECT 3509.485 2410.265 3509.765 2410.545 ;
        RECT 3500.255 2409.555 3500.535 2409.835 ;
        RECT 3500.965 2409.555 3501.245 2409.835 ;
        RECT 3501.675 2409.555 3501.955 2409.835 ;
        RECT 3502.385 2409.555 3502.665 2409.835 ;
        RECT 3503.095 2409.555 3503.375 2409.835 ;
        RECT 3503.805 2409.555 3504.085 2409.835 ;
        RECT 3504.515 2409.555 3504.795 2409.835 ;
        RECT 3505.225 2409.555 3505.505 2409.835 ;
        RECT 3505.935 2409.555 3506.215 2409.835 ;
        RECT 3506.645 2409.555 3506.925 2409.835 ;
        RECT 3507.355 2409.555 3507.635 2409.835 ;
        RECT 3508.065 2409.555 3508.345 2409.835 ;
        RECT 3508.775 2409.555 3509.055 2409.835 ;
        RECT 3509.485 2409.555 3509.765 2409.835 ;
        RECT 3500.255 2408.845 3500.535 2409.125 ;
        RECT 3500.965 2408.845 3501.245 2409.125 ;
        RECT 3501.675 2408.845 3501.955 2409.125 ;
        RECT 3502.385 2408.845 3502.665 2409.125 ;
        RECT 3503.095 2408.845 3503.375 2409.125 ;
        RECT 3503.805 2408.845 3504.085 2409.125 ;
        RECT 3504.515 2408.845 3504.795 2409.125 ;
        RECT 3505.225 2408.845 3505.505 2409.125 ;
        RECT 3505.935 2408.845 3506.215 2409.125 ;
        RECT 3506.645 2408.845 3506.925 2409.125 ;
        RECT 3507.355 2408.845 3507.635 2409.125 ;
        RECT 3508.065 2408.845 3508.345 2409.125 ;
        RECT 3508.775 2408.845 3509.055 2409.125 ;
        RECT 3509.485 2408.845 3509.765 2409.125 ;
        RECT 3500.255 2408.135 3500.535 2408.415 ;
        RECT 3500.965 2408.135 3501.245 2408.415 ;
        RECT 3501.675 2408.135 3501.955 2408.415 ;
        RECT 3502.385 2408.135 3502.665 2408.415 ;
        RECT 3503.095 2408.135 3503.375 2408.415 ;
        RECT 3503.805 2408.135 3504.085 2408.415 ;
        RECT 3504.515 2408.135 3504.795 2408.415 ;
        RECT 3505.225 2408.135 3505.505 2408.415 ;
        RECT 3505.935 2408.135 3506.215 2408.415 ;
        RECT 3506.645 2408.135 3506.925 2408.415 ;
        RECT 3507.355 2408.135 3507.635 2408.415 ;
        RECT 3508.065 2408.135 3508.345 2408.415 ;
        RECT 3508.775 2408.135 3509.055 2408.415 ;
        RECT 3509.485 2408.135 3509.765 2408.415 ;
        RECT 3500.255 2407.425 3500.535 2407.705 ;
        RECT 3500.965 2407.425 3501.245 2407.705 ;
        RECT 3501.675 2407.425 3501.955 2407.705 ;
        RECT 3502.385 2407.425 3502.665 2407.705 ;
        RECT 3503.095 2407.425 3503.375 2407.705 ;
        RECT 3503.805 2407.425 3504.085 2407.705 ;
        RECT 3504.515 2407.425 3504.795 2407.705 ;
        RECT 3505.225 2407.425 3505.505 2407.705 ;
        RECT 3505.935 2407.425 3506.215 2407.705 ;
        RECT 3506.645 2407.425 3506.925 2407.705 ;
        RECT 3507.355 2407.425 3507.635 2407.705 ;
        RECT 3508.065 2407.425 3508.345 2407.705 ;
        RECT 3508.775 2407.425 3509.055 2407.705 ;
        RECT 3509.485 2407.425 3509.765 2407.705 ;
        RECT 3500.255 2406.715 3500.535 2406.995 ;
        RECT 3500.965 2406.715 3501.245 2406.995 ;
        RECT 3501.675 2406.715 3501.955 2406.995 ;
        RECT 3502.385 2406.715 3502.665 2406.995 ;
        RECT 3503.095 2406.715 3503.375 2406.995 ;
        RECT 3503.805 2406.715 3504.085 2406.995 ;
        RECT 3504.515 2406.715 3504.795 2406.995 ;
        RECT 3505.225 2406.715 3505.505 2406.995 ;
        RECT 3505.935 2406.715 3506.215 2406.995 ;
        RECT 3506.645 2406.715 3506.925 2406.995 ;
        RECT 3507.355 2406.715 3507.635 2406.995 ;
        RECT 3508.065 2406.715 3508.345 2406.995 ;
        RECT 3508.775 2406.715 3509.055 2406.995 ;
        RECT 3509.485 2406.715 3509.765 2406.995 ;
        RECT 3500.255 2406.005 3500.535 2406.285 ;
        RECT 3500.965 2406.005 3501.245 2406.285 ;
        RECT 3501.675 2406.005 3501.955 2406.285 ;
        RECT 3502.385 2406.005 3502.665 2406.285 ;
        RECT 3503.095 2406.005 3503.375 2406.285 ;
        RECT 3503.805 2406.005 3504.085 2406.285 ;
        RECT 3504.515 2406.005 3504.795 2406.285 ;
        RECT 3505.225 2406.005 3505.505 2406.285 ;
        RECT 3505.935 2406.005 3506.215 2406.285 ;
        RECT 3506.645 2406.005 3506.925 2406.285 ;
        RECT 3507.355 2406.005 3507.635 2406.285 ;
        RECT 3508.065 2406.005 3508.345 2406.285 ;
        RECT 3508.775 2406.005 3509.055 2406.285 ;
        RECT 3509.485 2406.005 3509.765 2406.285 ;
        RECT 3500.255 2403.385 3500.535 2403.665 ;
        RECT 3500.965 2403.385 3501.245 2403.665 ;
        RECT 3501.675 2403.385 3501.955 2403.665 ;
        RECT 3502.385 2403.385 3502.665 2403.665 ;
        RECT 3503.095 2403.385 3503.375 2403.665 ;
        RECT 3503.805 2403.385 3504.085 2403.665 ;
        RECT 3504.515 2403.385 3504.795 2403.665 ;
        RECT 3505.225 2403.385 3505.505 2403.665 ;
        RECT 3505.935 2403.385 3506.215 2403.665 ;
        RECT 3506.645 2403.385 3506.925 2403.665 ;
        RECT 3507.355 2403.385 3507.635 2403.665 ;
        RECT 3508.065 2403.385 3508.345 2403.665 ;
        RECT 3508.775 2403.385 3509.055 2403.665 ;
        RECT 3509.485 2403.385 3509.765 2403.665 ;
        RECT 3500.255 2402.675 3500.535 2402.955 ;
        RECT 3500.965 2402.675 3501.245 2402.955 ;
        RECT 3501.675 2402.675 3501.955 2402.955 ;
        RECT 3502.385 2402.675 3502.665 2402.955 ;
        RECT 3503.095 2402.675 3503.375 2402.955 ;
        RECT 3503.805 2402.675 3504.085 2402.955 ;
        RECT 3504.515 2402.675 3504.795 2402.955 ;
        RECT 3505.225 2402.675 3505.505 2402.955 ;
        RECT 3505.935 2402.675 3506.215 2402.955 ;
        RECT 3506.645 2402.675 3506.925 2402.955 ;
        RECT 3507.355 2402.675 3507.635 2402.955 ;
        RECT 3508.065 2402.675 3508.345 2402.955 ;
        RECT 3508.775 2402.675 3509.055 2402.955 ;
        RECT 3509.485 2402.675 3509.765 2402.955 ;
        RECT 3500.255 2401.965 3500.535 2402.245 ;
        RECT 3500.965 2401.965 3501.245 2402.245 ;
        RECT 3501.675 2401.965 3501.955 2402.245 ;
        RECT 3502.385 2401.965 3502.665 2402.245 ;
        RECT 3503.095 2401.965 3503.375 2402.245 ;
        RECT 3503.805 2401.965 3504.085 2402.245 ;
        RECT 3504.515 2401.965 3504.795 2402.245 ;
        RECT 3505.225 2401.965 3505.505 2402.245 ;
        RECT 3505.935 2401.965 3506.215 2402.245 ;
        RECT 3506.645 2401.965 3506.925 2402.245 ;
        RECT 3507.355 2401.965 3507.635 2402.245 ;
        RECT 3508.065 2401.965 3508.345 2402.245 ;
        RECT 3508.775 2401.965 3509.055 2402.245 ;
        RECT 3509.485 2401.965 3509.765 2402.245 ;
        RECT 3500.255 2401.255 3500.535 2401.535 ;
        RECT 3500.965 2401.255 3501.245 2401.535 ;
        RECT 3501.675 2401.255 3501.955 2401.535 ;
        RECT 3502.385 2401.255 3502.665 2401.535 ;
        RECT 3503.095 2401.255 3503.375 2401.535 ;
        RECT 3503.805 2401.255 3504.085 2401.535 ;
        RECT 3504.515 2401.255 3504.795 2401.535 ;
        RECT 3505.225 2401.255 3505.505 2401.535 ;
        RECT 3505.935 2401.255 3506.215 2401.535 ;
        RECT 3506.645 2401.255 3506.925 2401.535 ;
        RECT 3507.355 2401.255 3507.635 2401.535 ;
        RECT 3508.065 2401.255 3508.345 2401.535 ;
        RECT 3508.775 2401.255 3509.055 2401.535 ;
        RECT 3509.485 2401.255 3509.765 2401.535 ;
        RECT 3500.255 2400.545 3500.535 2400.825 ;
        RECT 3500.965 2400.545 3501.245 2400.825 ;
        RECT 3501.675 2400.545 3501.955 2400.825 ;
        RECT 3502.385 2400.545 3502.665 2400.825 ;
        RECT 3503.095 2400.545 3503.375 2400.825 ;
        RECT 3503.805 2400.545 3504.085 2400.825 ;
        RECT 3504.515 2400.545 3504.795 2400.825 ;
        RECT 3505.225 2400.545 3505.505 2400.825 ;
        RECT 3505.935 2400.545 3506.215 2400.825 ;
        RECT 3506.645 2400.545 3506.925 2400.825 ;
        RECT 3507.355 2400.545 3507.635 2400.825 ;
        RECT 3508.065 2400.545 3508.345 2400.825 ;
        RECT 3508.775 2400.545 3509.055 2400.825 ;
        RECT 3509.485 2400.545 3509.765 2400.825 ;
        RECT 3500.255 2399.835 3500.535 2400.115 ;
        RECT 3500.965 2399.835 3501.245 2400.115 ;
        RECT 3501.675 2399.835 3501.955 2400.115 ;
        RECT 3502.385 2399.835 3502.665 2400.115 ;
        RECT 3503.095 2399.835 3503.375 2400.115 ;
        RECT 3503.805 2399.835 3504.085 2400.115 ;
        RECT 3504.515 2399.835 3504.795 2400.115 ;
        RECT 3505.225 2399.835 3505.505 2400.115 ;
        RECT 3505.935 2399.835 3506.215 2400.115 ;
        RECT 3506.645 2399.835 3506.925 2400.115 ;
        RECT 3507.355 2399.835 3507.635 2400.115 ;
        RECT 3508.065 2399.835 3508.345 2400.115 ;
        RECT 3508.775 2399.835 3509.055 2400.115 ;
        RECT 3509.485 2399.835 3509.765 2400.115 ;
        RECT 3500.255 2399.125 3500.535 2399.405 ;
        RECT 3500.965 2399.125 3501.245 2399.405 ;
        RECT 3501.675 2399.125 3501.955 2399.405 ;
        RECT 3502.385 2399.125 3502.665 2399.405 ;
        RECT 3503.095 2399.125 3503.375 2399.405 ;
        RECT 3503.805 2399.125 3504.085 2399.405 ;
        RECT 3504.515 2399.125 3504.795 2399.405 ;
        RECT 3505.225 2399.125 3505.505 2399.405 ;
        RECT 3505.935 2399.125 3506.215 2399.405 ;
        RECT 3506.645 2399.125 3506.925 2399.405 ;
        RECT 3507.355 2399.125 3507.635 2399.405 ;
        RECT 3508.065 2399.125 3508.345 2399.405 ;
        RECT 3508.775 2399.125 3509.055 2399.405 ;
        RECT 3509.485 2399.125 3509.765 2399.405 ;
        RECT 3500.255 2398.415 3500.535 2398.695 ;
        RECT 3500.965 2398.415 3501.245 2398.695 ;
        RECT 3501.675 2398.415 3501.955 2398.695 ;
        RECT 3502.385 2398.415 3502.665 2398.695 ;
        RECT 3503.095 2398.415 3503.375 2398.695 ;
        RECT 3503.805 2398.415 3504.085 2398.695 ;
        RECT 3504.515 2398.415 3504.795 2398.695 ;
        RECT 3505.225 2398.415 3505.505 2398.695 ;
        RECT 3505.935 2398.415 3506.215 2398.695 ;
        RECT 3506.645 2398.415 3506.925 2398.695 ;
        RECT 3507.355 2398.415 3507.635 2398.695 ;
        RECT 3508.065 2398.415 3508.345 2398.695 ;
        RECT 3508.775 2398.415 3509.055 2398.695 ;
        RECT 3509.485 2398.415 3509.765 2398.695 ;
        RECT 3500.255 2397.705 3500.535 2397.985 ;
        RECT 3500.965 2397.705 3501.245 2397.985 ;
        RECT 3501.675 2397.705 3501.955 2397.985 ;
        RECT 3502.385 2397.705 3502.665 2397.985 ;
        RECT 3503.095 2397.705 3503.375 2397.985 ;
        RECT 3503.805 2397.705 3504.085 2397.985 ;
        RECT 3504.515 2397.705 3504.795 2397.985 ;
        RECT 3505.225 2397.705 3505.505 2397.985 ;
        RECT 3505.935 2397.705 3506.215 2397.985 ;
        RECT 3506.645 2397.705 3506.925 2397.985 ;
        RECT 3507.355 2397.705 3507.635 2397.985 ;
        RECT 3508.065 2397.705 3508.345 2397.985 ;
        RECT 3508.775 2397.705 3509.055 2397.985 ;
        RECT 3509.485 2397.705 3509.765 2397.985 ;
        RECT 3500.255 2396.995 3500.535 2397.275 ;
        RECT 3500.965 2396.995 3501.245 2397.275 ;
        RECT 3501.675 2396.995 3501.955 2397.275 ;
        RECT 3502.385 2396.995 3502.665 2397.275 ;
        RECT 3503.095 2396.995 3503.375 2397.275 ;
        RECT 3503.805 2396.995 3504.085 2397.275 ;
        RECT 3504.515 2396.995 3504.795 2397.275 ;
        RECT 3505.225 2396.995 3505.505 2397.275 ;
        RECT 3505.935 2396.995 3506.215 2397.275 ;
        RECT 3506.645 2396.995 3506.925 2397.275 ;
        RECT 3507.355 2396.995 3507.635 2397.275 ;
        RECT 3508.065 2396.995 3508.345 2397.275 ;
        RECT 3508.775 2396.995 3509.055 2397.275 ;
        RECT 3509.485 2396.995 3509.765 2397.275 ;
        RECT 3500.255 2396.285 3500.535 2396.565 ;
        RECT 3500.965 2396.285 3501.245 2396.565 ;
        RECT 3501.675 2396.285 3501.955 2396.565 ;
        RECT 3502.385 2396.285 3502.665 2396.565 ;
        RECT 3503.095 2396.285 3503.375 2396.565 ;
        RECT 3503.805 2396.285 3504.085 2396.565 ;
        RECT 3504.515 2396.285 3504.795 2396.565 ;
        RECT 3505.225 2396.285 3505.505 2396.565 ;
        RECT 3505.935 2396.285 3506.215 2396.565 ;
        RECT 3506.645 2396.285 3506.925 2396.565 ;
        RECT 3507.355 2396.285 3507.635 2396.565 ;
        RECT 3508.065 2396.285 3508.345 2396.565 ;
        RECT 3508.775 2396.285 3509.055 2396.565 ;
        RECT 3509.485 2396.285 3509.765 2396.565 ;
        RECT 3500.255 2395.575 3500.535 2395.855 ;
        RECT 3500.965 2395.575 3501.245 2395.855 ;
        RECT 3501.675 2395.575 3501.955 2395.855 ;
        RECT 3502.385 2395.575 3502.665 2395.855 ;
        RECT 3503.095 2395.575 3503.375 2395.855 ;
        RECT 3503.805 2395.575 3504.085 2395.855 ;
        RECT 3504.515 2395.575 3504.795 2395.855 ;
        RECT 3505.225 2395.575 3505.505 2395.855 ;
        RECT 3505.935 2395.575 3506.215 2395.855 ;
        RECT 3506.645 2395.575 3506.925 2395.855 ;
        RECT 3507.355 2395.575 3507.635 2395.855 ;
        RECT 3508.065 2395.575 3508.345 2395.855 ;
        RECT 3508.775 2395.575 3509.055 2395.855 ;
        RECT 3509.485 2395.575 3509.765 2395.855 ;
        RECT 3500.255 2394.865 3500.535 2395.145 ;
        RECT 3500.965 2394.865 3501.245 2395.145 ;
        RECT 3501.675 2394.865 3501.955 2395.145 ;
        RECT 3502.385 2394.865 3502.665 2395.145 ;
        RECT 3503.095 2394.865 3503.375 2395.145 ;
        RECT 3503.805 2394.865 3504.085 2395.145 ;
        RECT 3504.515 2394.865 3504.795 2395.145 ;
        RECT 3505.225 2394.865 3505.505 2395.145 ;
        RECT 3505.935 2394.865 3506.215 2395.145 ;
        RECT 3506.645 2394.865 3506.925 2395.145 ;
        RECT 3507.355 2394.865 3507.635 2395.145 ;
        RECT 3508.065 2394.865 3508.345 2395.145 ;
        RECT 3508.775 2394.865 3509.055 2395.145 ;
        RECT 3509.485 2394.865 3509.765 2395.145 ;
        RECT 3500.255 2394.155 3500.535 2394.435 ;
        RECT 3500.965 2394.155 3501.245 2394.435 ;
        RECT 3501.675 2394.155 3501.955 2394.435 ;
        RECT 3502.385 2394.155 3502.665 2394.435 ;
        RECT 3503.095 2394.155 3503.375 2394.435 ;
        RECT 3503.805 2394.155 3504.085 2394.435 ;
        RECT 3504.515 2394.155 3504.795 2394.435 ;
        RECT 3505.225 2394.155 3505.505 2394.435 ;
        RECT 3505.935 2394.155 3506.215 2394.435 ;
        RECT 3506.645 2394.155 3506.925 2394.435 ;
        RECT 3507.355 2394.155 3507.635 2394.435 ;
        RECT 3508.065 2394.155 3508.345 2394.435 ;
        RECT 3508.775 2394.155 3509.055 2394.435 ;
        RECT 3509.485 2394.155 3509.765 2394.435 ;
        RECT 3500.200 2390.270 3500.480 2390.550 ;
        RECT 3500.910 2390.270 3501.190 2390.550 ;
        RECT 3501.620 2390.270 3501.900 2390.550 ;
        RECT 3502.330 2390.270 3502.610 2390.550 ;
        RECT 3503.040 2390.270 3503.320 2390.550 ;
        RECT 3503.750 2390.270 3504.030 2390.550 ;
        RECT 3504.460 2390.270 3504.740 2390.550 ;
        RECT 3505.170 2390.270 3505.450 2390.550 ;
        RECT 3505.880 2390.270 3506.160 2390.550 ;
        RECT 3506.590 2390.270 3506.870 2390.550 ;
        RECT 3507.300 2390.270 3507.580 2390.550 ;
        RECT 3508.010 2390.270 3508.290 2390.550 ;
        RECT 3508.720 2390.270 3509.000 2390.550 ;
        RECT 3509.430 2390.270 3509.710 2390.550 ;
        RECT 3500.200 2389.560 3500.480 2389.840 ;
        RECT 3500.910 2389.560 3501.190 2389.840 ;
        RECT 3501.620 2389.560 3501.900 2389.840 ;
        RECT 3502.330 2389.560 3502.610 2389.840 ;
        RECT 3503.040 2389.560 3503.320 2389.840 ;
        RECT 3503.750 2389.560 3504.030 2389.840 ;
        RECT 3504.460 2389.560 3504.740 2389.840 ;
        RECT 3505.170 2389.560 3505.450 2389.840 ;
        RECT 3505.880 2389.560 3506.160 2389.840 ;
        RECT 3506.590 2389.560 3506.870 2389.840 ;
        RECT 3507.300 2389.560 3507.580 2389.840 ;
        RECT 3508.010 2389.560 3508.290 2389.840 ;
        RECT 3508.720 2389.560 3509.000 2389.840 ;
        RECT 3509.430 2389.560 3509.710 2389.840 ;
        RECT 3500.200 2388.850 3500.480 2389.130 ;
        RECT 3500.910 2388.850 3501.190 2389.130 ;
        RECT 3501.620 2388.850 3501.900 2389.130 ;
        RECT 3502.330 2388.850 3502.610 2389.130 ;
        RECT 3503.040 2388.850 3503.320 2389.130 ;
        RECT 3503.750 2388.850 3504.030 2389.130 ;
        RECT 3504.460 2388.850 3504.740 2389.130 ;
        RECT 3505.170 2388.850 3505.450 2389.130 ;
        RECT 3505.880 2388.850 3506.160 2389.130 ;
        RECT 3506.590 2388.850 3506.870 2389.130 ;
        RECT 3507.300 2388.850 3507.580 2389.130 ;
        RECT 3508.010 2388.850 3508.290 2389.130 ;
        RECT 3508.720 2388.850 3509.000 2389.130 ;
        RECT 3509.430 2388.850 3509.710 2389.130 ;
        RECT 3500.200 2388.140 3500.480 2388.420 ;
        RECT 3500.910 2388.140 3501.190 2388.420 ;
        RECT 3501.620 2388.140 3501.900 2388.420 ;
        RECT 3502.330 2388.140 3502.610 2388.420 ;
        RECT 3503.040 2388.140 3503.320 2388.420 ;
        RECT 3503.750 2388.140 3504.030 2388.420 ;
        RECT 3504.460 2388.140 3504.740 2388.420 ;
        RECT 3505.170 2388.140 3505.450 2388.420 ;
        RECT 3505.880 2388.140 3506.160 2388.420 ;
        RECT 3506.590 2388.140 3506.870 2388.420 ;
        RECT 3507.300 2388.140 3507.580 2388.420 ;
        RECT 3508.010 2388.140 3508.290 2388.420 ;
        RECT 3508.720 2388.140 3509.000 2388.420 ;
        RECT 3509.430 2388.140 3509.710 2388.420 ;
        RECT 3500.200 2387.430 3500.480 2387.710 ;
        RECT 3500.910 2387.430 3501.190 2387.710 ;
        RECT 3501.620 2387.430 3501.900 2387.710 ;
        RECT 3502.330 2387.430 3502.610 2387.710 ;
        RECT 3503.040 2387.430 3503.320 2387.710 ;
        RECT 3503.750 2387.430 3504.030 2387.710 ;
        RECT 3504.460 2387.430 3504.740 2387.710 ;
        RECT 3505.170 2387.430 3505.450 2387.710 ;
        RECT 3505.880 2387.430 3506.160 2387.710 ;
        RECT 3506.590 2387.430 3506.870 2387.710 ;
        RECT 3507.300 2387.430 3507.580 2387.710 ;
        RECT 3508.010 2387.430 3508.290 2387.710 ;
        RECT 3508.720 2387.430 3509.000 2387.710 ;
        RECT 3509.430 2387.430 3509.710 2387.710 ;
        RECT 3500.200 2386.720 3500.480 2387.000 ;
        RECT 3500.910 2386.720 3501.190 2387.000 ;
        RECT 3501.620 2386.720 3501.900 2387.000 ;
        RECT 3502.330 2386.720 3502.610 2387.000 ;
        RECT 3503.040 2386.720 3503.320 2387.000 ;
        RECT 3503.750 2386.720 3504.030 2387.000 ;
        RECT 3504.460 2386.720 3504.740 2387.000 ;
        RECT 3505.170 2386.720 3505.450 2387.000 ;
        RECT 3505.880 2386.720 3506.160 2387.000 ;
        RECT 3506.590 2386.720 3506.870 2387.000 ;
        RECT 3507.300 2386.720 3507.580 2387.000 ;
        RECT 3508.010 2386.720 3508.290 2387.000 ;
        RECT 3508.720 2386.720 3509.000 2387.000 ;
        RECT 3509.430 2386.720 3509.710 2387.000 ;
        RECT 3500.200 2386.010 3500.480 2386.290 ;
        RECT 3500.910 2386.010 3501.190 2386.290 ;
        RECT 3501.620 2386.010 3501.900 2386.290 ;
        RECT 3502.330 2386.010 3502.610 2386.290 ;
        RECT 3503.040 2386.010 3503.320 2386.290 ;
        RECT 3503.750 2386.010 3504.030 2386.290 ;
        RECT 3504.460 2386.010 3504.740 2386.290 ;
        RECT 3505.170 2386.010 3505.450 2386.290 ;
        RECT 3505.880 2386.010 3506.160 2386.290 ;
        RECT 3506.590 2386.010 3506.870 2386.290 ;
        RECT 3507.300 2386.010 3507.580 2386.290 ;
        RECT 3508.010 2386.010 3508.290 2386.290 ;
        RECT 3508.720 2386.010 3509.000 2386.290 ;
        RECT 3509.430 2386.010 3509.710 2386.290 ;
        RECT 3500.200 2385.300 3500.480 2385.580 ;
        RECT 3500.910 2385.300 3501.190 2385.580 ;
        RECT 3501.620 2385.300 3501.900 2385.580 ;
        RECT 3502.330 2385.300 3502.610 2385.580 ;
        RECT 3503.040 2385.300 3503.320 2385.580 ;
        RECT 3503.750 2385.300 3504.030 2385.580 ;
        RECT 3504.460 2385.300 3504.740 2385.580 ;
        RECT 3505.170 2385.300 3505.450 2385.580 ;
        RECT 3505.880 2385.300 3506.160 2385.580 ;
        RECT 3506.590 2385.300 3506.870 2385.580 ;
        RECT 3507.300 2385.300 3507.580 2385.580 ;
        RECT 3508.010 2385.300 3508.290 2385.580 ;
        RECT 3508.720 2385.300 3509.000 2385.580 ;
        RECT 3509.430 2385.300 3509.710 2385.580 ;
        RECT 3500.200 2384.590 3500.480 2384.870 ;
        RECT 3500.910 2384.590 3501.190 2384.870 ;
        RECT 3501.620 2384.590 3501.900 2384.870 ;
        RECT 3502.330 2384.590 3502.610 2384.870 ;
        RECT 3503.040 2384.590 3503.320 2384.870 ;
        RECT 3503.750 2384.590 3504.030 2384.870 ;
        RECT 3504.460 2384.590 3504.740 2384.870 ;
        RECT 3505.170 2384.590 3505.450 2384.870 ;
        RECT 3505.880 2384.590 3506.160 2384.870 ;
        RECT 3506.590 2384.590 3506.870 2384.870 ;
        RECT 3507.300 2384.590 3507.580 2384.870 ;
        RECT 3508.010 2384.590 3508.290 2384.870 ;
        RECT 3508.720 2384.590 3509.000 2384.870 ;
        RECT 3509.430 2384.590 3509.710 2384.870 ;
        RECT 3500.200 2383.880 3500.480 2384.160 ;
        RECT 3500.910 2383.880 3501.190 2384.160 ;
        RECT 3501.620 2383.880 3501.900 2384.160 ;
        RECT 3502.330 2383.880 3502.610 2384.160 ;
        RECT 3503.040 2383.880 3503.320 2384.160 ;
        RECT 3503.750 2383.880 3504.030 2384.160 ;
        RECT 3504.460 2383.880 3504.740 2384.160 ;
        RECT 3505.170 2383.880 3505.450 2384.160 ;
        RECT 3505.880 2383.880 3506.160 2384.160 ;
        RECT 3506.590 2383.880 3506.870 2384.160 ;
        RECT 3507.300 2383.880 3507.580 2384.160 ;
        RECT 3508.010 2383.880 3508.290 2384.160 ;
        RECT 3508.720 2383.880 3509.000 2384.160 ;
        RECT 3509.430 2383.880 3509.710 2384.160 ;
        RECT 3500.200 2383.170 3500.480 2383.450 ;
        RECT 3500.910 2383.170 3501.190 2383.450 ;
        RECT 3501.620 2383.170 3501.900 2383.450 ;
        RECT 3502.330 2383.170 3502.610 2383.450 ;
        RECT 3503.040 2383.170 3503.320 2383.450 ;
        RECT 3503.750 2383.170 3504.030 2383.450 ;
        RECT 3504.460 2383.170 3504.740 2383.450 ;
        RECT 3505.170 2383.170 3505.450 2383.450 ;
        RECT 3505.880 2383.170 3506.160 2383.450 ;
        RECT 3506.590 2383.170 3506.870 2383.450 ;
        RECT 3507.300 2383.170 3507.580 2383.450 ;
        RECT 3508.010 2383.170 3508.290 2383.450 ;
        RECT 3508.720 2383.170 3509.000 2383.450 ;
        RECT 3509.430 2383.170 3509.710 2383.450 ;
        RECT 3500.200 2382.460 3500.480 2382.740 ;
        RECT 3500.910 2382.460 3501.190 2382.740 ;
        RECT 3501.620 2382.460 3501.900 2382.740 ;
        RECT 3502.330 2382.460 3502.610 2382.740 ;
        RECT 3503.040 2382.460 3503.320 2382.740 ;
        RECT 3503.750 2382.460 3504.030 2382.740 ;
        RECT 3504.460 2382.460 3504.740 2382.740 ;
        RECT 3505.170 2382.460 3505.450 2382.740 ;
        RECT 3505.880 2382.460 3506.160 2382.740 ;
        RECT 3506.590 2382.460 3506.870 2382.740 ;
        RECT 3507.300 2382.460 3507.580 2382.740 ;
        RECT 3508.010 2382.460 3508.290 2382.740 ;
        RECT 3508.720 2382.460 3509.000 2382.740 ;
        RECT 3509.430 2382.460 3509.710 2382.740 ;
        RECT 3500.200 2381.750 3500.480 2382.030 ;
        RECT 3500.910 2381.750 3501.190 2382.030 ;
        RECT 3501.620 2381.750 3501.900 2382.030 ;
        RECT 3502.330 2381.750 3502.610 2382.030 ;
        RECT 3503.040 2381.750 3503.320 2382.030 ;
        RECT 3503.750 2381.750 3504.030 2382.030 ;
        RECT 3504.460 2381.750 3504.740 2382.030 ;
        RECT 3505.170 2381.750 3505.450 2382.030 ;
        RECT 3505.880 2381.750 3506.160 2382.030 ;
        RECT 3506.590 2381.750 3506.870 2382.030 ;
        RECT 3507.300 2381.750 3507.580 2382.030 ;
        RECT 3508.010 2381.750 3508.290 2382.030 ;
        RECT 3508.720 2381.750 3509.000 2382.030 ;
        RECT 3509.430 2381.750 3509.710 2382.030 ;
        RECT 369.330 2342.970 369.610 2343.250 ;
        RECT 370.040 2342.970 370.320 2343.250 ;
        RECT 370.750 2342.970 371.030 2343.250 ;
        RECT 371.460 2342.970 371.740 2343.250 ;
        RECT 372.170 2342.970 372.450 2343.250 ;
        RECT 372.880 2342.970 373.160 2343.250 ;
        RECT 373.590 2342.970 373.870 2343.250 ;
        RECT 374.300 2342.970 374.580 2343.250 ;
        RECT 375.010 2342.970 375.290 2343.250 ;
        RECT 375.720 2342.970 376.000 2343.250 ;
        RECT 376.430 2342.970 376.710 2343.250 ;
        RECT 369.330 2342.260 369.610 2342.540 ;
        RECT 370.040 2342.260 370.320 2342.540 ;
        RECT 370.750 2342.260 371.030 2342.540 ;
        RECT 371.460 2342.260 371.740 2342.540 ;
        RECT 372.170 2342.260 372.450 2342.540 ;
        RECT 372.880 2342.260 373.160 2342.540 ;
        RECT 373.590 2342.260 373.870 2342.540 ;
        RECT 374.300 2342.260 374.580 2342.540 ;
        RECT 375.010 2342.260 375.290 2342.540 ;
        RECT 375.720 2342.260 376.000 2342.540 ;
        RECT 376.430 2342.260 376.710 2342.540 ;
        RECT 369.330 2341.550 369.610 2341.830 ;
        RECT 370.040 2341.550 370.320 2341.830 ;
        RECT 370.750 2341.550 371.030 2341.830 ;
        RECT 371.460 2341.550 371.740 2341.830 ;
        RECT 372.170 2341.550 372.450 2341.830 ;
        RECT 372.880 2341.550 373.160 2341.830 ;
        RECT 373.590 2341.550 373.870 2341.830 ;
        RECT 374.300 2341.550 374.580 2341.830 ;
        RECT 375.010 2341.550 375.290 2341.830 ;
        RECT 375.720 2341.550 376.000 2341.830 ;
        RECT 376.430 2341.550 376.710 2341.830 ;
        RECT 369.330 2340.840 369.610 2341.120 ;
        RECT 370.040 2340.840 370.320 2341.120 ;
        RECT 370.750 2340.840 371.030 2341.120 ;
        RECT 371.460 2340.840 371.740 2341.120 ;
        RECT 372.170 2340.840 372.450 2341.120 ;
        RECT 372.880 2340.840 373.160 2341.120 ;
        RECT 373.590 2340.840 373.870 2341.120 ;
        RECT 374.300 2340.840 374.580 2341.120 ;
        RECT 375.010 2340.840 375.290 2341.120 ;
        RECT 375.720 2340.840 376.000 2341.120 ;
        RECT 376.430 2340.840 376.710 2341.120 ;
        RECT 369.330 2340.130 369.610 2340.410 ;
        RECT 370.040 2340.130 370.320 2340.410 ;
        RECT 370.750 2340.130 371.030 2340.410 ;
        RECT 371.460 2340.130 371.740 2340.410 ;
        RECT 372.170 2340.130 372.450 2340.410 ;
        RECT 372.880 2340.130 373.160 2340.410 ;
        RECT 373.590 2340.130 373.870 2340.410 ;
        RECT 374.300 2340.130 374.580 2340.410 ;
        RECT 375.010 2340.130 375.290 2340.410 ;
        RECT 375.720 2340.130 376.000 2340.410 ;
        RECT 376.430 2340.130 376.710 2340.410 ;
        RECT 369.330 2339.420 369.610 2339.700 ;
        RECT 370.040 2339.420 370.320 2339.700 ;
        RECT 370.750 2339.420 371.030 2339.700 ;
        RECT 371.460 2339.420 371.740 2339.700 ;
        RECT 372.170 2339.420 372.450 2339.700 ;
        RECT 372.880 2339.420 373.160 2339.700 ;
        RECT 373.590 2339.420 373.870 2339.700 ;
        RECT 374.300 2339.420 374.580 2339.700 ;
        RECT 375.010 2339.420 375.290 2339.700 ;
        RECT 375.720 2339.420 376.000 2339.700 ;
        RECT 376.430 2339.420 376.710 2339.700 ;
        RECT 369.330 2338.710 369.610 2338.990 ;
        RECT 370.040 2338.710 370.320 2338.990 ;
        RECT 370.750 2338.710 371.030 2338.990 ;
        RECT 371.460 2338.710 371.740 2338.990 ;
        RECT 372.170 2338.710 372.450 2338.990 ;
        RECT 372.880 2338.710 373.160 2338.990 ;
        RECT 373.590 2338.710 373.870 2338.990 ;
        RECT 374.300 2338.710 374.580 2338.990 ;
        RECT 375.010 2338.710 375.290 2338.990 ;
        RECT 375.720 2338.710 376.000 2338.990 ;
        RECT 376.430 2338.710 376.710 2338.990 ;
        RECT 369.330 2338.000 369.610 2338.280 ;
        RECT 370.040 2338.000 370.320 2338.280 ;
        RECT 370.750 2338.000 371.030 2338.280 ;
        RECT 371.460 2338.000 371.740 2338.280 ;
        RECT 372.170 2338.000 372.450 2338.280 ;
        RECT 372.880 2338.000 373.160 2338.280 ;
        RECT 373.590 2338.000 373.870 2338.280 ;
        RECT 374.300 2338.000 374.580 2338.280 ;
        RECT 375.010 2338.000 375.290 2338.280 ;
        RECT 375.720 2338.000 376.000 2338.280 ;
        RECT 376.430 2338.000 376.710 2338.280 ;
        RECT 369.330 2337.290 369.610 2337.570 ;
        RECT 370.040 2337.290 370.320 2337.570 ;
        RECT 370.750 2337.290 371.030 2337.570 ;
        RECT 371.460 2337.290 371.740 2337.570 ;
        RECT 372.170 2337.290 372.450 2337.570 ;
        RECT 372.880 2337.290 373.160 2337.570 ;
        RECT 373.590 2337.290 373.870 2337.570 ;
        RECT 374.300 2337.290 374.580 2337.570 ;
        RECT 375.010 2337.290 375.290 2337.570 ;
        RECT 375.720 2337.290 376.000 2337.570 ;
        RECT 376.430 2337.290 376.710 2337.570 ;
        RECT 369.330 2336.580 369.610 2336.860 ;
        RECT 370.040 2336.580 370.320 2336.860 ;
        RECT 370.750 2336.580 371.030 2336.860 ;
        RECT 371.460 2336.580 371.740 2336.860 ;
        RECT 372.170 2336.580 372.450 2336.860 ;
        RECT 372.880 2336.580 373.160 2336.860 ;
        RECT 373.590 2336.580 373.870 2336.860 ;
        RECT 374.300 2336.580 374.580 2336.860 ;
        RECT 375.010 2336.580 375.290 2336.860 ;
        RECT 375.720 2336.580 376.000 2336.860 ;
        RECT 376.430 2336.580 376.710 2336.860 ;
        RECT 369.330 2335.870 369.610 2336.150 ;
        RECT 370.040 2335.870 370.320 2336.150 ;
        RECT 370.750 2335.870 371.030 2336.150 ;
        RECT 371.460 2335.870 371.740 2336.150 ;
        RECT 372.170 2335.870 372.450 2336.150 ;
        RECT 372.880 2335.870 373.160 2336.150 ;
        RECT 373.590 2335.870 373.870 2336.150 ;
        RECT 374.300 2335.870 374.580 2336.150 ;
        RECT 375.010 2335.870 375.290 2336.150 ;
        RECT 375.720 2335.870 376.000 2336.150 ;
        RECT 376.430 2335.870 376.710 2336.150 ;
        RECT 369.330 2335.160 369.610 2335.440 ;
        RECT 370.040 2335.160 370.320 2335.440 ;
        RECT 370.750 2335.160 371.030 2335.440 ;
        RECT 371.460 2335.160 371.740 2335.440 ;
        RECT 372.170 2335.160 372.450 2335.440 ;
        RECT 372.880 2335.160 373.160 2335.440 ;
        RECT 373.590 2335.160 373.870 2335.440 ;
        RECT 374.300 2335.160 374.580 2335.440 ;
        RECT 375.010 2335.160 375.290 2335.440 ;
        RECT 375.720 2335.160 376.000 2335.440 ;
        RECT 376.430 2335.160 376.710 2335.440 ;
        RECT 369.330 2334.450 369.610 2334.730 ;
        RECT 370.040 2334.450 370.320 2334.730 ;
        RECT 370.750 2334.450 371.030 2334.730 ;
        RECT 371.460 2334.450 371.740 2334.730 ;
        RECT 372.170 2334.450 372.450 2334.730 ;
        RECT 372.880 2334.450 373.160 2334.730 ;
        RECT 373.590 2334.450 373.870 2334.730 ;
        RECT 374.300 2334.450 374.580 2334.730 ;
        RECT 375.010 2334.450 375.290 2334.730 ;
        RECT 375.720 2334.450 376.000 2334.730 ;
        RECT 376.430 2334.450 376.710 2334.730 ;
        RECT 369.275 2330.565 369.555 2330.845 ;
        RECT 369.985 2330.565 370.265 2330.845 ;
        RECT 370.695 2330.565 370.975 2330.845 ;
        RECT 371.405 2330.565 371.685 2330.845 ;
        RECT 372.115 2330.565 372.395 2330.845 ;
        RECT 372.825 2330.565 373.105 2330.845 ;
        RECT 373.535 2330.565 373.815 2330.845 ;
        RECT 374.245 2330.565 374.525 2330.845 ;
        RECT 374.955 2330.565 375.235 2330.845 ;
        RECT 375.665 2330.565 375.945 2330.845 ;
        RECT 376.375 2330.565 376.655 2330.845 ;
        RECT 369.275 2329.855 369.555 2330.135 ;
        RECT 369.985 2329.855 370.265 2330.135 ;
        RECT 370.695 2329.855 370.975 2330.135 ;
        RECT 371.405 2329.855 371.685 2330.135 ;
        RECT 372.115 2329.855 372.395 2330.135 ;
        RECT 372.825 2329.855 373.105 2330.135 ;
        RECT 373.535 2329.855 373.815 2330.135 ;
        RECT 374.245 2329.855 374.525 2330.135 ;
        RECT 374.955 2329.855 375.235 2330.135 ;
        RECT 375.665 2329.855 375.945 2330.135 ;
        RECT 376.375 2329.855 376.655 2330.135 ;
        RECT 369.275 2329.145 369.555 2329.425 ;
        RECT 369.985 2329.145 370.265 2329.425 ;
        RECT 370.695 2329.145 370.975 2329.425 ;
        RECT 371.405 2329.145 371.685 2329.425 ;
        RECT 372.115 2329.145 372.395 2329.425 ;
        RECT 372.825 2329.145 373.105 2329.425 ;
        RECT 373.535 2329.145 373.815 2329.425 ;
        RECT 374.245 2329.145 374.525 2329.425 ;
        RECT 374.955 2329.145 375.235 2329.425 ;
        RECT 375.665 2329.145 375.945 2329.425 ;
        RECT 376.375 2329.145 376.655 2329.425 ;
        RECT 369.275 2328.435 369.555 2328.715 ;
        RECT 369.985 2328.435 370.265 2328.715 ;
        RECT 370.695 2328.435 370.975 2328.715 ;
        RECT 371.405 2328.435 371.685 2328.715 ;
        RECT 372.115 2328.435 372.395 2328.715 ;
        RECT 372.825 2328.435 373.105 2328.715 ;
        RECT 373.535 2328.435 373.815 2328.715 ;
        RECT 374.245 2328.435 374.525 2328.715 ;
        RECT 374.955 2328.435 375.235 2328.715 ;
        RECT 375.665 2328.435 375.945 2328.715 ;
        RECT 376.375 2328.435 376.655 2328.715 ;
        RECT 369.275 2327.725 369.555 2328.005 ;
        RECT 369.985 2327.725 370.265 2328.005 ;
        RECT 370.695 2327.725 370.975 2328.005 ;
        RECT 371.405 2327.725 371.685 2328.005 ;
        RECT 372.115 2327.725 372.395 2328.005 ;
        RECT 372.825 2327.725 373.105 2328.005 ;
        RECT 373.535 2327.725 373.815 2328.005 ;
        RECT 374.245 2327.725 374.525 2328.005 ;
        RECT 374.955 2327.725 375.235 2328.005 ;
        RECT 375.665 2327.725 375.945 2328.005 ;
        RECT 376.375 2327.725 376.655 2328.005 ;
        RECT 369.275 2327.015 369.555 2327.295 ;
        RECT 369.985 2327.015 370.265 2327.295 ;
        RECT 370.695 2327.015 370.975 2327.295 ;
        RECT 371.405 2327.015 371.685 2327.295 ;
        RECT 372.115 2327.015 372.395 2327.295 ;
        RECT 372.825 2327.015 373.105 2327.295 ;
        RECT 373.535 2327.015 373.815 2327.295 ;
        RECT 374.245 2327.015 374.525 2327.295 ;
        RECT 374.955 2327.015 375.235 2327.295 ;
        RECT 375.665 2327.015 375.945 2327.295 ;
        RECT 376.375 2327.015 376.655 2327.295 ;
        RECT 369.275 2326.305 369.555 2326.585 ;
        RECT 369.985 2326.305 370.265 2326.585 ;
        RECT 370.695 2326.305 370.975 2326.585 ;
        RECT 371.405 2326.305 371.685 2326.585 ;
        RECT 372.115 2326.305 372.395 2326.585 ;
        RECT 372.825 2326.305 373.105 2326.585 ;
        RECT 373.535 2326.305 373.815 2326.585 ;
        RECT 374.245 2326.305 374.525 2326.585 ;
        RECT 374.955 2326.305 375.235 2326.585 ;
        RECT 375.665 2326.305 375.945 2326.585 ;
        RECT 376.375 2326.305 376.655 2326.585 ;
        RECT 369.275 2325.595 369.555 2325.875 ;
        RECT 369.985 2325.595 370.265 2325.875 ;
        RECT 370.695 2325.595 370.975 2325.875 ;
        RECT 371.405 2325.595 371.685 2325.875 ;
        RECT 372.115 2325.595 372.395 2325.875 ;
        RECT 372.825 2325.595 373.105 2325.875 ;
        RECT 373.535 2325.595 373.815 2325.875 ;
        RECT 374.245 2325.595 374.525 2325.875 ;
        RECT 374.955 2325.595 375.235 2325.875 ;
        RECT 375.665 2325.595 375.945 2325.875 ;
        RECT 376.375 2325.595 376.655 2325.875 ;
        RECT 369.275 2324.885 369.555 2325.165 ;
        RECT 369.985 2324.885 370.265 2325.165 ;
        RECT 370.695 2324.885 370.975 2325.165 ;
        RECT 371.405 2324.885 371.685 2325.165 ;
        RECT 372.115 2324.885 372.395 2325.165 ;
        RECT 372.825 2324.885 373.105 2325.165 ;
        RECT 373.535 2324.885 373.815 2325.165 ;
        RECT 374.245 2324.885 374.525 2325.165 ;
        RECT 374.955 2324.885 375.235 2325.165 ;
        RECT 375.665 2324.885 375.945 2325.165 ;
        RECT 376.375 2324.885 376.655 2325.165 ;
        RECT 369.275 2324.175 369.555 2324.455 ;
        RECT 369.985 2324.175 370.265 2324.455 ;
        RECT 370.695 2324.175 370.975 2324.455 ;
        RECT 371.405 2324.175 371.685 2324.455 ;
        RECT 372.115 2324.175 372.395 2324.455 ;
        RECT 372.825 2324.175 373.105 2324.455 ;
        RECT 373.535 2324.175 373.815 2324.455 ;
        RECT 374.245 2324.175 374.525 2324.455 ;
        RECT 374.955 2324.175 375.235 2324.455 ;
        RECT 375.665 2324.175 375.945 2324.455 ;
        RECT 376.375 2324.175 376.655 2324.455 ;
        RECT 369.275 2323.465 369.555 2323.745 ;
        RECT 369.985 2323.465 370.265 2323.745 ;
        RECT 370.695 2323.465 370.975 2323.745 ;
        RECT 371.405 2323.465 371.685 2323.745 ;
        RECT 372.115 2323.465 372.395 2323.745 ;
        RECT 372.825 2323.465 373.105 2323.745 ;
        RECT 373.535 2323.465 373.815 2323.745 ;
        RECT 374.245 2323.465 374.525 2323.745 ;
        RECT 374.955 2323.465 375.235 2323.745 ;
        RECT 375.665 2323.465 375.945 2323.745 ;
        RECT 376.375 2323.465 376.655 2323.745 ;
        RECT 369.275 2322.755 369.555 2323.035 ;
        RECT 369.985 2322.755 370.265 2323.035 ;
        RECT 370.695 2322.755 370.975 2323.035 ;
        RECT 371.405 2322.755 371.685 2323.035 ;
        RECT 372.115 2322.755 372.395 2323.035 ;
        RECT 372.825 2322.755 373.105 2323.035 ;
        RECT 373.535 2322.755 373.815 2323.035 ;
        RECT 374.245 2322.755 374.525 2323.035 ;
        RECT 374.955 2322.755 375.235 2323.035 ;
        RECT 375.665 2322.755 375.945 2323.035 ;
        RECT 376.375 2322.755 376.655 2323.035 ;
        RECT 369.275 2322.045 369.555 2322.325 ;
        RECT 369.985 2322.045 370.265 2322.325 ;
        RECT 370.695 2322.045 370.975 2322.325 ;
        RECT 371.405 2322.045 371.685 2322.325 ;
        RECT 372.115 2322.045 372.395 2322.325 ;
        RECT 372.825 2322.045 373.105 2322.325 ;
        RECT 373.535 2322.045 373.815 2322.325 ;
        RECT 374.245 2322.045 374.525 2322.325 ;
        RECT 374.955 2322.045 375.235 2322.325 ;
        RECT 375.665 2322.045 375.945 2322.325 ;
        RECT 376.375 2322.045 376.655 2322.325 ;
        RECT 369.275 2321.335 369.555 2321.615 ;
        RECT 369.985 2321.335 370.265 2321.615 ;
        RECT 370.695 2321.335 370.975 2321.615 ;
        RECT 371.405 2321.335 371.685 2321.615 ;
        RECT 372.115 2321.335 372.395 2321.615 ;
        RECT 372.825 2321.335 373.105 2321.615 ;
        RECT 373.535 2321.335 373.815 2321.615 ;
        RECT 374.245 2321.335 374.525 2321.615 ;
        RECT 374.955 2321.335 375.235 2321.615 ;
        RECT 375.665 2321.335 375.945 2321.615 ;
        RECT 376.375 2321.335 376.655 2321.615 ;
        RECT 369.275 2318.715 369.555 2318.995 ;
        RECT 369.985 2318.715 370.265 2318.995 ;
        RECT 370.695 2318.715 370.975 2318.995 ;
        RECT 371.405 2318.715 371.685 2318.995 ;
        RECT 372.115 2318.715 372.395 2318.995 ;
        RECT 372.825 2318.715 373.105 2318.995 ;
        RECT 373.535 2318.715 373.815 2318.995 ;
        RECT 374.245 2318.715 374.525 2318.995 ;
        RECT 374.955 2318.715 375.235 2318.995 ;
        RECT 375.665 2318.715 375.945 2318.995 ;
        RECT 376.375 2318.715 376.655 2318.995 ;
        RECT 369.275 2318.005 369.555 2318.285 ;
        RECT 369.985 2318.005 370.265 2318.285 ;
        RECT 370.695 2318.005 370.975 2318.285 ;
        RECT 371.405 2318.005 371.685 2318.285 ;
        RECT 372.115 2318.005 372.395 2318.285 ;
        RECT 372.825 2318.005 373.105 2318.285 ;
        RECT 373.535 2318.005 373.815 2318.285 ;
        RECT 374.245 2318.005 374.525 2318.285 ;
        RECT 374.955 2318.005 375.235 2318.285 ;
        RECT 375.665 2318.005 375.945 2318.285 ;
        RECT 376.375 2318.005 376.655 2318.285 ;
        RECT 369.275 2317.295 369.555 2317.575 ;
        RECT 369.985 2317.295 370.265 2317.575 ;
        RECT 370.695 2317.295 370.975 2317.575 ;
        RECT 371.405 2317.295 371.685 2317.575 ;
        RECT 372.115 2317.295 372.395 2317.575 ;
        RECT 372.825 2317.295 373.105 2317.575 ;
        RECT 373.535 2317.295 373.815 2317.575 ;
        RECT 374.245 2317.295 374.525 2317.575 ;
        RECT 374.955 2317.295 375.235 2317.575 ;
        RECT 375.665 2317.295 375.945 2317.575 ;
        RECT 376.375 2317.295 376.655 2317.575 ;
        RECT 369.275 2316.585 369.555 2316.865 ;
        RECT 369.985 2316.585 370.265 2316.865 ;
        RECT 370.695 2316.585 370.975 2316.865 ;
        RECT 371.405 2316.585 371.685 2316.865 ;
        RECT 372.115 2316.585 372.395 2316.865 ;
        RECT 372.825 2316.585 373.105 2316.865 ;
        RECT 373.535 2316.585 373.815 2316.865 ;
        RECT 374.245 2316.585 374.525 2316.865 ;
        RECT 374.955 2316.585 375.235 2316.865 ;
        RECT 375.665 2316.585 375.945 2316.865 ;
        RECT 376.375 2316.585 376.655 2316.865 ;
        RECT 369.275 2315.875 369.555 2316.155 ;
        RECT 369.985 2315.875 370.265 2316.155 ;
        RECT 370.695 2315.875 370.975 2316.155 ;
        RECT 371.405 2315.875 371.685 2316.155 ;
        RECT 372.115 2315.875 372.395 2316.155 ;
        RECT 372.825 2315.875 373.105 2316.155 ;
        RECT 373.535 2315.875 373.815 2316.155 ;
        RECT 374.245 2315.875 374.525 2316.155 ;
        RECT 374.955 2315.875 375.235 2316.155 ;
        RECT 375.665 2315.875 375.945 2316.155 ;
        RECT 376.375 2315.875 376.655 2316.155 ;
        RECT 369.275 2315.165 369.555 2315.445 ;
        RECT 369.985 2315.165 370.265 2315.445 ;
        RECT 370.695 2315.165 370.975 2315.445 ;
        RECT 371.405 2315.165 371.685 2315.445 ;
        RECT 372.115 2315.165 372.395 2315.445 ;
        RECT 372.825 2315.165 373.105 2315.445 ;
        RECT 373.535 2315.165 373.815 2315.445 ;
        RECT 374.245 2315.165 374.525 2315.445 ;
        RECT 374.955 2315.165 375.235 2315.445 ;
        RECT 375.665 2315.165 375.945 2315.445 ;
        RECT 376.375 2315.165 376.655 2315.445 ;
        RECT 369.275 2314.455 369.555 2314.735 ;
        RECT 369.985 2314.455 370.265 2314.735 ;
        RECT 370.695 2314.455 370.975 2314.735 ;
        RECT 371.405 2314.455 371.685 2314.735 ;
        RECT 372.115 2314.455 372.395 2314.735 ;
        RECT 372.825 2314.455 373.105 2314.735 ;
        RECT 373.535 2314.455 373.815 2314.735 ;
        RECT 374.245 2314.455 374.525 2314.735 ;
        RECT 374.955 2314.455 375.235 2314.735 ;
        RECT 375.665 2314.455 375.945 2314.735 ;
        RECT 376.375 2314.455 376.655 2314.735 ;
        RECT 369.275 2313.745 369.555 2314.025 ;
        RECT 369.985 2313.745 370.265 2314.025 ;
        RECT 370.695 2313.745 370.975 2314.025 ;
        RECT 371.405 2313.745 371.685 2314.025 ;
        RECT 372.115 2313.745 372.395 2314.025 ;
        RECT 372.825 2313.745 373.105 2314.025 ;
        RECT 373.535 2313.745 373.815 2314.025 ;
        RECT 374.245 2313.745 374.525 2314.025 ;
        RECT 374.955 2313.745 375.235 2314.025 ;
        RECT 375.665 2313.745 375.945 2314.025 ;
        RECT 376.375 2313.745 376.655 2314.025 ;
        RECT 369.275 2313.035 369.555 2313.315 ;
        RECT 369.985 2313.035 370.265 2313.315 ;
        RECT 370.695 2313.035 370.975 2313.315 ;
        RECT 371.405 2313.035 371.685 2313.315 ;
        RECT 372.115 2313.035 372.395 2313.315 ;
        RECT 372.825 2313.035 373.105 2313.315 ;
        RECT 373.535 2313.035 373.815 2313.315 ;
        RECT 374.245 2313.035 374.525 2313.315 ;
        RECT 374.955 2313.035 375.235 2313.315 ;
        RECT 375.665 2313.035 375.945 2313.315 ;
        RECT 376.375 2313.035 376.655 2313.315 ;
        RECT 369.275 2312.325 369.555 2312.605 ;
        RECT 369.985 2312.325 370.265 2312.605 ;
        RECT 370.695 2312.325 370.975 2312.605 ;
        RECT 371.405 2312.325 371.685 2312.605 ;
        RECT 372.115 2312.325 372.395 2312.605 ;
        RECT 372.825 2312.325 373.105 2312.605 ;
        RECT 373.535 2312.325 373.815 2312.605 ;
        RECT 374.245 2312.325 374.525 2312.605 ;
        RECT 374.955 2312.325 375.235 2312.605 ;
        RECT 375.665 2312.325 375.945 2312.605 ;
        RECT 376.375 2312.325 376.655 2312.605 ;
        RECT 369.275 2311.615 369.555 2311.895 ;
        RECT 369.985 2311.615 370.265 2311.895 ;
        RECT 370.695 2311.615 370.975 2311.895 ;
        RECT 371.405 2311.615 371.685 2311.895 ;
        RECT 372.115 2311.615 372.395 2311.895 ;
        RECT 372.825 2311.615 373.105 2311.895 ;
        RECT 373.535 2311.615 373.815 2311.895 ;
        RECT 374.245 2311.615 374.525 2311.895 ;
        RECT 374.955 2311.615 375.235 2311.895 ;
        RECT 375.665 2311.615 375.945 2311.895 ;
        RECT 376.375 2311.615 376.655 2311.895 ;
        RECT 369.275 2310.905 369.555 2311.185 ;
        RECT 369.985 2310.905 370.265 2311.185 ;
        RECT 370.695 2310.905 370.975 2311.185 ;
        RECT 371.405 2310.905 371.685 2311.185 ;
        RECT 372.115 2310.905 372.395 2311.185 ;
        RECT 372.825 2310.905 373.105 2311.185 ;
        RECT 373.535 2310.905 373.815 2311.185 ;
        RECT 374.245 2310.905 374.525 2311.185 ;
        RECT 374.955 2310.905 375.235 2311.185 ;
        RECT 375.665 2310.905 375.945 2311.185 ;
        RECT 376.375 2310.905 376.655 2311.185 ;
        RECT 369.275 2310.195 369.555 2310.475 ;
        RECT 369.985 2310.195 370.265 2310.475 ;
        RECT 370.695 2310.195 370.975 2310.475 ;
        RECT 371.405 2310.195 371.685 2310.475 ;
        RECT 372.115 2310.195 372.395 2310.475 ;
        RECT 372.825 2310.195 373.105 2310.475 ;
        RECT 373.535 2310.195 373.815 2310.475 ;
        RECT 374.245 2310.195 374.525 2310.475 ;
        RECT 374.955 2310.195 375.235 2310.475 ;
        RECT 375.665 2310.195 375.945 2310.475 ;
        RECT 376.375 2310.195 376.655 2310.475 ;
        RECT 369.275 2309.485 369.555 2309.765 ;
        RECT 369.985 2309.485 370.265 2309.765 ;
        RECT 370.695 2309.485 370.975 2309.765 ;
        RECT 371.405 2309.485 371.685 2309.765 ;
        RECT 372.115 2309.485 372.395 2309.765 ;
        RECT 372.825 2309.485 373.105 2309.765 ;
        RECT 373.535 2309.485 373.815 2309.765 ;
        RECT 374.245 2309.485 374.525 2309.765 ;
        RECT 374.955 2309.485 375.235 2309.765 ;
        RECT 375.665 2309.485 375.945 2309.765 ;
        RECT 376.375 2309.485 376.655 2309.765 ;
        RECT 369.275 2305.185 369.555 2305.465 ;
        RECT 369.985 2305.185 370.265 2305.465 ;
        RECT 370.695 2305.185 370.975 2305.465 ;
        RECT 371.405 2305.185 371.685 2305.465 ;
        RECT 372.115 2305.185 372.395 2305.465 ;
        RECT 372.825 2305.185 373.105 2305.465 ;
        RECT 373.535 2305.185 373.815 2305.465 ;
        RECT 374.245 2305.185 374.525 2305.465 ;
        RECT 374.955 2305.185 375.235 2305.465 ;
        RECT 375.665 2305.185 375.945 2305.465 ;
        RECT 376.375 2305.185 376.655 2305.465 ;
        RECT 369.275 2304.475 369.555 2304.755 ;
        RECT 369.985 2304.475 370.265 2304.755 ;
        RECT 370.695 2304.475 370.975 2304.755 ;
        RECT 371.405 2304.475 371.685 2304.755 ;
        RECT 372.115 2304.475 372.395 2304.755 ;
        RECT 372.825 2304.475 373.105 2304.755 ;
        RECT 373.535 2304.475 373.815 2304.755 ;
        RECT 374.245 2304.475 374.525 2304.755 ;
        RECT 374.955 2304.475 375.235 2304.755 ;
        RECT 375.665 2304.475 375.945 2304.755 ;
        RECT 376.375 2304.475 376.655 2304.755 ;
        RECT 369.275 2303.765 369.555 2304.045 ;
        RECT 369.985 2303.765 370.265 2304.045 ;
        RECT 370.695 2303.765 370.975 2304.045 ;
        RECT 371.405 2303.765 371.685 2304.045 ;
        RECT 372.115 2303.765 372.395 2304.045 ;
        RECT 372.825 2303.765 373.105 2304.045 ;
        RECT 373.535 2303.765 373.815 2304.045 ;
        RECT 374.245 2303.765 374.525 2304.045 ;
        RECT 374.955 2303.765 375.235 2304.045 ;
        RECT 375.665 2303.765 375.945 2304.045 ;
        RECT 376.375 2303.765 376.655 2304.045 ;
        RECT 369.275 2303.055 369.555 2303.335 ;
        RECT 369.985 2303.055 370.265 2303.335 ;
        RECT 370.695 2303.055 370.975 2303.335 ;
        RECT 371.405 2303.055 371.685 2303.335 ;
        RECT 372.115 2303.055 372.395 2303.335 ;
        RECT 372.825 2303.055 373.105 2303.335 ;
        RECT 373.535 2303.055 373.815 2303.335 ;
        RECT 374.245 2303.055 374.525 2303.335 ;
        RECT 374.955 2303.055 375.235 2303.335 ;
        RECT 375.665 2303.055 375.945 2303.335 ;
        RECT 376.375 2303.055 376.655 2303.335 ;
        RECT 369.275 2302.345 369.555 2302.625 ;
        RECT 369.985 2302.345 370.265 2302.625 ;
        RECT 370.695 2302.345 370.975 2302.625 ;
        RECT 371.405 2302.345 371.685 2302.625 ;
        RECT 372.115 2302.345 372.395 2302.625 ;
        RECT 372.825 2302.345 373.105 2302.625 ;
        RECT 373.535 2302.345 373.815 2302.625 ;
        RECT 374.245 2302.345 374.525 2302.625 ;
        RECT 374.955 2302.345 375.235 2302.625 ;
        RECT 375.665 2302.345 375.945 2302.625 ;
        RECT 376.375 2302.345 376.655 2302.625 ;
        RECT 369.275 2301.635 369.555 2301.915 ;
        RECT 369.985 2301.635 370.265 2301.915 ;
        RECT 370.695 2301.635 370.975 2301.915 ;
        RECT 371.405 2301.635 371.685 2301.915 ;
        RECT 372.115 2301.635 372.395 2301.915 ;
        RECT 372.825 2301.635 373.105 2301.915 ;
        RECT 373.535 2301.635 373.815 2301.915 ;
        RECT 374.245 2301.635 374.525 2301.915 ;
        RECT 374.955 2301.635 375.235 2301.915 ;
        RECT 375.665 2301.635 375.945 2301.915 ;
        RECT 376.375 2301.635 376.655 2301.915 ;
        RECT 369.275 2300.925 369.555 2301.205 ;
        RECT 369.985 2300.925 370.265 2301.205 ;
        RECT 370.695 2300.925 370.975 2301.205 ;
        RECT 371.405 2300.925 371.685 2301.205 ;
        RECT 372.115 2300.925 372.395 2301.205 ;
        RECT 372.825 2300.925 373.105 2301.205 ;
        RECT 373.535 2300.925 373.815 2301.205 ;
        RECT 374.245 2300.925 374.525 2301.205 ;
        RECT 374.955 2300.925 375.235 2301.205 ;
        RECT 375.665 2300.925 375.945 2301.205 ;
        RECT 376.375 2300.925 376.655 2301.205 ;
        RECT 369.275 2300.215 369.555 2300.495 ;
        RECT 369.985 2300.215 370.265 2300.495 ;
        RECT 370.695 2300.215 370.975 2300.495 ;
        RECT 371.405 2300.215 371.685 2300.495 ;
        RECT 372.115 2300.215 372.395 2300.495 ;
        RECT 372.825 2300.215 373.105 2300.495 ;
        RECT 373.535 2300.215 373.815 2300.495 ;
        RECT 374.245 2300.215 374.525 2300.495 ;
        RECT 374.955 2300.215 375.235 2300.495 ;
        RECT 375.665 2300.215 375.945 2300.495 ;
        RECT 376.375 2300.215 376.655 2300.495 ;
        RECT 369.275 2299.505 369.555 2299.785 ;
        RECT 369.985 2299.505 370.265 2299.785 ;
        RECT 370.695 2299.505 370.975 2299.785 ;
        RECT 371.405 2299.505 371.685 2299.785 ;
        RECT 372.115 2299.505 372.395 2299.785 ;
        RECT 372.825 2299.505 373.105 2299.785 ;
        RECT 373.535 2299.505 373.815 2299.785 ;
        RECT 374.245 2299.505 374.525 2299.785 ;
        RECT 374.955 2299.505 375.235 2299.785 ;
        RECT 375.665 2299.505 375.945 2299.785 ;
        RECT 376.375 2299.505 376.655 2299.785 ;
        RECT 369.275 2298.795 369.555 2299.075 ;
        RECT 369.985 2298.795 370.265 2299.075 ;
        RECT 370.695 2298.795 370.975 2299.075 ;
        RECT 371.405 2298.795 371.685 2299.075 ;
        RECT 372.115 2298.795 372.395 2299.075 ;
        RECT 372.825 2298.795 373.105 2299.075 ;
        RECT 373.535 2298.795 373.815 2299.075 ;
        RECT 374.245 2298.795 374.525 2299.075 ;
        RECT 374.955 2298.795 375.235 2299.075 ;
        RECT 375.665 2298.795 375.945 2299.075 ;
        RECT 376.375 2298.795 376.655 2299.075 ;
        RECT 369.275 2298.085 369.555 2298.365 ;
        RECT 369.985 2298.085 370.265 2298.365 ;
        RECT 370.695 2298.085 370.975 2298.365 ;
        RECT 371.405 2298.085 371.685 2298.365 ;
        RECT 372.115 2298.085 372.395 2298.365 ;
        RECT 372.825 2298.085 373.105 2298.365 ;
        RECT 373.535 2298.085 373.815 2298.365 ;
        RECT 374.245 2298.085 374.525 2298.365 ;
        RECT 374.955 2298.085 375.235 2298.365 ;
        RECT 375.665 2298.085 375.945 2298.365 ;
        RECT 376.375 2298.085 376.655 2298.365 ;
        RECT 369.275 2297.375 369.555 2297.655 ;
        RECT 369.985 2297.375 370.265 2297.655 ;
        RECT 370.695 2297.375 370.975 2297.655 ;
        RECT 371.405 2297.375 371.685 2297.655 ;
        RECT 372.115 2297.375 372.395 2297.655 ;
        RECT 372.825 2297.375 373.105 2297.655 ;
        RECT 373.535 2297.375 373.815 2297.655 ;
        RECT 374.245 2297.375 374.525 2297.655 ;
        RECT 374.955 2297.375 375.235 2297.655 ;
        RECT 375.665 2297.375 375.945 2297.655 ;
        RECT 376.375 2297.375 376.655 2297.655 ;
        RECT 369.275 2296.665 369.555 2296.945 ;
        RECT 369.985 2296.665 370.265 2296.945 ;
        RECT 370.695 2296.665 370.975 2296.945 ;
        RECT 371.405 2296.665 371.685 2296.945 ;
        RECT 372.115 2296.665 372.395 2296.945 ;
        RECT 372.825 2296.665 373.105 2296.945 ;
        RECT 373.535 2296.665 373.815 2296.945 ;
        RECT 374.245 2296.665 374.525 2296.945 ;
        RECT 374.955 2296.665 375.235 2296.945 ;
        RECT 375.665 2296.665 375.945 2296.945 ;
        RECT 376.375 2296.665 376.655 2296.945 ;
        RECT 369.275 2295.955 369.555 2296.235 ;
        RECT 369.985 2295.955 370.265 2296.235 ;
        RECT 370.695 2295.955 370.975 2296.235 ;
        RECT 371.405 2295.955 371.685 2296.235 ;
        RECT 372.115 2295.955 372.395 2296.235 ;
        RECT 372.825 2295.955 373.105 2296.235 ;
        RECT 373.535 2295.955 373.815 2296.235 ;
        RECT 374.245 2295.955 374.525 2296.235 ;
        RECT 374.955 2295.955 375.235 2296.235 ;
        RECT 375.665 2295.955 375.945 2296.235 ;
        RECT 376.375 2295.955 376.655 2296.235 ;
        RECT 369.275 2293.335 369.555 2293.615 ;
        RECT 369.985 2293.335 370.265 2293.615 ;
        RECT 370.695 2293.335 370.975 2293.615 ;
        RECT 371.405 2293.335 371.685 2293.615 ;
        RECT 372.115 2293.335 372.395 2293.615 ;
        RECT 372.825 2293.335 373.105 2293.615 ;
        RECT 373.535 2293.335 373.815 2293.615 ;
        RECT 374.245 2293.335 374.525 2293.615 ;
        RECT 374.955 2293.335 375.235 2293.615 ;
        RECT 375.665 2293.335 375.945 2293.615 ;
        RECT 376.375 2293.335 376.655 2293.615 ;
        RECT 369.275 2292.625 369.555 2292.905 ;
        RECT 369.985 2292.625 370.265 2292.905 ;
        RECT 370.695 2292.625 370.975 2292.905 ;
        RECT 371.405 2292.625 371.685 2292.905 ;
        RECT 372.115 2292.625 372.395 2292.905 ;
        RECT 372.825 2292.625 373.105 2292.905 ;
        RECT 373.535 2292.625 373.815 2292.905 ;
        RECT 374.245 2292.625 374.525 2292.905 ;
        RECT 374.955 2292.625 375.235 2292.905 ;
        RECT 375.665 2292.625 375.945 2292.905 ;
        RECT 376.375 2292.625 376.655 2292.905 ;
        RECT 369.275 2291.915 369.555 2292.195 ;
        RECT 369.985 2291.915 370.265 2292.195 ;
        RECT 370.695 2291.915 370.975 2292.195 ;
        RECT 371.405 2291.915 371.685 2292.195 ;
        RECT 372.115 2291.915 372.395 2292.195 ;
        RECT 372.825 2291.915 373.105 2292.195 ;
        RECT 373.535 2291.915 373.815 2292.195 ;
        RECT 374.245 2291.915 374.525 2292.195 ;
        RECT 374.955 2291.915 375.235 2292.195 ;
        RECT 375.665 2291.915 375.945 2292.195 ;
        RECT 376.375 2291.915 376.655 2292.195 ;
        RECT 369.275 2291.205 369.555 2291.485 ;
        RECT 369.985 2291.205 370.265 2291.485 ;
        RECT 370.695 2291.205 370.975 2291.485 ;
        RECT 371.405 2291.205 371.685 2291.485 ;
        RECT 372.115 2291.205 372.395 2291.485 ;
        RECT 372.825 2291.205 373.105 2291.485 ;
        RECT 373.535 2291.205 373.815 2291.485 ;
        RECT 374.245 2291.205 374.525 2291.485 ;
        RECT 374.955 2291.205 375.235 2291.485 ;
        RECT 375.665 2291.205 375.945 2291.485 ;
        RECT 376.375 2291.205 376.655 2291.485 ;
        RECT 369.275 2290.495 369.555 2290.775 ;
        RECT 369.985 2290.495 370.265 2290.775 ;
        RECT 370.695 2290.495 370.975 2290.775 ;
        RECT 371.405 2290.495 371.685 2290.775 ;
        RECT 372.115 2290.495 372.395 2290.775 ;
        RECT 372.825 2290.495 373.105 2290.775 ;
        RECT 373.535 2290.495 373.815 2290.775 ;
        RECT 374.245 2290.495 374.525 2290.775 ;
        RECT 374.955 2290.495 375.235 2290.775 ;
        RECT 375.665 2290.495 375.945 2290.775 ;
        RECT 376.375 2290.495 376.655 2290.775 ;
        RECT 369.275 2289.785 369.555 2290.065 ;
        RECT 369.985 2289.785 370.265 2290.065 ;
        RECT 370.695 2289.785 370.975 2290.065 ;
        RECT 371.405 2289.785 371.685 2290.065 ;
        RECT 372.115 2289.785 372.395 2290.065 ;
        RECT 372.825 2289.785 373.105 2290.065 ;
        RECT 373.535 2289.785 373.815 2290.065 ;
        RECT 374.245 2289.785 374.525 2290.065 ;
        RECT 374.955 2289.785 375.235 2290.065 ;
        RECT 375.665 2289.785 375.945 2290.065 ;
        RECT 376.375 2289.785 376.655 2290.065 ;
        RECT 369.275 2289.075 369.555 2289.355 ;
        RECT 369.985 2289.075 370.265 2289.355 ;
        RECT 370.695 2289.075 370.975 2289.355 ;
        RECT 371.405 2289.075 371.685 2289.355 ;
        RECT 372.115 2289.075 372.395 2289.355 ;
        RECT 372.825 2289.075 373.105 2289.355 ;
        RECT 373.535 2289.075 373.815 2289.355 ;
        RECT 374.245 2289.075 374.525 2289.355 ;
        RECT 374.955 2289.075 375.235 2289.355 ;
        RECT 375.665 2289.075 375.945 2289.355 ;
        RECT 376.375 2289.075 376.655 2289.355 ;
        RECT 369.275 2288.365 369.555 2288.645 ;
        RECT 369.985 2288.365 370.265 2288.645 ;
        RECT 370.695 2288.365 370.975 2288.645 ;
        RECT 371.405 2288.365 371.685 2288.645 ;
        RECT 372.115 2288.365 372.395 2288.645 ;
        RECT 372.825 2288.365 373.105 2288.645 ;
        RECT 373.535 2288.365 373.815 2288.645 ;
        RECT 374.245 2288.365 374.525 2288.645 ;
        RECT 374.955 2288.365 375.235 2288.645 ;
        RECT 375.665 2288.365 375.945 2288.645 ;
        RECT 376.375 2288.365 376.655 2288.645 ;
        RECT 369.275 2287.655 369.555 2287.935 ;
        RECT 369.985 2287.655 370.265 2287.935 ;
        RECT 370.695 2287.655 370.975 2287.935 ;
        RECT 371.405 2287.655 371.685 2287.935 ;
        RECT 372.115 2287.655 372.395 2287.935 ;
        RECT 372.825 2287.655 373.105 2287.935 ;
        RECT 373.535 2287.655 373.815 2287.935 ;
        RECT 374.245 2287.655 374.525 2287.935 ;
        RECT 374.955 2287.655 375.235 2287.935 ;
        RECT 375.665 2287.655 375.945 2287.935 ;
        RECT 376.375 2287.655 376.655 2287.935 ;
        RECT 369.275 2286.945 369.555 2287.225 ;
        RECT 369.985 2286.945 370.265 2287.225 ;
        RECT 370.695 2286.945 370.975 2287.225 ;
        RECT 371.405 2286.945 371.685 2287.225 ;
        RECT 372.115 2286.945 372.395 2287.225 ;
        RECT 372.825 2286.945 373.105 2287.225 ;
        RECT 373.535 2286.945 373.815 2287.225 ;
        RECT 374.245 2286.945 374.525 2287.225 ;
        RECT 374.955 2286.945 375.235 2287.225 ;
        RECT 375.665 2286.945 375.945 2287.225 ;
        RECT 376.375 2286.945 376.655 2287.225 ;
        RECT 369.275 2286.235 369.555 2286.515 ;
        RECT 369.985 2286.235 370.265 2286.515 ;
        RECT 370.695 2286.235 370.975 2286.515 ;
        RECT 371.405 2286.235 371.685 2286.515 ;
        RECT 372.115 2286.235 372.395 2286.515 ;
        RECT 372.825 2286.235 373.105 2286.515 ;
        RECT 373.535 2286.235 373.815 2286.515 ;
        RECT 374.245 2286.235 374.525 2286.515 ;
        RECT 374.955 2286.235 375.235 2286.515 ;
        RECT 375.665 2286.235 375.945 2286.515 ;
        RECT 376.375 2286.235 376.655 2286.515 ;
        RECT 369.275 2285.525 369.555 2285.805 ;
        RECT 369.985 2285.525 370.265 2285.805 ;
        RECT 370.695 2285.525 370.975 2285.805 ;
        RECT 371.405 2285.525 371.685 2285.805 ;
        RECT 372.115 2285.525 372.395 2285.805 ;
        RECT 372.825 2285.525 373.105 2285.805 ;
        RECT 373.535 2285.525 373.815 2285.805 ;
        RECT 374.245 2285.525 374.525 2285.805 ;
        RECT 374.955 2285.525 375.235 2285.805 ;
        RECT 375.665 2285.525 375.945 2285.805 ;
        RECT 376.375 2285.525 376.655 2285.805 ;
        RECT 369.275 2284.815 369.555 2285.095 ;
        RECT 369.985 2284.815 370.265 2285.095 ;
        RECT 370.695 2284.815 370.975 2285.095 ;
        RECT 371.405 2284.815 371.685 2285.095 ;
        RECT 372.115 2284.815 372.395 2285.095 ;
        RECT 372.825 2284.815 373.105 2285.095 ;
        RECT 373.535 2284.815 373.815 2285.095 ;
        RECT 374.245 2284.815 374.525 2285.095 ;
        RECT 374.955 2284.815 375.235 2285.095 ;
        RECT 375.665 2284.815 375.945 2285.095 ;
        RECT 376.375 2284.815 376.655 2285.095 ;
        RECT 369.275 2284.105 369.555 2284.385 ;
        RECT 369.985 2284.105 370.265 2284.385 ;
        RECT 370.695 2284.105 370.975 2284.385 ;
        RECT 371.405 2284.105 371.685 2284.385 ;
        RECT 372.115 2284.105 372.395 2284.385 ;
        RECT 372.825 2284.105 373.105 2284.385 ;
        RECT 373.535 2284.105 373.815 2284.385 ;
        RECT 374.245 2284.105 374.525 2284.385 ;
        RECT 374.955 2284.105 375.235 2284.385 ;
        RECT 375.665 2284.105 375.945 2284.385 ;
        RECT 376.375 2284.105 376.655 2284.385 ;
        RECT 369.330 2280.190 369.610 2280.470 ;
        RECT 370.040 2280.190 370.320 2280.470 ;
        RECT 370.750 2280.190 371.030 2280.470 ;
        RECT 371.460 2280.190 371.740 2280.470 ;
        RECT 372.170 2280.190 372.450 2280.470 ;
        RECT 372.880 2280.190 373.160 2280.470 ;
        RECT 373.590 2280.190 373.870 2280.470 ;
        RECT 374.300 2280.190 374.580 2280.470 ;
        RECT 375.010 2280.190 375.290 2280.470 ;
        RECT 375.720 2280.190 376.000 2280.470 ;
        RECT 376.430 2280.190 376.710 2280.470 ;
        RECT 369.330 2279.480 369.610 2279.760 ;
        RECT 370.040 2279.480 370.320 2279.760 ;
        RECT 370.750 2279.480 371.030 2279.760 ;
        RECT 371.460 2279.480 371.740 2279.760 ;
        RECT 372.170 2279.480 372.450 2279.760 ;
        RECT 372.880 2279.480 373.160 2279.760 ;
        RECT 373.590 2279.480 373.870 2279.760 ;
        RECT 374.300 2279.480 374.580 2279.760 ;
        RECT 375.010 2279.480 375.290 2279.760 ;
        RECT 375.720 2279.480 376.000 2279.760 ;
        RECT 376.430 2279.480 376.710 2279.760 ;
        RECT 369.330 2278.770 369.610 2279.050 ;
        RECT 370.040 2278.770 370.320 2279.050 ;
        RECT 370.750 2278.770 371.030 2279.050 ;
        RECT 371.460 2278.770 371.740 2279.050 ;
        RECT 372.170 2278.770 372.450 2279.050 ;
        RECT 372.880 2278.770 373.160 2279.050 ;
        RECT 373.590 2278.770 373.870 2279.050 ;
        RECT 374.300 2278.770 374.580 2279.050 ;
        RECT 375.010 2278.770 375.290 2279.050 ;
        RECT 375.720 2278.770 376.000 2279.050 ;
        RECT 376.430 2278.770 376.710 2279.050 ;
        RECT 369.330 2278.060 369.610 2278.340 ;
        RECT 370.040 2278.060 370.320 2278.340 ;
        RECT 370.750 2278.060 371.030 2278.340 ;
        RECT 371.460 2278.060 371.740 2278.340 ;
        RECT 372.170 2278.060 372.450 2278.340 ;
        RECT 372.880 2278.060 373.160 2278.340 ;
        RECT 373.590 2278.060 373.870 2278.340 ;
        RECT 374.300 2278.060 374.580 2278.340 ;
        RECT 375.010 2278.060 375.290 2278.340 ;
        RECT 375.720 2278.060 376.000 2278.340 ;
        RECT 376.430 2278.060 376.710 2278.340 ;
        RECT 369.330 2277.350 369.610 2277.630 ;
        RECT 370.040 2277.350 370.320 2277.630 ;
        RECT 370.750 2277.350 371.030 2277.630 ;
        RECT 371.460 2277.350 371.740 2277.630 ;
        RECT 372.170 2277.350 372.450 2277.630 ;
        RECT 372.880 2277.350 373.160 2277.630 ;
        RECT 373.590 2277.350 373.870 2277.630 ;
        RECT 374.300 2277.350 374.580 2277.630 ;
        RECT 375.010 2277.350 375.290 2277.630 ;
        RECT 375.720 2277.350 376.000 2277.630 ;
        RECT 376.430 2277.350 376.710 2277.630 ;
        RECT 369.330 2276.640 369.610 2276.920 ;
        RECT 370.040 2276.640 370.320 2276.920 ;
        RECT 370.750 2276.640 371.030 2276.920 ;
        RECT 371.460 2276.640 371.740 2276.920 ;
        RECT 372.170 2276.640 372.450 2276.920 ;
        RECT 372.880 2276.640 373.160 2276.920 ;
        RECT 373.590 2276.640 373.870 2276.920 ;
        RECT 374.300 2276.640 374.580 2276.920 ;
        RECT 375.010 2276.640 375.290 2276.920 ;
        RECT 375.720 2276.640 376.000 2276.920 ;
        RECT 376.430 2276.640 376.710 2276.920 ;
        RECT 369.330 2275.930 369.610 2276.210 ;
        RECT 370.040 2275.930 370.320 2276.210 ;
        RECT 370.750 2275.930 371.030 2276.210 ;
        RECT 371.460 2275.930 371.740 2276.210 ;
        RECT 372.170 2275.930 372.450 2276.210 ;
        RECT 372.880 2275.930 373.160 2276.210 ;
        RECT 373.590 2275.930 373.870 2276.210 ;
        RECT 374.300 2275.930 374.580 2276.210 ;
        RECT 375.010 2275.930 375.290 2276.210 ;
        RECT 375.720 2275.930 376.000 2276.210 ;
        RECT 376.430 2275.930 376.710 2276.210 ;
        RECT 369.330 2275.220 369.610 2275.500 ;
        RECT 370.040 2275.220 370.320 2275.500 ;
        RECT 370.750 2275.220 371.030 2275.500 ;
        RECT 371.460 2275.220 371.740 2275.500 ;
        RECT 372.170 2275.220 372.450 2275.500 ;
        RECT 372.880 2275.220 373.160 2275.500 ;
        RECT 373.590 2275.220 373.870 2275.500 ;
        RECT 374.300 2275.220 374.580 2275.500 ;
        RECT 375.010 2275.220 375.290 2275.500 ;
        RECT 375.720 2275.220 376.000 2275.500 ;
        RECT 376.430 2275.220 376.710 2275.500 ;
        RECT 369.330 2274.510 369.610 2274.790 ;
        RECT 370.040 2274.510 370.320 2274.790 ;
        RECT 370.750 2274.510 371.030 2274.790 ;
        RECT 371.460 2274.510 371.740 2274.790 ;
        RECT 372.170 2274.510 372.450 2274.790 ;
        RECT 372.880 2274.510 373.160 2274.790 ;
        RECT 373.590 2274.510 373.870 2274.790 ;
        RECT 374.300 2274.510 374.580 2274.790 ;
        RECT 375.010 2274.510 375.290 2274.790 ;
        RECT 375.720 2274.510 376.000 2274.790 ;
        RECT 376.430 2274.510 376.710 2274.790 ;
        RECT 369.330 2273.800 369.610 2274.080 ;
        RECT 370.040 2273.800 370.320 2274.080 ;
        RECT 370.750 2273.800 371.030 2274.080 ;
        RECT 371.460 2273.800 371.740 2274.080 ;
        RECT 372.170 2273.800 372.450 2274.080 ;
        RECT 372.880 2273.800 373.160 2274.080 ;
        RECT 373.590 2273.800 373.870 2274.080 ;
        RECT 374.300 2273.800 374.580 2274.080 ;
        RECT 375.010 2273.800 375.290 2274.080 ;
        RECT 375.720 2273.800 376.000 2274.080 ;
        RECT 376.430 2273.800 376.710 2274.080 ;
        RECT 369.330 2273.090 369.610 2273.370 ;
        RECT 370.040 2273.090 370.320 2273.370 ;
        RECT 370.750 2273.090 371.030 2273.370 ;
        RECT 371.460 2273.090 371.740 2273.370 ;
        RECT 372.170 2273.090 372.450 2273.370 ;
        RECT 372.880 2273.090 373.160 2273.370 ;
        RECT 373.590 2273.090 373.870 2273.370 ;
        RECT 374.300 2273.090 374.580 2273.370 ;
        RECT 375.010 2273.090 375.290 2273.370 ;
        RECT 375.720 2273.090 376.000 2273.370 ;
        RECT 376.430 2273.090 376.710 2273.370 ;
        RECT 369.330 2272.380 369.610 2272.660 ;
        RECT 370.040 2272.380 370.320 2272.660 ;
        RECT 370.750 2272.380 371.030 2272.660 ;
        RECT 371.460 2272.380 371.740 2272.660 ;
        RECT 372.170 2272.380 372.450 2272.660 ;
        RECT 372.880 2272.380 373.160 2272.660 ;
        RECT 373.590 2272.380 373.870 2272.660 ;
        RECT 374.300 2272.380 374.580 2272.660 ;
        RECT 375.010 2272.380 375.290 2272.660 ;
        RECT 375.720 2272.380 376.000 2272.660 ;
        RECT 376.430 2272.380 376.710 2272.660 ;
        RECT 369.330 2271.670 369.610 2271.950 ;
        RECT 370.040 2271.670 370.320 2271.950 ;
        RECT 370.750 2271.670 371.030 2271.950 ;
        RECT 371.460 2271.670 371.740 2271.950 ;
        RECT 372.170 2271.670 372.450 2271.950 ;
        RECT 372.880 2271.670 373.160 2271.950 ;
        RECT 373.590 2271.670 373.870 2271.950 ;
        RECT 374.300 2271.670 374.580 2271.950 ;
        RECT 375.010 2271.670 375.290 2271.950 ;
        RECT 375.720 2271.670 376.000 2271.950 ;
        RECT 376.430 2271.670 376.710 2271.950 ;
        RECT 3512.200 2238.050 3512.480 2238.330 ;
        RECT 3512.910 2238.050 3513.190 2238.330 ;
        RECT 3513.620 2238.050 3513.900 2238.330 ;
        RECT 3514.330 2238.050 3514.610 2238.330 ;
        RECT 3515.040 2238.050 3515.320 2238.330 ;
        RECT 3515.750 2238.050 3516.030 2238.330 ;
        RECT 3516.460 2238.050 3516.740 2238.330 ;
        RECT 3517.170 2238.050 3517.450 2238.330 ;
        RECT 3517.880 2238.050 3518.160 2238.330 ;
        RECT 3518.590 2238.050 3518.870 2238.330 ;
        RECT 3519.300 2238.050 3519.580 2238.330 ;
        RECT 3520.010 2238.050 3520.290 2238.330 ;
        RECT 3520.720 2238.050 3521.000 2238.330 ;
        RECT 3521.430 2238.050 3521.710 2238.330 ;
        RECT 3512.200 2237.340 3512.480 2237.620 ;
        RECT 3512.910 2237.340 3513.190 2237.620 ;
        RECT 3513.620 2237.340 3513.900 2237.620 ;
        RECT 3514.330 2237.340 3514.610 2237.620 ;
        RECT 3515.040 2237.340 3515.320 2237.620 ;
        RECT 3515.750 2237.340 3516.030 2237.620 ;
        RECT 3516.460 2237.340 3516.740 2237.620 ;
        RECT 3517.170 2237.340 3517.450 2237.620 ;
        RECT 3517.880 2237.340 3518.160 2237.620 ;
        RECT 3518.590 2237.340 3518.870 2237.620 ;
        RECT 3519.300 2237.340 3519.580 2237.620 ;
        RECT 3520.010 2237.340 3520.290 2237.620 ;
        RECT 3520.720 2237.340 3521.000 2237.620 ;
        RECT 3521.430 2237.340 3521.710 2237.620 ;
        RECT 3512.200 2236.630 3512.480 2236.910 ;
        RECT 3512.910 2236.630 3513.190 2236.910 ;
        RECT 3513.620 2236.630 3513.900 2236.910 ;
        RECT 3514.330 2236.630 3514.610 2236.910 ;
        RECT 3515.040 2236.630 3515.320 2236.910 ;
        RECT 3515.750 2236.630 3516.030 2236.910 ;
        RECT 3516.460 2236.630 3516.740 2236.910 ;
        RECT 3517.170 2236.630 3517.450 2236.910 ;
        RECT 3517.880 2236.630 3518.160 2236.910 ;
        RECT 3518.590 2236.630 3518.870 2236.910 ;
        RECT 3519.300 2236.630 3519.580 2236.910 ;
        RECT 3520.010 2236.630 3520.290 2236.910 ;
        RECT 3520.720 2236.630 3521.000 2236.910 ;
        RECT 3521.430 2236.630 3521.710 2236.910 ;
        RECT 3512.200 2235.920 3512.480 2236.200 ;
        RECT 3512.910 2235.920 3513.190 2236.200 ;
        RECT 3513.620 2235.920 3513.900 2236.200 ;
        RECT 3514.330 2235.920 3514.610 2236.200 ;
        RECT 3515.040 2235.920 3515.320 2236.200 ;
        RECT 3515.750 2235.920 3516.030 2236.200 ;
        RECT 3516.460 2235.920 3516.740 2236.200 ;
        RECT 3517.170 2235.920 3517.450 2236.200 ;
        RECT 3517.880 2235.920 3518.160 2236.200 ;
        RECT 3518.590 2235.920 3518.870 2236.200 ;
        RECT 3519.300 2235.920 3519.580 2236.200 ;
        RECT 3520.010 2235.920 3520.290 2236.200 ;
        RECT 3520.720 2235.920 3521.000 2236.200 ;
        RECT 3521.430 2235.920 3521.710 2236.200 ;
        RECT 3512.200 2235.210 3512.480 2235.490 ;
        RECT 3512.910 2235.210 3513.190 2235.490 ;
        RECT 3513.620 2235.210 3513.900 2235.490 ;
        RECT 3514.330 2235.210 3514.610 2235.490 ;
        RECT 3515.040 2235.210 3515.320 2235.490 ;
        RECT 3515.750 2235.210 3516.030 2235.490 ;
        RECT 3516.460 2235.210 3516.740 2235.490 ;
        RECT 3517.170 2235.210 3517.450 2235.490 ;
        RECT 3517.880 2235.210 3518.160 2235.490 ;
        RECT 3518.590 2235.210 3518.870 2235.490 ;
        RECT 3519.300 2235.210 3519.580 2235.490 ;
        RECT 3520.010 2235.210 3520.290 2235.490 ;
        RECT 3520.720 2235.210 3521.000 2235.490 ;
        RECT 3521.430 2235.210 3521.710 2235.490 ;
        RECT 3512.200 2234.500 3512.480 2234.780 ;
        RECT 3512.910 2234.500 3513.190 2234.780 ;
        RECT 3513.620 2234.500 3513.900 2234.780 ;
        RECT 3514.330 2234.500 3514.610 2234.780 ;
        RECT 3515.040 2234.500 3515.320 2234.780 ;
        RECT 3515.750 2234.500 3516.030 2234.780 ;
        RECT 3516.460 2234.500 3516.740 2234.780 ;
        RECT 3517.170 2234.500 3517.450 2234.780 ;
        RECT 3517.880 2234.500 3518.160 2234.780 ;
        RECT 3518.590 2234.500 3518.870 2234.780 ;
        RECT 3519.300 2234.500 3519.580 2234.780 ;
        RECT 3520.010 2234.500 3520.290 2234.780 ;
        RECT 3520.720 2234.500 3521.000 2234.780 ;
        RECT 3521.430 2234.500 3521.710 2234.780 ;
        RECT 3512.200 2233.790 3512.480 2234.070 ;
        RECT 3512.910 2233.790 3513.190 2234.070 ;
        RECT 3513.620 2233.790 3513.900 2234.070 ;
        RECT 3514.330 2233.790 3514.610 2234.070 ;
        RECT 3515.040 2233.790 3515.320 2234.070 ;
        RECT 3515.750 2233.790 3516.030 2234.070 ;
        RECT 3516.460 2233.790 3516.740 2234.070 ;
        RECT 3517.170 2233.790 3517.450 2234.070 ;
        RECT 3517.880 2233.790 3518.160 2234.070 ;
        RECT 3518.590 2233.790 3518.870 2234.070 ;
        RECT 3519.300 2233.790 3519.580 2234.070 ;
        RECT 3520.010 2233.790 3520.290 2234.070 ;
        RECT 3520.720 2233.790 3521.000 2234.070 ;
        RECT 3521.430 2233.790 3521.710 2234.070 ;
        RECT 3512.200 2233.080 3512.480 2233.360 ;
        RECT 3512.910 2233.080 3513.190 2233.360 ;
        RECT 3513.620 2233.080 3513.900 2233.360 ;
        RECT 3514.330 2233.080 3514.610 2233.360 ;
        RECT 3515.040 2233.080 3515.320 2233.360 ;
        RECT 3515.750 2233.080 3516.030 2233.360 ;
        RECT 3516.460 2233.080 3516.740 2233.360 ;
        RECT 3517.170 2233.080 3517.450 2233.360 ;
        RECT 3517.880 2233.080 3518.160 2233.360 ;
        RECT 3518.590 2233.080 3518.870 2233.360 ;
        RECT 3519.300 2233.080 3519.580 2233.360 ;
        RECT 3520.010 2233.080 3520.290 2233.360 ;
        RECT 3520.720 2233.080 3521.000 2233.360 ;
        RECT 3521.430 2233.080 3521.710 2233.360 ;
        RECT 3512.200 2232.370 3512.480 2232.650 ;
        RECT 3512.910 2232.370 3513.190 2232.650 ;
        RECT 3513.620 2232.370 3513.900 2232.650 ;
        RECT 3514.330 2232.370 3514.610 2232.650 ;
        RECT 3515.040 2232.370 3515.320 2232.650 ;
        RECT 3515.750 2232.370 3516.030 2232.650 ;
        RECT 3516.460 2232.370 3516.740 2232.650 ;
        RECT 3517.170 2232.370 3517.450 2232.650 ;
        RECT 3517.880 2232.370 3518.160 2232.650 ;
        RECT 3518.590 2232.370 3518.870 2232.650 ;
        RECT 3519.300 2232.370 3519.580 2232.650 ;
        RECT 3520.010 2232.370 3520.290 2232.650 ;
        RECT 3520.720 2232.370 3521.000 2232.650 ;
        RECT 3521.430 2232.370 3521.710 2232.650 ;
        RECT 3512.200 2231.660 3512.480 2231.940 ;
        RECT 3512.910 2231.660 3513.190 2231.940 ;
        RECT 3513.620 2231.660 3513.900 2231.940 ;
        RECT 3514.330 2231.660 3514.610 2231.940 ;
        RECT 3515.040 2231.660 3515.320 2231.940 ;
        RECT 3515.750 2231.660 3516.030 2231.940 ;
        RECT 3516.460 2231.660 3516.740 2231.940 ;
        RECT 3517.170 2231.660 3517.450 2231.940 ;
        RECT 3517.880 2231.660 3518.160 2231.940 ;
        RECT 3518.590 2231.660 3518.870 2231.940 ;
        RECT 3519.300 2231.660 3519.580 2231.940 ;
        RECT 3520.010 2231.660 3520.290 2231.940 ;
        RECT 3520.720 2231.660 3521.000 2231.940 ;
        RECT 3521.430 2231.660 3521.710 2231.940 ;
        RECT 3512.200 2230.950 3512.480 2231.230 ;
        RECT 3512.910 2230.950 3513.190 2231.230 ;
        RECT 3513.620 2230.950 3513.900 2231.230 ;
        RECT 3514.330 2230.950 3514.610 2231.230 ;
        RECT 3515.040 2230.950 3515.320 2231.230 ;
        RECT 3515.750 2230.950 3516.030 2231.230 ;
        RECT 3516.460 2230.950 3516.740 2231.230 ;
        RECT 3517.170 2230.950 3517.450 2231.230 ;
        RECT 3517.880 2230.950 3518.160 2231.230 ;
        RECT 3518.590 2230.950 3518.870 2231.230 ;
        RECT 3519.300 2230.950 3519.580 2231.230 ;
        RECT 3520.010 2230.950 3520.290 2231.230 ;
        RECT 3520.720 2230.950 3521.000 2231.230 ;
        RECT 3521.430 2230.950 3521.710 2231.230 ;
        RECT 3512.200 2230.240 3512.480 2230.520 ;
        RECT 3512.910 2230.240 3513.190 2230.520 ;
        RECT 3513.620 2230.240 3513.900 2230.520 ;
        RECT 3514.330 2230.240 3514.610 2230.520 ;
        RECT 3515.040 2230.240 3515.320 2230.520 ;
        RECT 3515.750 2230.240 3516.030 2230.520 ;
        RECT 3516.460 2230.240 3516.740 2230.520 ;
        RECT 3517.170 2230.240 3517.450 2230.520 ;
        RECT 3517.880 2230.240 3518.160 2230.520 ;
        RECT 3518.590 2230.240 3518.870 2230.520 ;
        RECT 3519.300 2230.240 3519.580 2230.520 ;
        RECT 3520.010 2230.240 3520.290 2230.520 ;
        RECT 3520.720 2230.240 3521.000 2230.520 ;
        RECT 3521.430 2230.240 3521.710 2230.520 ;
        RECT 3512.200 2229.530 3512.480 2229.810 ;
        RECT 3512.910 2229.530 3513.190 2229.810 ;
        RECT 3513.620 2229.530 3513.900 2229.810 ;
        RECT 3514.330 2229.530 3514.610 2229.810 ;
        RECT 3515.040 2229.530 3515.320 2229.810 ;
        RECT 3515.750 2229.530 3516.030 2229.810 ;
        RECT 3516.460 2229.530 3516.740 2229.810 ;
        RECT 3517.170 2229.530 3517.450 2229.810 ;
        RECT 3517.880 2229.530 3518.160 2229.810 ;
        RECT 3518.590 2229.530 3518.870 2229.810 ;
        RECT 3519.300 2229.530 3519.580 2229.810 ;
        RECT 3520.010 2229.530 3520.290 2229.810 ;
        RECT 3520.720 2229.530 3521.000 2229.810 ;
        RECT 3521.430 2229.530 3521.710 2229.810 ;
        RECT 3512.255 2225.615 3512.535 2225.895 ;
        RECT 3512.965 2225.615 3513.245 2225.895 ;
        RECT 3513.675 2225.615 3513.955 2225.895 ;
        RECT 3514.385 2225.615 3514.665 2225.895 ;
        RECT 3515.095 2225.615 3515.375 2225.895 ;
        RECT 3515.805 2225.615 3516.085 2225.895 ;
        RECT 3516.515 2225.615 3516.795 2225.895 ;
        RECT 3517.225 2225.615 3517.505 2225.895 ;
        RECT 3517.935 2225.615 3518.215 2225.895 ;
        RECT 3518.645 2225.615 3518.925 2225.895 ;
        RECT 3519.355 2225.615 3519.635 2225.895 ;
        RECT 3520.065 2225.615 3520.345 2225.895 ;
        RECT 3520.775 2225.615 3521.055 2225.895 ;
        RECT 3521.485 2225.615 3521.765 2225.895 ;
        RECT 3512.255 2224.905 3512.535 2225.185 ;
        RECT 3512.965 2224.905 3513.245 2225.185 ;
        RECT 3513.675 2224.905 3513.955 2225.185 ;
        RECT 3514.385 2224.905 3514.665 2225.185 ;
        RECT 3515.095 2224.905 3515.375 2225.185 ;
        RECT 3515.805 2224.905 3516.085 2225.185 ;
        RECT 3516.515 2224.905 3516.795 2225.185 ;
        RECT 3517.225 2224.905 3517.505 2225.185 ;
        RECT 3517.935 2224.905 3518.215 2225.185 ;
        RECT 3518.645 2224.905 3518.925 2225.185 ;
        RECT 3519.355 2224.905 3519.635 2225.185 ;
        RECT 3520.065 2224.905 3520.345 2225.185 ;
        RECT 3520.775 2224.905 3521.055 2225.185 ;
        RECT 3521.485 2224.905 3521.765 2225.185 ;
        RECT 3512.255 2224.195 3512.535 2224.475 ;
        RECT 3512.965 2224.195 3513.245 2224.475 ;
        RECT 3513.675 2224.195 3513.955 2224.475 ;
        RECT 3514.385 2224.195 3514.665 2224.475 ;
        RECT 3515.095 2224.195 3515.375 2224.475 ;
        RECT 3515.805 2224.195 3516.085 2224.475 ;
        RECT 3516.515 2224.195 3516.795 2224.475 ;
        RECT 3517.225 2224.195 3517.505 2224.475 ;
        RECT 3517.935 2224.195 3518.215 2224.475 ;
        RECT 3518.645 2224.195 3518.925 2224.475 ;
        RECT 3519.355 2224.195 3519.635 2224.475 ;
        RECT 3520.065 2224.195 3520.345 2224.475 ;
        RECT 3520.775 2224.195 3521.055 2224.475 ;
        RECT 3521.485 2224.195 3521.765 2224.475 ;
        RECT 3512.255 2223.485 3512.535 2223.765 ;
        RECT 3512.965 2223.485 3513.245 2223.765 ;
        RECT 3513.675 2223.485 3513.955 2223.765 ;
        RECT 3514.385 2223.485 3514.665 2223.765 ;
        RECT 3515.095 2223.485 3515.375 2223.765 ;
        RECT 3515.805 2223.485 3516.085 2223.765 ;
        RECT 3516.515 2223.485 3516.795 2223.765 ;
        RECT 3517.225 2223.485 3517.505 2223.765 ;
        RECT 3517.935 2223.485 3518.215 2223.765 ;
        RECT 3518.645 2223.485 3518.925 2223.765 ;
        RECT 3519.355 2223.485 3519.635 2223.765 ;
        RECT 3520.065 2223.485 3520.345 2223.765 ;
        RECT 3520.775 2223.485 3521.055 2223.765 ;
        RECT 3521.485 2223.485 3521.765 2223.765 ;
        RECT 3512.255 2222.775 3512.535 2223.055 ;
        RECT 3512.965 2222.775 3513.245 2223.055 ;
        RECT 3513.675 2222.775 3513.955 2223.055 ;
        RECT 3514.385 2222.775 3514.665 2223.055 ;
        RECT 3515.095 2222.775 3515.375 2223.055 ;
        RECT 3515.805 2222.775 3516.085 2223.055 ;
        RECT 3516.515 2222.775 3516.795 2223.055 ;
        RECT 3517.225 2222.775 3517.505 2223.055 ;
        RECT 3517.935 2222.775 3518.215 2223.055 ;
        RECT 3518.645 2222.775 3518.925 2223.055 ;
        RECT 3519.355 2222.775 3519.635 2223.055 ;
        RECT 3520.065 2222.775 3520.345 2223.055 ;
        RECT 3520.775 2222.775 3521.055 2223.055 ;
        RECT 3521.485 2222.775 3521.765 2223.055 ;
        RECT 3512.255 2222.065 3512.535 2222.345 ;
        RECT 3512.965 2222.065 3513.245 2222.345 ;
        RECT 3513.675 2222.065 3513.955 2222.345 ;
        RECT 3514.385 2222.065 3514.665 2222.345 ;
        RECT 3515.095 2222.065 3515.375 2222.345 ;
        RECT 3515.805 2222.065 3516.085 2222.345 ;
        RECT 3516.515 2222.065 3516.795 2222.345 ;
        RECT 3517.225 2222.065 3517.505 2222.345 ;
        RECT 3517.935 2222.065 3518.215 2222.345 ;
        RECT 3518.645 2222.065 3518.925 2222.345 ;
        RECT 3519.355 2222.065 3519.635 2222.345 ;
        RECT 3520.065 2222.065 3520.345 2222.345 ;
        RECT 3520.775 2222.065 3521.055 2222.345 ;
        RECT 3521.485 2222.065 3521.765 2222.345 ;
        RECT 3512.255 2221.355 3512.535 2221.635 ;
        RECT 3512.965 2221.355 3513.245 2221.635 ;
        RECT 3513.675 2221.355 3513.955 2221.635 ;
        RECT 3514.385 2221.355 3514.665 2221.635 ;
        RECT 3515.095 2221.355 3515.375 2221.635 ;
        RECT 3515.805 2221.355 3516.085 2221.635 ;
        RECT 3516.515 2221.355 3516.795 2221.635 ;
        RECT 3517.225 2221.355 3517.505 2221.635 ;
        RECT 3517.935 2221.355 3518.215 2221.635 ;
        RECT 3518.645 2221.355 3518.925 2221.635 ;
        RECT 3519.355 2221.355 3519.635 2221.635 ;
        RECT 3520.065 2221.355 3520.345 2221.635 ;
        RECT 3520.775 2221.355 3521.055 2221.635 ;
        RECT 3521.485 2221.355 3521.765 2221.635 ;
        RECT 3512.255 2220.645 3512.535 2220.925 ;
        RECT 3512.965 2220.645 3513.245 2220.925 ;
        RECT 3513.675 2220.645 3513.955 2220.925 ;
        RECT 3514.385 2220.645 3514.665 2220.925 ;
        RECT 3515.095 2220.645 3515.375 2220.925 ;
        RECT 3515.805 2220.645 3516.085 2220.925 ;
        RECT 3516.515 2220.645 3516.795 2220.925 ;
        RECT 3517.225 2220.645 3517.505 2220.925 ;
        RECT 3517.935 2220.645 3518.215 2220.925 ;
        RECT 3518.645 2220.645 3518.925 2220.925 ;
        RECT 3519.355 2220.645 3519.635 2220.925 ;
        RECT 3520.065 2220.645 3520.345 2220.925 ;
        RECT 3520.775 2220.645 3521.055 2220.925 ;
        RECT 3521.485 2220.645 3521.765 2220.925 ;
        RECT 3512.255 2219.935 3512.535 2220.215 ;
        RECT 3512.965 2219.935 3513.245 2220.215 ;
        RECT 3513.675 2219.935 3513.955 2220.215 ;
        RECT 3514.385 2219.935 3514.665 2220.215 ;
        RECT 3515.095 2219.935 3515.375 2220.215 ;
        RECT 3515.805 2219.935 3516.085 2220.215 ;
        RECT 3516.515 2219.935 3516.795 2220.215 ;
        RECT 3517.225 2219.935 3517.505 2220.215 ;
        RECT 3517.935 2219.935 3518.215 2220.215 ;
        RECT 3518.645 2219.935 3518.925 2220.215 ;
        RECT 3519.355 2219.935 3519.635 2220.215 ;
        RECT 3520.065 2219.935 3520.345 2220.215 ;
        RECT 3520.775 2219.935 3521.055 2220.215 ;
        RECT 3521.485 2219.935 3521.765 2220.215 ;
        RECT 3512.255 2219.225 3512.535 2219.505 ;
        RECT 3512.965 2219.225 3513.245 2219.505 ;
        RECT 3513.675 2219.225 3513.955 2219.505 ;
        RECT 3514.385 2219.225 3514.665 2219.505 ;
        RECT 3515.095 2219.225 3515.375 2219.505 ;
        RECT 3515.805 2219.225 3516.085 2219.505 ;
        RECT 3516.515 2219.225 3516.795 2219.505 ;
        RECT 3517.225 2219.225 3517.505 2219.505 ;
        RECT 3517.935 2219.225 3518.215 2219.505 ;
        RECT 3518.645 2219.225 3518.925 2219.505 ;
        RECT 3519.355 2219.225 3519.635 2219.505 ;
        RECT 3520.065 2219.225 3520.345 2219.505 ;
        RECT 3520.775 2219.225 3521.055 2219.505 ;
        RECT 3521.485 2219.225 3521.765 2219.505 ;
        RECT 3512.255 2218.515 3512.535 2218.795 ;
        RECT 3512.965 2218.515 3513.245 2218.795 ;
        RECT 3513.675 2218.515 3513.955 2218.795 ;
        RECT 3514.385 2218.515 3514.665 2218.795 ;
        RECT 3515.095 2218.515 3515.375 2218.795 ;
        RECT 3515.805 2218.515 3516.085 2218.795 ;
        RECT 3516.515 2218.515 3516.795 2218.795 ;
        RECT 3517.225 2218.515 3517.505 2218.795 ;
        RECT 3517.935 2218.515 3518.215 2218.795 ;
        RECT 3518.645 2218.515 3518.925 2218.795 ;
        RECT 3519.355 2218.515 3519.635 2218.795 ;
        RECT 3520.065 2218.515 3520.345 2218.795 ;
        RECT 3520.775 2218.515 3521.055 2218.795 ;
        RECT 3521.485 2218.515 3521.765 2218.795 ;
        RECT 3512.255 2217.805 3512.535 2218.085 ;
        RECT 3512.965 2217.805 3513.245 2218.085 ;
        RECT 3513.675 2217.805 3513.955 2218.085 ;
        RECT 3514.385 2217.805 3514.665 2218.085 ;
        RECT 3515.095 2217.805 3515.375 2218.085 ;
        RECT 3515.805 2217.805 3516.085 2218.085 ;
        RECT 3516.515 2217.805 3516.795 2218.085 ;
        RECT 3517.225 2217.805 3517.505 2218.085 ;
        RECT 3517.935 2217.805 3518.215 2218.085 ;
        RECT 3518.645 2217.805 3518.925 2218.085 ;
        RECT 3519.355 2217.805 3519.635 2218.085 ;
        RECT 3520.065 2217.805 3520.345 2218.085 ;
        RECT 3520.775 2217.805 3521.055 2218.085 ;
        RECT 3521.485 2217.805 3521.765 2218.085 ;
        RECT 3512.255 2217.095 3512.535 2217.375 ;
        RECT 3512.965 2217.095 3513.245 2217.375 ;
        RECT 3513.675 2217.095 3513.955 2217.375 ;
        RECT 3514.385 2217.095 3514.665 2217.375 ;
        RECT 3515.095 2217.095 3515.375 2217.375 ;
        RECT 3515.805 2217.095 3516.085 2217.375 ;
        RECT 3516.515 2217.095 3516.795 2217.375 ;
        RECT 3517.225 2217.095 3517.505 2217.375 ;
        RECT 3517.935 2217.095 3518.215 2217.375 ;
        RECT 3518.645 2217.095 3518.925 2217.375 ;
        RECT 3519.355 2217.095 3519.635 2217.375 ;
        RECT 3520.065 2217.095 3520.345 2217.375 ;
        RECT 3520.775 2217.095 3521.055 2217.375 ;
        RECT 3521.485 2217.095 3521.765 2217.375 ;
        RECT 3512.255 2216.385 3512.535 2216.665 ;
        RECT 3512.965 2216.385 3513.245 2216.665 ;
        RECT 3513.675 2216.385 3513.955 2216.665 ;
        RECT 3514.385 2216.385 3514.665 2216.665 ;
        RECT 3515.095 2216.385 3515.375 2216.665 ;
        RECT 3515.805 2216.385 3516.085 2216.665 ;
        RECT 3516.515 2216.385 3516.795 2216.665 ;
        RECT 3517.225 2216.385 3517.505 2216.665 ;
        RECT 3517.935 2216.385 3518.215 2216.665 ;
        RECT 3518.645 2216.385 3518.925 2216.665 ;
        RECT 3519.355 2216.385 3519.635 2216.665 ;
        RECT 3520.065 2216.385 3520.345 2216.665 ;
        RECT 3520.775 2216.385 3521.055 2216.665 ;
        RECT 3521.485 2216.385 3521.765 2216.665 ;
        RECT 3512.255 2213.765 3512.535 2214.045 ;
        RECT 3512.965 2213.765 3513.245 2214.045 ;
        RECT 3513.675 2213.765 3513.955 2214.045 ;
        RECT 3514.385 2213.765 3514.665 2214.045 ;
        RECT 3515.095 2213.765 3515.375 2214.045 ;
        RECT 3515.805 2213.765 3516.085 2214.045 ;
        RECT 3516.515 2213.765 3516.795 2214.045 ;
        RECT 3517.225 2213.765 3517.505 2214.045 ;
        RECT 3517.935 2213.765 3518.215 2214.045 ;
        RECT 3518.645 2213.765 3518.925 2214.045 ;
        RECT 3519.355 2213.765 3519.635 2214.045 ;
        RECT 3520.065 2213.765 3520.345 2214.045 ;
        RECT 3520.775 2213.765 3521.055 2214.045 ;
        RECT 3521.485 2213.765 3521.765 2214.045 ;
        RECT 3512.255 2213.055 3512.535 2213.335 ;
        RECT 3512.965 2213.055 3513.245 2213.335 ;
        RECT 3513.675 2213.055 3513.955 2213.335 ;
        RECT 3514.385 2213.055 3514.665 2213.335 ;
        RECT 3515.095 2213.055 3515.375 2213.335 ;
        RECT 3515.805 2213.055 3516.085 2213.335 ;
        RECT 3516.515 2213.055 3516.795 2213.335 ;
        RECT 3517.225 2213.055 3517.505 2213.335 ;
        RECT 3517.935 2213.055 3518.215 2213.335 ;
        RECT 3518.645 2213.055 3518.925 2213.335 ;
        RECT 3519.355 2213.055 3519.635 2213.335 ;
        RECT 3520.065 2213.055 3520.345 2213.335 ;
        RECT 3520.775 2213.055 3521.055 2213.335 ;
        RECT 3521.485 2213.055 3521.765 2213.335 ;
        RECT 3512.255 2212.345 3512.535 2212.625 ;
        RECT 3512.965 2212.345 3513.245 2212.625 ;
        RECT 3513.675 2212.345 3513.955 2212.625 ;
        RECT 3514.385 2212.345 3514.665 2212.625 ;
        RECT 3515.095 2212.345 3515.375 2212.625 ;
        RECT 3515.805 2212.345 3516.085 2212.625 ;
        RECT 3516.515 2212.345 3516.795 2212.625 ;
        RECT 3517.225 2212.345 3517.505 2212.625 ;
        RECT 3517.935 2212.345 3518.215 2212.625 ;
        RECT 3518.645 2212.345 3518.925 2212.625 ;
        RECT 3519.355 2212.345 3519.635 2212.625 ;
        RECT 3520.065 2212.345 3520.345 2212.625 ;
        RECT 3520.775 2212.345 3521.055 2212.625 ;
        RECT 3521.485 2212.345 3521.765 2212.625 ;
        RECT 3512.255 2211.635 3512.535 2211.915 ;
        RECT 3512.965 2211.635 3513.245 2211.915 ;
        RECT 3513.675 2211.635 3513.955 2211.915 ;
        RECT 3514.385 2211.635 3514.665 2211.915 ;
        RECT 3515.095 2211.635 3515.375 2211.915 ;
        RECT 3515.805 2211.635 3516.085 2211.915 ;
        RECT 3516.515 2211.635 3516.795 2211.915 ;
        RECT 3517.225 2211.635 3517.505 2211.915 ;
        RECT 3517.935 2211.635 3518.215 2211.915 ;
        RECT 3518.645 2211.635 3518.925 2211.915 ;
        RECT 3519.355 2211.635 3519.635 2211.915 ;
        RECT 3520.065 2211.635 3520.345 2211.915 ;
        RECT 3520.775 2211.635 3521.055 2211.915 ;
        RECT 3521.485 2211.635 3521.765 2211.915 ;
        RECT 3512.255 2210.925 3512.535 2211.205 ;
        RECT 3512.965 2210.925 3513.245 2211.205 ;
        RECT 3513.675 2210.925 3513.955 2211.205 ;
        RECT 3514.385 2210.925 3514.665 2211.205 ;
        RECT 3515.095 2210.925 3515.375 2211.205 ;
        RECT 3515.805 2210.925 3516.085 2211.205 ;
        RECT 3516.515 2210.925 3516.795 2211.205 ;
        RECT 3517.225 2210.925 3517.505 2211.205 ;
        RECT 3517.935 2210.925 3518.215 2211.205 ;
        RECT 3518.645 2210.925 3518.925 2211.205 ;
        RECT 3519.355 2210.925 3519.635 2211.205 ;
        RECT 3520.065 2210.925 3520.345 2211.205 ;
        RECT 3520.775 2210.925 3521.055 2211.205 ;
        RECT 3521.485 2210.925 3521.765 2211.205 ;
        RECT 3512.255 2210.215 3512.535 2210.495 ;
        RECT 3512.965 2210.215 3513.245 2210.495 ;
        RECT 3513.675 2210.215 3513.955 2210.495 ;
        RECT 3514.385 2210.215 3514.665 2210.495 ;
        RECT 3515.095 2210.215 3515.375 2210.495 ;
        RECT 3515.805 2210.215 3516.085 2210.495 ;
        RECT 3516.515 2210.215 3516.795 2210.495 ;
        RECT 3517.225 2210.215 3517.505 2210.495 ;
        RECT 3517.935 2210.215 3518.215 2210.495 ;
        RECT 3518.645 2210.215 3518.925 2210.495 ;
        RECT 3519.355 2210.215 3519.635 2210.495 ;
        RECT 3520.065 2210.215 3520.345 2210.495 ;
        RECT 3520.775 2210.215 3521.055 2210.495 ;
        RECT 3521.485 2210.215 3521.765 2210.495 ;
        RECT 3512.255 2209.505 3512.535 2209.785 ;
        RECT 3512.965 2209.505 3513.245 2209.785 ;
        RECT 3513.675 2209.505 3513.955 2209.785 ;
        RECT 3514.385 2209.505 3514.665 2209.785 ;
        RECT 3515.095 2209.505 3515.375 2209.785 ;
        RECT 3515.805 2209.505 3516.085 2209.785 ;
        RECT 3516.515 2209.505 3516.795 2209.785 ;
        RECT 3517.225 2209.505 3517.505 2209.785 ;
        RECT 3517.935 2209.505 3518.215 2209.785 ;
        RECT 3518.645 2209.505 3518.925 2209.785 ;
        RECT 3519.355 2209.505 3519.635 2209.785 ;
        RECT 3520.065 2209.505 3520.345 2209.785 ;
        RECT 3520.775 2209.505 3521.055 2209.785 ;
        RECT 3521.485 2209.505 3521.765 2209.785 ;
        RECT 3512.255 2208.795 3512.535 2209.075 ;
        RECT 3512.965 2208.795 3513.245 2209.075 ;
        RECT 3513.675 2208.795 3513.955 2209.075 ;
        RECT 3514.385 2208.795 3514.665 2209.075 ;
        RECT 3515.095 2208.795 3515.375 2209.075 ;
        RECT 3515.805 2208.795 3516.085 2209.075 ;
        RECT 3516.515 2208.795 3516.795 2209.075 ;
        RECT 3517.225 2208.795 3517.505 2209.075 ;
        RECT 3517.935 2208.795 3518.215 2209.075 ;
        RECT 3518.645 2208.795 3518.925 2209.075 ;
        RECT 3519.355 2208.795 3519.635 2209.075 ;
        RECT 3520.065 2208.795 3520.345 2209.075 ;
        RECT 3520.775 2208.795 3521.055 2209.075 ;
        RECT 3521.485 2208.795 3521.765 2209.075 ;
        RECT 3512.255 2208.085 3512.535 2208.365 ;
        RECT 3512.965 2208.085 3513.245 2208.365 ;
        RECT 3513.675 2208.085 3513.955 2208.365 ;
        RECT 3514.385 2208.085 3514.665 2208.365 ;
        RECT 3515.095 2208.085 3515.375 2208.365 ;
        RECT 3515.805 2208.085 3516.085 2208.365 ;
        RECT 3516.515 2208.085 3516.795 2208.365 ;
        RECT 3517.225 2208.085 3517.505 2208.365 ;
        RECT 3517.935 2208.085 3518.215 2208.365 ;
        RECT 3518.645 2208.085 3518.925 2208.365 ;
        RECT 3519.355 2208.085 3519.635 2208.365 ;
        RECT 3520.065 2208.085 3520.345 2208.365 ;
        RECT 3520.775 2208.085 3521.055 2208.365 ;
        RECT 3521.485 2208.085 3521.765 2208.365 ;
        RECT 3512.255 2207.375 3512.535 2207.655 ;
        RECT 3512.965 2207.375 3513.245 2207.655 ;
        RECT 3513.675 2207.375 3513.955 2207.655 ;
        RECT 3514.385 2207.375 3514.665 2207.655 ;
        RECT 3515.095 2207.375 3515.375 2207.655 ;
        RECT 3515.805 2207.375 3516.085 2207.655 ;
        RECT 3516.515 2207.375 3516.795 2207.655 ;
        RECT 3517.225 2207.375 3517.505 2207.655 ;
        RECT 3517.935 2207.375 3518.215 2207.655 ;
        RECT 3518.645 2207.375 3518.925 2207.655 ;
        RECT 3519.355 2207.375 3519.635 2207.655 ;
        RECT 3520.065 2207.375 3520.345 2207.655 ;
        RECT 3520.775 2207.375 3521.055 2207.655 ;
        RECT 3521.485 2207.375 3521.765 2207.655 ;
        RECT 3512.255 2206.665 3512.535 2206.945 ;
        RECT 3512.965 2206.665 3513.245 2206.945 ;
        RECT 3513.675 2206.665 3513.955 2206.945 ;
        RECT 3514.385 2206.665 3514.665 2206.945 ;
        RECT 3515.095 2206.665 3515.375 2206.945 ;
        RECT 3515.805 2206.665 3516.085 2206.945 ;
        RECT 3516.515 2206.665 3516.795 2206.945 ;
        RECT 3517.225 2206.665 3517.505 2206.945 ;
        RECT 3517.935 2206.665 3518.215 2206.945 ;
        RECT 3518.645 2206.665 3518.925 2206.945 ;
        RECT 3519.355 2206.665 3519.635 2206.945 ;
        RECT 3520.065 2206.665 3520.345 2206.945 ;
        RECT 3520.775 2206.665 3521.055 2206.945 ;
        RECT 3521.485 2206.665 3521.765 2206.945 ;
        RECT 3512.255 2205.955 3512.535 2206.235 ;
        RECT 3512.965 2205.955 3513.245 2206.235 ;
        RECT 3513.675 2205.955 3513.955 2206.235 ;
        RECT 3514.385 2205.955 3514.665 2206.235 ;
        RECT 3515.095 2205.955 3515.375 2206.235 ;
        RECT 3515.805 2205.955 3516.085 2206.235 ;
        RECT 3516.515 2205.955 3516.795 2206.235 ;
        RECT 3517.225 2205.955 3517.505 2206.235 ;
        RECT 3517.935 2205.955 3518.215 2206.235 ;
        RECT 3518.645 2205.955 3518.925 2206.235 ;
        RECT 3519.355 2205.955 3519.635 2206.235 ;
        RECT 3520.065 2205.955 3520.345 2206.235 ;
        RECT 3520.775 2205.955 3521.055 2206.235 ;
        RECT 3521.485 2205.955 3521.765 2206.235 ;
        RECT 3512.255 2205.245 3512.535 2205.525 ;
        RECT 3512.965 2205.245 3513.245 2205.525 ;
        RECT 3513.675 2205.245 3513.955 2205.525 ;
        RECT 3514.385 2205.245 3514.665 2205.525 ;
        RECT 3515.095 2205.245 3515.375 2205.525 ;
        RECT 3515.805 2205.245 3516.085 2205.525 ;
        RECT 3516.515 2205.245 3516.795 2205.525 ;
        RECT 3517.225 2205.245 3517.505 2205.525 ;
        RECT 3517.935 2205.245 3518.215 2205.525 ;
        RECT 3518.645 2205.245 3518.925 2205.525 ;
        RECT 3519.355 2205.245 3519.635 2205.525 ;
        RECT 3520.065 2205.245 3520.345 2205.525 ;
        RECT 3520.775 2205.245 3521.055 2205.525 ;
        RECT 3521.485 2205.245 3521.765 2205.525 ;
        RECT 3512.255 2204.535 3512.535 2204.815 ;
        RECT 3512.965 2204.535 3513.245 2204.815 ;
        RECT 3513.675 2204.535 3513.955 2204.815 ;
        RECT 3514.385 2204.535 3514.665 2204.815 ;
        RECT 3515.095 2204.535 3515.375 2204.815 ;
        RECT 3515.805 2204.535 3516.085 2204.815 ;
        RECT 3516.515 2204.535 3516.795 2204.815 ;
        RECT 3517.225 2204.535 3517.505 2204.815 ;
        RECT 3517.935 2204.535 3518.215 2204.815 ;
        RECT 3518.645 2204.535 3518.925 2204.815 ;
        RECT 3519.355 2204.535 3519.635 2204.815 ;
        RECT 3520.065 2204.535 3520.345 2204.815 ;
        RECT 3520.775 2204.535 3521.055 2204.815 ;
        RECT 3521.485 2204.535 3521.765 2204.815 ;
        RECT 3512.255 2200.235 3512.535 2200.515 ;
        RECT 3512.965 2200.235 3513.245 2200.515 ;
        RECT 3513.675 2200.235 3513.955 2200.515 ;
        RECT 3514.385 2200.235 3514.665 2200.515 ;
        RECT 3515.095 2200.235 3515.375 2200.515 ;
        RECT 3515.805 2200.235 3516.085 2200.515 ;
        RECT 3516.515 2200.235 3516.795 2200.515 ;
        RECT 3517.225 2200.235 3517.505 2200.515 ;
        RECT 3517.935 2200.235 3518.215 2200.515 ;
        RECT 3518.645 2200.235 3518.925 2200.515 ;
        RECT 3519.355 2200.235 3519.635 2200.515 ;
        RECT 3520.065 2200.235 3520.345 2200.515 ;
        RECT 3520.775 2200.235 3521.055 2200.515 ;
        RECT 3521.485 2200.235 3521.765 2200.515 ;
        RECT 3512.255 2199.525 3512.535 2199.805 ;
        RECT 3512.965 2199.525 3513.245 2199.805 ;
        RECT 3513.675 2199.525 3513.955 2199.805 ;
        RECT 3514.385 2199.525 3514.665 2199.805 ;
        RECT 3515.095 2199.525 3515.375 2199.805 ;
        RECT 3515.805 2199.525 3516.085 2199.805 ;
        RECT 3516.515 2199.525 3516.795 2199.805 ;
        RECT 3517.225 2199.525 3517.505 2199.805 ;
        RECT 3517.935 2199.525 3518.215 2199.805 ;
        RECT 3518.645 2199.525 3518.925 2199.805 ;
        RECT 3519.355 2199.525 3519.635 2199.805 ;
        RECT 3520.065 2199.525 3520.345 2199.805 ;
        RECT 3520.775 2199.525 3521.055 2199.805 ;
        RECT 3521.485 2199.525 3521.765 2199.805 ;
        RECT 3512.255 2198.815 3512.535 2199.095 ;
        RECT 3512.965 2198.815 3513.245 2199.095 ;
        RECT 3513.675 2198.815 3513.955 2199.095 ;
        RECT 3514.385 2198.815 3514.665 2199.095 ;
        RECT 3515.095 2198.815 3515.375 2199.095 ;
        RECT 3515.805 2198.815 3516.085 2199.095 ;
        RECT 3516.515 2198.815 3516.795 2199.095 ;
        RECT 3517.225 2198.815 3517.505 2199.095 ;
        RECT 3517.935 2198.815 3518.215 2199.095 ;
        RECT 3518.645 2198.815 3518.925 2199.095 ;
        RECT 3519.355 2198.815 3519.635 2199.095 ;
        RECT 3520.065 2198.815 3520.345 2199.095 ;
        RECT 3520.775 2198.815 3521.055 2199.095 ;
        RECT 3521.485 2198.815 3521.765 2199.095 ;
        RECT 3512.255 2198.105 3512.535 2198.385 ;
        RECT 3512.965 2198.105 3513.245 2198.385 ;
        RECT 3513.675 2198.105 3513.955 2198.385 ;
        RECT 3514.385 2198.105 3514.665 2198.385 ;
        RECT 3515.095 2198.105 3515.375 2198.385 ;
        RECT 3515.805 2198.105 3516.085 2198.385 ;
        RECT 3516.515 2198.105 3516.795 2198.385 ;
        RECT 3517.225 2198.105 3517.505 2198.385 ;
        RECT 3517.935 2198.105 3518.215 2198.385 ;
        RECT 3518.645 2198.105 3518.925 2198.385 ;
        RECT 3519.355 2198.105 3519.635 2198.385 ;
        RECT 3520.065 2198.105 3520.345 2198.385 ;
        RECT 3520.775 2198.105 3521.055 2198.385 ;
        RECT 3521.485 2198.105 3521.765 2198.385 ;
        RECT 3512.255 2197.395 3512.535 2197.675 ;
        RECT 3512.965 2197.395 3513.245 2197.675 ;
        RECT 3513.675 2197.395 3513.955 2197.675 ;
        RECT 3514.385 2197.395 3514.665 2197.675 ;
        RECT 3515.095 2197.395 3515.375 2197.675 ;
        RECT 3515.805 2197.395 3516.085 2197.675 ;
        RECT 3516.515 2197.395 3516.795 2197.675 ;
        RECT 3517.225 2197.395 3517.505 2197.675 ;
        RECT 3517.935 2197.395 3518.215 2197.675 ;
        RECT 3518.645 2197.395 3518.925 2197.675 ;
        RECT 3519.355 2197.395 3519.635 2197.675 ;
        RECT 3520.065 2197.395 3520.345 2197.675 ;
        RECT 3520.775 2197.395 3521.055 2197.675 ;
        RECT 3521.485 2197.395 3521.765 2197.675 ;
        RECT 3512.255 2196.685 3512.535 2196.965 ;
        RECT 3512.965 2196.685 3513.245 2196.965 ;
        RECT 3513.675 2196.685 3513.955 2196.965 ;
        RECT 3514.385 2196.685 3514.665 2196.965 ;
        RECT 3515.095 2196.685 3515.375 2196.965 ;
        RECT 3515.805 2196.685 3516.085 2196.965 ;
        RECT 3516.515 2196.685 3516.795 2196.965 ;
        RECT 3517.225 2196.685 3517.505 2196.965 ;
        RECT 3517.935 2196.685 3518.215 2196.965 ;
        RECT 3518.645 2196.685 3518.925 2196.965 ;
        RECT 3519.355 2196.685 3519.635 2196.965 ;
        RECT 3520.065 2196.685 3520.345 2196.965 ;
        RECT 3520.775 2196.685 3521.055 2196.965 ;
        RECT 3521.485 2196.685 3521.765 2196.965 ;
        RECT 3512.255 2195.975 3512.535 2196.255 ;
        RECT 3512.965 2195.975 3513.245 2196.255 ;
        RECT 3513.675 2195.975 3513.955 2196.255 ;
        RECT 3514.385 2195.975 3514.665 2196.255 ;
        RECT 3515.095 2195.975 3515.375 2196.255 ;
        RECT 3515.805 2195.975 3516.085 2196.255 ;
        RECT 3516.515 2195.975 3516.795 2196.255 ;
        RECT 3517.225 2195.975 3517.505 2196.255 ;
        RECT 3517.935 2195.975 3518.215 2196.255 ;
        RECT 3518.645 2195.975 3518.925 2196.255 ;
        RECT 3519.355 2195.975 3519.635 2196.255 ;
        RECT 3520.065 2195.975 3520.345 2196.255 ;
        RECT 3520.775 2195.975 3521.055 2196.255 ;
        RECT 3521.485 2195.975 3521.765 2196.255 ;
        RECT 3512.255 2195.265 3512.535 2195.545 ;
        RECT 3512.965 2195.265 3513.245 2195.545 ;
        RECT 3513.675 2195.265 3513.955 2195.545 ;
        RECT 3514.385 2195.265 3514.665 2195.545 ;
        RECT 3515.095 2195.265 3515.375 2195.545 ;
        RECT 3515.805 2195.265 3516.085 2195.545 ;
        RECT 3516.515 2195.265 3516.795 2195.545 ;
        RECT 3517.225 2195.265 3517.505 2195.545 ;
        RECT 3517.935 2195.265 3518.215 2195.545 ;
        RECT 3518.645 2195.265 3518.925 2195.545 ;
        RECT 3519.355 2195.265 3519.635 2195.545 ;
        RECT 3520.065 2195.265 3520.345 2195.545 ;
        RECT 3520.775 2195.265 3521.055 2195.545 ;
        RECT 3521.485 2195.265 3521.765 2195.545 ;
        RECT 3512.255 2194.555 3512.535 2194.835 ;
        RECT 3512.965 2194.555 3513.245 2194.835 ;
        RECT 3513.675 2194.555 3513.955 2194.835 ;
        RECT 3514.385 2194.555 3514.665 2194.835 ;
        RECT 3515.095 2194.555 3515.375 2194.835 ;
        RECT 3515.805 2194.555 3516.085 2194.835 ;
        RECT 3516.515 2194.555 3516.795 2194.835 ;
        RECT 3517.225 2194.555 3517.505 2194.835 ;
        RECT 3517.935 2194.555 3518.215 2194.835 ;
        RECT 3518.645 2194.555 3518.925 2194.835 ;
        RECT 3519.355 2194.555 3519.635 2194.835 ;
        RECT 3520.065 2194.555 3520.345 2194.835 ;
        RECT 3520.775 2194.555 3521.055 2194.835 ;
        RECT 3521.485 2194.555 3521.765 2194.835 ;
        RECT 3512.255 2193.845 3512.535 2194.125 ;
        RECT 3512.965 2193.845 3513.245 2194.125 ;
        RECT 3513.675 2193.845 3513.955 2194.125 ;
        RECT 3514.385 2193.845 3514.665 2194.125 ;
        RECT 3515.095 2193.845 3515.375 2194.125 ;
        RECT 3515.805 2193.845 3516.085 2194.125 ;
        RECT 3516.515 2193.845 3516.795 2194.125 ;
        RECT 3517.225 2193.845 3517.505 2194.125 ;
        RECT 3517.935 2193.845 3518.215 2194.125 ;
        RECT 3518.645 2193.845 3518.925 2194.125 ;
        RECT 3519.355 2193.845 3519.635 2194.125 ;
        RECT 3520.065 2193.845 3520.345 2194.125 ;
        RECT 3520.775 2193.845 3521.055 2194.125 ;
        RECT 3521.485 2193.845 3521.765 2194.125 ;
        RECT 3512.255 2193.135 3512.535 2193.415 ;
        RECT 3512.965 2193.135 3513.245 2193.415 ;
        RECT 3513.675 2193.135 3513.955 2193.415 ;
        RECT 3514.385 2193.135 3514.665 2193.415 ;
        RECT 3515.095 2193.135 3515.375 2193.415 ;
        RECT 3515.805 2193.135 3516.085 2193.415 ;
        RECT 3516.515 2193.135 3516.795 2193.415 ;
        RECT 3517.225 2193.135 3517.505 2193.415 ;
        RECT 3517.935 2193.135 3518.215 2193.415 ;
        RECT 3518.645 2193.135 3518.925 2193.415 ;
        RECT 3519.355 2193.135 3519.635 2193.415 ;
        RECT 3520.065 2193.135 3520.345 2193.415 ;
        RECT 3520.775 2193.135 3521.055 2193.415 ;
        RECT 3521.485 2193.135 3521.765 2193.415 ;
        RECT 3512.255 2192.425 3512.535 2192.705 ;
        RECT 3512.965 2192.425 3513.245 2192.705 ;
        RECT 3513.675 2192.425 3513.955 2192.705 ;
        RECT 3514.385 2192.425 3514.665 2192.705 ;
        RECT 3515.095 2192.425 3515.375 2192.705 ;
        RECT 3515.805 2192.425 3516.085 2192.705 ;
        RECT 3516.515 2192.425 3516.795 2192.705 ;
        RECT 3517.225 2192.425 3517.505 2192.705 ;
        RECT 3517.935 2192.425 3518.215 2192.705 ;
        RECT 3518.645 2192.425 3518.925 2192.705 ;
        RECT 3519.355 2192.425 3519.635 2192.705 ;
        RECT 3520.065 2192.425 3520.345 2192.705 ;
        RECT 3520.775 2192.425 3521.055 2192.705 ;
        RECT 3521.485 2192.425 3521.765 2192.705 ;
        RECT 3512.255 2191.715 3512.535 2191.995 ;
        RECT 3512.965 2191.715 3513.245 2191.995 ;
        RECT 3513.675 2191.715 3513.955 2191.995 ;
        RECT 3514.385 2191.715 3514.665 2191.995 ;
        RECT 3515.095 2191.715 3515.375 2191.995 ;
        RECT 3515.805 2191.715 3516.085 2191.995 ;
        RECT 3516.515 2191.715 3516.795 2191.995 ;
        RECT 3517.225 2191.715 3517.505 2191.995 ;
        RECT 3517.935 2191.715 3518.215 2191.995 ;
        RECT 3518.645 2191.715 3518.925 2191.995 ;
        RECT 3519.355 2191.715 3519.635 2191.995 ;
        RECT 3520.065 2191.715 3520.345 2191.995 ;
        RECT 3520.775 2191.715 3521.055 2191.995 ;
        RECT 3521.485 2191.715 3521.765 2191.995 ;
        RECT 3512.255 2191.005 3512.535 2191.285 ;
        RECT 3512.965 2191.005 3513.245 2191.285 ;
        RECT 3513.675 2191.005 3513.955 2191.285 ;
        RECT 3514.385 2191.005 3514.665 2191.285 ;
        RECT 3515.095 2191.005 3515.375 2191.285 ;
        RECT 3515.805 2191.005 3516.085 2191.285 ;
        RECT 3516.515 2191.005 3516.795 2191.285 ;
        RECT 3517.225 2191.005 3517.505 2191.285 ;
        RECT 3517.935 2191.005 3518.215 2191.285 ;
        RECT 3518.645 2191.005 3518.925 2191.285 ;
        RECT 3519.355 2191.005 3519.635 2191.285 ;
        RECT 3520.065 2191.005 3520.345 2191.285 ;
        RECT 3520.775 2191.005 3521.055 2191.285 ;
        RECT 3521.485 2191.005 3521.765 2191.285 ;
        RECT 3512.255 2188.385 3512.535 2188.665 ;
        RECT 3512.965 2188.385 3513.245 2188.665 ;
        RECT 3513.675 2188.385 3513.955 2188.665 ;
        RECT 3514.385 2188.385 3514.665 2188.665 ;
        RECT 3515.095 2188.385 3515.375 2188.665 ;
        RECT 3515.805 2188.385 3516.085 2188.665 ;
        RECT 3516.515 2188.385 3516.795 2188.665 ;
        RECT 3517.225 2188.385 3517.505 2188.665 ;
        RECT 3517.935 2188.385 3518.215 2188.665 ;
        RECT 3518.645 2188.385 3518.925 2188.665 ;
        RECT 3519.355 2188.385 3519.635 2188.665 ;
        RECT 3520.065 2188.385 3520.345 2188.665 ;
        RECT 3520.775 2188.385 3521.055 2188.665 ;
        RECT 3521.485 2188.385 3521.765 2188.665 ;
        RECT 3512.255 2187.675 3512.535 2187.955 ;
        RECT 3512.965 2187.675 3513.245 2187.955 ;
        RECT 3513.675 2187.675 3513.955 2187.955 ;
        RECT 3514.385 2187.675 3514.665 2187.955 ;
        RECT 3515.095 2187.675 3515.375 2187.955 ;
        RECT 3515.805 2187.675 3516.085 2187.955 ;
        RECT 3516.515 2187.675 3516.795 2187.955 ;
        RECT 3517.225 2187.675 3517.505 2187.955 ;
        RECT 3517.935 2187.675 3518.215 2187.955 ;
        RECT 3518.645 2187.675 3518.925 2187.955 ;
        RECT 3519.355 2187.675 3519.635 2187.955 ;
        RECT 3520.065 2187.675 3520.345 2187.955 ;
        RECT 3520.775 2187.675 3521.055 2187.955 ;
        RECT 3521.485 2187.675 3521.765 2187.955 ;
        RECT 3512.255 2186.965 3512.535 2187.245 ;
        RECT 3512.965 2186.965 3513.245 2187.245 ;
        RECT 3513.675 2186.965 3513.955 2187.245 ;
        RECT 3514.385 2186.965 3514.665 2187.245 ;
        RECT 3515.095 2186.965 3515.375 2187.245 ;
        RECT 3515.805 2186.965 3516.085 2187.245 ;
        RECT 3516.515 2186.965 3516.795 2187.245 ;
        RECT 3517.225 2186.965 3517.505 2187.245 ;
        RECT 3517.935 2186.965 3518.215 2187.245 ;
        RECT 3518.645 2186.965 3518.925 2187.245 ;
        RECT 3519.355 2186.965 3519.635 2187.245 ;
        RECT 3520.065 2186.965 3520.345 2187.245 ;
        RECT 3520.775 2186.965 3521.055 2187.245 ;
        RECT 3521.485 2186.965 3521.765 2187.245 ;
        RECT 3512.255 2186.255 3512.535 2186.535 ;
        RECT 3512.965 2186.255 3513.245 2186.535 ;
        RECT 3513.675 2186.255 3513.955 2186.535 ;
        RECT 3514.385 2186.255 3514.665 2186.535 ;
        RECT 3515.095 2186.255 3515.375 2186.535 ;
        RECT 3515.805 2186.255 3516.085 2186.535 ;
        RECT 3516.515 2186.255 3516.795 2186.535 ;
        RECT 3517.225 2186.255 3517.505 2186.535 ;
        RECT 3517.935 2186.255 3518.215 2186.535 ;
        RECT 3518.645 2186.255 3518.925 2186.535 ;
        RECT 3519.355 2186.255 3519.635 2186.535 ;
        RECT 3520.065 2186.255 3520.345 2186.535 ;
        RECT 3520.775 2186.255 3521.055 2186.535 ;
        RECT 3521.485 2186.255 3521.765 2186.535 ;
        RECT 3512.255 2185.545 3512.535 2185.825 ;
        RECT 3512.965 2185.545 3513.245 2185.825 ;
        RECT 3513.675 2185.545 3513.955 2185.825 ;
        RECT 3514.385 2185.545 3514.665 2185.825 ;
        RECT 3515.095 2185.545 3515.375 2185.825 ;
        RECT 3515.805 2185.545 3516.085 2185.825 ;
        RECT 3516.515 2185.545 3516.795 2185.825 ;
        RECT 3517.225 2185.545 3517.505 2185.825 ;
        RECT 3517.935 2185.545 3518.215 2185.825 ;
        RECT 3518.645 2185.545 3518.925 2185.825 ;
        RECT 3519.355 2185.545 3519.635 2185.825 ;
        RECT 3520.065 2185.545 3520.345 2185.825 ;
        RECT 3520.775 2185.545 3521.055 2185.825 ;
        RECT 3521.485 2185.545 3521.765 2185.825 ;
        RECT 3512.255 2184.835 3512.535 2185.115 ;
        RECT 3512.965 2184.835 3513.245 2185.115 ;
        RECT 3513.675 2184.835 3513.955 2185.115 ;
        RECT 3514.385 2184.835 3514.665 2185.115 ;
        RECT 3515.095 2184.835 3515.375 2185.115 ;
        RECT 3515.805 2184.835 3516.085 2185.115 ;
        RECT 3516.515 2184.835 3516.795 2185.115 ;
        RECT 3517.225 2184.835 3517.505 2185.115 ;
        RECT 3517.935 2184.835 3518.215 2185.115 ;
        RECT 3518.645 2184.835 3518.925 2185.115 ;
        RECT 3519.355 2184.835 3519.635 2185.115 ;
        RECT 3520.065 2184.835 3520.345 2185.115 ;
        RECT 3520.775 2184.835 3521.055 2185.115 ;
        RECT 3521.485 2184.835 3521.765 2185.115 ;
        RECT 3512.255 2184.125 3512.535 2184.405 ;
        RECT 3512.965 2184.125 3513.245 2184.405 ;
        RECT 3513.675 2184.125 3513.955 2184.405 ;
        RECT 3514.385 2184.125 3514.665 2184.405 ;
        RECT 3515.095 2184.125 3515.375 2184.405 ;
        RECT 3515.805 2184.125 3516.085 2184.405 ;
        RECT 3516.515 2184.125 3516.795 2184.405 ;
        RECT 3517.225 2184.125 3517.505 2184.405 ;
        RECT 3517.935 2184.125 3518.215 2184.405 ;
        RECT 3518.645 2184.125 3518.925 2184.405 ;
        RECT 3519.355 2184.125 3519.635 2184.405 ;
        RECT 3520.065 2184.125 3520.345 2184.405 ;
        RECT 3520.775 2184.125 3521.055 2184.405 ;
        RECT 3521.485 2184.125 3521.765 2184.405 ;
        RECT 3512.255 2183.415 3512.535 2183.695 ;
        RECT 3512.965 2183.415 3513.245 2183.695 ;
        RECT 3513.675 2183.415 3513.955 2183.695 ;
        RECT 3514.385 2183.415 3514.665 2183.695 ;
        RECT 3515.095 2183.415 3515.375 2183.695 ;
        RECT 3515.805 2183.415 3516.085 2183.695 ;
        RECT 3516.515 2183.415 3516.795 2183.695 ;
        RECT 3517.225 2183.415 3517.505 2183.695 ;
        RECT 3517.935 2183.415 3518.215 2183.695 ;
        RECT 3518.645 2183.415 3518.925 2183.695 ;
        RECT 3519.355 2183.415 3519.635 2183.695 ;
        RECT 3520.065 2183.415 3520.345 2183.695 ;
        RECT 3520.775 2183.415 3521.055 2183.695 ;
        RECT 3521.485 2183.415 3521.765 2183.695 ;
        RECT 3512.255 2182.705 3512.535 2182.985 ;
        RECT 3512.965 2182.705 3513.245 2182.985 ;
        RECT 3513.675 2182.705 3513.955 2182.985 ;
        RECT 3514.385 2182.705 3514.665 2182.985 ;
        RECT 3515.095 2182.705 3515.375 2182.985 ;
        RECT 3515.805 2182.705 3516.085 2182.985 ;
        RECT 3516.515 2182.705 3516.795 2182.985 ;
        RECT 3517.225 2182.705 3517.505 2182.985 ;
        RECT 3517.935 2182.705 3518.215 2182.985 ;
        RECT 3518.645 2182.705 3518.925 2182.985 ;
        RECT 3519.355 2182.705 3519.635 2182.985 ;
        RECT 3520.065 2182.705 3520.345 2182.985 ;
        RECT 3520.775 2182.705 3521.055 2182.985 ;
        RECT 3521.485 2182.705 3521.765 2182.985 ;
        RECT 3512.255 2181.995 3512.535 2182.275 ;
        RECT 3512.965 2181.995 3513.245 2182.275 ;
        RECT 3513.675 2181.995 3513.955 2182.275 ;
        RECT 3514.385 2181.995 3514.665 2182.275 ;
        RECT 3515.095 2181.995 3515.375 2182.275 ;
        RECT 3515.805 2181.995 3516.085 2182.275 ;
        RECT 3516.515 2181.995 3516.795 2182.275 ;
        RECT 3517.225 2181.995 3517.505 2182.275 ;
        RECT 3517.935 2181.995 3518.215 2182.275 ;
        RECT 3518.645 2181.995 3518.925 2182.275 ;
        RECT 3519.355 2181.995 3519.635 2182.275 ;
        RECT 3520.065 2181.995 3520.345 2182.275 ;
        RECT 3520.775 2181.995 3521.055 2182.275 ;
        RECT 3521.485 2181.995 3521.765 2182.275 ;
        RECT 3512.255 2181.285 3512.535 2181.565 ;
        RECT 3512.965 2181.285 3513.245 2181.565 ;
        RECT 3513.675 2181.285 3513.955 2181.565 ;
        RECT 3514.385 2181.285 3514.665 2181.565 ;
        RECT 3515.095 2181.285 3515.375 2181.565 ;
        RECT 3515.805 2181.285 3516.085 2181.565 ;
        RECT 3516.515 2181.285 3516.795 2181.565 ;
        RECT 3517.225 2181.285 3517.505 2181.565 ;
        RECT 3517.935 2181.285 3518.215 2181.565 ;
        RECT 3518.645 2181.285 3518.925 2181.565 ;
        RECT 3519.355 2181.285 3519.635 2181.565 ;
        RECT 3520.065 2181.285 3520.345 2181.565 ;
        RECT 3520.775 2181.285 3521.055 2181.565 ;
        RECT 3521.485 2181.285 3521.765 2181.565 ;
        RECT 3512.255 2180.575 3512.535 2180.855 ;
        RECT 3512.965 2180.575 3513.245 2180.855 ;
        RECT 3513.675 2180.575 3513.955 2180.855 ;
        RECT 3514.385 2180.575 3514.665 2180.855 ;
        RECT 3515.095 2180.575 3515.375 2180.855 ;
        RECT 3515.805 2180.575 3516.085 2180.855 ;
        RECT 3516.515 2180.575 3516.795 2180.855 ;
        RECT 3517.225 2180.575 3517.505 2180.855 ;
        RECT 3517.935 2180.575 3518.215 2180.855 ;
        RECT 3518.645 2180.575 3518.925 2180.855 ;
        RECT 3519.355 2180.575 3519.635 2180.855 ;
        RECT 3520.065 2180.575 3520.345 2180.855 ;
        RECT 3520.775 2180.575 3521.055 2180.855 ;
        RECT 3521.485 2180.575 3521.765 2180.855 ;
        RECT 3512.200 2175.270 3512.480 2175.550 ;
        RECT 3512.910 2175.270 3513.190 2175.550 ;
        RECT 3513.620 2175.270 3513.900 2175.550 ;
        RECT 3514.330 2175.270 3514.610 2175.550 ;
        RECT 3515.040 2175.270 3515.320 2175.550 ;
        RECT 3515.750 2175.270 3516.030 2175.550 ;
        RECT 3516.460 2175.270 3516.740 2175.550 ;
        RECT 3517.170 2175.270 3517.450 2175.550 ;
        RECT 3517.880 2175.270 3518.160 2175.550 ;
        RECT 3518.590 2175.270 3518.870 2175.550 ;
        RECT 3519.300 2175.270 3519.580 2175.550 ;
        RECT 3520.010 2175.270 3520.290 2175.550 ;
        RECT 3520.720 2175.270 3521.000 2175.550 ;
        RECT 3521.430 2175.270 3521.710 2175.550 ;
        RECT 3512.200 2174.560 3512.480 2174.840 ;
        RECT 3512.910 2174.560 3513.190 2174.840 ;
        RECT 3513.620 2174.560 3513.900 2174.840 ;
        RECT 3514.330 2174.560 3514.610 2174.840 ;
        RECT 3515.040 2174.560 3515.320 2174.840 ;
        RECT 3515.750 2174.560 3516.030 2174.840 ;
        RECT 3516.460 2174.560 3516.740 2174.840 ;
        RECT 3517.170 2174.560 3517.450 2174.840 ;
        RECT 3517.880 2174.560 3518.160 2174.840 ;
        RECT 3518.590 2174.560 3518.870 2174.840 ;
        RECT 3519.300 2174.560 3519.580 2174.840 ;
        RECT 3520.010 2174.560 3520.290 2174.840 ;
        RECT 3520.720 2174.560 3521.000 2174.840 ;
        RECT 3521.430 2174.560 3521.710 2174.840 ;
        RECT 3512.200 2173.850 3512.480 2174.130 ;
        RECT 3512.910 2173.850 3513.190 2174.130 ;
        RECT 3513.620 2173.850 3513.900 2174.130 ;
        RECT 3514.330 2173.850 3514.610 2174.130 ;
        RECT 3515.040 2173.850 3515.320 2174.130 ;
        RECT 3515.750 2173.850 3516.030 2174.130 ;
        RECT 3516.460 2173.850 3516.740 2174.130 ;
        RECT 3517.170 2173.850 3517.450 2174.130 ;
        RECT 3517.880 2173.850 3518.160 2174.130 ;
        RECT 3518.590 2173.850 3518.870 2174.130 ;
        RECT 3519.300 2173.850 3519.580 2174.130 ;
        RECT 3520.010 2173.850 3520.290 2174.130 ;
        RECT 3520.720 2173.850 3521.000 2174.130 ;
        RECT 3521.430 2173.850 3521.710 2174.130 ;
        RECT 3512.200 2173.140 3512.480 2173.420 ;
        RECT 3512.910 2173.140 3513.190 2173.420 ;
        RECT 3513.620 2173.140 3513.900 2173.420 ;
        RECT 3514.330 2173.140 3514.610 2173.420 ;
        RECT 3515.040 2173.140 3515.320 2173.420 ;
        RECT 3515.750 2173.140 3516.030 2173.420 ;
        RECT 3516.460 2173.140 3516.740 2173.420 ;
        RECT 3517.170 2173.140 3517.450 2173.420 ;
        RECT 3517.880 2173.140 3518.160 2173.420 ;
        RECT 3518.590 2173.140 3518.870 2173.420 ;
        RECT 3519.300 2173.140 3519.580 2173.420 ;
        RECT 3520.010 2173.140 3520.290 2173.420 ;
        RECT 3520.720 2173.140 3521.000 2173.420 ;
        RECT 3521.430 2173.140 3521.710 2173.420 ;
        RECT 3512.200 2172.430 3512.480 2172.710 ;
        RECT 3512.910 2172.430 3513.190 2172.710 ;
        RECT 3513.620 2172.430 3513.900 2172.710 ;
        RECT 3514.330 2172.430 3514.610 2172.710 ;
        RECT 3515.040 2172.430 3515.320 2172.710 ;
        RECT 3515.750 2172.430 3516.030 2172.710 ;
        RECT 3516.460 2172.430 3516.740 2172.710 ;
        RECT 3517.170 2172.430 3517.450 2172.710 ;
        RECT 3517.880 2172.430 3518.160 2172.710 ;
        RECT 3518.590 2172.430 3518.870 2172.710 ;
        RECT 3519.300 2172.430 3519.580 2172.710 ;
        RECT 3520.010 2172.430 3520.290 2172.710 ;
        RECT 3520.720 2172.430 3521.000 2172.710 ;
        RECT 3521.430 2172.430 3521.710 2172.710 ;
        RECT 3512.200 2171.720 3512.480 2172.000 ;
        RECT 3512.910 2171.720 3513.190 2172.000 ;
        RECT 3513.620 2171.720 3513.900 2172.000 ;
        RECT 3514.330 2171.720 3514.610 2172.000 ;
        RECT 3515.040 2171.720 3515.320 2172.000 ;
        RECT 3515.750 2171.720 3516.030 2172.000 ;
        RECT 3516.460 2171.720 3516.740 2172.000 ;
        RECT 3517.170 2171.720 3517.450 2172.000 ;
        RECT 3517.880 2171.720 3518.160 2172.000 ;
        RECT 3518.590 2171.720 3518.870 2172.000 ;
        RECT 3519.300 2171.720 3519.580 2172.000 ;
        RECT 3520.010 2171.720 3520.290 2172.000 ;
        RECT 3520.720 2171.720 3521.000 2172.000 ;
        RECT 3521.430 2171.720 3521.710 2172.000 ;
        RECT 3512.200 2171.010 3512.480 2171.290 ;
        RECT 3512.910 2171.010 3513.190 2171.290 ;
        RECT 3513.620 2171.010 3513.900 2171.290 ;
        RECT 3514.330 2171.010 3514.610 2171.290 ;
        RECT 3515.040 2171.010 3515.320 2171.290 ;
        RECT 3515.750 2171.010 3516.030 2171.290 ;
        RECT 3516.460 2171.010 3516.740 2171.290 ;
        RECT 3517.170 2171.010 3517.450 2171.290 ;
        RECT 3517.880 2171.010 3518.160 2171.290 ;
        RECT 3518.590 2171.010 3518.870 2171.290 ;
        RECT 3519.300 2171.010 3519.580 2171.290 ;
        RECT 3520.010 2171.010 3520.290 2171.290 ;
        RECT 3520.720 2171.010 3521.000 2171.290 ;
        RECT 3521.430 2171.010 3521.710 2171.290 ;
        RECT 3512.200 2170.300 3512.480 2170.580 ;
        RECT 3512.910 2170.300 3513.190 2170.580 ;
        RECT 3513.620 2170.300 3513.900 2170.580 ;
        RECT 3514.330 2170.300 3514.610 2170.580 ;
        RECT 3515.040 2170.300 3515.320 2170.580 ;
        RECT 3515.750 2170.300 3516.030 2170.580 ;
        RECT 3516.460 2170.300 3516.740 2170.580 ;
        RECT 3517.170 2170.300 3517.450 2170.580 ;
        RECT 3517.880 2170.300 3518.160 2170.580 ;
        RECT 3518.590 2170.300 3518.870 2170.580 ;
        RECT 3519.300 2170.300 3519.580 2170.580 ;
        RECT 3520.010 2170.300 3520.290 2170.580 ;
        RECT 3520.720 2170.300 3521.000 2170.580 ;
        RECT 3521.430 2170.300 3521.710 2170.580 ;
        RECT 3512.200 2169.590 3512.480 2169.870 ;
        RECT 3512.910 2169.590 3513.190 2169.870 ;
        RECT 3513.620 2169.590 3513.900 2169.870 ;
        RECT 3514.330 2169.590 3514.610 2169.870 ;
        RECT 3515.040 2169.590 3515.320 2169.870 ;
        RECT 3515.750 2169.590 3516.030 2169.870 ;
        RECT 3516.460 2169.590 3516.740 2169.870 ;
        RECT 3517.170 2169.590 3517.450 2169.870 ;
        RECT 3517.880 2169.590 3518.160 2169.870 ;
        RECT 3518.590 2169.590 3518.870 2169.870 ;
        RECT 3519.300 2169.590 3519.580 2169.870 ;
        RECT 3520.010 2169.590 3520.290 2169.870 ;
        RECT 3520.720 2169.590 3521.000 2169.870 ;
        RECT 3521.430 2169.590 3521.710 2169.870 ;
        RECT 3512.200 2168.880 3512.480 2169.160 ;
        RECT 3512.910 2168.880 3513.190 2169.160 ;
        RECT 3513.620 2168.880 3513.900 2169.160 ;
        RECT 3514.330 2168.880 3514.610 2169.160 ;
        RECT 3515.040 2168.880 3515.320 2169.160 ;
        RECT 3515.750 2168.880 3516.030 2169.160 ;
        RECT 3516.460 2168.880 3516.740 2169.160 ;
        RECT 3517.170 2168.880 3517.450 2169.160 ;
        RECT 3517.880 2168.880 3518.160 2169.160 ;
        RECT 3518.590 2168.880 3518.870 2169.160 ;
        RECT 3519.300 2168.880 3519.580 2169.160 ;
        RECT 3520.010 2168.880 3520.290 2169.160 ;
        RECT 3520.720 2168.880 3521.000 2169.160 ;
        RECT 3521.430 2168.880 3521.710 2169.160 ;
        RECT 3512.200 2168.170 3512.480 2168.450 ;
        RECT 3512.910 2168.170 3513.190 2168.450 ;
        RECT 3513.620 2168.170 3513.900 2168.450 ;
        RECT 3514.330 2168.170 3514.610 2168.450 ;
        RECT 3515.040 2168.170 3515.320 2168.450 ;
        RECT 3515.750 2168.170 3516.030 2168.450 ;
        RECT 3516.460 2168.170 3516.740 2168.450 ;
        RECT 3517.170 2168.170 3517.450 2168.450 ;
        RECT 3517.880 2168.170 3518.160 2168.450 ;
        RECT 3518.590 2168.170 3518.870 2168.450 ;
        RECT 3519.300 2168.170 3519.580 2168.450 ;
        RECT 3520.010 2168.170 3520.290 2168.450 ;
        RECT 3520.720 2168.170 3521.000 2168.450 ;
        RECT 3521.430 2168.170 3521.710 2168.450 ;
        RECT 3512.200 2167.460 3512.480 2167.740 ;
        RECT 3512.910 2167.460 3513.190 2167.740 ;
        RECT 3513.620 2167.460 3513.900 2167.740 ;
        RECT 3514.330 2167.460 3514.610 2167.740 ;
        RECT 3515.040 2167.460 3515.320 2167.740 ;
        RECT 3515.750 2167.460 3516.030 2167.740 ;
        RECT 3516.460 2167.460 3516.740 2167.740 ;
        RECT 3517.170 2167.460 3517.450 2167.740 ;
        RECT 3517.880 2167.460 3518.160 2167.740 ;
        RECT 3518.590 2167.460 3518.870 2167.740 ;
        RECT 3519.300 2167.460 3519.580 2167.740 ;
        RECT 3520.010 2167.460 3520.290 2167.740 ;
        RECT 3520.720 2167.460 3521.000 2167.740 ;
        RECT 3521.430 2167.460 3521.710 2167.740 ;
        RECT 3512.200 2166.750 3512.480 2167.030 ;
        RECT 3512.910 2166.750 3513.190 2167.030 ;
        RECT 3513.620 2166.750 3513.900 2167.030 ;
        RECT 3514.330 2166.750 3514.610 2167.030 ;
        RECT 3515.040 2166.750 3515.320 2167.030 ;
        RECT 3515.750 2166.750 3516.030 2167.030 ;
        RECT 3516.460 2166.750 3516.740 2167.030 ;
        RECT 3517.170 2166.750 3517.450 2167.030 ;
        RECT 3517.880 2166.750 3518.160 2167.030 ;
        RECT 3518.590 2166.750 3518.870 2167.030 ;
        RECT 3519.300 2166.750 3519.580 2167.030 ;
        RECT 3520.010 2166.750 3520.290 2167.030 ;
        RECT 3520.720 2166.750 3521.000 2167.030 ;
        RECT 3521.430 2166.750 3521.710 2167.030 ;
        RECT 357.330 2137.970 357.610 2138.250 ;
        RECT 358.040 2137.970 358.320 2138.250 ;
        RECT 358.750 2137.970 359.030 2138.250 ;
        RECT 359.460 2137.970 359.740 2138.250 ;
        RECT 360.170 2137.970 360.450 2138.250 ;
        RECT 360.880 2137.970 361.160 2138.250 ;
        RECT 361.590 2137.970 361.870 2138.250 ;
        RECT 362.300 2137.970 362.580 2138.250 ;
        RECT 363.010 2137.970 363.290 2138.250 ;
        RECT 363.720 2137.970 364.000 2138.250 ;
        RECT 364.430 2137.970 364.710 2138.250 ;
        RECT 365.140 2137.970 365.420 2138.250 ;
        RECT 365.850 2137.970 366.130 2138.250 ;
        RECT 366.560 2137.970 366.840 2138.250 ;
        RECT 357.330 2137.260 357.610 2137.540 ;
        RECT 358.040 2137.260 358.320 2137.540 ;
        RECT 358.750 2137.260 359.030 2137.540 ;
        RECT 359.460 2137.260 359.740 2137.540 ;
        RECT 360.170 2137.260 360.450 2137.540 ;
        RECT 360.880 2137.260 361.160 2137.540 ;
        RECT 361.590 2137.260 361.870 2137.540 ;
        RECT 362.300 2137.260 362.580 2137.540 ;
        RECT 363.010 2137.260 363.290 2137.540 ;
        RECT 363.720 2137.260 364.000 2137.540 ;
        RECT 364.430 2137.260 364.710 2137.540 ;
        RECT 365.140 2137.260 365.420 2137.540 ;
        RECT 365.850 2137.260 366.130 2137.540 ;
        RECT 366.560 2137.260 366.840 2137.540 ;
        RECT 357.330 2136.550 357.610 2136.830 ;
        RECT 358.040 2136.550 358.320 2136.830 ;
        RECT 358.750 2136.550 359.030 2136.830 ;
        RECT 359.460 2136.550 359.740 2136.830 ;
        RECT 360.170 2136.550 360.450 2136.830 ;
        RECT 360.880 2136.550 361.160 2136.830 ;
        RECT 361.590 2136.550 361.870 2136.830 ;
        RECT 362.300 2136.550 362.580 2136.830 ;
        RECT 363.010 2136.550 363.290 2136.830 ;
        RECT 363.720 2136.550 364.000 2136.830 ;
        RECT 364.430 2136.550 364.710 2136.830 ;
        RECT 365.140 2136.550 365.420 2136.830 ;
        RECT 365.850 2136.550 366.130 2136.830 ;
        RECT 366.560 2136.550 366.840 2136.830 ;
        RECT 357.330 2135.840 357.610 2136.120 ;
        RECT 358.040 2135.840 358.320 2136.120 ;
        RECT 358.750 2135.840 359.030 2136.120 ;
        RECT 359.460 2135.840 359.740 2136.120 ;
        RECT 360.170 2135.840 360.450 2136.120 ;
        RECT 360.880 2135.840 361.160 2136.120 ;
        RECT 361.590 2135.840 361.870 2136.120 ;
        RECT 362.300 2135.840 362.580 2136.120 ;
        RECT 363.010 2135.840 363.290 2136.120 ;
        RECT 363.720 2135.840 364.000 2136.120 ;
        RECT 364.430 2135.840 364.710 2136.120 ;
        RECT 365.140 2135.840 365.420 2136.120 ;
        RECT 365.850 2135.840 366.130 2136.120 ;
        RECT 366.560 2135.840 366.840 2136.120 ;
        RECT 357.330 2135.130 357.610 2135.410 ;
        RECT 358.040 2135.130 358.320 2135.410 ;
        RECT 358.750 2135.130 359.030 2135.410 ;
        RECT 359.460 2135.130 359.740 2135.410 ;
        RECT 360.170 2135.130 360.450 2135.410 ;
        RECT 360.880 2135.130 361.160 2135.410 ;
        RECT 361.590 2135.130 361.870 2135.410 ;
        RECT 362.300 2135.130 362.580 2135.410 ;
        RECT 363.010 2135.130 363.290 2135.410 ;
        RECT 363.720 2135.130 364.000 2135.410 ;
        RECT 364.430 2135.130 364.710 2135.410 ;
        RECT 365.140 2135.130 365.420 2135.410 ;
        RECT 365.850 2135.130 366.130 2135.410 ;
        RECT 366.560 2135.130 366.840 2135.410 ;
        RECT 357.330 2134.420 357.610 2134.700 ;
        RECT 358.040 2134.420 358.320 2134.700 ;
        RECT 358.750 2134.420 359.030 2134.700 ;
        RECT 359.460 2134.420 359.740 2134.700 ;
        RECT 360.170 2134.420 360.450 2134.700 ;
        RECT 360.880 2134.420 361.160 2134.700 ;
        RECT 361.590 2134.420 361.870 2134.700 ;
        RECT 362.300 2134.420 362.580 2134.700 ;
        RECT 363.010 2134.420 363.290 2134.700 ;
        RECT 363.720 2134.420 364.000 2134.700 ;
        RECT 364.430 2134.420 364.710 2134.700 ;
        RECT 365.140 2134.420 365.420 2134.700 ;
        RECT 365.850 2134.420 366.130 2134.700 ;
        RECT 366.560 2134.420 366.840 2134.700 ;
        RECT 357.330 2133.710 357.610 2133.990 ;
        RECT 358.040 2133.710 358.320 2133.990 ;
        RECT 358.750 2133.710 359.030 2133.990 ;
        RECT 359.460 2133.710 359.740 2133.990 ;
        RECT 360.170 2133.710 360.450 2133.990 ;
        RECT 360.880 2133.710 361.160 2133.990 ;
        RECT 361.590 2133.710 361.870 2133.990 ;
        RECT 362.300 2133.710 362.580 2133.990 ;
        RECT 363.010 2133.710 363.290 2133.990 ;
        RECT 363.720 2133.710 364.000 2133.990 ;
        RECT 364.430 2133.710 364.710 2133.990 ;
        RECT 365.140 2133.710 365.420 2133.990 ;
        RECT 365.850 2133.710 366.130 2133.990 ;
        RECT 366.560 2133.710 366.840 2133.990 ;
        RECT 357.330 2133.000 357.610 2133.280 ;
        RECT 358.040 2133.000 358.320 2133.280 ;
        RECT 358.750 2133.000 359.030 2133.280 ;
        RECT 359.460 2133.000 359.740 2133.280 ;
        RECT 360.170 2133.000 360.450 2133.280 ;
        RECT 360.880 2133.000 361.160 2133.280 ;
        RECT 361.590 2133.000 361.870 2133.280 ;
        RECT 362.300 2133.000 362.580 2133.280 ;
        RECT 363.010 2133.000 363.290 2133.280 ;
        RECT 363.720 2133.000 364.000 2133.280 ;
        RECT 364.430 2133.000 364.710 2133.280 ;
        RECT 365.140 2133.000 365.420 2133.280 ;
        RECT 365.850 2133.000 366.130 2133.280 ;
        RECT 366.560 2133.000 366.840 2133.280 ;
        RECT 357.330 2132.290 357.610 2132.570 ;
        RECT 358.040 2132.290 358.320 2132.570 ;
        RECT 358.750 2132.290 359.030 2132.570 ;
        RECT 359.460 2132.290 359.740 2132.570 ;
        RECT 360.170 2132.290 360.450 2132.570 ;
        RECT 360.880 2132.290 361.160 2132.570 ;
        RECT 361.590 2132.290 361.870 2132.570 ;
        RECT 362.300 2132.290 362.580 2132.570 ;
        RECT 363.010 2132.290 363.290 2132.570 ;
        RECT 363.720 2132.290 364.000 2132.570 ;
        RECT 364.430 2132.290 364.710 2132.570 ;
        RECT 365.140 2132.290 365.420 2132.570 ;
        RECT 365.850 2132.290 366.130 2132.570 ;
        RECT 366.560 2132.290 366.840 2132.570 ;
        RECT 357.330 2131.580 357.610 2131.860 ;
        RECT 358.040 2131.580 358.320 2131.860 ;
        RECT 358.750 2131.580 359.030 2131.860 ;
        RECT 359.460 2131.580 359.740 2131.860 ;
        RECT 360.170 2131.580 360.450 2131.860 ;
        RECT 360.880 2131.580 361.160 2131.860 ;
        RECT 361.590 2131.580 361.870 2131.860 ;
        RECT 362.300 2131.580 362.580 2131.860 ;
        RECT 363.010 2131.580 363.290 2131.860 ;
        RECT 363.720 2131.580 364.000 2131.860 ;
        RECT 364.430 2131.580 364.710 2131.860 ;
        RECT 365.140 2131.580 365.420 2131.860 ;
        RECT 365.850 2131.580 366.130 2131.860 ;
        RECT 366.560 2131.580 366.840 2131.860 ;
        RECT 357.330 2130.870 357.610 2131.150 ;
        RECT 358.040 2130.870 358.320 2131.150 ;
        RECT 358.750 2130.870 359.030 2131.150 ;
        RECT 359.460 2130.870 359.740 2131.150 ;
        RECT 360.170 2130.870 360.450 2131.150 ;
        RECT 360.880 2130.870 361.160 2131.150 ;
        RECT 361.590 2130.870 361.870 2131.150 ;
        RECT 362.300 2130.870 362.580 2131.150 ;
        RECT 363.010 2130.870 363.290 2131.150 ;
        RECT 363.720 2130.870 364.000 2131.150 ;
        RECT 364.430 2130.870 364.710 2131.150 ;
        RECT 365.140 2130.870 365.420 2131.150 ;
        RECT 365.850 2130.870 366.130 2131.150 ;
        RECT 366.560 2130.870 366.840 2131.150 ;
        RECT 357.330 2130.160 357.610 2130.440 ;
        RECT 358.040 2130.160 358.320 2130.440 ;
        RECT 358.750 2130.160 359.030 2130.440 ;
        RECT 359.460 2130.160 359.740 2130.440 ;
        RECT 360.170 2130.160 360.450 2130.440 ;
        RECT 360.880 2130.160 361.160 2130.440 ;
        RECT 361.590 2130.160 361.870 2130.440 ;
        RECT 362.300 2130.160 362.580 2130.440 ;
        RECT 363.010 2130.160 363.290 2130.440 ;
        RECT 363.720 2130.160 364.000 2130.440 ;
        RECT 364.430 2130.160 364.710 2130.440 ;
        RECT 365.140 2130.160 365.420 2130.440 ;
        RECT 365.850 2130.160 366.130 2130.440 ;
        RECT 366.560 2130.160 366.840 2130.440 ;
        RECT 357.330 2129.450 357.610 2129.730 ;
        RECT 358.040 2129.450 358.320 2129.730 ;
        RECT 358.750 2129.450 359.030 2129.730 ;
        RECT 359.460 2129.450 359.740 2129.730 ;
        RECT 360.170 2129.450 360.450 2129.730 ;
        RECT 360.880 2129.450 361.160 2129.730 ;
        RECT 361.590 2129.450 361.870 2129.730 ;
        RECT 362.300 2129.450 362.580 2129.730 ;
        RECT 363.010 2129.450 363.290 2129.730 ;
        RECT 363.720 2129.450 364.000 2129.730 ;
        RECT 364.430 2129.450 364.710 2129.730 ;
        RECT 365.140 2129.450 365.420 2129.730 ;
        RECT 365.850 2129.450 366.130 2129.730 ;
        RECT 366.560 2129.450 366.840 2129.730 ;
        RECT 357.275 2125.565 357.555 2125.845 ;
        RECT 357.985 2125.565 358.265 2125.845 ;
        RECT 358.695 2125.565 358.975 2125.845 ;
        RECT 359.405 2125.565 359.685 2125.845 ;
        RECT 360.115 2125.565 360.395 2125.845 ;
        RECT 360.825 2125.565 361.105 2125.845 ;
        RECT 361.535 2125.565 361.815 2125.845 ;
        RECT 362.245 2125.565 362.525 2125.845 ;
        RECT 362.955 2125.565 363.235 2125.845 ;
        RECT 363.665 2125.565 363.945 2125.845 ;
        RECT 364.375 2125.565 364.655 2125.845 ;
        RECT 365.085 2125.565 365.365 2125.845 ;
        RECT 365.795 2125.565 366.075 2125.845 ;
        RECT 366.505 2125.565 366.785 2125.845 ;
        RECT 357.275 2124.855 357.555 2125.135 ;
        RECT 357.985 2124.855 358.265 2125.135 ;
        RECT 358.695 2124.855 358.975 2125.135 ;
        RECT 359.405 2124.855 359.685 2125.135 ;
        RECT 360.115 2124.855 360.395 2125.135 ;
        RECT 360.825 2124.855 361.105 2125.135 ;
        RECT 361.535 2124.855 361.815 2125.135 ;
        RECT 362.245 2124.855 362.525 2125.135 ;
        RECT 362.955 2124.855 363.235 2125.135 ;
        RECT 363.665 2124.855 363.945 2125.135 ;
        RECT 364.375 2124.855 364.655 2125.135 ;
        RECT 365.085 2124.855 365.365 2125.135 ;
        RECT 365.795 2124.855 366.075 2125.135 ;
        RECT 366.505 2124.855 366.785 2125.135 ;
        RECT 357.275 2124.145 357.555 2124.425 ;
        RECT 357.985 2124.145 358.265 2124.425 ;
        RECT 358.695 2124.145 358.975 2124.425 ;
        RECT 359.405 2124.145 359.685 2124.425 ;
        RECT 360.115 2124.145 360.395 2124.425 ;
        RECT 360.825 2124.145 361.105 2124.425 ;
        RECT 361.535 2124.145 361.815 2124.425 ;
        RECT 362.245 2124.145 362.525 2124.425 ;
        RECT 362.955 2124.145 363.235 2124.425 ;
        RECT 363.665 2124.145 363.945 2124.425 ;
        RECT 364.375 2124.145 364.655 2124.425 ;
        RECT 365.085 2124.145 365.365 2124.425 ;
        RECT 365.795 2124.145 366.075 2124.425 ;
        RECT 366.505 2124.145 366.785 2124.425 ;
        RECT 357.275 2123.435 357.555 2123.715 ;
        RECT 357.985 2123.435 358.265 2123.715 ;
        RECT 358.695 2123.435 358.975 2123.715 ;
        RECT 359.405 2123.435 359.685 2123.715 ;
        RECT 360.115 2123.435 360.395 2123.715 ;
        RECT 360.825 2123.435 361.105 2123.715 ;
        RECT 361.535 2123.435 361.815 2123.715 ;
        RECT 362.245 2123.435 362.525 2123.715 ;
        RECT 362.955 2123.435 363.235 2123.715 ;
        RECT 363.665 2123.435 363.945 2123.715 ;
        RECT 364.375 2123.435 364.655 2123.715 ;
        RECT 365.085 2123.435 365.365 2123.715 ;
        RECT 365.795 2123.435 366.075 2123.715 ;
        RECT 366.505 2123.435 366.785 2123.715 ;
        RECT 357.275 2122.725 357.555 2123.005 ;
        RECT 357.985 2122.725 358.265 2123.005 ;
        RECT 358.695 2122.725 358.975 2123.005 ;
        RECT 359.405 2122.725 359.685 2123.005 ;
        RECT 360.115 2122.725 360.395 2123.005 ;
        RECT 360.825 2122.725 361.105 2123.005 ;
        RECT 361.535 2122.725 361.815 2123.005 ;
        RECT 362.245 2122.725 362.525 2123.005 ;
        RECT 362.955 2122.725 363.235 2123.005 ;
        RECT 363.665 2122.725 363.945 2123.005 ;
        RECT 364.375 2122.725 364.655 2123.005 ;
        RECT 365.085 2122.725 365.365 2123.005 ;
        RECT 365.795 2122.725 366.075 2123.005 ;
        RECT 366.505 2122.725 366.785 2123.005 ;
        RECT 357.275 2122.015 357.555 2122.295 ;
        RECT 357.985 2122.015 358.265 2122.295 ;
        RECT 358.695 2122.015 358.975 2122.295 ;
        RECT 359.405 2122.015 359.685 2122.295 ;
        RECT 360.115 2122.015 360.395 2122.295 ;
        RECT 360.825 2122.015 361.105 2122.295 ;
        RECT 361.535 2122.015 361.815 2122.295 ;
        RECT 362.245 2122.015 362.525 2122.295 ;
        RECT 362.955 2122.015 363.235 2122.295 ;
        RECT 363.665 2122.015 363.945 2122.295 ;
        RECT 364.375 2122.015 364.655 2122.295 ;
        RECT 365.085 2122.015 365.365 2122.295 ;
        RECT 365.795 2122.015 366.075 2122.295 ;
        RECT 366.505 2122.015 366.785 2122.295 ;
        RECT 357.275 2121.305 357.555 2121.585 ;
        RECT 357.985 2121.305 358.265 2121.585 ;
        RECT 358.695 2121.305 358.975 2121.585 ;
        RECT 359.405 2121.305 359.685 2121.585 ;
        RECT 360.115 2121.305 360.395 2121.585 ;
        RECT 360.825 2121.305 361.105 2121.585 ;
        RECT 361.535 2121.305 361.815 2121.585 ;
        RECT 362.245 2121.305 362.525 2121.585 ;
        RECT 362.955 2121.305 363.235 2121.585 ;
        RECT 363.665 2121.305 363.945 2121.585 ;
        RECT 364.375 2121.305 364.655 2121.585 ;
        RECT 365.085 2121.305 365.365 2121.585 ;
        RECT 365.795 2121.305 366.075 2121.585 ;
        RECT 366.505 2121.305 366.785 2121.585 ;
        RECT 357.275 2120.595 357.555 2120.875 ;
        RECT 357.985 2120.595 358.265 2120.875 ;
        RECT 358.695 2120.595 358.975 2120.875 ;
        RECT 359.405 2120.595 359.685 2120.875 ;
        RECT 360.115 2120.595 360.395 2120.875 ;
        RECT 360.825 2120.595 361.105 2120.875 ;
        RECT 361.535 2120.595 361.815 2120.875 ;
        RECT 362.245 2120.595 362.525 2120.875 ;
        RECT 362.955 2120.595 363.235 2120.875 ;
        RECT 363.665 2120.595 363.945 2120.875 ;
        RECT 364.375 2120.595 364.655 2120.875 ;
        RECT 365.085 2120.595 365.365 2120.875 ;
        RECT 365.795 2120.595 366.075 2120.875 ;
        RECT 366.505 2120.595 366.785 2120.875 ;
        RECT 357.275 2119.885 357.555 2120.165 ;
        RECT 357.985 2119.885 358.265 2120.165 ;
        RECT 358.695 2119.885 358.975 2120.165 ;
        RECT 359.405 2119.885 359.685 2120.165 ;
        RECT 360.115 2119.885 360.395 2120.165 ;
        RECT 360.825 2119.885 361.105 2120.165 ;
        RECT 361.535 2119.885 361.815 2120.165 ;
        RECT 362.245 2119.885 362.525 2120.165 ;
        RECT 362.955 2119.885 363.235 2120.165 ;
        RECT 363.665 2119.885 363.945 2120.165 ;
        RECT 364.375 2119.885 364.655 2120.165 ;
        RECT 365.085 2119.885 365.365 2120.165 ;
        RECT 365.795 2119.885 366.075 2120.165 ;
        RECT 366.505 2119.885 366.785 2120.165 ;
        RECT 357.275 2119.175 357.555 2119.455 ;
        RECT 357.985 2119.175 358.265 2119.455 ;
        RECT 358.695 2119.175 358.975 2119.455 ;
        RECT 359.405 2119.175 359.685 2119.455 ;
        RECT 360.115 2119.175 360.395 2119.455 ;
        RECT 360.825 2119.175 361.105 2119.455 ;
        RECT 361.535 2119.175 361.815 2119.455 ;
        RECT 362.245 2119.175 362.525 2119.455 ;
        RECT 362.955 2119.175 363.235 2119.455 ;
        RECT 363.665 2119.175 363.945 2119.455 ;
        RECT 364.375 2119.175 364.655 2119.455 ;
        RECT 365.085 2119.175 365.365 2119.455 ;
        RECT 365.795 2119.175 366.075 2119.455 ;
        RECT 366.505 2119.175 366.785 2119.455 ;
        RECT 357.275 2118.465 357.555 2118.745 ;
        RECT 357.985 2118.465 358.265 2118.745 ;
        RECT 358.695 2118.465 358.975 2118.745 ;
        RECT 359.405 2118.465 359.685 2118.745 ;
        RECT 360.115 2118.465 360.395 2118.745 ;
        RECT 360.825 2118.465 361.105 2118.745 ;
        RECT 361.535 2118.465 361.815 2118.745 ;
        RECT 362.245 2118.465 362.525 2118.745 ;
        RECT 362.955 2118.465 363.235 2118.745 ;
        RECT 363.665 2118.465 363.945 2118.745 ;
        RECT 364.375 2118.465 364.655 2118.745 ;
        RECT 365.085 2118.465 365.365 2118.745 ;
        RECT 365.795 2118.465 366.075 2118.745 ;
        RECT 366.505 2118.465 366.785 2118.745 ;
        RECT 357.275 2117.755 357.555 2118.035 ;
        RECT 357.985 2117.755 358.265 2118.035 ;
        RECT 358.695 2117.755 358.975 2118.035 ;
        RECT 359.405 2117.755 359.685 2118.035 ;
        RECT 360.115 2117.755 360.395 2118.035 ;
        RECT 360.825 2117.755 361.105 2118.035 ;
        RECT 361.535 2117.755 361.815 2118.035 ;
        RECT 362.245 2117.755 362.525 2118.035 ;
        RECT 362.955 2117.755 363.235 2118.035 ;
        RECT 363.665 2117.755 363.945 2118.035 ;
        RECT 364.375 2117.755 364.655 2118.035 ;
        RECT 365.085 2117.755 365.365 2118.035 ;
        RECT 365.795 2117.755 366.075 2118.035 ;
        RECT 366.505 2117.755 366.785 2118.035 ;
        RECT 357.275 2117.045 357.555 2117.325 ;
        RECT 357.985 2117.045 358.265 2117.325 ;
        RECT 358.695 2117.045 358.975 2117.325 ;
        RECT 359.405 2117.045 359.685 2117.325 ;
        RECT 360.115 2117.045 360.395 2117.325 ;
        RECT 360.825 2117.045 361.105 2117.325 ;
        RECT 361.535 2117.045 361.815 2117.325 ;
        RECT 362.245 2117.045 362.525 2117.325 ;
        RECT 362.955 2117.045 363.235 2117.325 ;
        RECT 363.665 2117.045 363.945 2117.325 ;
        RECT 364.375 2117.045 364.655 2117.325 ;
        RECT 365.085 2117.045 365.365 2117.325 ;
        RECT 365.795 2117.045 366.075 2117.325 ;
        RECT 366.505 2117.045 366.785 2117.325 ;
        RECT 357.275 2116.335 357.555 2116.615 ;
        RECT 357.985 2116.335 358.265 2116.615 ;
        RECT 358.695 2116.335 358.975 2116.615 ;
        RECT 359.405 2116.335 359.685 2116.615 ;
        RECT 360.115 2116.335 360.395 2116.615 ;
        RECT 360.825 2116.335 361.105 2116.615 ;
        RECT 361.535 2116.335 361.815 2116.615 ;
        RECT 362.245 2116.335 362.525 2116.615 ;
        RECT 362.955 2116.335 363.235 2116.615 ;
        RECT 363.665 2116.335 363.945 2116.615 ;
        RECT 364.375 2116.335 364.655 2116.615 ;
        RECT 365.085 2116.335 365.365 2116.615 ;
        RECT 365.795 2116.335 366.075 2116.615 ;
        RECT 366.505 2116.335 366.785 2116.615 ;
        RECT 357.275 2113.715 357.555 2113.995 ;
        RECT 357.985 2113.715 358.265 2113.995 ;
        RECT 358.695 2113.715 358.975 2113.995 ;
        RECT 359.405 2113.715 359.685 2113.995 ;
        RECT 360.115 2113.715 360.395 2113.995 ;
        RECT 360.825 2113.715 361.105 2113.995 ;
        RECT 361.535 2113.715 361.815 2113.995 ;
        RECT 362.245 2113.715 362.525 2113.995 ;
        RECT 362.955 2113.715 363.235 2113.995 ;
        RECT 363.665 2113.715 363.945 2113.995 ;
        RECT 364.375 2113.715 364.655 2113.995 ;
        RECT 365.085 2113.715 365.365 2113.995 ;
        RECT 365.795 2113.715 366.075 2113.995 ;
        RECT 366.505 2113.715 366.785 2113.995 ;
        RECT 357.275 2113.005 357.555 2113.285 ;
        RECT 357.985 2113.005 358.265 2113.285 ;
        RECT 358.695 2113.005 358.975 2113.285 ;
        RECT 359.405 2113.005 359.685 2113.285 ;
        RECT 360.115 2113.005 360.395 2113.285 ;
        RECT 360.825 2113.005 361.105 2113.285 ;
        RECT 361.535 2113.005 361.815 2113.285 ;
        RECT 362.245 2113.005 362.525 2113.285 ;
        RECT 362.955 2113.005 363.235 2113.285 ;
        RECT 363.665 2113.005 363.945 2113.285 ;
        RECT 364.375 2113.005 364.655 2113.285 ;
        RECT 365.085 2113.005 365.365 2113.285 ;
        RECT 365.795 2113.005 366.075 2113.285 ;
        RECT 366.505 2113.005 366.785 2113.285 ;
        RECT 357.275 2112.295 357.555 2112.575 ;
        RECT 357.985 2112.295 358.265 2112.575 ;
        RECT 358.695 2112.295 358.975 2112.575 ;
        RECT 359.405 2112.295 359.685 2112.575 ;
        RECT 360.115 2112.295 360.395 2112.575 ;
        RECT 360.825 2112.295 361.105 2112.575 ;
        RECT 361.535 2112.295 361.815 2112.575 ;
        RECT 362.245 2112.295 362.525 2112.575 ;
        RECT 362.955 2112.295 363.235 2112.575 ;
        RECT 363.665 2112.295 363.945 2112.575 ;
        RECT 364.375 2112.295 364.655 2112.575 ;
        RECT 365.085 2112.295 365.365 2112.575 ;
        RECT 365.795 2112.295 366.075 2112.575 ;
        RECT 366.505 2112.295 366.785 2112.575 ;
        RECT 357.275 2111.585 357.555 2111.865 ;
        RECT 357.985 2111.585 358.265 2111.865 ;
        RECT 358.695 2111.585 358.975 2111.865 ;
        RECT 359.405 2111.585 359.685 2111.865 ;
        RECT 360.115 2111.585 360.395 2111.865 ;
        RECT 360.825 2111.585 361.105 2111.865 ;
        RECT 361.535 2111.585 361.815 2111.865 ;
        RECT 362.245 2111.585 362.525 2111.865 ;
        RECT 362.955 2111.585 363.235 2111.865 ;
        RECT 363.665 2111.585 363.945 2111.865 ;
        RECT 364.375 2111.585 364.655 2111.865 ;
        RECT 365.085 2111.585 365.365 2111.865 ;
        RECT 365.795 2111.585 366.075 2111.865 ;
        RECT 366.505 2111.585 366.785 2111.865 ;
        RECT 357.275 2110.875 357.555 2111.155 ;
        RECT 357.985 2110.875 358.265 2111.155 ;
        RECT 358.695 2110.875 358.975 2111.155 ;
        RECT 359.405 2110.875 359.685 2111.155 ;
        RECT 360.115 2110.875 360.395 2111.155 ;
        RECT 360.825 2110.875 361.105 2111.155 ;
        RECT 361.535 2110.875 361.815 2111.155 ;
        RECT 362.245 2110.875 362.525 2111.155 ;
        RECT 362.955 2110.875 363.235 2111.155 ;
        RECT 363.665 2110.875 363.945 2111.155 ;
        RECT 364.375 2110.875 364.655 2111.155 ;
        RECT 365.085 2110.875 365.365 2111.155 ;
        RECT 365.795 2110.875 366.075 2111.155 ;
        RECT 366.505 2110.875 366.785 2111.155 ;
        RECT 357.275 2110.165 357.555 2110.445 ;
        RECT 357.985 2110.165 358.265 2110.445 ;
        RECT 358.695 2110.165 358.975 2110.445 ;
        RECT 359.405 2110.165 359.685 2110.445 ;
        RECT 360.115 2110.165 360.395 2110.445 ;
        RECT 360.825 2110.165 361.105 2110.445 ;
        RECT 361.535 2110.165 361.815 2110.445 ;
        RECT 362.245 2110.165 362.525 2110.445 ;
        RECT 362.955 2110.165 363.235 2110.445 ;
        RECT 363.665 2110.165 363.945 2110.445 ;
        RECT 364.375 2110.165 364.655 2110.445 ;
        RECT 365.085 2110.165 365.365 2110.445 ;
        RECT 365.795 2110.165 366.075 2110.445 ;
        RECT 366.505 2110.165 366.785 2110.445 ;
        RECT 357.275 2109.455 357.555 2109.735 ;
        RECT 357.985 2109.455 358.265 2109.735 ;
        RECT 358.695 2109.455 358.975 2109.735 ;
        RECT 359.405 2109.455 359.685 2109.735 ;
        RECT 360.115 2109.455 360.395 2109.735 ;
        RECT 360.825 2109.455 361.105 2109.735 ;
        RECT 361.535 2109.455 361.815 2109.735 ;
        RECT 362.245 2109.455 362.525 2109.735 ;
        RECT 362.955 2109.455 363.235 2109.735 ;
        RECT 363.665 2109.455 363.945 2109.735 ;
        RECT 364.375 2109.455 364.655 2109.735 ;
        RECT 365.085 2109.455 365.365 2109.735 ;
        RECT 365.795 2109.455 366.075 2109.735 ;
        RECT 366.505 2109.455 366.785 2109.735 ;
        RECT 357.275 2108.745 357.555 2109.025 ;
        RECT 357.985 2108.745 358.265 2109.025 ;
        RECT 358.695 2108.745 358.975 2109.025 ;
        RECT 359.405 2108.745 359.685 2109.025 ;
        RECT 360.115 2108.745 360.395 2109.025 ;
        RECT 360.825 2108.745 361.105 2109.025 ;
        RECT 361.535 2108.745 361.815 2109.025 ;
        RECT 362.245 2108.745 362.525 2109.025 ;
        RECT 362.955 2108.745 363.235 2109.025 ;
        RECT 363.665 2108.745 363.945 2109.025 ;
        RECT 364.375 2108.745 364.655 2109.025 ;
        RECT 365.085 2108.745 365.365 2109.025 ;
        RECT 365.795 2108.745 366.075 2109.025 ;
        RECT 366.505 2108.745 366.785 2109.025 ;
        RECT 357.275 2108.035 357.555 2108.315 ;
        RECT 357.985 2108.035 358.265 2108.315 ;
        RECT 358.695 2108.035 358.975 2108.315 ;
        RECT 359.405 2108.035 359.685 2108.315 ;
        RECT 360.115 2108.035 360.395 2108.315 ;
        RECT 360.825 2108.035 361.105 2108.315 ;
        RECT 361.535 2108.035 361.815 2108.315 ;
        RECT 362.245 2108.035 362.525 2108.315 ;
        RECT 362.955 2108.035 363.235 2108.315 ;
        RECT 363.665 2108.035 363.945 2108.315 ;
        RECT 364.375 2108.035 364.655 2108.315 ;
        RECT 365.085 2108.035 365.365 2108.315 ;
        RECT 365.795 2108.035 366.075 2108.315 ;
        RECT 366.505 2108.035 366.785 2108.315 ;
        RECT 357.275 2107.325 357.555 2107.605 ;
        RECT 357.985 2107.325 358.265 2107.605 ;
        RECT 358.695 2107.325 358.975 2107.605 ;
        RECT 359.405 2107.325 359.685 2107.605 ;
        RECT 360.115 2107.325 360.395 2107.605 ;
        RECT 360.825 2107.325 361.105 2107.605 ;
        RECT 361.535 2107.325 361.815 2107.605 ;
        RECT 362.245 2107.325 362.525 2107.605 ;
        RECT 362.955 2107.325 363.235 2107.605 ;
        RECT 363.665 2107.325 363.945 2107.605 ;
        RECT 364.375 2107.325 364.655 2107.605 ;
        RECT 365.085 2107.325 365.365 2107.605 ;
        RECT 365.795 2107.325 366.075 2107.605 ;
        RECT 366.505 2107.325 366.785 2107.605 ;
        RECT 357.275 2106.615 357.555 2106.895 ;
        RECT 357.985 2106.615 358.265 2106.895 ;
        RECT 358.695 2106.615 358.975 2106.895 ;
        RECT 359.405 2106.615 359.685 2106.895 ;
        RECT 360.115 2106.615 360.395 2106.895 ;
        RECT 360.825 2106.615 361.105 2106.895 ;
        RECT 361.535 2106.615 361.815 2106.895 ;
        RECT 362.245 2106.615 362.525 2106.895 ;
        RECT 362.955 2106.615 363.235 2106.895 ;
        RECT 363.665 2106.615 363.945 2106.895 ;
        RECT 364.375 2106.615 364.655 2106.895 ;
        RECT 365.085 2106.615 365.365 2106.895 ;
        RECT 365.795 2106.615 366.075 2106.895 ;
        RECT 366.505 2106.615 366.785 2106.895 ;
        RECT 357.275 2105.905 357.555 2106.185 ;
        RECT 357.985 2105.905 358.265 2106.185 ;
        RECT 358.695 2105.905 358.975 2106.185 ;
        RECT 359.405 2105.905 359.685 2106.185 ;
        RECT 360.115 2105.905 360.395 2106.185 ;
        RECT 360.825 2105.905 361.105 2106.185 ;
        RECT 361.535 2105.905 361.815 2106.185 ;
        RECT 362.245 2105.905 362.525 2106.185 ;
        RECT 362.955 2105.905 363.235 2106.185 ;
        RECT 363.665 2105.905 363.945 2106.185 ;
        RECT 364.375 2105.905 364.655 2106.185 ;
        RECT 365.085 2105.905 365.365 2106.185 ;
        RECT 365.795 2105.905 366.075 2106.185 ;
        RECT 366.505 2105.905 366.785 2106.185 ;
        RECT 357.275 2105.195 357.555 2105.475 ;
        RECT 357.985 2105.195 358.265 2105.475 ;
        RECT 358.695 2105.195 358.975 2105.475 ;
        RECT 359.405 2105.195 359.685 2105.475 ;
        RECT 360.115 2105.195 360.395 2105.475 ;
        RECT 360.825 2105.195 361.105 2105.475 ;
        RECT 361.535 2105.195 361.815 2105.475 ;
        RECT 362.245 2105.195 362.525 2105.475 ;
        RECT 362.955 2105.195 363.235 2105.475 ;
        RECT 363.665 2105.195 363.945 2105.475 ;
        RECT 364.375 2105.195 364.655 2105.475 ;
        RECT 365.085 2105.195 365.365 2105.475 ;
        RECT 365.795 2105.195 366.075 2105.475 ;
        RECT 366.505 2105.195 366.785 2105.475 ;
        RECT 357.275 2104.485 357.555 2104.765 ;
        RECT 357.985 2104.485 358.265 2104.765 ;
        RECT 358.695 2104.485 358.975 2104.765 ;
        RECT 359.405 2104.485 359.685 2104.765 ;
        RECT 360.115 2104.485 360.395 2104.765 ;
        RECT 360.825 2104.485 361.105 2104.765 ;
        RECT 361.535 2104.485 361.815 2104.765 ;
        RECT 362.245 2104.485 362.525 2104.765 ;
        RECT 362.955 2104.485 363.235 2104.765 ;
        RECT 363.665 2104.485 363.945 2104.765 ;
        RECT 364.375 2104.485 364.655 2104.765 ;
        RECT 365.085 2104.485 365.365 2104.765 ;
        RECT 365.795 2104.485 366.075 2104.765 ;
        RECT 366.505 2104.485 366.785 2104.765 ;
        RECT 357.275 2100.185 357.555 2100.465 ;
        RECT 357.985 2100.185 358.265 2100.465 ;
        RECT 358.695 2100.185 358.975 2100.465 ;
        RECT 359.405 2100.185 359.685 2100.465 ;
        RECT 360.115 2100.185 360.395 2100.465 ;
        RECT 360.825 2100.185 361.105 2100.465 ;
        RECT 361.535 2100.185 361.815 2100.465 ;
        RECT 362.245 2100.185 362.525 2100.465 ;
        RECT 362.955 2100.185 363.235 2100.465 ;
        RECT 363.665 2100.185 363.945 2100.465 ;
        RECT 364.375 2100.185 364.655 2100.465 ;
        RECT 365.085 2100.185 365.365 2100.465 ;
        RECT 365.795 2100.185 366.075 2100.465 ;
        RECT 366.505 2100.185 366.785 2100.465 ;
        RECT 357.275 2099.475 357.555 2099.755 ;
        RECT 357.985 2099.475 358.265 2099.755 ;
        RECT 358.695 2099.475 358.975 2099.755 ;
        RECT 359.405 2099.475 359.685 2099.755 ;
        RECT 360.115 2099.475 360.395 2099.755 ;
        RECT 360.825 2099.475 361.105 2099.755 ;
        RECT 361.535 2099.475 361.815 2099.755 ;
        RECT 362.245 2099.475 362.525 2099.755 ;
        RECT 362.955 2099.475 363.235 2099.755 ;
        RECT 363.665 2099.475 363.945 2099.755 ;
        RECT 364.375 2099.475 364.655 2099.755 ;
        RECT 365.085 2099.475 365.365 2099.755 ;
        RECT 365.795 2099.475 366.075 2099.755 ;
        RECT 366.505 2099.475 366.785 2099.755 ;
        RECT 357.275 2098.765 357.555 2099.045 ;
        RECT 357.985 2098.765 358.265 2099.045 ;
        RECT 358.695 2098.765 358.975 2099.045 ;
        RECT 359.405 2098.765 359.685 2099.045 ;
        RECT 360.115 2098.765 360.395 2099.045 ;
        RECT 360.825 2098.765 361.105 2099.045 ;
        RECT 361.535 2098.765 361.815 2099.045 ;
        RECT 362.245 2098.765 362.525 2099.045 ;
        RECT 362.955 2098.765 363.235 2099.045 ;
        RECT 363.665 2098.765 363.945 2099.045 ;
        RECT 364.375 2098.765 364.655 2099.045 ;
        RECT 365.085 2098.765 365.365 2099.045 ;
        RECT 365.795 2098.765 366.075 2099.045 ;
        RECT 366.505 2098.765 366.785 2099.045 ;
        RECT 357.275 2098.055 357.555 2098.335 ;
        RECT 357.985 2098.055 358.265 2098.335 ;
        RECT 358.695 2098.055 358.975 2098.335 ;
        RECT 359.405 2098.055 359.685 2098.335 ;
        RECT 360.115 2098.055 360.395 2098.335 ;
        RECT 360.825 2098.055 361.105 2098.335 ;
        RECT 361.535 2098.055 361.815 2098.335 ;
        RECT 362.245 2098.055 362.525 2098.335 ;
        RECT 362.955 2098.055 363.235 2098.335 ;
        RECT 363.665 2098.055 363.945 2098.335 ;
        RECT 364.375 2098.055 364.655 2098.335 ;
        RECT 365.085 2098.055 365.365 2098.335 ;
        RECT 365.795 2098.055 366.075 2098.335 ;
        RECT 366.505 2098.055 366.785 2098.335 ;
        RECT 357.275 2097.345 357.555 2097.625 ;
        RECT 357.985 2097.345 358.265 2097.625 ;
        RECT 358.695 2097.345 358.975 2097.625 ;
        RECT 359.405 2097.345 359.685 2097.625 ;
        RECT 360.115 2097.345 360.395 2097.625 ;
        RECT 360.825 2097.345 361.105 2097.625 ;
        RECT 361.535 2097.345 361.815 2097.625 ;
        RECT 362.245 2097.345 362.525 2097.625 ;
        RECT 362.955 2097.345 363.235 2097.625 ;
        RECT 363.665 2097.345 363.945 2097.625 ;
        RECT 364.375 2097.345 364.655 2097.625 ;
        RECT 365.085 2097.345 365.365 2097.625 ;
        RECT 365.795 2097.345 366.075 2097.625 ;
        RECT 366.505 2097.345 366.785 2097.625 ;
        RECT 357.275 2096.635 357.555 2096.915 ;
        RECT 357.985 2096.635 358.265 2096.915 ;
        RECT 358.695 2096.635 358.975 2096.915 ;
        RECT 359.405 2096.635 359.685 2096.915 ;
        RECT 360.115 2096.635 360.395 2096.915 ;
        RECT 360.825 2096.635 361.105 2096.915 ;
        RECT 361.535 2096.635 361.815 2096.915 ;
        RECT 362.245 2096.635 362.525 2096.915 ;
        RECT 362.955 2096.635 363.235 2096.915 ;
        RECT 363.665 2096.635 363.945 2096.915 ;
        RECT 364.375 2096.635 364.655 2096.915 ;
        RECT 365.085 2096.635 365.365 2096.915 ;
        RECT 365.795 2096.635 366.075 2096.915 ;
        RECT 366.505 2096.635 366.785 2096.915 ;
        RECT 357.275 2095.925 357.555 2096.205 ;
        RECT 357.985 2095.925 358.265 2096.205 ;
        RECT 358.695 2095.925 358.975 2096.205 ;
        RECT 359.405 2095.925 359.685 2096.205 ;
        RECT 360.115 2095.925 360.395 2096.205 ;
        RECT 360.825 2095.925 361.105 2096.205 ;
        RECT 361.535 2095.925 361.815 2096.205 ;
        RECT 362.245 2095.925 362.525 2096.205 ;
        RECT 362.955 2095.925 363.235 2096.205 ;
        RECT 363.665 2095.925 363.945 2096.205 ;
        RECT 364.375 2095.925 364.655 2096.205 ;
        RECT 365.085 2095.925 365.365 2096.205 ;
        RECT 365.795 2095.925 366.075 2096.205 ;
        RECT 366.505 2095.925 366.785 2096.205 ;
        RECT 357.275 2095.215 357.555 2095.495 ;
        RECT 357.985 2095.215 358.265 2095.495 ;
        RECT 358.695 2095.215 358.975 2095.495 ;
        RECT 359.405 2095.215 359.685 2095.495 ;
        RECT 360.115 2095.215 360.395 2095.495 ;
        RECT 360.825 2095.215 361.105 2095.495 ;
        RECT 361.535 2095.215 361.815 2095.495 ;
        RECT 362.245 2095.215 362.525 2095.495 ;
        RECT 362.955 2095.215 363.235 2095.495 ;
        RECT 363.665 2095.215 363.945 2095.495 ;
        RECT 364.375 2095.215 364.655 2095.495 ;
        RECT 365.085 2095.215 365.365 2095.495 ;
        RECT 365.795 2095.215 366.075 2095.495 ;
        RECT 366.505 2095.215 366.785 2095.495 ;
        RECT 357.275 2094.505 357.555 2094.785 ;
        RECT 357.985 2094.505 358.265 2094.785 ;
        RECT 358.695 2094.505 358.975 2094.785 ;
        RECT 359.405 2094.505 359.685 2094.785 ;
        RECT 360.115 2094.505 360.395 2094.785 ;
        RECT 360.825 2094.505 361.105 2094.785 ;
        RECT 361.535 2094.505 361.815 2094.785 ;
        RECT 362.245 2094.505 362.525 2094.785 ;
        RECT 362.955 2094.505 363.235 2094.785 ;
        RECT 363.665 2094.505 363.945 2094.785 ;
        RECT 364.375 2094.505 364.655 2094.785 ;
        RECT 365.085 2094.505 365.365 2094.785 ;
        RECT 365.795 2094.505 366.075 2094.785 ;
        RECT 366.505 2094.505 366.785 2094.785 ;
        RECT 357.275 2093.795 357.555 2094.075 ;
        RECT 357.985 2093.795 358.265 2094.075 ;
        RECT 358.695 2093.795 358.975 2094.075 ;
        RECT 359.405 2093.795 359.685 2094.075 ;
        RECT 360.115 2093.795 360.395 2094.075 ;
        RECT 360.825 2093.795 361.105 2094.075 ;
        RECT 361.535 2093.795 361.815 2094.075 ;
        RECT 362.245 2093.795 362.525 2094.075 ;
        RECT 362.955 2093.795 363.235 2094.075 ;
        RECT 363.665 2093.795 363.945 2094.075 ;
        RECT 364.375 2093.795 364.655 2094.075 ;
        RECT 365.085 2093.795 365.365 2094.075 ;
        RECT 365.795 2093.795 366.075 2094.075 ;
        RECT 366.505 2093.795 366.785 2094.075 ;
        RECT 357.275 2093.085 357.555 2093.365 ;
        RECT 357.985 2093.085 358.265 2093.365 ;
        RECT 358.695 2093.085 358.975 2093.365 ;
        RECT 359.405 2093.085 359.685 2093.365 ;
        RECT 360.115 2093.085 360.395 2093.365 ;
        RECT 360.825 2093.085 361.105 2093.365 ;
        RECT 361.535 2093.085 361.815 2093.365 ;
        RECT 362.245 2093.085 362.525 2093.365 ;
        RECT 362.955 2093.085 363.235 2093.365 ;
        RECT 363.665 2093.085 363.945 2093.365 ;
        RECT 364.375 2093.085 364.655 2093.365 ;
        RECT 365.085 2093.085 365.365 2093.365 ;
        RECT 365.795 2093.085 366.075 2093.365 ;
        RECT 366.505 2093.085 366.785 2093.365 ;
        RECT 357.275 2092.375 357.555 2092.655 ;
        RECT 357.985 2092.375 358.265 2092.655 ;
        RECT 358.695 2092.375 358.975 2092.655 ;
        RECT 359.405 2092.375 359.685 2092.655 ;
        RECT 360.115 2092.375 360.395 2092.655 ;
        RECT 360.825 2092.375 361.105 2092.655 ;
        RECT 361.535 2092.375 361.815 2092.655 ;
        RECT 362.245 2092.375 362.525 2092.655 ;
        RECT 362.955 2092.375 363.235 2092.655 ;
        RECT 363.665 2092.375 363.945 2092.655 ;
        RECT 364.375 2092.375 364.655 2092.655 ;
        RECT 365.085 2092.375 365.365 2092.655 ;
        RECT 365.795 2092.375 366.075 2092.655 ;
        RECT 366.505 2092.375 366.785 2092.655 ;
        RECT 357.275 2091.665 357.555 2091.945 ;
        RECT 357.985 2091.665 358.265 2091.945 ;
        RECT 358.695 2091.665 358.975 2091.945 ;
        RECT 359.405 2091.665 359.685 2091.945 ;
        RECT 360.115 2091.665 360.395 2091.945 ;
        RECT 360.825 2091.665 361.105 2091.945 ;
        RECT 361.535 2091.665 361.815 2091.945 ;
        RECT 362.245 2091.665 362.525 2091.945 ;
        RECT 362.955 2091.665 363.235 2091.945 ;
        RECT 363.665 2091.665 363.945 2091.945 ;
        RECT 364.375 2091.665 364.655 2091.945 ;
        RECT 365.085 2091.665 365.365 2091.945 ;
        RECT 365.795 2091.665 366.075 2091.945 ;
        RECT 366.505 2091.665 366.785 2091.945 ;
        RECT 357.275 2090.955 357.555 2091.235 ;
        RECT 357.985 2090.955 358.265 2091.235 ;
        RECT 358.695 2090.955 358.975 2091.235 ;
        RECT 359.405 2090.955 359.685 2091.235 ;
        RECT 360.115 2090.955 360.395 2091.235 ;
        RECT 360.825 2090.955 361.105 2091.235 ;
        RECT 361.535 2090.955 361.815 2091.235 ;
        RECT 362.245 2090.955 362.525 2091.235 ;
        RECT 362.955 2090.955 363.235 2091.235 ;
        RECT 363.665 2090.955 363.945 2091.235 ;
        RECT 364.375 2090.955 364.655 2091.235 ;
        RECT 365.085 2090.955 365.365 2091.235 ;
        RECT 365.795 2090.955 366.075 2091.235 ;
        RECT 366.505 2090.955 366.785 2091.235 ;
        RECT 357.275 2088.335 357.555 2088.615 ;
        RECT 357.985 2088.335 358.265 2088.615 ;
        RECT 358.695 2088.335 358.975 2088.615 ;
        RECT 359.405 2088.335 359.685 2088.615 ;
        RECT 360.115 2088.335 360.395 2088.615 ;
        RECT 360.825 2088.335 361.105 2088.615 ;
        RECT 361.535 2088.335 361.815 2088.615 ;
        RECT 362.245 2088.335 362.525 2088.615 ;
        RECT 362.955 2088.335 363.235 2088.615 ;
        RECT 363.665 2088.335 363.945 2088.615 ;
        RECT 364.375 2088.335 364.655 2088.615 ;
        RECT 365.085 2088.335 365.365 2088.615 ;
        RECT 365.795 2088.335 366.075 2088.615 ;
        RECT 366.505 2088.335 366.785 2088.615 ;
        RECT 357.275 2087.625 357.555 2087.905 ;
        RECT 357.985 2087.625 358.265 2087.905 ;
        RECT 358.695 2087.625 358.975 2087.905 ;
        RECT 359.405 2087.625 359.685 2087.905 ;
        RECT 360.115 2087.625 360.395 2087.905 ;
        RECT 360.825 2087.625 361.105 2087.905 ;
        RECT 361.535 2087.625 361.815 2087.905 ;
        RECT 362.245 2087.625 362.525 2087.905 ;
        RECT 362.955 2087.625 363.235 2087.905 ;
        RECT 363.665 2087.625 363.945 2087.905 ;
        RECT 364.375 2087.625 364.655 2087.905 ;
        RECT 365.085 2087.625 365.365 2087.905 ;
        RECT 365.795 2087.625 366.075 2087.905 ;
        RECT 366.505 2087.625 366.785 2087.905 ;
        RECT 357.275 2086.915 357.555 2087.195 ;
        RECT 357.985 2086.915 358.265 2087.195 ;
        RECT 358.695 2086.915 358.975 2087.195 ;
        RECT 359.405 2086.915 359.685 2087.195 ;
        RECT 360.115 2086.915 360.395 2087.195 ;
        RECT 360.825 2086.915 361.105 2087.195 ;
        RECT 361.535 2086.915 361.815 2087.195 ;
        RECT 362.245 2086.915 362.525 2087.195 ;
        RECT 362.955 2086.915 363.235 2087.195 ;
        RECT 363.665 2086.915 363.945 2087.195 ;
        RECT 364.375 2086.915 364.655 2087.195 ;
        RECT 365.085 2086.915 365.365 2087.195 ;
        RECT 365.795 2086.915 366.075 2087.195 ;
        RECT 366.505 2086.915 366.785 2087.195 ;
        RECT 357.275 2086.205 357.555 2086.485 ;
        RECT 357.985 2086.205 358.265 2086.485 ;
        RECT 358.695 2086.205 358.975 2086.485 ;
        RECT 359.405 2086.205 359.685 2086.485 ;
        RECT 360.115 2086.205 360.395 2086.485 ;
        RECT 360.825 2086.205 361.105 2086.485 ;
        RECT 361.535 2086.205 361.815 2086.485 ;
        RECT 362.245 2086.205 362.525 2086.485 ;
        RECT 362.955 2086.205 363.235 2086.485 ;
        RECT 363.665 2086.205 363.945 2086.485 ;
        RECT 364.375 2086.205 364.655 2086.485 ;
        RECT 365.085 2086.205 365.365 2086.485 ;
        RECT 365.795 2086.205 366.075 2086.485 ;
        RECT 366.505 2086.205 366.785 2086.485 ;
        RECT 357.275 2085.495 357.555 2085.775 ;
        RECT 357.985 2085.495 358.265 2085.775 ;
        RECT 358.695 2085.495 358.975 2085.775 ;
        RECT 359.405 2085.495 359.685 2085.775 ;
        RECT 360.115 2085.495 360.395 2085.775 ;
        RECT 360.825 2085.495 361.105 2085.775 ;
        RECT 361.535 2085.495 361.815 2085.775 ;
        RECT 362.245 2085.495 362.525 2085.775 ;
        RECT 362.955 2085.495 363.235 2085.775 ;
        RECT 363.665 2085.495 363.945 2085.775 ;
        RECT 364.375 2085.495 364.655 2085.775 ;
        RECT 365.085 2085.495 365.365 2085.775 ;
        RECT 365.795 2085.495 366.075 2085.775 ;
        RECT 366.505 2085.495 366.785 2085.775 ;
        RECT 357.275 2084.785 357.555 2085.065 ;
        RECT 357.985 2084.785 358.265 2085.065 ;
        RECT 358.695 2084.785 358.975 2085.065 ;
        RECT 359.405 2084.785 359.685 2085.065 ;
        RECT 360.115 2084.785 360.395 2085.065 ;
        RECT 360.825 2084.785 361.105 2085.065 ;
        RECT 361.535 2084.785 361.815 2085.065 ;
        RECT 362.245 2084.785 362.525 2085.065 ;
        RECT 362.955 2084.785 363.235 2085.065 ;
        RECT 363.665 2084.785 363.945 2085.065 ;
        RECT 364.375 2084.785 364.655 2085.065 ;
        RECT 365.085 2084.785 365.365 2085.065 ;
        RECT 365.795 2084.785 366.075 2085.065 ;
        RECT 366.505 2084.785 366.785 2085.065 ;
        RECT 357.275 2084.075 357.555 2084.355 ;
        RECT 357.985 2084.075 358.265 2084.355 ;
        RECT 358.695 2084.075 358.975 2084.355 ;
        RECT 359.405 2084.075 359.685 2084.355 ;
        RECT 360.115 2084.075 360.395 2084.355 ;
        RECT 360.825 2084.075 361.105 2084.355 ;
        RECT 361.535 2084.075 361.815 2084.355 ;
        RECT 362.245 2084.075 362.525 2084.355 ;
        RECT 362.955 2084.075 363.235 2084.355 ;
        RECT 363.665 2084.075 363.945 2084.355 ;
        RECT 364.375 2084.075 364.655 2084.355 ;
        RECT 365.085 2084.075 365.365 2084.355 ;
        RECT 365.795 2084.075 366.075 2084.355 ;
        RECT 366.505 2084.075 366.785 2084.355 ;
        RECT 357.275 2083.365 357.555 2083.645 ;
        RECT 357.985 2083.365 358.265 2083.645 ;
        RECT 358.695 2083.365 358.975 2083.645 ;
        RECT 359.405 2083.365 359.685 2083.645 ;
        RECT 360.115 2083.365 360.395 2083.645 ;
        RECT 360.825 2083.365 361.105 2083.645 ;
        RECT 361.535 2083.365 361.815 2083.645 ;
        RECT 362.245 2083.365 362.525 2083.645 ;
        RECT 362.955 2083.365 363.235 2083.645 ;
        RECT 363.665 2083.365 363.945 2083.645 ;
        RECT 364.375 2083.365 364.655 2083.645 ;
        RECT 365.085 2083.365 365.365 2083.645 ;
        RECT 365.795 2083.365 366.075 2083.645 ;
        RECT 366.505 2083.365 366.785 2083.645 ;
        RECT 357.275 2082.655 357.555 2082.935 ;
        RECT 357.985 2082.655 358.265 2082.935 ;
        RECT 358.695 2082.655 358.975 2082.935 ;
        RECT 359.405 2082.655 359.685 2082.935 ;
        RECT 360.115 2082.655 360.395 2082.935 ;
        RECT 360.825 2082.655 361.105 2082.935 ;
        RECT 361.535 2082.655 361.815 2082.935 ;
        RECT 362.245 2082.655 362.525 2082.935 ;
        RECT 362.955 2082.655 363.235 2082.935 ;
        RECT 363.665 2082.655 363.945 2082.935 ;
        RECT 364.375 2082.655 364.655 2082.935 ;
        RECT 365.085 2082.655 365.365 2082.935 ;
        RECT 365.795 2082.655 366.075 2082.935 ;
        RECT 366.505 2082.655 366.785 2082.935 ;
        RECT 357.275 2081.945 357.555 2082.225 ;
        RECT 357.985 2081.945 358.265 2082.225 ;
        RECT 358.695 2081.945 358.975 2082.225 ;
        RECT 359.405 2081.945 359.685 2082.225 ;
        RECT 360.115 2081.945 360.395 2082.225 ;
        RECT 360.825 2081.945 361.105 2082.225 ;
        RECT 361.535 2081.945 361.815 2082.225 ;
        RECT 362.245 2081.945 362.525 2082.225 ;
        RECT 362.955 2081.945 363.235 2082.225 ;
        RECT 363.665 2081.945 363.945 2082.225 ;
        RECT 364.375 2081.945 364.655 2082.225 ;
        RECT 365.085 2081.945 365.365 2082.225 ;
        RECT 365.795 2081.945 366.075 2082.225 ;
        RECT 366.505 2081.945 366.785 2082.225 ;
        RECT 357.275 2081.235 357.555 2081.515 ;
        RECT 357.985 2081.235 358.265 2081.515 ;
        RECT 358.695 2081.235 358.975 2081.515 ;
        RECT 359.405 2081.235 359.685 2081.515 ;
        RECT 360.115 2081.235 360.395 2081.515 ;
        RECT 360.825 2081.235 361.105 2081.515 ;
        RECT 361.535 2081.235 361.815 2081.515 ;
        RECT 362.245 2081.235 362.525 2081.515 ;
        RECT 362.955 2081.235 363.235 2081.515 ;
        RECT 363.665 2081.235 363.945 2081.515 ;
        RECT 364.375 2081.235 364.655 2081.515 ;
        RECT 365.085 2081.235 365.365 2081.515 ;
        RECT 365.795 2081.235 366.075 2081.515 ;
        RECT 366.505 2081.235 366.785 2081.515 ;
        RECT 357.275 2080.525 357.555 2080.805 ;
        RECT 357.985 2080.525 358.265 2080.805 ;
        RECT 358.695 2080.525 358.975 2080.805 ;
        RECT 359.405 2080.525 359.685 2080.805 ;
        RECT 360.115 2080.525 360.395 2080.805 ;
        RECT 360.825 2080.525 361.105 2080.805 ;
        RECT 361.535 2080.525 361.815 2080.805 ;
        RECT 362.245 2080.525 362.525 2080.805 ;
        RECT 362.955 2080.525 363.235 2080.805 ;
        RECT 363.665 2080.525 363.945 2080.805 ;
        RECT 364.375 2080.525 364.655 2080.805 ;
        RECT 365.085 2080.525 365.365 2080.805 ;
        RECT 365.795 2080.525 366.075 2080.805 ;
        RECT 366.505 2080.525 366.785 2080.805 ;
        RECT 357.275 2079.815 357.555 2080.095 ;
        RECT 357.985 2079.815 358.265 2080.095 ;
        RECT 358.695 2079.815 358.975 2080.095 ;
        RECT 359.405 2079.815 359.685 2080.095 ;
        RECT 360.115 2079.815 360.395 2080.095 ;
        RECT 360.825 2079.815 361.105 2080.095 ;
        RECT 361.535 2079.815 361.815 2080.095 ;
        RECT 362.245 2079.815 362.525 2080.095 ;
        RECT 362.955 2079.815 363.235 2080.095 ;
        RECT 363.665 2079.815 363.945 2080.095 ;
        RECT 364.375 2079.815 364.655 2080.095 ;
        RECT 365.085 2079.815 365.365 2080.095 ;
        RECT 365.795 2079.815 366.075 2080.095 ;
        RECT 366.505 2079.815 366.785 2080.095 ;
        RECT 357.275 2079.105 357.555 2079.385 ;
        RECT 357.985 2079.105 358.265 2079.385 ;
        RECT 358.695 2079.105 358.975 2079.385 ;
        RECT 359.405 2079.105 359.685 2079.385 ;
        RECT 360.115 2079.105 360.395 2079.385 ;
        RECT 360.825 2079.105 361.105 2079.385 ;
        RECT 361.535 2079.105 361.815 2079.385 ;
        RECT 362.245 2079.105 362.525 2079.385 ;
        RECT 362.955 2079.105 363.235 2079.385 ;
        RECT 363.665 2079.105 363.945 2079.385 ;
        RECT 364.375 2079.105 364.655 2079.385 ;
        RECT 365.085 2079.105 365.365 2079.385 ;
        RECT 365.795 2079.105 366.075 2079.385 ;
        RECT 366.505 2079.105 366.785 2079.385 ;
        RECT 357.330 2075.190 357.610 2075.470 ;
        RECT 358.040 2075.190 358.320 2075.470 ;
        RECT 358.750 2075.190 359.030 2075.470 ;
        RECT 359.460 2075.190 359.740 2075.470 ;
        RECT 360.170 2075.190 360.450 2075.470 ;
        RECT 360.880 2075.190 361.160 2075.470 ;
        RECT 361.590 2075.190 361.870 2075.470 ;
        RECT 362.300 2075.190 362.580 2075.470 ;
        RECT 363.010 2075.190 363.290 2075.470 ;
        RECT 363.720 2075.190 364.000 2075.470 ;
        RECT 364.430 2075.190 364.710 2075.470 ;
        RECT 365.140 2075.190 365.420 2075.470 ;
        RECT 365.850 2075.190 366.130 2075.470 ;
        RECT 366.560 2075.190 366.840 2075.470 ;
        RECT 357.330 2074.480 357.610 2074.760 ;
        RECT 358.040 2074.480 358.320 2074.760 ;
        RECT 358.750 2074.480 359.030 2074.760 ;
        RECT 359.460 2074.480 359.740 2074.760 ;
        RECT 360.170 2074.480 360.450 2074.760 ;
        RECT 360.880 2074.480 361.160 2074.760 ;
        RECT 361.590 2074.480 361.870 2074.760 ;
        RECT 362.300 2074.480 362.580 2074.760 ;
        RECT 363.010 2074.480 363.290 2074.760 ;
        RECT 363.720 2074.480 364.000 2074.760 ;
        RECT 364.430 2074.480 364.710 2074.760 ;
        RECT 365.140 2074.480 365.420 2074.760 ;
        RECT 365.850 2074.480 366.130 2074.760 ;
        RECT 366.560 2074.480 366.840 2074.760 ;
        RECT 357.330 2073.770 357.610 2074.050 ;
        RECT 358.040 2073.770 358.320 2074.050 ;
        RECT 358.750 2073.770 359.030 2074.050 ;
        RECT 359.460 2073.770 359.740 2074.050 ;
        RECT 360.170 2073.770 360.450 2074.050 ;
        RECT 360.880 2073.770 361.160 2074.050 ;
        RECT 361.590 2073.770 361.870 2074.050 ;
        RECT 362.300 2073.770 362.580 2074.050 ;
        RECT 363.010 2073.770 363.290 2074.050 ;
        RECT 363.720 2073.770 364.000 2074.050 ;
        RECT 364.430 2073.770 364.710 2074.050 ;
        RECT 365.140 2073.770 365.420 2074.050 ;
        RECT 365.850 2073.770 366.130 2074.050 ;
        RECT 366.560 2073.770 366.840 2074.050 ;
        RECT 357.330 2073.060 357.610 2073.340 ;
        RECT 358.040 2073.060 358.320 2073.340 ;
        RECT 358.750 2073.060 359.030 2073.340 ;
        RECT 359.460 2073.060 359.740 2073.340 ;
        RECT 360.170 2073.060 360.450 2073.340 ;
        RECT 360.880 2073.060 361.160 2073.340 ;
        RECT 361.590 2073.060 361.870 2073.340 ;
        RECT 362.300 2073.060 362.580 2073.340 ;
        RECT 363.010 2073.060 363.290 2073.340 ;
        RECT 363.720 2073.060 364.000 2073.340 ;
        RECT 364.430 2073.060 364.710 2073.340 ;
        RECT 365.140 2073.060 365.420 2073.340 ;
        RECT 365.850 2073.060 366.130 2073.340 ;
        RECT 366.560 2073.060 366.840 2073.340 ;
        RECT 357.330 2072.350 357.610 2072.630 ;
        RECT 358.040 2072.350 358.320 2072.630 ;
        RECT 358.750 2072.350 359.030 2072.630 ;
        RECT 359.460 2072.350 359.740 2072.630 ;
        RECT 360.170 2072.350 360.450 2072.630 ;
        RECT 360.880 2072.350 361.160 2072.630 ;
        RECT 361.590 2072.350 361.870 2072.630 ;
        RECT 362.300 2072.350 362.580 2072.630 ;
        RECT 363.010 2072.350 363.290 2072.630 ;
        RECT 363.720 2072.350 364.000 2072.630 ;
        RECT 364.430 2072.350 364.710 2072.630 ;
        RECT 365.140 2072.350 365.420 2072.630 ;
        RECT 365.850 2072.350 366.130 2072.630 ;
        RECT 366.560 2072.350 366.840 2072.630 ;
        RECT 357.330 2071.640 357.610 2071.920 ;
        RECT 358.040 2071.640 358.320 2071.920 ;
        RECT 358.750 2071.640 359.030 2071.920 ;
        RECT 359.460 2071.640 359.740 2071.920 ;
        RECT 360.170 2071.640 360.450 2071.920 ;
        RECT 360.880 2071.640 361.160 2071.920 ;
        RECT 361.590 2071.640 361.870 2071.920 ;
        RECT 362.300 2071.640 362.580 2071.920 ;
        RECT 363.010 2071.640 363.290 2071.920 ;
        RECT 363.720 2071.640 364.000 2071.920 ;
        RECT 364.430 2071.640 364.710 2071.920 ;
        RECT 365.140 2071.640 365.420 2071.920 ;
        RECT 365.850 2071.640 366.130 2071.920 ;
        RECT 366.560 2071.640 366.840 2071.920 ;
        RECT 357.330 2070.930 357.610 2071.210 ;
        RECT 358.040 2070.930 358.320 2071.210 ;
        RECT 358.750 2070.930 359.030 2071.210 ;
        RECT 359.460 2070.930 359.740 2071.210 ;
        RECT 360.170 2070.930 360.450 2071.210 ;
        RECT 360.880 2070.930 361.160 2071.210 ;
        RECT 361.590 2070.930 361.870 2071.210 ;
        RECT 362.300 2070.930 362.580 2071.210 ;
        RECT 363.010 2070.930 363.290 2071.210 ;
        RECT 363.720 2070.930 364.000 2071.210 ;
        RECT 364.430 2070.930 364.710 2071.210 ;
        RECT 365.140 2070.930 365.420 2071.210 ;
        RECT 365.850 2070.930 366.130 2071.210 ;
        RECT 366.560 2070.930 366.840 2071.210 ;
        RECT 357.330 2070.220 357.610 2070.500 ;
        RECT 358.040 2070.220 358.320 2070.500 ;
        RECT 358.750 2070.220 359.030 2070.500 ;
        RECT 359.460 2070.220 359.740 2070.500 ;
        RECT 360.170 2070.220 360.450 2070.500 ;
        RECT 360.880 2070.220 361.160 2070.500 ;
        RECT 361.590 2070.220 361.870 2070.500 ;
        RECT 362.300 2070.220 362.580 2070.500 ;
        RECT 363.010 2070.220 363.290 2070.500 ;
        RECT 363.720 2070.220 364.000 2070.500 ;
        RECT 364.430 2070.220 364.710 2070.500 ;
        RECT 365.140 2070.220 365.420 2070.500 ;
        RECT 365.850 2070.220 366.130 2070.500 ;
        RECT 366.560 2070.220 366.840 2070.500 ;
        RECT 357.330 2069.510 357.610 2069.790 ;
        RECT 358.040 2069.510 358.320 2069.790 ;
        RECT 358.750 2069.510 359.030 2069.790 ;
        RECT 359.460 2069.510 359.740 2069.790 ;
        RECT 360.170 2069.510 360.450 2069.790 ;
        RECT 360.880 2069.510 361.160 2069.790 ;
        RECT 361.590 2069.510 361.870 2069.790 ;
        RECT 362.300 2069.510 362.580 2069.790 ;
        RECT 363.010 2069.510 363.290 2069.790 ;
        RECT 363.720 2069.510 364.000 2069.790 ;
        RECT 364.430 2069.510 364.710 2069.790 ;
        RECT 365.140 2069.510 365.420 2069.790 ;
        RECT 365.850 2069.510 366.130 2069.790 ;
        RECT 366.560 2069.510 366.840 2069.790 ;
        RECT 357.330 2068.800 357.610 2069.080 ;
        RECT 358.040 2068.800 358.320 2069.080 ;
        RECT 358.750 2068.800 359.030 2069.080 ;
        RECT 359.460 2068.800 359.740 2069.080 ;
        RECT 360.170 2068.800 360.450 2069.080 ;
        RECT 360.880 2068.800 361.160 2069.080 ;
        RECT 361.590 2068.800 361.870 2069.080 ;
        RECT 362.300 2068.800 362.580 2069.080 ;
        RECT 363.010 2068.800 363.290 2069.080 ;
        RECT 363.720 2068.800 364.000 2069.080 ;
        RECT 364.430 2068.800 364.710 2069.080 ;
        RECT 365.140 2068.800 365.420 2069.080 ;
        RECT 365.850 2068.800 366.130 2069.080 ;
        RECT 366.560 2068.800 366.840 2069.080 ;
        RECT 357.330 2068.090 357.610 2068.370 ;
        RECT 358.040 2068.090 358.320 2068.370 ;
        RECT 358.750 2068.090 359.030 2068.370 ;
        RECT 359.460 2068.090 359.740 2068.370 ;
        RECT 360.170 2068.090 360.450 2068.370 ;
        RECT 360.880 2068.090 361.160 2068.370 ;
        RECT 361.590 2068.090 361.870 2068.370 ;
        RECT 362.300 2068.090 362.580 2068.370 ;
        RECT 363.010 2068.090 363.290 2068.370 ;
        RECT 363.720 2068.090 364.000 2068.370 ;
        RECT 364.430 2068.090 364.710 2068.370 ;
        RECT 365.140 2068.090 365.420 2068.370 ;
        RECT 365.850 2068.090 366.130 2068.370 ;
        RECT 366.560 2068.090 366.840 2068.370 ;
        RECT 357.330 2067.380 357.610 2067.660 ;
        RECT 358.040 2067.380 358.320 2067.660 ;
        RECT 358.750 2067.380 359.030 2067.660 ;
        RECT 359.460 2067.380 359.740 2067.660 ;
        RECT 360.170 2067.380 360.450 2067.660 ;
        RECT 360.880 2067.380 361.160 2067.660 ;
        RECT 361.590 2067.380 361.870 2067.660 ;
        RECT 362.300 2067.380 362.580 2067.660 ;
        RECT 363.010 2067.380 363.290 2067.660 ;
        RECT 363.720 2067.380 364.000 2067.660 ;
        RECT 364.430 2067.380 364.710 2067.660 ;
        RECT 365.140 2067.380 365.420 2067.660 ;
        RECT 365.850 2067.380 366.130 2067.660 ;
        RECT 366.560 2067.380 366.840 2067.660 ;
        RECT 357.330 2066.670 357.610 2066.950 ;
        RECT 358.040 2066.670 358.320 2066.950 ;
        RECT 358.750 2066.670 359.030 2066.950 ;
        RECT 359.460 2066.670 359.740 2066.950 ;
        RECT 360.170 2066.670 360.450 2066.950 ;
        RECT 360.880 2066.670 361.160 2066.950 ;
        RECT 361.590 2066.670 361.870 2066.950 ;
        RECT 362.300 2066.670 362.580 2066.950 ;
        RECT 363.010 2066.670 363.290 2066.950 ;
        RECT 363.720 2066.670 364.000 2066.950 ;
        RECT 364.430 2066.670 364.710 2066.950 ;
        RECT 365.140 2066.670 365.420 2066.950 ;
        RECT 365.850 2066.670 366.130 2066.950 ;
        RECT 366.560 2066.670 366.840 2066.950 ;
        RECT 3512.200 2023.050 3512.480 2023.330 ;
        RECT 3512.910 2023.050 3513.190 2023.330 ;
        RECT 3513.620 2023.050 3513.900 2023.330 ;
        RECT 3514.330 2023.050 3514.610 2023.330 ;
        RECT 3515.040 2023.050 3515.320 2023.330 ;
        RECT 3515.750 2023.050 3516.030 2023.330 ;
        RECT 3516.460 2023.050 3516.740 2023.330 ;
        RECT 3517.170 2023.050 3517.450 2023.330 ;
        RECT 3517.880 2023.050 3518.160 2023.330 ;
        RECT 3518.590 2023.050 3518.870 2023.330 ;
        RECT 3519.300 2023.050 3519.580 2023.330 ;
        RECT 3520.010 2023.050 3520.290 2023.330 ;
        RECT 3520.720 2023.050 3521.000 2023.330 ;
        RECT 3521.430 2023.050 3521.710 2023.330 ;
        RECT 3512.200 2022.340 3512.480 2022.620 ;
        RECT 3512.910 2022.340 3513.190 2022.620 ;
        RECT 3513.620 2022.340 3513.900 2022.620 ;
        RECT 3514.330 2022.340 3514.610 2022.620 ;
        RECT 3515.040 2022.340 3515.320 2022.620 ;
        RECT 3515.750 2022.340 3516.030 2022.620 ;
        RECT 3516.460 2022.340 3516.740 2022.620 ;
        RECT 3517.170 2022.340 3517.450 2022.620 ;
        RECT 3517.880 2022.340 3518.160 2022.620 ;
        RECT 3518.590 2022.340 3518.870 2022.620 ;
        RECT 3519.300 2022.340 3519.580 2022.620 ;
        RECT 3520.010 2022.340 3520.290 2022.620 ;
        RECT 3520.720 2022.340 3521.000 2022.620 ;
        RECT 3521.430 2022.340 3521.710 2022.620 ;
        RECT 3512.200 2021.630 3512.480 2021.910 ;
        RECT 3512.910 2021.630 3513.190 2021.910 ;
        RECT 3513.620 2021.630 3513.900 2021.910 ;
        RECT 3514.330 2021.630 3514.610 2021.910 ;
        RECT 3515.040 2021.630 3515.320 2021.910 ;
        RECT 3515.750 2021.630 3516.030 2021.910 ;
        RECT 3516.460 2021.630 3516.740 2021.910 ;
        RECT 3517.170 2021.630 3517.450 2021.910 ;
        RECT 3517.880 2021.630 3518.160 2021.910 ;
        RECT 3518.590 2021.630 3518.870 2021.910 ;
        RECT 3519.300 2021.630 3519.580 2021.910 ;
        RECT 3520.010 2021.630 3520.290 2021.910 ;
        RECT 3520.720 2021.630 3521.000 2021.910 ;
        RECT 3521.430 2021.630 3521.710 2021.910 ;
        RECT 3512.200 2020.920 3512.480 2021.200 ;
        RECT 3512.910 2020.920 3513.190 2021.200 ;
        RECT 3513.620 2020.920 3513.900 2021.200 ;
        RECT 3514.330 2020.920 3514.610 2021.200 ;
        RECT 3515.040 2020.920 3515.320 2021.200 ;
        RECT 3515.750 2020.920 3516.030 2021.200 ;
        RECT 3516.460 2020.920 3516.740 2021.200 ;
        RECT 3517.170 2020.920 3517.450 2021.200 ;
        RECT 3517.880 2020.920 3518.160 2021.200 ;
        RECT 3518.590 2020.920 3518.870 2021.200 ;
        RECT 3519.300 2020.920 3519.580 2021.200 ;
        RECT 3520.010 2020.920 3520.290 2021.200 ;
        RECT 3520.720 2020.920 3521.000 2021.200 ;
        RECT 3521.430 2020.920 3521.710 2021.200 ;
        RECT 3512.200 2020.210 3512.480 2020.490 ;
        RECT 3512.910 2020.210 3513.190 2020.490 ;
        RECT 3513.620 2020.210 3513.900 2020.490 ;
        RECT 3514.330 2020.210 3514.610 2020.490 ;
        RECT 3515.040 2020.210 3515.320 2020.490 ;
        RECT 3515.750 2020.210 3516.030 2020.490 ;
        RECT 3516.460 2020.210 3516.740 2020.490 ;
        RECT 3517.170 2020.210 3517.450 2020.490 ;
        RECT 3517.880 2020.210 3518.160 2020.490 ;
        RECT 3518.590 2020.210 3518.870 2020.490 ;
        RECT 3519.300 2020.210 3519.580 2020.490 ;
        RECT 3520.010 2020.210 3520.290 2020.490 ;
        RECT 3520.720 2020.210 3521.000 2020.490 ;
        RECT 3521.430 2020.210 3521.710 2020.490 ;
        RECT 3512.200 2019.500 3512.480 2019.780 ;
        RECT 3512.910 2019.500 3513.190 2019.780 ;
        RECT 3513.620 2019.500 3513.900 2019.780 ;
        RECT 3514.330 2019.500 3514.610 2019.780 ;
        RECT 3515.040 2019.500 3515.320 2019.780 ;
        RECT 3515.750 2019.500 3516.030 2019.780 ;
        RECT 3516.460 2019.500 3516.740 2019.780 ;
        RECT 3517.170 2019.500 3517.450 2019.780 ;
        RECT 3517.880 2019.500 3518.160 2019.780 ;
        RECT 3518.590 2019.500 3518.870 2019.780 ;
        RECT 3519.300 2019.500 3519.580 2019.780 ;
        RECT 3520.010 2019.500 3520.290 2019.780 ;
        RECT 3520.720 2019.500 3521.000 2019.780 ;
        RECT 3521.430 2019.500 3521.710 2019.780 ;
        RECT 3512.200 2018.790 3512.480 2019.070 ;
        RECT 3512.910 2018.790 3513.190 2019.070 ;
        RECT 3513.620 2018.790 3513.900 2019.070 ;
        RECT 3514.330 2018.790 3514.610 2019.070 ;
        RECT 3515.040 2018.790 3515.320 2019.070 ;
        RECT 3515.750 2018.790 3516.030 2019.070 ;
        RECT 3516.460 2018.790 3516.740 2019.070 ;
        RECT 3517.170 2018.790 3517.450 2019.070 ;
        RECT 3517.880 2018.790 3518.160 2019.070 ;
        RECT 3518.590 2018.790 3518.870 2019.070 ;
        RECT 3519.300 2018.790 3519.580 2019.070 ;
        RECT 3520.010 2018.790 3520.290 2019.070 ;
        RECT 3520.720 2018.790 3521.000 2019.070 ;
        RECT 3521.430 2018.790 3521.710 2019.070 ;
        RECT 3512.200 2018.080 3512.480 2018.360 ;
        RECT 3512.910 2018.080 3513.190 2018.360 ;
        RECT 3513.620 2018.080 3513.900 2018.360 ;
        RECT 3514.330 2018.080 3514.610 2018.360 ;
        RECT 3515.040 2018.080 3515.320 2018.360 ;
        RECT 3515.750 2018.080 3516.030 2018.360 ;
        RECT 3516.460 2018.080 3516.740 2018.360 ;
        RECT 3517.170 2018.080 3517.450 2018.360 ;
        RECT 3517.880 2018.080 3518.160 2018.360 ;
        RECT 3518.590 2018.080 3518.870 2018.360 ;
        RECT 3519.300 2018.080 3519.580 2018.360 ;
        RECT 3520.010 2018.080 3520.290 2018.360 ;
        RECT 3520.720 2018.080 3521.000 2018.360 ;
        RECT 3521.430 2018.080 3521.710 2018.360 ;
        RECT 3512.200 2017.370 3512.480 2017.650 ;
        RECT 3512.910 2017.370 3513.190 2017.650 ;
        RECT 3513.620 2017.370 3513.900 2017.650 ;
        RECT 3514.330 2017.370 3514.610 2017.650 ;
        RECT 3515.040 2017.370 3515.320 2017.650 ;
        RECT 3515.750 2017.370 3516.030 2017.650 ;
        RECT 3516.460 2017.370 3516.740 2017.650 ;
        RECT 3517.170 2017.370 3517.450 2017.650 ;
        RECT 3517.880 2017.370 3518.160 2017.650 ;
        RECT 3518.590 2017.370 3518.870 2017.650 ;
        RECT 3519.300 2017.370 3519.580 2017.650 ;
        RECT 3520.010 2017.370 3520.290 2017.650 ;
        RECT 3520.720 2017.370 3521.000 2017.650 ;
        RECT 3521.430 2017.370 3521.710 2017.650 ;
        RECT 3512.200 2016.660 3512.480 2016.940 ;
        RECT 3512.910 2016.660 3513.190 2016.940 ;
        RECT 3513.620 2016.660 3513.900 2016.940 ;
        RECT 3514.330 2016.660 3514.610 2016.940 ;
        RECT 3515.040 2016.660 3515.320 2016.940 ;
        RECT 3515.750 2016.660 3516.030 2016.940 ;
        RECT 3516.460 2016.660 3516.740 2016.940 ;
        RECT 3517.170 2016.660 3517.450 2016.940 ;
        RECT 3517.880 2016.660 3518.160 2016.940 ;
        RECT 3518.590 2016.660 3518.870 2016.940 ;
        RECT 3519.300 2016.660 3519.580 2016.940 ;
        RECT 3520.010 2016.660 3520.290 2016.940 ;
        RECT 3520.720 2016.660 3521.000 2016.940 ;
        RECT 3521.430 2016.660 3521.710 2016.940 ;
        RECT 3512.200 2015.950 3512.480 2016.230 ;
        RECT 3512.910 2015.950 3513.190 2016.230 ;
        RECT 3513.620 2015.950 3513.900 2016.230 ;
        RECT 3514.330 2015.950 3514.610 2016.230 ;
        RECT 3515.040 2015.950 3515.320 2016.230 ;
        RECT 3515.750 2015.950 3516.030 2016.230 ;
        RECT 3516.460 2015.950 3516.740 2016.230 ;
        RECT 3517.170 2015.950 3517.450 2016.230 ;
        RECT 3517.880 2015.950 3518.160 2016.230 ;
        RECT 3518.590 2015.950 3518.870 2016.230 ;
        RECT 3519.300 2015.950 3519.580 2016.230 ;
        RECT 3520.010 2015.950 3520.290 2016.230 ;
        RECT 3520.720 2015.950 3521.000 2016.230 ;
        RECT 3521.430 2015.950 3521.710 2016.230 ;
        RECT 3512.200 2015.240 3512.480 2015.520 ;
        RECT 3512.910 2015.240 3513.190 2015.520 ;
        RECT 3513.620 2015.240 3513.900 2015.520 ;
        RECT 3514.330 2015.240 3514.610 2015.520 ;
        RECT 3515.040 2015.240 3515.320 2015.520 ;
        RECT 3515.750 2015.240 3516.030 2015.520 ;
        RECT 3516.460 2015.240 3516.740 2015.520 ;
        RECT 3517.170 2015.240 3517.450 2015.520 ;
        RECT 3517.880 2015.240 3518.160 2015.520 ;
        RECT 3518.590 2015.240 3518.870 2015.520 ;
        RECT 3519.300 2015.240 3519.580 2015.520 ;
        RECT 3520.010 2015.240 3520.290 2015.520 ;
        RECT 3520.720 2015.240 3521.000 2015.520 ;
        RECT 3521.430 2015.240 3521.710 2015.520 ;
        RECT 3512.200 2014.530 3512.480 2014.810 ;
        RECT 3512.910 2014.530 3513.190 2014.810 ;
        RECT 3513.620 2014.530 3513.900 2014.810 ;
        RECT 3514.330 2014.530 3514.610 2014.810 ;
        RECT 3515.040 2014.530 3515.320 2014.810 ;
        RECT 3515.750 2014.530 3516.030 2014.810 ;
        RECT 3516.460 2014.530 3516.740 2014.810 ;
        RECT 3517.170 2014.530 3517.450 2014.810 ;
        RECT 3517.880 2014.530 3518.160 2014.810 ;
        RECT 3518.590 2014.530 3518.870 2014.810 ;
        RECT 3519.300 2014.530 3519.580 2014.810 ;
        RECT 3520.010 2014.530 3520.290 2014.810 ;
        RECT 3520.720 2014.530 3521.000 2014.810 ;
        RECT 3521.430 2014.530 3521.710 2014.810 ;
        RECT 3512.255 2010.615 3512.535 2010.895 ;
        RECT 3512.965 2010.615 3513.245 2010.895 ;
        RECT 3513.675 2010.615 3513.955 2010.895 ;
        RECT 3514.385 2010.615 3514.665 2010.895 ;
        RECT 3515.095 2010.615 3515.375 2010.895 ;
        RECT 3515.805 2010.615 3516.085 2010.895 ;
        RECT 3516.515 2010.615 3516.795 2010.895 ;
        RECT 3517.225 2010.615 3517.505 2010.895 ;
        RECT 3517.935 2010.615 3518.215 2010.895 ;
        RECT 3518.645 2010.615 3518.925 2010.895 ;
        RECT 3519.355 2010.615 3519.635 2010.895 ;
        RECT 3520.065 2010.615 3520.345 2010.895 ;
        RECT 3520.775 2010.615 3521.055 2010.895 ;
        RECT 3521.485 2010.615 3521.765 2010.895 ;
        RECT 3512.255 2009.905 3512.535 2010.185 ;
        RECT 3512.965 2009.905 3513.245 2010.185 ;
        RECT 3513.675 2009.905 3513.955 2010.185 ;
        RECT 3514.385 2009.905 3514.665 2010.185 ;
        RECT 3515.095 2009.905 3515.375 2010.185 ;
        RECT 3515.805 2009.905 3516.085 2010.185 ;
        RECT 3516.515 2009.905 3516.795 2010.185 ;
        RECT 3517.225 2009.905 3517.505 2010.185 ;
        RECT 3517.935 2009.905 3518.215 2010.185 ;
        RECT 3518.645 2009.905 3518.925 2010.185 ;
        RECT 3519.355 2009.905 3519.635 2010.185 ;
        RECT 3520.065 2009.905 3520.345 2010.185 ;
        RECT 3520.775 2009.905 3521.055 2010.185 ;
        RECT 3521.485 2009.905 3521.765 2010.185 ;
        RECT 3512.255 2009.195 3512.535 2009.475 ;
        RECT 3512.965 2009.195 3513.245 2009.475 ;
        RECT 3513.675 2009.195 3513.955 2009.475 ;
        RECT 3514.385 2009.195 3514.665 2009.475 ;
        RECT 3515.095 2009.195 3515.375 2009.475 ;
        RECT 3515.805 2009.195 3516.085 2009.475 ;
        RECT 3516.515 2009.195 3516.795 2009.475 ;
        RECT 3517.225 2009.195 3517.505 2009.475 ;
        RECT 3517.935 2009.195 3518.215 2009.475 ;
        RECT 3518.645 2009.195 3518.925 2009.475 ;
        RECT 3519.355 2009.195 3519.635 2009.475 ;
        RECT 3520.065 2009.195 3520.345 2009.475 ;
        RECT 3520.775 2009.195 3521.055 2009.475 ;
        RECT 3521.485 2009.195 3521.765 2009.475 ;
        RECT 3512.255 2008.485 3512.535 2008.765 ;
        RECT 3512.965 2008.485 3513.245 2008.765 ;
        RECT 3513.675 2008.485 3513.955 2008.765 ;
        RECT 3514.385 2008.485 3514.665 2008.765 ;
        RECT 3515.095 2008.485 3515.375 2008.765 ;
        RECT 3515.805 2008.485 3516.085 2008.765 ;
        RECT 3516.515 2008.485 3516.795 2008.765 ;
        RECT 3517.225 2008.485 3517.505 2008.765 ;
        RECT 3517.935 2008.485 3518.215 2008.765 ;
        RECT 3518.645 2008.485 3518.925 2008.765 ;
        RECT 3519.355 2008.485 3519.635 2008.765 ;
        RECT 3520.065 2008.485 3520.345 2008.765 ;
        RECT 3520.775 2008.485 3521.055 2008.765 ;
        RECT 3521.485 2008.485 3521.765 2008.765 ;
        RECT 3512.255 2007.775 3512.535 2008.055 ;
        RECT 3512.965 2007.775 3513.245 2008.055 ;
        RECT 3513.675 2007.775 3513.955 2008.055 ;
        RECT 3514.385 2007.775 3514.665 2008.055 ;
        RECT 3515.095 2007.775 3515.375 2008.055 ;
        RECT 3515.805 2007.775 3516.085 2008.055 ;
        RECT 3516.515 2007.775 3516.795 2008.055 ;
        RECT 3517.225 2007.775 3517.505 2008.055 ;
        RECT 3517.935 2007.775 3518.215 2008.055 ;
        RECT 3518.645 2007.775 3518.925 2008.055 ;
        RECT 3519.355 2007.775 3519.635 2008.055 ;
        RECT 3520.065 2007.775 3520.345 2008.055 ;
        RECT 3520.775 2007.775 3521.055 2008.055 ;
        RECT 3521.485 2007.775 3521.765 2008.055 ;
        RECT 3512.255 2007.065 3512.535 2007.345 ;
        RECT 3512.965 2007.065 3513.245 2007.345 ;
        RECT 3513.675 2007.065 3513.955 2007.345 ;
        RECT 3514.385 2007.065 3514.665 2007.345 ;
        RECT 3515.095 2007.065 3515.375 2007.345 ;
        RECT 3515.805 2007.065 3516.085 2007.345 ;
        RECT 3516.515 2007.065 3516.795 2007.345 ;
        RECT 3517.225 2007.065 3517.505 2007.345 ;
        RECT 3517.935 2007.065 3518.215 2007.345 ;
        RECT 3518.645 2007.065 3518.925 2007.345 ;
        RECT 3519.355 2007.065 3519.635 2007.345 ;
        RECT 3520.065 2007.065 3520.345 2007.345 ;
        RECT 3520.775 2007.065 3521.055 2007.345 ;
        RECT 3521.485 2007.065 3521.765 2007.345 ;
        RECT 3512.255 2006.355 3512.535 2006.635 ;
        RECT 3512.965 2006.355 3513.245 2006.635 ;
        RECT 3513.675 2006.355 3513.955 2006.635 ;
        RECT 3514.385 2006.355 3514.665 2006.635 ;
        RECT 3515.095 2006.355 3515.375 2006.635 ;
        RECT 3515.805 2006.355 3516.085 2006.635 ;
        RECT 3516.515 2006.355 3516.795 2006.635 ;
        RECT 3517.225 2006.355 3517.505 2006.635 ;
        RECT 3517.935 2006.355 3518.215 2006.635 ;
        RECT 3518.645 2006.355 3518.925 2006.635 ;
        RECT 3519.355 2006.355 3519.635 2006.635 ;
        RECT 3520.065 2006.355 3520.345 2006.635 ;
        RECT 3520.775 2006.355 3521.055 2006.635 ;
        RECT 3521.485 2006.355 3521.765 2006.635 ;
        RECT 3512.255 2005.645 3512.535 2005.925 ;
        RECT 3512.965 2005.645 3513.245 2005.925 ;
        RECT 3513.675 2005.645 3513.955 2005.925 ;
        RECT 3514.385 2005.645 3514.665 2005.925 ;
        RECT 3515.095 2005.645 3515.375 2005.925 ;
        RECT 3515.805 2005.645 3516.085 2005.925 ;
        RECT 3516.515 2005.645 3516.795 2005.925 ;
        RECT 3517.225 2005.645 3517.505 2005.925 ;
        RECT 3517.935 2005.645 3518.215 2005.925 ;
        RECT 3518.645 2005.645 3518.925 2005.925 ;
        RECT 3519.355 2005.645 3519.635 2005.925 ;
        RECT 3520.065 2005.645 3520.345 2005.925 ;
        RECT 3520.775 2005.645 3521.055 2005.925 ;
        RECT 3521.485 2005.645 3521.765 2005.925 ;
        RECT 3512.255 2004.935 3512.535 2005.215 ;
        RECT 3512.965 2004.935 3513.245 2005.215 ;
        RECT 3513.675 2004.935 3513.955 2005.215 ;
        RECT 3514.385 2004.935 3514.665 2005.215 ;
        RECT 3515.095 2004.935 3515.375 2005.215 ;
        RECT 3515.805 2004.935 3516.085 2005.215 ;
        RECT 3516.515 2004.935 3516.795 2005.215 ;
        RECT 3517.225 2004.935 3517.505 2005.215 ;
        RECT 3517.935 2004.935 3518.215 2005.215 ;
        RECT 3518.645 2004.935 3518.925 2005.215 ;
        RECT 3519.355 2004.935 3519.635 2005.215 ;
        RECT 3520.065 2004.935 3520.345 2005.215 ;
        RECT 3520.775 2004.935 3521.055 2005.215 ;
        RECT 3521.485 2004.935 3521.765 2005.215 ;
        RECT 3512.255 2004.225 3512.535 2004.505 ;
        RECT 3512.965 2004.225 3513.245 2004.505 ;
        RECT 3513.675 2004.225 3513.955 2004.505 ;
        RECT 3514.385 2004.225 3514.665 2004.505 ;
        RECT 3515.095 2004.225 3515.375 2004.505 ;
        RECT 3515.805 2004.225 3516.085 2004.505 ;
        RECT 3516.515 2004.225 3516.795 2004.505 ;
        RECT 3517.225 2004.225 3517.505 2004.505 ;
        RECT 3517.935 2004.225 3518.215 2004.505 ;
        RECT 3518.645 2004.225 3518.925 2004.505 ;
        RECT 3519.355 2004.225 3519.635 2004.505 ;
        RECT 3520.065 2004.225 3520.345 2004.505 ;
        RECT 3520.775 2004.225 3521.055 2004.505 ;
        RECT 3521.485 2004.225 3521.765 2004.505 ;
        RECT 3512.255 2003.515 3512.535 2003.795 ;
        RECT 3512.965 2003.515 3513.245 2003.795 ;
        RECT 3513.675 2003.515 3513.955 2003.795 ;
        RECT 3514.385 2003.515 3514.665 2003.795 ;
        RECT 3515.095 2003.515 3515.375 2003.795 ;
        RECT 3515.805 2003.515 3516.085 2003.795 ;
        RECT 3516.515 2003.515 3516.795 2003.795 ;
        RECT 3517.225 2003.515 3517.505 2003.795 ;
        RECT 3517.935 2003.515 3518.215 2003.795 ;
        RECT 3518.645 2003.515 3518.925 2003.795 ;
        RECT 3519.355 2003.515 3519.635 2003.795 ;
        RECT 3520.065 2003.515 3520.345 2003.795 ;
        RECT 3520.775 2003.515 3521.055 2003.795 ;
        RECT 3521.485 2003.515 3521.765 2003.795 ;
        RECT 3512.255 2002.805 3512.535 2003.085 ;
        RECT 3512.965 2002.805 3513.245 2003.085 ;
        RECT 3513.675 2002.805 3513.955 2003.085 ;
        RECT 3514.385 2002.805 3514.665 2003.085 ;
        RECT 3515.095 2002.805 3515.375 2003.085 ;
        RECT 3515.805 2002.805 3516.085 2003.085 ;
        RECT 3516.515 2002.805 3516.795 2003.085 ;
        RECT 3517.225 2002.805 3517.505 2003.085 ;
        RECT 3517.935 2002.805 3518.215 2003.085 ;
        RECT 3518.645 2002.805 3518.925 2003.085 ;
        RECT 3519.355 2002.805 3519.635 2003.085 ;
        RECT 3520.065 2002.805 3520.345 2003.085 ;
        RECT 3520.775 2002.805 3521.055 2003.085 ;
        RECT 3521.485 2002.805 3521.765 2003.085 ;
        RECT 3512.255 2002.095 3512.535 2002.375 ;
        RECT 3512.965 2002.095 3513.245 2002.375 ;
        RECT 3513.675 2002.095 3513.955 2002.375 ;
        RECT 3514.385 2002.095 3514.665 2002.375 ;
        RECT 3515.095 2002.095 3515.375 2002.375 ;
        RECT 3515.805 2002.095 3516.085 2002.375 ;
        RECT 3516.515 2002.095 3516.795 2002.375 ;
        RECT 3517.225 2002.095 3517.505 2002.375 ;
        RECT 3517.935 2002.095 3518.215 2002.375 ;
        RECT 3518.645 2002.095 3518.925 2002.375 ;
        RECT 3519.355 2002.095 3519.635 2002.375 ;
        RECT 3520.065 2002.095 3520.345 2002.375 ;
        RECT 3520.775 2002.095 3521.055 2002.375 ;
        RECT 3521.485 2002.095 3521.765 2002.375 ;
        RECT 3512.255 2001.385 3512.535 2001.665 ;
        RECT 3512.965 2001.385 3513.245 2001.665 ;
        RECT 3513.675 2001.385 3513.955 2001.665 ;
        RECT 3514.385 2001.385 3514.665 2001.665 ;
        RECT 3515.095 2001.385 3515.375 2001.665 ;
        RECT 3515.805 2001.385 3516.085 2001.665 ;
        RECT 3516.515 2001.385 3516.795 2001.665 ;
        RECT 3517.225 2001.385 3517.505 2001.665 ;
        RECT 3517.935 2001.385 3518.215 2001.665 ;
        RECT 3518.645 2001.385 3518.925 2001.665 ;
        RECT 3519.355 2001.385 3519.635 2001.665 ;
        RECT 3520.065 2001.385 3520.345 2001.665 ;
        RECT 3520.775 2001.385 3521.055 2001.665 ;
        RECT 3521.485 2001.385 3521.765 2001.665 ;
        RECT 3512.255 1998.765 3512.535 1999.045 ;
        RECT 3512.965 1998.765 3513.245 1999.045 ;
        RECT 3513.675 1998.765 3513.955 1999.045 ;
        RECT 3514.385 1998.765 3514.665 1999.045 ;
        RECT 3515.095 1998.765 3515.375 1999.045 ;
        RECT 3515.805 1998.765 3516.085 1999.045 ;
        RECT 3516.515 1998.765 3516.795 1999.045 ;
        RECT 3517.225 1998.765 3517.505 1999.045 ;
        RECT 3517.935 1998.765 3518.215 1999.045 ;
        RECT 3518.645 1998.765 3518.925 1999.045 ;
        RECT 3519.355 1998.765 3519.635 1999.045 ;
        RECT 3520.065 1998.765 3520.345 1999.045 ;
        RECT 3520.775 1998.765 3521.055 1999.045 ;
        RECT 3521.485 1998.765 3521.765 1999.045 ;
        RECT 3512.255 1998.055 3512.535 1998.335 ;
        RECT 3512.965 1998.055 3513.245 1998.335 ;
        RECT 3513.675 1998.055 3513.955 1998.335 ;
        RECT 3514.385 1998.055 3514.665 1998.335 ;
        RECT 3515.095 1998.055 3515.375 1998.335 ;
        RECT 3515.805 1998.055 3516.085 1998.335 ;
        RECT 3516.515 1998.055 3516.795 1998.335 ;
        RECT 3517.225 1998.055 3517.505 1998.335 ;
        RECT 3517.935 1998.055 3518.215 1998.335 ;
        RECT 3518.645 1998.055 3518.925 1998.335 ;
        RECT 3519.355 1998.055 3519.635 1998.335 ;
        RECT 3520.065 1998.055 3520.345 1998.335 ;
        RECT 3520.775 1998.055 3521.055 1998.335 ;
        RECT 3521.485 1998.055 3521.765 1998.335 ;
        RECT 3512.255 1997.345 3512.535 1997.625 ;
        RECT 3512.965 1997.345 3513.245 1997.625 ;
        RECT 3513.675 1997.345 3513.955 1997.625 ;
        RECT 3514.385 1997.345 3514.665 1997.625 ;
        RECT 3515.095 1997.345 3515.375 1997.625 ;
        RECT 3515.805 1997.345 3516.085 1997.625 ;
        RECT 3516.515 1997.345 3516.795 1997.625 ;
        RECT 3517.225 1997.345 3517.505 1997.625 ;
        RECT 3517.935 1997.345 3518.215 1997.625 ;
        RECT 3518.645 1997.345 3518.925 1997.625 ;
        RECT 3519.355 1997.345 3519.635 1997.625 ;
        RECT 3520.065 1997.345 3520.345 1997.625 ;
        RECT 3520.775 1997.345 3521.055 1997.625 ;
        RECT 3521.485 1997.345 3521.765 1997.625 ;
        RECT 3512.255 1996.635 3512.535 1996.915 ;
        RECT 3512.965 1996.635 3513.245 1996.915 ;
        RECT 3513.675 1996.635 3513.955 1996.915 ;
        RECT 3514.385 1996.635 3514.665 1996.915 ;
        RECT 3515.095 1996.635 3515.375 1996.915 ;
        RECT 3515.805 1996.635 3516.085 1996.915 ;
        RECT 3516.515 1996.635 3516.795 1996.915 ;
        RECT 3517.225 1996.635 3517.505 1996.915 ;
        RECT 3517.935 1996.635 3518.215 1996.915 ;
        RECT 3518.645 1996.635 3518.925 1996.915 ;
        RECT 3519.355 1996.635 3519.635 1996.915 ;
        RECT 3520.065 1996.635 3520.345 1996.915 ;
        RECT 3520.775 1996.635 3521.055 1996.915 ;
        RECT 3521.485 1996.635 3521.765 1996.915 ;
        RECT 3512.255 1995.925 3512.535 1996.205 ;
        RECT 3512.965 1995.925 3513.245 1996.205 ;
        RECT 3513.675 1995.925 3513.955 1996.205 ;
        RECT 3514.385 1995.925 3514.665 1996.205 ;
        RECT 3515.095 1995.925 3515.375 1996.205 ;
        RECT 3515.805 1995.925 3516.085 1996.205 ;
        RECT 3516.515 1995.925 3516.795 1996.205 ;
        RECT 3517.225 1995.925 3517.505 1996.205 ;
        RECT 3517.935 1995.925 3518.215 1996.205 ;
        RECT 3518.645 1995.925 3518.925 1996.205 ;
        RECT 3519.355 1995.925 3519.635 1996.205 ;
        RECT 3520.065 1995.925 3520.345 1996.205 ;
        RECT 3520.775 1995.925 3521.055 1996.205 ;
        RECT 3521.485 1995.925 3521.765 1996.205 ;
        RECT 3512.255 1995.215 3512.535 1995.495 ;
        RECT 3512.965 1995.215 3513.245 1995.495 ;
        RECT 3513.675 1995.215 3513.955 1995.495 ;
        RECT 3514.385 1995.215 3514.665 1995.495 ;
        RECT 3515.095 1995.215 3515.375 1995.495 ;
        RECT 3515.805 1995.215 3516.085 1995.495 ;
        RECT 3516.515 1995.215 3516.795 1995.495 ;
        RECT 3517.225 1995.215 3517.505 1995.495 ;
        RECT 3517.935 1995.215 3518.215 1995.495 ;
        RECT 3518.645 1995.215 3518.925 1995.495 ;
        RECT 3519.355 1995.215 3519.635 1995.495 ;
        RECT 3520.065 1995.215 3520.345 1995.495 ;
        RECT 3520.775 1995.215 3521.055 1995.495 ;
        RECT 3521.485 1995.215 3521.765 1995.495 ;
        RECT 3512.255 1994.505 3512.535 1994.785 ;
        RECT 3512.965 1994.505 3513.245 1994.785 ;
        RECT 3513.675 1994.505 3513.955 1994.785 ;
        RECT 3514.385 1994.505 3514.665 1994.785 ;
        RECT 3515.095 1994.505 3515.375 1994.785 ;
        RECT 3515.805 1994.505 3516.085 1994.785 ;
        RECT 3516.515 1994.505 3516.795 1994.785 ;
        RECT 3517.225 1994.505 3517.505 1994.785 ;
        RECT 3517.935 1994.505 3518.215 1994.785 ;
        RECT 3518.645 1994.505 3518.925 1994.785 ;
        RECT 3519.355 1994.505 3519.635 1994.785 ;
        RECT 3520.065 1994.505 3520.345 1994.785 ;
        RECT 3520.775 1994.505 3521.055 1994.785 ;
        RECT 3521.485 1994.505 3521.765 1994.785 ;
        RECT 3512.255 1993.795 3512.535 1994.075 ;
        RECT 3512.965 1993.795 3513.245 1994.075 ;
        RECT 3513.675 1993.795 3513.955 1994.075 ;
        RECT 3514.385 1993.795 3514.665 1994.075 ;
        RECT 3515.095 1993.795 3515.375 1994.075 ;
        RECT 3515.805 1993.795 3516.085 1994.075 ;
        RECT 3516.515 1993.795 3516.795 1994.075 ;
        RECT 3517.225 1993.795 3517.505 1994.075 ;
        RECT 3517.935 1993.795 3518.215 1994.075 ;
        RECT 3518.645 1993.795 3518.925 1994.075 ;
        RECT 3519.355 1993.795 3519.635 1994.075 ;
        RECT 3520.065 1993.795 3520.345 1994.075 ;
        RECT 3520.775 1993.795 3521.055 1994.075 ;
        RECT 3521.485 1993.795 3521.765 1994.075 ;
        RECT 3512.255 1993.085 3512.535 1993.365 ;
        RECT 3512.965 1993.085 3513.245 1993.365 ;
        RECT 3513.675 1993.085 3513.955 1993.365 ;
        RECT 3514.385 1993.085 3514.665 1993.365 ;
        RECT 3515.095 1993.085 3515.375 1993.365 ;
        RECT 3515.805 1993.085 3516.085 1993.365 ;
        RECT 3516.515 1993.085 3516.795 1993.365 ;
        RECT 3517.225 1993.085 3517.505 1993.365 ;
        RECT 3517.935 1993.085 3518.215 1993.365 ;
        RECT 3518.645 1993.085 3518.925 1993.365 ;
        RECT 3519.355 1993.085 3519.635 1993.365 ;
        RECT 3520.065 1993.085 3520.345 1993.365 ;
        RECT 3520.775 1993.085 3521.055 1993.365 ;
        RECT 3521.485 1993.085 3521.765 1993.365 ;
        RECT 3512.255 1992.375 3512.535 1992.655 ;
        RECT 3512.965 1992.375 3513.245 1992.655 ;
        RECT 3513.675 1992.375 3513.955 1992.655 ;
        RECT 3514.385 1992.375 3514.665 1992.655 ;
        RECT 3515.095 1992.375 3515.375 1992.655 ;
        RECT 3515.805 1992.375 3516.085 1992.655 ;
        RECT 3516.515 1992.375 3516.795 1992.655 ;
        RECT 3517.225 1992.375 3517.505 1992.655 ;
        RECT 3517.935 1992.375 3518.215 1992.655 ;
        RECT 3518.645 1992.375 3518.925 1992.655 ;
        RECT 3519.355 1992.375 3519.635 1992.655 ;
        RECT 3520.065 1992.375 3520.345 1992.655 ;
        RECT 3520.775 1992.375 3521.055 1992.655 ;
        RECT 3521.485 1992.375 3521.765 1992.655 ;
        RECT 3512.255 1991.665 3512.535 1991.945 ;
        RECT 3512.965 1991.665 3513.245 1991.945 ;
        RECT 3513.675 1991.665 3513.955 1991.945 ;
        RECT 3514.385 1991.665 3514.665 1991.945 ;
        RECT 3515.095 1991.665 3515.375 1991.945 ;
        RECT 3515.805 1991.665 3516.085 1991.945 ;
        RECT 3516.515 1991.665 3516.795 1991.945 ;
        RECT 3517.225 1991.665 3517.505 1991.945 ;
        RECT 3517.935 1991.665 3518.215 1991.945 ;
        RECT 3518.645 1991.665 3518.925 1991.945 ;
        RECT 3519.355 1991.665 3519.635 1991.945 ;
        RECT 3520.065 1991.665 3520.345 1991.945 ;
        RECT 3520.775 1991.665 3521.055 1991.945 ;
        RECT 3521.485 1991.665 3521.765 1991.945 ;
        RECT 3512.255 1990.955 3512.535 1991.235 ;
        RECT 3512.965 1990.955 3513.245 1991.235 ;
        RECT 3513.675 1990.955 3513.955 1991.235 ;
        RECT 3514.385 1990.955 3514.665 1991.235 ;
        RECT 3515.095 1990.955 3515.375 1991.235 ;
        RECT 3515.805 1990.955 3516.085 1991.235 ;
        RECT 3516.515 1990.955 3516.795 1991.235 ;
        RECT 3517.225 1990.955 3517.505 1991.235 ;
        RECT 3517.935 1990.955 3518.215 1991.235 ;
        RECT 3518.645 1990.955 3518.925 1991.235 ;
        RECT 3519.355 1990.955 3519.635 1991.235 ;
        RECT 3520.065 1990.955 3520.345 1991.235 ;
        RECT 3520.775 1990.955 3521.055 1991.235 ;
        RECT 3521.485 1990.955 3521.765 1991.235 ;
        RECT 3512.255 1990.245 3512.535 1990.525 ;
        RECT 3512.965 1990.245 3513.245 1990.525 ;
        RECT 3513.675 1990.245 3513.955 1990.525 ;
        RECT 3514.385 1990.245 3514.665 1990.525 ;
        RECT 3515.095 1990.245 3515.375 1990.525 ;
        RECT 3515.805 1990.245 3516.085 1990.525 ;
        RECT 3516.515 1990.245 3516.795 1990.525 ;
        RECT 3517.225 1990.245 3517.505 1990.525 ;
        RECT 3517.935 1990.245 3518.215 1990.525 ;
        RECT 3518.645 1990.245 3518.925 1990.525 ;
        RECT 3519.355 1990.245 3519.635 1990.525 ;
        RECT 3520.065 1990.245 3520.345 1990.525 ;
        RECT 3520.775 1990.245 3521.055 1990.525 ;
        RECT 3521.485 1990.245 3521.765 1990.525 ;
        RECT 3512.255 1989.535 3512.535 1989.815 ;
        RECT 3512.965 1989.535 3513.245 1989.815 ;
        RECT 3513.675 1989.535 3513.955 1989.815 ;
        RECT 3514.385 1989.535 3514.665 1989.815 ;
        RECT 3515.095 1989.535 3515.375 1989.815 ;
        RECT 3515.805 1989.535 3516.085 1989.815 ;
        RECT 3516.515 1989.535 3516.795 1989.815 ;
        RECT 3517.225 1989.535 3517.505 1989.815 ;
        RECT 3517.935 1989.535 3518.215 1989.815 ;
        RECT 3518.645 1989.535 3518.925 1989.815 ;
        RECT 3519.355 1989.535 3519.635 1989.815 ;
        RECT 3520.065 1989.535 3520.345 1989.815 ;
        RECT 3520.775 1989.535 3521.055 1989.815 ;
        RECT 3521.485 1989.535 3521.765 1989.815 ;
        RECT 3512.255 1985.235 3512.535 1985.515 ;
        RECT 3512.965 1985.235 3513.245 1985.515 ;
        RECT 3513.675 1985.235 3513.955 1985.515 ;
        RECT 3514.385 1985.235 3514.665 1985.515 ;
        RECT 3515.095 1985.235 3515.375 1985.515 ;
        RECT 3515.805 1985.235 3516.085 1985.515 ;
        RECT 3516.515 1985.235 3516.795 1985.515 ;
        RECT 3517.225 1985.235 3517.505 1985.515 ;
        RECT 3517.935 1985.235 3518.215 1985.515 ;
        RECT 3518.645 1985.235 3518.925 1985.515 ;
        RECT 3519.355 1985.235 3519.635 1985.515 ;
        RECT 3520.065 1985.235 3520.345 1985.515 ;
        RECT 3520.775 1985.235 3521.055 1985.515 ;
        RECT 3521.485 1985.235 3521.765 1985.515 ;
        RECT 3512.255 1984.525 3512.535 1984.805 ;
        RECT 3512.965 1984.525 3513.245 1984.805 ;
        RECT 3513.675 1984.525 3513.955 1984.805 ;
        RECT 3514.385 1984.525 3514.665 1984.805 ;
        RECT 3515.095 1984.525 3515.375 1984.805 ;
        RECT 3515.805 1984.525 3516.085 1984.805 ;
        RECT 3516.515 1984.525 3516.795 1984.805 ;
        RECT 3517.225 1984.525 3517.505 1984.805 ;
        RECT 3517.935 1984.525 3518.215 1984.805 ;
        RECT 3518.645 1984.525 3518.925 1984.805 ;
        RECT 3519.355 1984.525 3519.635 1984.805 ;
        RECT 3520.065 1984.525 3520.345 1984.805 ;
        RECT 3520.775 1984.525 3521.055 1984.805 ;
        RECT 3521.485 1984.525 3521.765 1984.805 ;
        RECT 3512.255 1983.815 3512.535 1984.095 ;
        RECT 3512.965 1983.815 3513.245 1984.095 ;
        RECT 3513.675 1983.815 3513.955 1984.095 ;
        RECT 3514.385 1983.815 3514.665 1984.095 ;
        RECT 3515.095 1983.815 3515.375 1984.095 ;
        RECT 3515.805 1983.815 3516.085 1984.095 ;
        RECT 3516.515 1983.815 3516.795 1984.095 ;
        RECT 3517.225 1983.815 3517.505 1984.095 ;
        RECT 3517.935 1983.815 3518.215 1984.095 ;
        RECT 3518.645 1983.815 3518.925 1984.095 ;
        RECT 3519.355 1983.815 3519.635 1984.095 ;
        RECT 3520.065 1983.815 3520.345 1984.095 ;
        RECT 3520.775 1983.815 3521.055 1984.095 ;
        RECT 3521.485 1983.815 3521.765 1984.095 ;
        RECT 3512.255 1983.105 3512.535 1983.385 ;
        RECT 3512.965 1983.105 3513.245 1983.385 ;
        RECT 3513.675 1983.105 3513.955 1983.385 ;
        RECT 3514.385 1983.105 3514.665 1983.385 ;
        RECT 3515.095 1983.105 3515.375 1983.385 ;
        RECT 3515.805 1983.105 3516.085 1983.385 ;
        RECT 3516.515 1983.105 3516.795 1983.385 ;
        RECT 3517.225 1983.105 3517.505 1983.385 ;
        RECT 3517.935 1983.105 3518.215 1983.385 ;
        RECT 3518.645 1983.105 3518.925 1983.385 ;
        RECT 3519.355 1983.105 3519.635 1983.385 ;
        RECT 3520.065 1983.105 3520.345 1983.385 ;
        RECT 3520.775 1983.105 3521.055 1983.385 ;
        RECT 3521.485 1983.105 3521.765 1983.385 ;
        RECT 3512.255 1982.395 3512.535 1982.675 ;
        RECT 3512.965 1982.395 3513.245 1982.675 ;
        RECT 3513.675 1982.395 3513.955 1982.675 ;
        RECT 3514.385 1982.395 3514.665 1982.675 ;
        RECT 3515.095 1982.395 3515.375 1982.675 ;
        RECT 3515.805 1982.395 3516.085 1982.675 ;
        RECT 3516.515 1982.395 3516.795 1982.675 ;
        RECT 3517.225 1982.395 3517.505 1982.675 ;
        RECT 3517.935 1982.395 3518.215 1982.675 ;
        RECT 3518.645 1982.395 3518.925 1982.675 ;
        RECT 3519.355 1982.395 3519.635 1982.675 ;
        RECT 3520.065 1982.395 3520.345 1982.675 ;
        RECT 3520.775 1982.395 3521.055 1982.675 ;
        RECT 3521.485 1982.395 3521.765 1982.675 ;
        RECT 3512.255 1981.685 3512.535 1981.965 ;
        RECT 3512.965 1981.685 3513.245 1981.965 ;
        RECT 3513.675 1981.685 3513.955 1981.965 ;
        RECT 3514.385 1981.685 3514.665 1981.965 ;
        RECT 3515.095 1981.685 3515.375 1981.965 ;
        RECT 3515.805 1981.685 3516.085 1981.965 ;
        RECT 3516.515 1981.685 3516.795 1981.965 ;
        RECT 3517.225 1981.685 3517.505 1981.965 ;
        RECT 3517.935 1981.685 3518.215 1981.965 ;
        RECT 3518.645 1981.685 3518.925 1981.965 ;
        RECT 3519.355 1981.685 3519.635 1981.965 ;
        RECT 3520.065 1981.685 3520.345 1981.965 ;
        RECT 3520.775 1981.685 3521.055 1981.965 ;
        RECT 3521.485 1981.685 3521.765 1981.965 ;
        RECT 3512.255 1980.975 3512.535 1981.255 ;
        RECT 3512.965 1980.975 3513.245 1981.255 ;
        RECT 3513.675 1980.975 3513.955 1981.255 ;
        RECT 3514.385 1980.975 3514.665 1981.255 ;
        RECT 3515.095 1980.975 3515.375 1981.255 ;
        RECT 3515.805 1980.975 3516.085 1981.255 ;
        RECT 3516.515 1980.975 3516.795 1981.255 ;
        RECT 3517.225 1980.975 3517.505 1981.255 ;
        RECT 3517.935 1980.975 3518.215 1981.255 ;
        RECT 3518.645 1980.975 3518.925 1981.255 ;
        RECT 3519.355 1980.975 3519.635 1981.255 ;
        RECT 3520.065 1980.975 3520.345 1981.255 ;
        RECT 3520.775 1980.975 3521.055 1981.255 ;
        RECT 3521.485 1980.975 3521.765 1981.255 ;
        RECT 3512.255 1980.265 3512.535 1980.545 ;
        RECT 3512.965 1980.265 3513.245 1980.545 ;
        RECT 3513.675 1980.265 3513.955 1980.545 ;
        RECT 3514.385 1980.265 3514.665 1980.545 ;
        RECT 3515.095 1980.265 3515.375 1980.545 ;
        RECT 3515.805 1980.265 3516.085 1980.545 ;
        RECT 3516.515 1980.265 3516.795 1980.545 ;
        RECT 3517.225 1980.265 3517.505 1980.545 ;
        RECT 3517.935 1980.265 3518.215 1980.545 ;
        RECT 3518.645 1980.265 3518.925 1980.545 ;
        RECT 3519.355 1980.265 3519.635 1980.545 ;
        RECT 3520.065 1980.265 3520.345 1980.545 ;
        RECT 3520.775 1980.265 3521.055 1980.545 ;
        RECT 3521.485 1980.265 3521.765 1980.545 ;
        RECT 3512.255 1979.555 3512.535 1979.835 ;
        RECT 3512.965 1979.555 3513.245 1979.835 ;
        RECT 3513.675 1979.555 3513.955 1979.835 ;
        RECT 3514.385 1979.555 3514.665 1979.835 ;
        RECT 3515.095 1979.555 3515.375 1979.835 ;
        RECT 3515.805 1979.555 3516.085 1979.835 ;
        RECT 3516.515 1979.555 3516.795 1979.835 ;
        RECT 3517.225 1979.555 3517.505 1979.835 ;
        RECT 3517.935 1979.555 3518.215 1979.835 ;
        RECT 3518.645 1979.555 3518.925 1979.835 ;
        RECT 3519.355 1979.555 3519.635 1979.835 ;
        RECT 3520.065 1979.555 3520.345 1979.835 ;
        RECT 3520.775 1979.555 3521.055 1979.835 ;
        RECT 3521.485 1979.555 3521.765 1979.835 ;
        RECT 3512.255 1978.845 3512.535 1979.125 ;
        RECT 3512.965 1978.845 3513.245 1979.125 ;
        RECT 3513.675 1978.845 3513.955 1979.125 ;
        RECT 3514.385 1978.845 3514.665 1979.125 ;
        RECT 3515.095 1978.845 3515.375 1979.125 ;
        RECT 3515.805 1978.845 3516.085 1979.125 ;
        RECT 3516.515 1978.845 3516.795 1979.125 ;
        RECT 3517.225 1978.845 3517.505 1979.125 ;
        RECT 3517.935 1978.845 3518.215 1979.125 ;
        RECT 3518.645 1978.845 3518.925 1979.125 ;
        RECT 3519.355 1978.845 3519.635 1979.125 ;
        RECT 3520.065 1978.845 3520.345 1979.125 ;
        RECT 3520.775 1978.845 3521.055 1979.125 ;
        RECT 3521.485 1978.845 3521.765 1979.125 ;
        RECT 3512.255 1978.135 3512.535 1978.415 ;
        RECT 3512.965 1978.135 3513.245 1978.415 ;
        RECT 3513.675 1978.135 3513.955 1978.415 ;
        RECT 3514.385 1978.135 3514.665 1978.415 ;
        RECT 3515.095 1978.135 3515.375 1978.415 ;
        RECT 3515.805 1978.135 3516.085 1978.415 ;
        RECT 3516.515 1978.135 3516.795 1978.415 ;
        RECT 3517.225 1978.135 3517.505 1978.415 ;
        RECT 3517.935 1978.135 3518.215 1978.415 ;
        RECT 3518.645 1978.135 3518.925 1978.415 ;
        RECT 3519.355 1978.135 3519.635 1978.415 ;
        RECT 3520.065 1978.135 3520.345 1978.415 ;
        RECT 3520.775 1978.135 3521.055 1978.415 ;
        RECT 3521.485 1978.135 3521.765 1978.415 ;
        RECT 3512.255 1977.425 3512.535 1977.705 ;
        RECT 3512.965 1977.425 3513.245 1977.705 ;
        RECT 3513.675 1977.425 3513.955 1977.705 ;
        RECT 3514.385 1977.425 3514.665 1977.705 ;
        RECT 3515.095 1977.425 3515.375 1977.705 ;
        RECT 3515.805 1977.425 3516.085 1977.705 ;
        RECT 3516.515 1977.425 3516.795 1977.705 ;
        RECT 3517.225 1977.425 3517.505 1977.705 ;
        RECT 3517.935 1977.425 3518.215 1977.705 ;
        RECT 3518.645 1977.425 3518.925 1977.705 ;
        RECT 3519.355 1977.425 3519.635 1977.705 ;
        RECT 3520.065 1977.425 3520.345 1977.705 ;
        RECT 3520.775 1977.425 3521.055 1977.705 ;
        RECT 3521.485 1977.425 3521.765 1977.705 ;
        RECT 3512.255 1976.715 3512.535 1976.995 ;
        RECT 3512.965 1976.715 3513.245 1976.995 ;
        RECT 3513.675 1976.715 3513.955 1976.995 ;
        RECT 3514.385 1976.715 3514.665 1976.995 ;
        RECT 3515.095 1976.715 3515.375 1976.995 ;
        RECT 3515.805 1976.715 3516.085 1976.995 ;
        RECT 3516.515 1976.715 3516.795 1976.995 ;
        RECT 3517.225 1976.715 3517.505 1976.995 ;
        RECT 3517.935 1976.715 3518.215 1976.995 ;
        RECT 3518.645 1976.715 3518.925 1976.995 ;
        RECT 3519.355 1976.715 3519.635 1976.995 ;
        RECT 3520.065 1976.715 3520.345 1976.995 ;
        RECT 3520.775 1976.715 3521.055 1976.995 ;
        RECT 3521.485 1976.715 3521.765 1976.995 ;
        RECT 3512.255 1976.005 3512.535 1976.285 ;
        RECT 3512.965 1976.005 3513.245 1976.285 ;
        RECT 3513.675 1976.005 3513.955 1976.285 ;
        RECT 3514.385 1976.005 3514.665 1976.285 ;
        RECT 3515.095 1976.005 3515.375 1976.285 ;
        RECT 3515.805 1976.005 3516.085 1976.285 ;
        RECT 3516.515 1976.005 3516.795 1976.285 ;
        RECT 3517.225 1976.005 3517.505 1976.285 ;
        RECT 3517.935 1976.005 3518.215 1976.285 ;
        RECT 3518.645 1976.005 3518.925 1976.285 ;
        RECT 3519.355 1976.005 3519.635 1976.285 ;
        RECT 3520.065 1976.005 3520.345 1976.285 ;
        RECT 3520.775 1976.005 3521.055 1976.285 ;
        RECT 3521.485 1976.005 3521.765 1976.285 ;
        RECT 3512.255 1973.385 3512.535 1973.665 ;
        RECT 3512.965 1973.385 3513.245 1973.665 ;
        RECT 3513.675 1973.385 3513.955 1973.665 ;
        RECT 3514.385 1973.385 3514.665 1973.665 ;
        RECT 3515.095 1973.385 3515.375 1973.665 ;
        RECT 3515.805 1973.385 3516.085 1973.665 ;
        RECT 3516.515 1973.385 3516.795 1973.665 ;
        RECT 3517.225 1973.385 3517.505 1973.665 ;
        RECT 3517.935 1973.385 3518.215 1973.665 ;
        RECT 3518.645 1973.385 3518.925 1973.665 ;
        RECT 3519.355 1973.385 3519.635 1973.665 ;
        RECT 3520.065 1973.385 3520.345 1973.665 ;
        RECT 3520.775 1973.385 3521.055 1973.665 ;
        RECT 3521.485 1973.385 3521.765 1973.665 ;
        RECT 3512.255 1972.675 3512.535 1972.955 ;
        RECT 3512.965 1972.675 3513.245 1972.955 ;
        RECT 3513.675 1972.675 3513.955 1972.955 ;
        RECT 3514.385 1972.675 3514.665 1972.955 ;
        RECT 3515.095 1972.675 3515.375 1972.955 ;
        RECT 3515.805 1972.675 3516.085 1972.955 ;
        RECT 3516.515 1972.675 3516.795 1972.955 ;
        RECT 3517.225 1972.675 3517.505 1972.955 ;
        RECT 3517.935 1972.675 3518.215 1972.955 ;
        RECT 3518.645 1972.675 3518.925 1972.955 ;
        RECT 3519.355 1972.675 3519.635 1972.955 ;
        RECT 3520.065 1972.675 3520.345 1972.955 ;
        RECT 3520.775 1972.675 3521.055 1972.955 ;
        RECT 3521.485 1972.675 3521.765 1972.955 ;
        RECT 3512.255 1971.965 3512.535 1972.245 ;
        RECT 3512.965 1971.965 3513.245 1972.245 ;
        RECT 3513.675 1971.965 3513.955 1972.245 ;
        RECT 3514.385 1971.965 3514.665 1972.245 ;
        RECT 3515.095 1971.965 3515.375 1972.245 ;
        RECT 3515.805 1971.965 3516.085 1972.245 ;
        RECT 3516.515 1971.965 3516.795 1972.245 ;
        RECT 3517.225 1971.965 3517.505 1972.245 ;
        RECT 3517.935 1971.965 3518.215 1972.245 ;
        RECT 3518.645 1971.965 3518.925 1972.245 ;
        RECT 3519.355 1971.965 3519.635 1972.245 ;
        RECT 3520.065 1971.965 3520.345 1972.245 ;
        RECT 3520.775 1971.965 3521.055 1972.245 ;
        RECT 3521.485 1971.965 3521.765 1972.245 ;
        RECT 3512.255 1971.255 3512.535 1971.535 ;
        RECT 3512.965 1971.255 3513.245 1971.535 ;
        RECT 3513.675 1971.255 3513.955 1971.535 ;
        RECT 3514.385 1971.255 3514.665 1971.535 ;
        RECT 3515.095 1971.255 3515.375 1971.535 ;
        RECT 3515.805 1971.255 3516.085 1971.535 ;
        RECT 3516.515 1971.255 3516.795 1971.535 ;
        RECT 3517.225 1971.255 3517.505 1971.535 ;
        RECT 3517.935 1971.255 3518.215 1971.535 ;
        RECT 3518.645 1971.255 3518.925 1971.535 ;
        RECT 3519.355 1971.255 3519.635 1971.535 ;
        RECT 3520.065 1971.255 3520.345 1971.535 ;
        RECT 3520.775 1971.255 3521.055 1971.535 ;
        RECT 3521.485 1971.255 3521.765 1971.535 ;
        RECT 3512.255 1970.545 3512.535 1970.825 ;
        RECT 3512.965 1970.545 3513.245 1970.825 ;
        RECT 3513.675 1970.545 3513.955 1970.825 ;
        RECT 3514.385 1970.545 3514.665 1970.825 ;
        RECT 3515.095 1970.545 3515.375 1970.825 ;
        RECT 3515.805 1970.545 3516.085 1970.825 ;
        RECT 3516.515 1970.545 3516.795 1970.825 ;
        RECT 3517.225 1970.545 3517.505 1970.825 ;
        RECT 3517.935 1970.545 3518.215 1970.825 ;
        RECT 3518.645 1970.545 3518.925 1970.825 ;
        RECT 3519.355 1970.545 3519.635 1970.825 ;
        RECT 3520.065 1970.545 3520.345 1970.825 ;
        RECT 3520.775 1970.545 3521.055 1970.825 ;
        RECT 3521.485 1970.545 3521.765 1970.825 ;
        RECT 3512.255 1969.835 3512.535 1970.115 ;
        RECT 3512.965 1969.835 3513.245 1970.115 ;
        RECT 3513.675 1969.835 3513.955 1970.115 ;
        RECT 3514.385 1969.835 3514.665 1970.115 ;
        RECT 3515.095 1969.835 3515.375 1970.115 ;
        RECT 3515.805 1969.835 3516.085 1970.115 ;
        RECT 3516.515 1969.835 3516.795 1970.115 ;
        RECT 3517.225 1969.835 3517.505 1970.115 ;
        RECT 3517.935 1969.835 3518.215 1970.115 ;
        RECT 3518.645 1969.835 3518.925 1970.115 ;
        RECT 3519.355 1969.835 3519.635 1970.115 ;
        RECT 3520.065 1969.835 3520.345 1970.115 ;
        RECT 3520.775 1969.835 3521.055 1970.115 ;
        RECT 3521.485 1969.835 3521.765 1970.115 ;
        RECT 3512.255 1969.125 3512.535 1969.405 ;
        RECT 3512.965 1969.125 3513.245 1969.405 ;
        RECT 3513.675 1969.125 3513.955 1969.405 ;
        RECT 3514.385 1969.125 3514.665 1969.405 ;
        RECT 3515.095 1969.125 3515.375 1969.405 ;
        RECT 3515.805 1969.125 3516.085 1969.405 ;
        RECT 3516.515 1969.125 3516.795 1969.405 ;
        RECT 3517.225 1969.125 3517.505 1969.405 ;
        RECT 3517.935 1969.125 3518.215 1969.405 ;
        RECT 3518.645 1969.125 3518.925 1969.405 ;
        RECT 3519.355 1969.125 3519.635 1969.405 ;
        RECT 3520.065 1969.125 3520.345 1969.405 ;
        RECT 3520.775 1969.125 3521.055 1969.405 ;
        RECT 3521.485 1969.125 3521.765 1969.405 ;
        RECT 3512.255 1968.415 3512.535 1968.695 ;
        RECT 3512.965 1968.415 3513.245 1968.695 ;
        RECT 3513.675 1968.415 3513.955 1968.695 ;
        RECT 3514.385 1968.415 3514.665 1968.695 ;
        RECT 3515.095 1968.415 3515.375 1968.695 ;
        RECT 3515.805 1968.415 3516.085 1968.695 ;
        RECT 3516.515 1968.415 3516.795 1968.695 ;
        RECT 3517.225 1968.415 3517.505 1968.695 ;
        RECT 3517.935 1968.415 3518.215 1968.695 ;
        RECT 3518.645 1968.415 3518.925 1968.695 ;
        RECT 3519.355 1968.415 3519.635 1968.695 ;
        RECT 3520.065 1968.415 3520.345 1968.695 ;
        RECT 3520.775 1968.415 3521.055 1968.695 ;
        RECT 3521.485 1968.415 3521.765 1968.695 ;
        RECT 3512.255 1967.705 3512.535 1967.985 ;
        RECT 3512.965 1967.705 3513.245 1967.985 ;
        RECT 3513.675 1967.705 3513.955 1967.985 ;
        RECT 3514.385 1967.705 3514.665 1967.985 ;
        RECT 3515.095 1967.705 3515.375 1967.985 ;
        RECT 3515.805 1967.705 3516.085 1967.985 ;
        RECT 3516.515 1967.705 3516.795 1967.985 ;
        RECT 3517.225 1967.705 3517.505 1967.985 ;
        RECT 3517.935 1967.705 3518.215 1967.985 ;
        RECT 3518.645 1967.705 3518.925 1967.985 ;
        RECT 3519.355 1967.705 3519.635 1967.985 ;
        RECT 3520.065 1967.705 3520.345 1967.985 ;
        RECT 3520.775 1967.705 3521.055 1967.985 ;
        RECT 3521.485 1967.705 3521.765 1967.985 ;
        RECT 3512.255 1966.995 3512.535 1967.275 ;
        RECT 3512.965 1966.995 3513.245 1967.275 ;
        RECT 3513.675 1966.995 3513.955 1967.275 ;
        RECT 3514.385 1966.995 3514.665 1967.275 ;
        RECT 3515.095 1966.995 3515.375 1967.275 ;
        RECT 3515.805 1966.995 3516.085 1967.275 ;
        RECT 3516.515 1966.995 3516.795 1967.275 ;
        RECT 3517.225 1966.995 3517.505 1967.275 ;
        RECT 3517.935 1966.995 3518.215 1967.275 ;
        RECT 3518.645 1966.995 3518.925 1967.275 ;
        RECT 3519.355 1966.995 3519.635 1967.275 ;
        RECT 3520.065 1966.995 3520.345 1967.275 ;
        RECT 3520.775 1966.995 3521.055 1967.275 ;
        RECT 3521.485 1966.995 3521.765 1967.275 ;
        RECT 3512.255 1966.285 3512.535 1966.565 ;
        RECT 3512.965 1966.285 3513.245 1966.565 ;
        RECT 3513.675 1966.285 3513.955 1966.565 ;
        RECT 3514.385 1966.285 3514.665 1966.565 ;
        RECT 3515.095 1966.285 3515.375 1966.565 ;
        RECT 3515.805 1966.285 3516.085 1966.565 ;
        RECT 3516.515 1966.285 3516.795 1966.565 ;
        RECT 3517.225 1966.285 3517.505 1966.565 ;
        RECT 3517.935 1966.285 3518.215 1966.565 ;
        RECT 3518.645 1966.285 3518.925 1966.565 ;
        RECT 3519.355 1966.285 3519.635 1966.565 ;
        RECT 3520.065 1966.285 3520.345 1966.565 ;
        RECT 3520.775 1966.285 3521.055 1966.565 ;
        RECT 3521.485 1966.285 3521.765 1966.565 ;
        RECT 3512.255 1965.575 3512.535 1965.855 ;
        RECT 3512.965 1965.575 3513.245 1965.855 ;
        RECT 3513.675 1965.575 3513.955 1965.855 ;
        RECT 3514.385 1965.575 3514.665 1965.855 ;
        RECT 3515.095 1965.575 3515.375 1965.855 ;
        RECT 3515.805 1965.575 3516.085 1965.855 ;
        RECT 3516.515 1965.575 3516.795 1965.855 ;
        RECT 3517.225 1965.575 3517.505 1965.855 ;
        RECT 3517.935 1965.575 3518.215 1965.855 ;
        RECT 3518.645 1965.575 3518.925 1965.855 ;
        RECT 3519.355 1965.575 3519.635 1965.855 ;
        RECT 3520.065 1965.575 3520.345 1965.855 ;
        RECT 3520.775 1965.575 3521.055 1965.855 ;
        RECT 3521.485 1965.575 3521.765 1965.855 ;
        RECT 3512.255 1964.865 3512.535 1965.145 ;
        RECT 3512.965 1964.865 3513.245 1965.145 ;
        RECT 3513.675 1964.865 3513.955 1965.145 ;
        RECT 3514.385 1964.865 3514.665 1965.145 ;
        RECT 3515.095 1964.865 3515.375 1965.145 ;
        RECT 3515.805 1964.865 3516.085 1965.145 ;
        RECT 3516.515 1964.865 3516.795 1965.145 ;
        RECT 3517.225 1964.865 3517.505 1965.145 ;
        RECT 3517.935 1964.865 3518.215 1965.145 ;
        RECT 3518.645 1964.865 3518.925 1965.145 ;
        RECT 3519.355 1964.865 3519.635 1965.145 ;
        RECT 3520.065 1964.865 3520.345 1965.145 ;
        RECT 3520.775 1964.865 3521.055 1965.145 ;
        RECT 3521.485 1964.865 3521.765 1965.145 ;
        RECT 3512.255 1964.155 3512.535 1964.435 ;
        RECT 3512.965 1964.155 3513.245 1964.435 ;
        RECT 3513.675 1964.155 3513.955 1964.435 ;
        RECT 3514.385 1964.155 3514.665 1964.435 ;
        RECT 3515.095 1964.155 3515.375 1964.435 ;
        RECT 3515.805 1964.155 3516.085 1964.435 ;
        RECT 3516.515 1964.155 3516.795 1964.435 ;
        RECT 3517.225 1964.155 3517.505 1964.435 ;
        RECT 3517.935 1964.155 3518.215 1964.435 ;
        RECT 3518.645 1964.155 3518.925 1964.435 ;
        RECT 3519.355 1964.155 3519.635 1964.435 ;
        RECT 3520.065 1964.155 3520.345 1964.435 ;
        RECT 3520.775 1964.155 3521.055 1964.435 ;
        RECT 3521.485 1964.155 3521.765 1964.435 ;
        RECT 3512.200 1960.270 3512.480 1960.550 ;
        RECT 3512.910 1960.270 3513.190 1960.550 ;
        RECT 3513.620 1960.270 3513.900 1960.550 ;
        RECT 3514.330 1960.270 3514.610 1960.550 ;
        RECT 3515.040 1960.270 3515.320 1960.550 ;
        RECT 3515.750 1960.270 3516.030 1960.550 ;
        RECT 3516.460 1960.270 3516.740 1960.550 ;
        RECT 3517.170 1960.270 3517.450 1960.550 ;
        RECT 3517.880 1960.270 3518.160 1960.550 ;
        RECT 3518.590 1960.270 3518.870 1960.550 ;
        RECT 3519.300 1960.270 3519.580 1960.550 ;
        RECT 3520.010 1960.270 3520.290 1960.550 ;
        RECT 3520.720 1960.270 3521.000 1960.550 ;
        RECT 3521.430 1960.270 3521.710 1960.550 ;
        RECT 3512.200 1959.560 3512.480 1959.840 ;
        RECT 3512.910 1959.560 3513.190 1959.840 ;
        RECT 3513.620 1959.560 3513.900 1959.840 ;
        RECT 3514.330 1959.560 3514.610 1959.840 ;
        RECT 3515.040 1959.560 3515.320 1959.840 ;
        RECT 3515.750 1959.560 3516.030 1959.840 ;
        RECT 3516.460 1959.560 3516.740 1959.840 ;
        RECT 3517.170 1959.560 3517.450 1959.840 ;
        RECT 3517.880 1959.560 3518.160 1959.840 ;
        RECT 3518.590 1959.560 3518.870 1959.840 ;
        RECT 3519.300 1959.560 3519.580 1959.840 ;
        RECT 3520.010 1959.560 3520.290 1959.840 ;
        RECT 3520.720 1959.560 3521.000 1959.840 ;
        RECT 3521.430 1959.560 3521.710 1959.840 ;
        RECT 3512.200 1958.850 3512.480 1959.130 ;
        RECT 3512.910 1958.850 3513.190 1959.130 ;
        RECT 3513.620 1958.850 3513.900 1959.130 ;
        RECT 3514.330 1958.850 3514.610 1959.130 ;
        RECT 3515.040 1958.850 3515.320 1959.130 ;
        RECT 3515.750 1958.850 3516.030 1959.130 ;
        RECT 3516.460 1958.850 3516.740 1959.130 ;
        RECT 3517.170 1958.850 3517.450 1959.130 ;
        RECT 3517.880 1958.850 3518.160 1959.130 ;
        RECT 3518.590 1958.850 3518.870 1959.130 ;
        RECT 3519.300 1958.850 3519.580 1959.130 ;
        RECT 3520.010 1958.850 3520.290 1959.130 ;
        RECT 3520.720 1958.850 3521.000 1959.130 ;
        RECT 3521.430 1958.850 3521.710 1959.130 ;
        RECT 3512.200 1958.140 3512.480 1958.420 ;
        RECT 3512.910 1958.140 3513.190 1958.420 ;
        RECT 3513.620 1958.140 3513.900 1958.420 ;
        RECT 3514.330 1958.140 3514.610 1958.420 ;
        RECT 3515.040 1958.140 3515.320 1958.420 ;
        RECT 3515.750 1958.140 3516.030 1958.420 ;
        RECT 3516.460 1958.140 3516.740 1958.420 ;
        RECT 3517.170 1958.140 3517.450 1958.420 ;
        RECT 3517.880 1958.140 3518.160 1958.420 ;
        RECT 3518.590 1958.140 3518.870 1958.420 ;
        RECT 3519.300 1958.140 3519.580 1958.420 ;
        RECT 3520.010 1958.140 3520.290 1958.420 ;
        RECT 3520.720 1958.140 3521.000 1958.420 ;
        RECT 3521.430 1958.140 3521.710 1958.420 ;
        RECT 3512.200 1957.430 3512.480 1957.710 ;
        RECT 3512.910 1957.430 3513.190 1957.710 ;
        RECT 3513.620 1957.430 3513.900 1957.710 ;
        RECT 3514.330 1957.430 3514.610 1957.710 ;
        RECT 3515.040 1957.430 3515.320 1957.710 ;
        RECT 3515.750 1957.430 3516.030 1957.710 ;
        RECT 3516.460 1957.430 3516.740 1957.710 ;
        RECT 3517.170 1957.430 3517.450 1957.710 ;
        RECT 3517.880 1957.430 3518.160 1957.710 ;
        RECT 3518.590 1957.430 3518.870 1957.710 ;
        RECT 3519.300 1957.430 3519.580 1957.710 ;
        RECT 3520.010 1957.430 3520.290 1957.710 ;
        RECT 3520.720 1957.430 3521.000 1957.710 ;
        RECT 3521.430 1957.430 3521.710 1957.710 ;
        RECT 3512.200 1956.720 3512.480 1957.000 ;
        RECT 3512.910 1956.720 3513.190 1957.000 ;
        RECT 3513.620 1956.720 3513.900 1957.000 ;
        RECT 3514.330 1956.720 3514.610 1957.000 ;
        RECT 3515.040 1956.720 3515.320 1957.000 ;
        RECT 3515.750 1956.720 3516.030 1957.000 ;
        RECT 3516.460 1956.720 3516.740 1957.000 ;
        RECT 3517.170 1956.720 3517.450 1957.000 ;
        RECT 3517.880 1956.720 3518.160 1957.000 ;
        RECT 3518.590 1956.720 3518.870 1957.000 ;
        RECT 3519.300 1956.720 3519.580 1957.000 ;
        RECT 3520.010 1956.720 3520.290 1957.000 ;
        RECT 3520.720 1956.720 3521.000 1957.000 ;
        RECT 3521.430 1956.720 3521.710 1957.000 ;
        RECT 3512.200 1956.010 3512.480 1956.290 ;
        RECT 3512.910 1956.010 3513.190 1956.290 ;
        RECT 3513.620 1956.010 3513.900 1956.290 ;
        RECT 3514.330 1956.010 3514.610 1956.290 ;
        RECT 3515.040 1956.010 3515.320 1956.290 ;
        RECT 3515.750 1956.010 3516.030 1956.290 ;
        RECT 3516.460 1956.010 3516.740 1956.290 ;
        RECT 3517.170 1956.010 3517.450 1956.290 ;
        RECT 3517.880 1956.010 3518.160 1956.290 ;
        RECT 3518.590 1956.010 3518.870 1956.290 ;
        RECT 3519.300 1956.010 3519.580 1956.290 ;
        RECT 3520.010 1956.010 3520.290 1956.290 ;
        RECT 3520.720 1956.010 3521.000 1956.290 ;
        RECT 3521.430 1956.010 3521.710 1956.290 ;
        RECT 3512.200 1955.300 3512.480 1955.580 ;
        RECT 3512.910 1955.300 3513.190 1955.580 ;
        RECT 3513.620 1955.300 3513.900 1955.580 ;
        RECT 3514.330 1955.300 3514.610 1955.580 ;
        RECT 3515.040 1955.300 3515.320 1955.580 ;
        RECT 3515.750 1955.300 3516.030 1955.580 ;
        RECT 3516.460 1955.300 3516.740 1955.580 ;
        RECT 3517.170 1955.300 3517.450 1955.580 ;
        RECT 3517.880 1955.300 3518.160 1955.580 ;
        RECT 3518.590 1955.300 3518.870 1955.580 ;
        RECT 3519.300 1955.300 3519.580 1955.580 ;
        RECT 3520.010 1955.300 3520.290 1955.580 ;
        RECT 3520.720 1955.300 3521.000 1955.580 ;
        RECT 3521.430 1955.300 3521.710 1955.580 ;
        RECT 3512.200 1954.590 3512.480 1954.870 ;
        RECT 3512.910 1954.590 3513.190 1954.870 ;
        RECT 3513.620 1954.590 3513.900 1954.870 ;
        RECT 3514.330 1954.590 3514.610 1954.870 ;
        RECT 3515.040 1954.590 3515.320 1954.870 ;
        RECT 3515.750 1954.590 3516.030 1954.870 ;
        RECT 3516.460 1954.590 3516.740 1954.870 ;
        RECT 3517.170 1954.590 3517.450 1954.870 ;
        RECT 3517.880 1954.590 3518.160 1954.870 ;
        RECT 3518.590 1954.590 3518.870 1954.870 ;
        RECT 3519.300 1954.590 3519.580 1954.870 ;
        RECT 3520.010 1954.590 3520.290 1954.870 ;
        RECT 3520.720 1954.590 3521.000 1954.870 ;
        RECT 3521.430 1954.590 3521.710 1954.870 ;
        RECT 3512.200 1953.880 3512.480 1954.160 ;
        RECT 3512.910 1953.880 3513.190 1954.160 ;
        RECT 3513.620 1953.880 3513.900 1954.160 ;
        RECT 3514.330 1953.880 3514.610 1954.160 ;
        RECT 3515.040 1953.880 3515.320 1954.160 ;
        RECT 3515.750 1953.880 3516.030 1954.160 ;
        RECT 3516.460 1953.880 3516.740 1954.160 ;
        RECT 3517.170 1953.880 3517.450 1954.160 ;
        RECT 3517.880 1953.880 3518.160 1954.160 ;
        RECT 3518.590 1953.880 3518.870 1954.160 ;
        RECT 3519.300 1953.880 3519.580 1954.160 ;
        RECT 3520.010 1953.880 3520.290 1954.160 ;
        RECT 3520.720 1953.880 3521.000 1954.160 ;
        RECT 3521.430 1953.880 3521.710 1954.160 ;
        RECT 3512.200 1953.170 3512.480 1953.450 ;
        RECT 3512.910 1953.170 3513.190 1953.450 ;
        RECT 3513.620 1953.170 3513.900 1953.450 ;
        RECT 3514.330 1953.170 3514.610 1953.450 ;
        RECT 3515.040 1953.170 3515.320 1953.450 ;
        RECT 3515.750 1953.170 3516.030 1953.450 ;
        RECT 3516.460 1953.170 3516.740 1953.450 ;
        RECT 3517.170 1953.170 3517.450 1953.450 ;
        RECT 3517.880 1953.170 3518.160 1953.450 ;
        RECT 3518.590 1953.170 3518.870 1953.450 ;
        RECT 3519.300 1953.170 3519.580 1953.450 ;
        RECT 3520.010 1953.170 3520.290 1953.450 ;
        RECT 3520.720 1953.170 3521.000 1953.450 ;
        RECT 3521.430 1953.170 3521.710 1953.450 ;
        RECT 3512.200 1952.460 3512.480 1952.740 ;
        RECT 3512.910 1952.460 3513.190 1952.740 ;
        RECT 3513.620 1952.460 3513.900 1952.740 ;
        RECT 3514.330 1952.460 3514.610 1952.740 ;
        RECT 3515.040 1952.460 3515.320 1952.740 ;
        RECT 3515.750 1952.460 3516.030 1952.740 ;
        RECT 3516.460 1952.460 3516.740 1952.740 ;
        RECT 3517.170 1952.460 3517.450 1952.740 ;
        RECT 3517.880 1952.460 3518.160 1952.740 ;
        RECT 3518.590 1952.460 3518.870 1952.740 ;
        RECT 3519.300 1952.460 3519.580 1952.740 ;
        RECT 3520.010 1952.460 3520.290 1952.740 ;
        RECT 3520.720 1952.460 3521.000 1952.740 ;
        RECT 3521.430 1952.460 3521.710 1952.740 ;
        RECT 3512.200 1951.750 3512.480 1952.030 ;
        RECT 3512.910 1951.750 3513.190 1952.030 ;
        RECT 3513.620 1951.750 3513.900 1952.030 ;
        RECT 3514.330 1951.750 3514.610 1952.030 ;
        RECT 3515.040 1951.750 3515.320 1952.030 ;
        RECT 3515.750 1951.750 3516.030 1952.030 ;
        RECT 3516.460 1951.750 3516.740 1952.030 ;
        RECT 3517.170 1951.750 3517.450 1952.030 ;
        RECT 3517.880 1951.750 3518.160 1952.030 ;
        RECT 3518.590 1951.750 3518.870 1952.030 ;
        RECT 3519.300 1951.750 3519.580 1952.030 ;
        RECT 3520.010 1951.750 3520.290 1952.030 ;
        RECT 3520.720 1951.750 3521.000 1952.030 ;
        RECT 3521.430 1951.750 3521.710 1952.030 ;
        RECT 369.330 702.970 369.610 703.250 ;
        RECT 370.040 702.970 370.320 703.250 ;
        RECT 370.750 702.970 371.030 703.250 ;
        RECT 371.460 702.970 371.740 703.250 ;
        RECT 372.170 702.970 372.450 703.250 ;
        RECT 372.880 702.970 373.160 703.250 ;
        RECT 373.590 702.970 373.870 703.250 ;
        RECT 374.300 702.970 374.580 703.250 ;
        RECT 375.010 702.970 375.290 703.250 ;
        RECT 375.720 702.970 376.000 703.250 ;
        RECT 376.430 702.970 376.710 703.250 ;
        RECT 369.330 702.260 369.610 702.540 ;
        RECT 370.040 702.260 370.320 702.540 ;
        RECT 370.750 702.260 371.030 702.540 ;
        RECT 371.460 702.260 371.740 702.540 ;
        RECT 372.170 702.260 372.450 702.540 ;
        RECT 372.880 702.260 373.160 702.540 ;
        RECT 373.590 702.260 373.870 702.540 ;
        RECT 374.300 702.260 374.580 702.540 ;
        RECT 375.010 702.260 375.290 702.540 ;
        RECT 375.720 702.260 376.000 702.540 ;
        RECT 376.430 702.260 376.710 702.540 ;
        RECT 369.330 701.550 369.610 701.830 ;
        RECT 370.040 701.550 370.320 701.830 ;
        RECT 370.750 701.550 371.030 701.830 ;
        RECT 371.460 701.550 371.740 701.830 ;
        RECT 372.170 701.550 372.450 701.830 ;
        RECT 372.880 701.550 373.160 701.830 ;
        RECT 373.590 701.550 373.870 701.830 ;
        RECT 374.300 701.550 374.580 701.830 ;
        RECT 375.010 701.550 375.290 701.830 ;
        RECT 375.720 701.550 376.000 701.830 ;
        RECT 376.430 701.550 376.710 701.830 ;
        RECT 369.330 700.840 369.610 701.120 ;
        RECT 370.040 700.840 370.320 701.120 ;
        RECT 370.750 700.840 371.030 701.120 ;
        RECT 371.460 700.840 371.740 701.120 ;
        RECT 372.170 700.840 372.450 701.120 ;
        RECT 372.880 700.840 373.160 701.120 ;
        RECT 373.590 700.840 373.870 701.120 ;
        RECT 374.300 700.840 374.580 701.120 ;
        RECT 375.010 700.840 375.290 701.120 ;
        RECT 375.720 700.840 376.000 701.120 ;
        RECT 376.430 700.840 376.710 701.120 ;
        RECT 369.330 700.130 369.610 700.410 ;
        RECT 370.040 700.130 370.320 700.410 ;
        RECT 370.750 700.130 371.030 700.410 ;
        RECT 371.460 700.130 371.740 700.410 ;
        RECT 372.170 700.130 372.450 700.410 ;
        RECT 372.880 700.130 373.160 700.410 ;
        RECT 373.590 700.130 373.870 700.410 ;
        RECT 374.300 700.130 374.580 700.410 ;
        RECT 375.010 700.130 375.290 700.410 ;
        RECT 375.720 700.130 376.000 700.410 ;
        RECT 376.430 700.130 376.710 700.410 ;
        RECT 369.330 699.420 369.610 699.700 ;
        RECT 370.040 699.420 370.320 699.700 ;
        RECT 370.750 699.420 371.030 699.700 ;
        RECT 371.460 699.420 371.740 699.700 ;
        RECT 372.170 699.420 372.450 699.700 ;
        RECT 372.880 699.420 373.160 699.700 ;
        RECT 373.590 699.420 373.870 699.700 ;
        RECT 374.300 699.420 374.580 699.700 ;
        RECT 375.010 699.420 375.290 699.700 ;
        RECT 375.720 699.420 376.000 699.700 ;
        RECT 376.430 699.420 376.710 699.700 ;
        RECT 369.330 698.710 369.610 698.990 ;
        RECT 370.040 698.710 370.320 698.990 ;
        RECT 370.750 698.710 371.030 698.990 ;
        RECT 371.460 698.710 371.740 698.990 ;
        RECT 372.170 698.710 372.450 698.990 ;
        RECT 372.880 698.710 373.160 698.990 ;
        RECT 373.590 698.710 373.870 698.990 ;
        RECT 374.300 698.710 374.580 698.990 ;
        RECT 375.010 698.710 375.290 698.990 ;
        RECT 375.720 698.710 376.000 698.990 ;
        RECT 376.430 698.710 376.710 698.990 ;
        RECT 369.330 698.000 369.610 698.280 ;
        RECT 370.040 698.000 370.320 698.280 ;
        RECT 370.750 698.000 371.030 698.280 ;
        RECT 371.460 698.000 371.740 698.280 ;
        RECT 372.170 698.000 372.450 698.280 ;
        RECT 372.880 698.000 373.160 698.280 ;
        RECT 373.590 698.000 373.870 698.280 ;
        RECT 374.300 698.000 374.580 698.280 ;
        RECT 375.010 698.000 375.290 698.280 ;
        RECT 375.720 698.000 376.000 698.280 ;
        RECT 376.430 698.000 376.710 698.280 ;
        RECT 369.330 697.290 369.610 697.570 ;
        RECT 370.040 697.290 370.320 697.570 ;
        RECT 370.750 697.290 371.030 697.570 ;
        RECT 371.460 697.290 371.740 697.570 ;
        RECT 372.170 697.290 372.450 697.570 ;
        RECT 372.880 697.290 373.160 697.570 ;
        RECT 373.590 697.290 373.870 697.570 ;
        RECT 374.300 697.290 374.580 697.570 ;
        RECT 375.010 697.290 375.290 697.570 ;
        RECT 375.720 697.290 376.000 697.570 ;
        RECT 376.430 697.290 376.710 697.570 ;
        RECT 369.330 696.580 369.610 696.860 ;
        RECT 370.040 696.580 370.320 696.860 ;
        RECT 370.750 696.580 371.030 696.860 ;
        RECT 371.460 696.580 371.740 696.860 ;
        RECT 372.170 696.580 372.450 696.860 ;
        RECT 372.880 696.580 373.160 696.860 ;
        RECT 373.590 696.580 373.870 696.860 ;
        RECT 374.300 696.580 374.580 696.860 ;
        RECT 375.010 696.580 375.290 696.860 ;
        RECT 375.720 696.580 376.000 696.860 ;
        RECT 376.430 696.580 376.710 696.860 ;
        RECT 369.330 695.870 369.610 696.150 ;
        RECT 370.040 695.870 370.320 696.150 ;
        RECT 370.750 695.870 371.030 696.150 ;
        RECT 371.460 695.870 371.740 696.150 ;
        RECT 372.170 695.870 372.450 696.150 ;
        RECT 372.880 695.870 373.160 696.150 ;
        RECT 373.590 695.870 373.870 696.150 ;
        RECT 374.300 695.870 374.580 696.150 ;
        RECT 375.010 695.870 375.290 696.150 ;
        RECT 375.720 695.870 376.000 696.150 ;
        RECT 376.430 695.870 376.710 696.150 ;
        RECT 369.330 695.160 369.610 695.440 ;
        RECT 370.040 695.160 370.320 695.440 ;
        RECT 370.750 695.160 371.030 695.440 ;
        RECT 371.460 695.160 371.740 695.440 ;
        RECT 372.170 695.160 372.450 695.440 ;
        RECT 372.880 695.160 373.160 695.440 ;
        RECT 373.590 695.160 373.870 695.440 ;
        RECT 374.300 695.160 374.580 695.440 ;
        RECT 375.010 695.160 375.290 695.440 ;
        RECT 375.720 695.160 376.000 695.440 ;
        RECT 376.430 695.160 376.710 695.440 ;
        RECT 369.330 694.450 369.610 694.730 ;
        RECT 370.040 694.450 370.320 694.730 ;
        RECT 370.750 694.450 371.030 694.730 ;
        RECT 371.460 694.450 371.740 694.730 ;
        RECT 372.170 694.450 372.450 694.730 ;
        RECT 372.880 694.450 373.160 694.730 ;
        RECT 373.590 694.450 373.870 694.730 ;
        RECT 374.300 694.450 374.580 694.730 ;
        RECT 375.010 694.450 375.290 694.730 ;
        RECT 375.720 694.450 376.000 694.730 ;
        RECT 376.430 694.450 376.710 694.730 ;
        RECT 369.275 690.565 369.555 690.845 ;
        RECT 369.985 690.565 370.265 690.845 ;
        RECT 370.695 690.565 370.975 690.845 ;
        RECT 371.405 690.565 371.685 690.845 ;
        RECT 372.115 690.565 372.395 690.845 ;
        RECT 372.825 690.565 373.105 690.845 ;
        RECT 373.535 690.565 373.815 690.845 ;
        RECT 374.245 690.565 374.525 690.845 ;
        RECT 374.955 690.565 375.235 690.845 ;
        RECT 375.665 690.565 375.945 690.845 ;
        RECT 376.375 690.565 376.655 690.845 ;
        RECT 369.275 689.855 369.555 690.135 ;
        RECT 369.985 689.855 370.265 690.135 ;
        RECT 370.695 689.855 370.975 690.135 ;
        RECT 371.405 689.855 371.685 690.135 ;
        RECT 372.115 689.855 372.395 690.135 ;
        RECT 372.825 689.855 373.105 690.135 ;
        RECT 373.535 689.855 373.815 690.135 ;
        RECT 374.245 689.855 374.525 690.135 ;
        RECT 374.955 689.855 375.235 690.135 ;
        RECT 375.665 689.855 375.945 690.135 ;
        RECT 376.375 689.855 376.655 690.135 ;
        RECT 369.275 689.145 369.555 689.425 ;
        RECT 369.985 689.145 370.265 689.425 ;
        RECT 370.695 689.145 370.975 689.425 ;
        RECT 371.405 689.145 371.685 689.425 ;
        RECT 372.115 689.145 372.395 689.425 ;
        RECT 372.825 689.145 373.105 689.425 ;
        RECT 373.535 689.145 373.815 689.425 ;
        RECT 374.245 689.145 374.525 689.425 ;
        RECT 374.955 689.145 375.235 689.425 ;
        RECT 375.665 689.145 375.945 689.425 ;
        RECT 376.375 689.145 376.655 689.425 ;
        RECT 369.275 688.435 369.555 688.715 ;
        RECT 369.985 688.435 370.265 688.715 ;
        RECT 370.695 688.435 370.975 688.715 ;
        RECT 371.405 688.435 371.685 688.715 ;
        RECT 372.115 688.435 372.395 688.715 ;
        RECT 372.825 688.435 373.105 688.715 ;
        RECT 373.535 688.435 373.815 688.715 ;
        RECT 374.245 688.435 374.525 688.715 ;
        RECT 374.955 688.435 375.235 688.715 ;
        RECT 375.665 688.435 375.945 688.715 ;
        RECT 376.375 688.435 376.655 688.715 ;
        RECT 369.275 687.725 369.555 688.005 ;
        RECT 369.985 687.725 370.265 688.005 ;
        RECT 370.695 687.725 370.975 688.005 ;
        RECT 371.405 687.725 371.685 688.005 ;
        RECT 372.115 687.725 372.395 688.005 ;
        RECT 372.825 687.725 373.105 688.005 ;
        RECT 373.535 687.725 373.815 688.005 ;
        RECT 374.245 687.725 374.525 688.005 ;
        RECT 374.955 687.725 375.235 688.005 ;
        RECT 375.665 687.725 375.945 688.005 ;
        RECT 376.375 687.725 376.655 688.005 ;
        RECT 369.275 687.015 369.555 687.295 ;
        RECT 369.985 687.015 370.265 687.295 ;
        RECT 370.695 687.015 370.975 687.295 ;
        RECT 371.405 687.015 371.685 687.295 ;
        RECT 372.115 687.015 372.395 687.295 ;
        RECT 372.825 687.015 373.105 687.295 ;
        RECT 373.535 687.015 373.815 687.295 ;
        RECT 374.245 687.015 374.525 687.295 ;
        RECT 374.955 687.015 375.235 687.295 ;
        RECT 375.665 687.015 375.945 687.295 ;
        RECT 376.375 687.015 376.655 687.295 ;
        RECT 369.275 686.305 369.555 686.585 ;
        RECT 369.985 686.305 370.265 686.585 ;
        RECT 370.695 686.305 370.975 686.585 ;
        RECT 371.405 686.305 371.685 686.585 ;
        RECT 372.115 686.305 372.395 686.585 ;
        RECT 372.825 686.305 373.105 686.585 ;
        RECT 373.535 686.305 373.815 686.585 ;
        RECT 374.245 686.305 374.525 686.585 ;
        RECT 374.955 686.305 375.235 686.585 ;
        RECT 375.665 686.305 375.945 686.585 ;
        RECT 376.375 686.305 376.655 686.585 ;
        RECT 369.275 685.595 369.555 685.875 ;
        RECT 369.985 685.595 370.265 685.875 ;
        RECT 370.695 685.595 370.975 685.875 ;
        RECT 371.405 685.595 371.685 685.875 ;
        RECT 372.115 685.595 372.395 685.875 ;
        RECT 372.825 685.595 373.105 685.875 ;
        RECT 373.535 685.595 373.815 685.875 ;
        RECT 374.245 685.595 374.525 685.875 ;
        RECT 374.955 685.595 375.235 685.875 ;
        RECT 375.665 685.595 375.945 685.875 ;
        RECT 376.375 685.595 376.655 685.875 ;
        RECT 369.275 684.885 369.555 685.165 ;
        RECT 369.985 684.885 370.265 685.165 ;
        RECT 370.695 684.885 370.975 685.165 ;
        RECT 371.405 684.885 371.685 685.165 ;
        RECT 372.115 684.885 372.395 685.165 ;
        RECT 372.825 684.885 373.105 685.165 ;
        RECT 373.535 684.885 373.815 685.165 ;
        RECT 374.245 684.885 374.525 685.165 ;
        RECT 374.955 684.885 375.235 685.165 ;
        RECT 375.665 684.885 375.945 685.165 ;
        RECT 376.375 684.885 376.655 685.165 ;
        RECT 369.275 684.175 369.555 684.455 ;
        RECT 369.985 684.175 370.265 684.455 ;
        RECT 370.695 684.175 370.975 684.455 ;
        RECT 371.405 684.175 371.685 684.455 ;
        RECT 372.115 684.175 372.395 684.455 ;
        RECT 372.825 684.175 373.105 684.455 ;
        RECT 373.535 684.175 373.815 684.455 ;
        RECT 374.245 684.175 374.525 684.455 ;
        RECT 374.955 684.175 375.235 684.455 ;
        RECT 375.665 684.175 375.945 684.455 ;
        RECT 376.375 684.175 376.655 684.455 ;
        RECT 369.275 683.465 369.555 683.745 ;
        RECT 369.985 683.465 370.265 683.745 ;
        RECT 370.695 683.465 370.975 683.745 ;
        RECT 371.405 683.465 371.685 683.745 ;
        RECT 372.115 683.465 372.395 683.745 ;
        RECT 372.825 683.465 373.105 683.745 ;
        RECT 373.535 683.465 373.815 683.745 ;
        RECT 374.245 683.465 374.525 683.745 ;
        RECT 374.955 683.465 375.235 683.745 ;
        RECT 375.665 683.465 375.945 683.745 ;
        RECT 376.375 683.465 376.655 683.745 ;
        RECT 369.275 682.755 369.555 683.035 ;
        RECT 369.985 682.755 370.265 683.035 ;
        RECT 370.695 682.755 370.975 683.035 ;
        RECT 371.405 682.755 371.685 683.035 ;
        RECT 372.115 682.755 372.395 683.035 ;
        RECT 372.825 682.755 373.105 683.035 ;
        RECT 373.535 682.755 373.815 683.035 ;
        RECT 374.245 682.755 374.525 683.035 ;
        RECT 374.955 682.755 375.235 683.035 ;
        RECT 375.665 682.755 375.945 683.035 ;
        RECT 376.375 682.755 376.655 683.035 ;
        RECT 369.275 682.045 369.555 682.325 ;
        RECT 369.985 682.045 370.265 682.325 ;
        RECT 370.695 682.045 370.975 682.325 ;
        RECT 371.405 682.045 371.685 682.325 ;
        RECT 372.115 682.045 372.395 682.325 ;
        RECT 372.825 682.045 373.105 682.325 ;
        RECT 373.535 682.045 373.815 682.325 ;
        RECT 374.245 682.045 374.525 682.325 ;
        RECT 374.955 682.045 375.235 682.325 ;
        RECT 375.665 682.045 375.945 682.325 ;
        RECT 376.375 682.045 376.655 682.325 ;
        RECT 369.275 681.335 369.555 681.615 ;
        RECT 369.985 681.335 370.265 681.615 ;
        RECT 370.695 681.335 370.975 681.615 ;
        RECT 371.405 681.335 371.685 681.615 ;
        RECT 372.115 681.335 372.395 681.615 ;
        RECT 372.825 681.335 373.105 681.615 ;
        RECT 373.535 681.335 373.815 681.615 ;
        RECT 374.245 681.335 374.525 681.615 ;
        RECT 374.955 681.335 375.235 681.615 ;
        RECT 375.665 681.335 375.945 681.615 ;
        RECT 376.375 681.335 376.655 681.615 ;
        RECT 369.275 678.715 369.555 678.995 ;
        RECT 369.985 678.715 370.265 678.995 ;
        RECT 370.695 678.715 370.975 678.995 ;
        RECT 371.405 678.715 371.685 678.995 ;
        RECT 372.115 678.715 372.395 678.995 ;
        RECT 372.825 678.715 373.105 678.995 ;
        RECT 373.535 678.715 373.815 678.995 ;
        RECT 374.245 678.715 374.525 678.995 ;
        RECT 374.955 678.715 375.235 678.995 ;
        RECT 375.665 678.715 375.945 678.995 ;
        RECT 376.375 678.715 376.655 678.995 ;
        RECT 369.275 678.005 369.555 678.285 ;
        RECT 369.985 678.005 370.265 678.285 ;
        RECT 370.695 678.005 370.975 678.285 ;
        RECT 371.405 678.005 371.685 678.285 ;
        RECT 372.115 678.005 372.395 678.285 ;
        RECT 372.825 678.005 373.105 678.285 ;
        RECT 373.535 678.005 373.815 678.285 ;
        RECT 374.245 678.005 374.525 678.285 ;
        RECT 374.955 678.005 375.235 678.285 ;
        RECT 375.665 678.005 375.945 678.285 ;
        RECT 376.375 678.005 376.655 678.285 ;
        RECT 369.275 677.295 369.555 677.575 ;
        RECT 369.985 677.295 370.265 677.575 ;
        RECT 370.695 677.295 370.975 677.575 ;
        RECT 371.405 677.295 371.685 677.575 ;
        RECT 372.115 677.295 372.395 677.575 ;
        RECT 372.825 677.295 373.105 677.575 ;
        RECT 373.535 677.295 373.815 677.575 ;
        RECT 374.245 677.295 374.525 677.575 ;
        RECT 374.955 677.295 375.235 677.575 ;
        RECT 375.665 677.295 375.945 677.575 ;
        RECT 376.375 677.295 376.655 677.575 ;
        RECT 369.275 676.585 369.555 676.865 ;
        RECT 369.985 676.585 370.265 676.865 ;
        RECT 370.695 676.585 370.975 676.865 ;
        RECT 371.405 676.585 371.685 676.865 ;
        RECT 372.115 676.585 372.395 676.865 ;
        RECT 372.825 676.585 373.105 676.865 ;
        RECT 373.535 676.585 373.815 676.865 ;
        RECT 374.245 676.585 374.525 676.865 ;
        RECT 374.955 676.585 375.235 676.865 ;
        RECT 375.665 676.585 375.945 676.865 ;
        RECT 376.375 676.585 376.655 676.865 ;
        RECT 369.275 675.875 369.555 676.155 ;
        RECT 369.985 675.875 370.265 676.155 ;
        RECT 370.695 675.875 370.975 676.155 ;
        RECT 371.405 675.875 371.685 676.155 ;
        RECT 372.115 675.875 372.395 676.155 ;
        RECT 372.825 675.875 373.105 676.155 ;
        RECT 373.535 675.875 373.815 676.155 ;
        RECT 374.245 675.875 374.525 676.155 ;
        RECT 374.955 675.875 375.235 676.155 ;
        RECT 375.665 675.875 375.945 676.155 ;
        RECT 376.375 675.875 376.655 676.155 ;
        RECT 369.275 675.165 369.555 675.445 ;
        RECT 369.985 675.165 370.265 675.445 ;
        RECT 370.695 675.165 370.975 675.445 ;
        RECT 371.405 675.165 371.685 675.445 ;
        RECT 372.115 675.165 372.395 675.445 ;
        RECT 372.825 675.165 373.105 675.445 ;
        RECT 373.535 675.165 373.815 675.445 ;
        RECT 374.245 675.165 374.525 675.445 ;
        RECT 374.955 675.165 375.235 675.445 ;
        RECT 375.665 675.165 375.945 675.445 ;
        RECT 376.375 675.165 376.655 675.445 ;
        RECT 369.275 674.455 369.555 674.735 ;
        RECT 369.985 674.455 370.265 674.735 ;
        RECT 370.695 674.455 370.975 674.735 ;
        RECT 371.405 674.455 371.685 674.735 ;
        RECT 372.115 674.455 372.395 674.735 ;
        RECT 372.825 674.455 373.105 674.735 ;
        RECT 373.535 674.455 373.815 674.735 ;
        RECT 374.245 674.455 374.525 674.735 ;
        RECT 374.955 674.455 375.235 674.735 ;
        RECT 375.665 674.455 375.945 674.735 ;
        RECT 376.375 674.455 376.655 674.735 ;
        RECT 369.275 673.745 369.555 674.025 ;
        RECT 369.985 673.745 370.265 674.025 ;
        RECT 370.695 673.745 370.975 674.025 ;
        RECT 371.405 673.745 371.685 674.025 ;
        RECT 372.115 673.745 372.395 674.025 ;
        RECT 372.825 673.745 373.105 674.025 ;
        RECT 373.535 673.745 373.815 674.025 ;
        RECT 374.245 673.745 374.525 674.025 ;
        RECT 374.955 673.745 375.235 674.025 ;
        RECT 375.665 673.745 375.945 674.025 ;
        RECT 376.375 673.745 376.655 674.025 ;
        RECT 369.275 673.035 369.555 673.315 ;
        RECT 369.985 673.035 370.265 673.315 ;
        RECT 370.695 673.035 370.975 673.315 ;
        RECT 371.405 673.035 371.685 673.315 ;
        RECT 372.115 673.035 372.395 673.315 ;
        RECT 372.825 673.035 373.105 673.315 ;
        RECT 373.535 673.035 373.815 673.315 ;
        RECT 374.245 673.035 374.525 673.315 ;
        RECT 374.955 673.035 375.235 673.315 ;
        RECT 375.665 673.035 375.945 673.315 ;
        RECT 376.375 673.035 376.655 673.315 ;
        RECT 369.275 672.325 369.555 672.605 ;
        RECT 369.985 672.325 370.265 672.605 ;
        RECT 370.695 672.325 370.975 672.605 ;
        RECT 371.405 672.325 371.685 672.605 ;
        RECT 372.115 672.325 372.395 672.605 ;
        RECT 372.825 672.325 373.105 672.605 ;
        RECT 373.535 672.325 373.815 672.605 ;
        RECT 374.245 672.325 374.525 672.605 ;
        RECT 374.955 672.325 375.235 672.605 ;
        RECT 375.665 672.325 375.945 672.605 ;
        RECT 376.375 672.325 376.655 672.605 ;
        RECT 369.275 671.615 369.555 671.895 ;
        RECT 369.985 671.615 370.265 671.895 ;
        RECT 370.695 671.615 370.975 671.895 ;
        RECT 371.405 671.615 371.685 671.895 ;
        RECT 372.115 671.615 372.395 671.895 ;
        RECT 372.825 671.615 373.105 671.895 ;
        RECT 373.535 671.615 373.815 671.895 ;
        RECT 374.245 671.615 374.525 671.895 ;
        RECT 374.955 671.615 375.235 671.895 ;
        RECT 375.665 671.615 375.945 671.895 ;
        RECT 376.375 671.615 376.655 671.895 ;
        RECT 369.275 670.905 369.555 671.185 ;
        RECT 369.985 670.905 370.265 671.185 ;
        RECT 370.695 670.905 370.975 671.185 ;
        RECT 371.405 670.905 371.685 671.185 ;
        RECT 372.115 670.905 372.395 671.185 ;
        RECT 372.825 670.905 373.105 671.185 ;
        RECT 373.535 670.905 373.815 671.185 ;
        RECT 374.245 670.905 374.525 671.185 ;
        RECT 374.955 670.905 375.235 671.185 ;
        RECT 375.665 670.905 375.945 671.185 ;
        RECT 376.375 670.905 376.655 671.185 ;
        RECT 369.275 670.195 369.555 670.475 ;
        RECT 369.985 670.195 370.265 670.475 ;
        RECT 370.695 670.195 370.975 670.475 ;
        RECT 371.405 670.195 371.685 670.475 ;
        RECT 372.115 670.195 372.395 670.475 ;
        RECT 372.825 670.195 373.105 670.475 ;
        RECT 373.535 670.195 373.815 670.475 ;
        RECT 374.245 670.195 374.525 670.475 ;
        RECT 374.955 670.195 375.235 670.475 ;
        RECT 375.665 670.195 375.945 670.475 ;
        RECT 376.375 670.195 376.655 670.475 ;
        RECT 369.275 669.485 369.555 669.765 ;
        RECT 369.985 669.485 370.265 669.765 ;
        RECT 370.695 669.485 370.975 669.765 ;
        RECT 371.405 669.485 371.685 669.765 ;
        RECT 372.115 669.485 372.395 669.765 ;
        RECT 372.825 669.485 373.105 669.765 ;
        RECT 373.535 669.485 373.815 669.765 ;
        RECT 374.245 669.485 374.525 669.765 ;
        RECT 374.955 669.485 375.235 669.765 ;
        RECT 375.665 669.485 375.945 669.765 ;
        RECT 376.375 669.485 376.655 669.765 ;
        RECT 369.275 665.185 369.555 665.465 ;
        RECT 369.985 665.185 370.265 665.465 ;
        RECT 370.695 665.185 370.975 665.465 ;
        RECT 371.405 665.185 371.685 665.465 ;
        RECT 372.115 665.185 372.395 665.465 ;
        RECT 372.825 665.185 373.105 665.465 ;
        RECT 373.535 665.185 373.815 665.465 ;
        RECT 374.245 665.185 374.525 665.465 ;
        RECT 374.955 665.185 375.235 665.465 ;
        RECT 375.665 665.185 375.945 665.465 ;
        RECT 376.375 665.185 376.655 665.465 ;
        RECT 369.275 664.475 369.555 664.755 ;
        RECT 369.985 664.475 370.265 664.755 ;
        RECT 370.695 664.475 370.975 664.755 ;
        RECT 371.405 664.475 371.685 664.755 ;
        RECT 372.115 664.475 372.395 664.755 ;
        RECT 372.825 664.475 373.105 664.755 ;
        RECT 373.535 664.475 373.815 664.755 ;
        RECT 374.245 664.475 374.525 664.755 ;
        RECT 374.955 664.475 375.235 664.755 ;
        RECT 375.665 664.475 375.945 664.755 ;
        RECT 376.375 664.475 376.655 664.755 ;
        RECT 369.275 663.765 369.555 664.045 ;
        RECT 369.985 663.765 370.265 664.045 ;
        RECT 370.695 663.765 370.975 664.045 ;
        RECT 371.405 663.765 371.685 664.045 ;
        RECT 372.115 663.765 372.395 664.045 ;
        RECT 372.825 663.765 373.105 664.045 ;
        RECT 373.535 663.765 373.815 664.045 ;
        RECT 374.245 663.765 374.525 664.045 ;
        RECT 374.955 663.765 375.235 664.045 ;
        RECT 375.665 663.765 375.945 664.045 ;
        RECT 376.375 663.765 376.655 664.045 ;
        RECT 369.275 663.055 369.555 663.335 ;
        RECT 369.985 663.055 370.265 663.335 ;
        RECT 370.695 663.055 370.975 663.335 ;
        RECT 371.405 663.055 371.685 663.335 ;
        RECT 372.115 663.055 372.395 663.335 ;
        RECT 372.825 663.055 373.105 663.335 ;
        RECT 373.535 663.055 373.815 663.335 ;
        RECT 374.245 663.055 374.525 663.335 ;
        RECT 374.955 663.055 375.235 663.335 ;
        RECT 375.665 663.055 375.945 663.335 ;
        RECT 376.375 663.055 376.655 663.335 ;
        RECT 369.275 662.345 369.555 662.625 ;
        RECT 369.985 662.345 370.265 662.625 ;
        RECT 370.695 662.345 370.975 662.625 ;
        RECT 371.405 662.345 371.685 662.625 ;
        RECT 372.115 662.345 372.395 662.625 ;
        RECT 372.825 662.345 373.105 662.625 ;
        RECT 373.535 662.345 373.815 662.625 ;
        RECT 374.245 662.345 374.525 662.625 ;
        RECT 374.955 662.345 375.235 662.625 ;
        RECT 375.665 662.345 375.945 662.625 ;
        RECT 376.375 662.345 376.655 662.625 ;
        RECT 369.275 661.635 369.555 661.915 ;
        RECT 369.985 661.635 370.265 661.915 ;
        RECT 370.695 661.635 370.975 661.915 ;
        RECT 371.405 661.635 371.685 661.915 ;
        RECT 372.115 661.635 372.395 661.915 ;
        RECT 372.825 661.635 373.105 661.915 ;
        RECT 373.535 661.635 373.815 661.915 ;
        RECT 374.245 661.635 374.525 661.915 ;
        RECT 374.955 661.635 375.235 661.915 ;
        RECT 375.665 661.635 375.945 661.915 ;
        RECT 376.375 661.635 376.655 661.915 ;
        RECT 369.275 660.925 369.555 661.205 ;
        RECT 369.985 660.925 370.265 661.205 ;
        RECT 370.695 660.925 370.975 661.205 ;
        RECT 371.405 660.925 371.685 661.205 ;
        RECT 372.115 660.925 372.395 661.205 ;
        RECT 372.825 660.925 373.105 661.205 ;
        RECT 373.535 660.925 373.815 661.205 ;
        RECT 374.245 660.925 374.525 661.205 ;
        RECT 374.955 660.925 375.235 661.205 ;
        RECT 375.665 660.925 375.945 661.205 ;
        RECT 376.375 660.925 376.655 661.205 ;
        RECT 369.275 660.215 369.555 660.495 ;
        RECT 369.985 660.215 370.265 660.495 ;
        RECT 370.695 660.215 370.975 660.495 ;
        RECT 371.405 660.215 371.685 660.495 ;
        RECT 372.115 660.215 372.395 660.495 ;
        RECT 372.825 660.215 373.105 660.495 ;
        RECT 373.535 660.215 373.815 660.495 ;
        RECT 374.245 660.215 374.525 660.495 ;
        RECT 374.955 660.215 375.235 660.495 ;
        RECT 375.665 660.215 375.945 660.495 ;
        RECT 376.375 660.215 376.655 660.495 ;
        RECT 369.275 659.505 369.555 659.785 ;
        RECT 369.985 659.505 370.265 659.785 ;
        RECT 370.695 659.505 370.975 659.785 ;
        RECT 371.405 659.505 371.685 659.785 ;
        RECT 372.115 659.505 372.395 659.785 ;
        RECT 372.825 659.505 373.105 659.785 ;
        RECT 373.535 659.505 373.815 659.785 ;
        RECT 374.245 659.505 374.525 659.785 ;
        RECT 374.955 659.505 375.235 659.785 ;
        RECT 375.665 659.505 375.945 659.785 ;
        RECT 376.375 659.505 376.655 659.785 ;
        RECT 369.275 658.795 369.555 659.075 ;
        RECT 369.985 658.795 370.265 659.075 ;
        RECT 370.695 658.795 370.975 659.075 ;
        RECT 371.405 658.795 371.685 659.075 ;
        RECT 372.115 658.795 372.395 659.075 ;
        RECT 372.825 658.795 373.105 659.075 ;
        RECT 373.535 658.795 373.815 659.075 ;
        RECT 374.245 658.795 374.525 659.075 ;
        RECT 374.955 658.795 375.235 659.075 ;
        RECT 375.665 658.795 375.945 659.075 ;
        RECT 376.375 658.795 376.655 659.075 ;
        RECT 369.275 658.085 369.555 658.365 ;
        RECT 369.985 658.085 370.265 658.365 ;
        RECT 370.695 658.085 370.975 658.365 ;
        RECT 371.405 658.085 371.685 658.365 ;
        RECT 372.115 658.085 372.395 658.365 ;
        RECT 372.825 658.085 373.105 658.365 ;
        RECT 373.535 658.085 373.815 658.365 ;
        RECT 374.245 658.085 374.525 658.365 ;
        RECT 374.955 658.085 375.235 658.365 ;
        RECT 375.665 658.085 375.945 658.365 ;
        RECT 376.375 658.085 376.655 658.365 ;
        RECT 369.275 657.375 369.555 657.655 ;
        RECT 369.985 657.375 370.265 657.655 ;
        RECT 370.695 657.375 370.975 657.655 ;
        RECT 371.405 657.375 371.685 657.655 ;
        RECT 372.115 657.375 372.395 657.655 ;
        RECT 372.825 657.375 373.105 657.655 ;
        RECT 373.535 657.375 373.815 657.655 ;
        RECT 374.245 657.375 374.525 657.655 ;
        RECT 374.955 657.375 375.235 657.655 ;
        RECT 375.665 657.375 375.945 657.655 ;
        RECT 376.375 657.375 376.655 657.655 ;
        RECT 369.275 656.665 369.555 656.945 ;
        RECT 369.985 656.665 370.265 656.945 ;
        RECT 370.695 656.665 370.975 656.945 ;
        RECT 371.405 656.665 371.685 656.945 ;
        RECT 372.115 656.665 372.395 656.945 ;
        RECT 372.825 656.665 373.105 656.945 ;
        RECT 373.535 656.665 373.815 656.945 ;
        RECT 374.245 656.665 374.525 656.945 ;
        RECT 374.955 656.665 375.235 656.945 ;
        RECT 375.665 656.665 375.945 656.945 ;
        RECT 376.375 656.665 376.655 656.945 ;
        RECT 369.275 655.955 369.555 656.235 ;
        RECT 369.985 655.955 370.265 656.235 ;
        RECT 370.695 655.955 370.975 656.235 ;
        RECT 371.405 655.955 371.685 656.235 ;
        RECT 372.115 655.955 372.395 656.235 ;
        RECT 372.825 655.955 373.105 656.235 ;
        RECT 373.535 655.955 373.815 656.235 ;
        RECT 374.245 655.955 374.525 656.235 ;
        RECT 374.955 655.955 375.235 656.235 ;
        RECT 375.665 655.955 375.945 656.235 ;
        RECT 376.375 655.955 376.655 656.235 ;
        RECT 369.275 653.335 369.555 653.615 ;
        RECT 369.985 653.335 370.265 653.615 ;
        RECT 370.695 653.335 370.975 653.615 ;
        RECT 371.405 653.335 371.685 653.615 ;
        RECT 372.115 653.335 372.395 653.615 ;
        RECT 372.825 653.335 373.105 653.615 ;
        RECT 373.535 653.335 373.815 653.615 ;
        RECT 374.245 653.335 374.525 653.615 ;
        RECT 374.955 653.335 375.235 653.615 ;
        RECT 375.665 653.335 375.945 653.615 ;
        RECT 376.375 653.335 376.655 653.615 ;
        RECT 369.275 652.625 369.555 652.905 ;
        RECT 369.985 652.625 370.265 652.905 ;
        RECT 370.695 652.625 370.975 652.905 ;
        RECT 371.405 652.625 371.685 652.905 ;
        RECT 372.115 652.625 372.395 652.905 ;
        RECT 372.825 652.625 373.105 652.905 ;
        RECT 373.535 652.625 373.815 652.905 ;
        RECT 374.245 652.625 374.525 652.905 ;
        RECT 374.955 652.625 375.235 652.905 ;
        RECT 375.665 652.625 375.945 652.905 ;
        RECT 376.375 652.625 376.655 652.905 ;
        RECT 369.275 651.915 369.555 652.195 ;
        RECT 369.985 651.915 370.265 652.195 ;
        RECT 370.695 651.915 370.975 652.195 ;
        RECT 371.405 651.915 371.685 652.195 ;
        RECT 372.115 651.915 372.395 652.195 ;
        RECT 372.825 651.915 373.105 652.195 ;
        RECT 373.535 651.915 373.815 652.195 ;
        RECT 374.245 651.915 374.525 652.195 ;
        RECT 374.955 651.915 375.235 652.195 ;
        RECT 375.665 651.915 375.945 652.195 ;
        RECT 376.375 651.915 376.655 652.195 ;
        RECT 369.275 651.205 369.555 651.485 ;
        RECT 369.985 651.205 370.265 651.485 ;
        RECT 370.695 651.205 370.975 651.485 ;
        RECT 371.405 651.205 371.685 651.485 ;
        RECT 372.115 651.205 372.395 651.485 ;
        RECT 372.825 651.205 373.105 651.485 ;
        RECT 373.535 651.205 373.815 651.485 ;
        RECT 374.245 651.205 374.525 651.485 ;
        RECT 374.955 651.205 375.235 651.485 ;
        RECT 375.665 651.205 375.945 651.485 ;
        RECT 376.375 651.205 376.655 651.485 ;
        RECT 369.275 650.495 369.555 650.775 ;
        RECT 369.985 650.495 370.265 650.775 ;
        RECT 370.695 650.495 370.975 650.775 ;
        RECT 371.405 650.495 371.685 650.775 ;
        RECT 372.115 650.495 372.395 650.775 ;
        RECT 372.825 650.495 373.105 650.775 ;
        RECT 373.535 650.495 373.815 650.775 ;
        RECT 374.245 650.495 374.525 650.775 ;
        RECT 374.955 650.495 375.235 650.775 ;
        RECT 375.665 650.495 375.945 650.775 ;
        RECT 376.375 650.495 376.655 650.775 ;
        RECT 369.275 649.785 369.555 650.065 ;
        RECT 369.985 649.785 370.265 650.065 ;
        RECT 370.695 649.785 370.975 650.065 ;
        RECT 371.405 649.785 371.685 650.065 ;
        RECT 372.115 649.785 372.395 650.065 ;
        RECT 372.825 649.785 373.105 650.065 ;
        RECT 373.535 649.785 373.815 650.065 ;
        RECT 374.245 649.785 374.525 650.065 ;
        RECT 374.955 649.785 375.235 650.065 ;
        RECT 375.665 649.785 375.945 650.065 ;
        RECT 376.375 649.785 376.655 650.065 ;
        RECT 369.275 649.075 369.555 649.355 ;
        RECT 369.985 649.075 370.265 649.355 ;
        RECT 370.695 649.075 370.975 649.355 ;
        RECT 371.405 649.075 371.685 649.355 ;
        RECT 372.115 649.075 372.395 649.355 ;
        RECT 372.825 649.075 373.105 649.355 ;
        RECT 373.535 649.075 373.815 649.355 ;
        RECT 374.245 649.075 374.525 649.355 ;
        RECT 374.955 649.075 375.235 649.355 ;
        RECT 375.665 649.075 375.945 649.355 ;
        RECT 376.375 649.075 376.655 649.355 ;
        RECT 369.275 648.365 369.555 648.645 ;
        RECT 369.985 648.365 370.265 648.645 ;
        RECT 370.695 648.365 370.975 648.645 ;
        RECT 371.405 648.365 371.685 648.645 ;
        RECT 372.115 648.365 372.395 648.645 ;
        RECT 372.825 648.365 373.105 648.645 ;
        RECT 373.535 648.365 373.815 648.645 ;
        RECT 374.245 648.365 374.525 648.645 ;
        RECT 374.955 648.365 375.235 648.645 ;
        RECT 375.665 648.365 375.945 648.645 ;
        RECT 376.375 648.365 376.655 648.645 ;
        RECT 369.275 647.655 369.555 647.935 ;
        RECT 369.985 647.655 370.265 647.935 ;
        RECT 370.695 647.655 370.975 647.935 ;
        RECT 371.405 647.655 371.685 647.935 ;
        RECT 372.115 647.655 372.395 647.935 ;
        RECT 372.825 647.655 373.105 647.935 ;
        RECT 373.535 647.655 373.815 647.935 ;
        RECT 374.245 647.655 374.525 647.935 ;
        RECT 374.955 647.655 375.235 647.935 ;
        RECT 375.665 647.655 375.945 647.935 ;
        RECT 376.375 647.655 376.655 647.935 ;
        RECT 369.275 646.945 369.555 647.225 ;
        RECT 369.985 646.945 370.265 647.225 ;
        RECT 370.695 646.945 370.975 647.225 ;
        RECT 371.405 646.945 371.685 647.225 ;
        RECT 372.115 646.945 372.395 647.225 ;
        RECT 372.825 646.945 373.105 647.225 ;
        RECT 373.535 646.945 373.815 647.225 ;
        RECT 374.245 646.945 374.525 647.225 ;
        RECT 374.955 646.945 375.235 647.225 ;
        RECT 375.665 646.945 375.945 647.225 ;
        RECT 376.375 646.945 376.655 647.225 ;
        RECT 369.275 646.235 369.555 646.515 ;
        RECT 369.985 646.235 370.265 646.515 ;
        RECT 370.695 646.235 370.975 646.515 ;
        RECT 371.405 646.235 371.685 646.515 ;
        RECT 372.115 646.235 372.395 646.515 ;
        RECT 372.825 646.235 373.105 646.515 ;
        RECT 373.535 646.235 373.815 646.515 ;
        RECT 374.245 646.235 374.525 646.515 ;
        RECT 374.955 646.235 375.235 646.515 ;
        RECT 375.665 646.235 375.945 646.515 ;
        RECT 376.375 646.235 376.655 646.515 ;
        RECT 369.275 645.525 369.555 645.805 ;
        RECT 369.985 645.525 370.265 645.805 ;
        RECT 370.695 645.525 370.975 645.805 ;
        RECT 371.405 645.525 371.685 645.805 ;
        RECT 372.115 645.525 372.395 645.805 ;
        RECT 372.825 645.525 373.105 645.805 ;
        RECT 373.535 645.525 373.815 645.805 ;
        RECT 374.245 645.525 374.525 645.805 ;
        RECT 374.955 645.525 375.235 645.805 ;
        RECT 375.665 645.525 375.945 645.805 ;
        RECT 376.375 645.525 376.655 645.805 ;
        RECT 369.275 644.815 369.555 645.095 ;
        RECT 369.985 644.815 370.265 645.095 ;
        RECT 370.695 644.815 370.975 645.095 ;
        RECT 371.405 644.815 371.685 645.095 ;
        RECT 372.115 644.815 372.395 645.095 ;
        RECT 372.825 644.815 373.105 645.095 ;
        RECT 373.535 644.815 373.815 645.095 ;
        RECT 374.245 644.815 374.525 645.095 ;
        RECT 374.955 644.815 375.235 645.095 ;
        RECT 375.665 644.815 375.945 645.095 ;
        RECT 376.375 644.815 376.655 645.095 ;
        RECT 369.275 644.105 369.555 644.385 ;
        RECT 369.985 644.105 370.265 644.385 ;
        RECT 370.695 644.105 370.975 644.385 ;
        RECT 371.405 644.105 371.685 644.385 ;
        RECT 372.115 644.105 372.395 644.385 ;
        RECT 372.825 644.105 373.105 644.385 ;
        RECT 373.535 644.105 373.815 644.385 ;
        RECT 374.245 644.105 374.525 644.385 ;
        RECT 374.955 644.105 375.235 644.385 ;
        RECT 375.665 644.105 375.945 644.385 ;
        RECT 376.375 644.105 376.655 644.385 ;
        RECT 369.330 640.190 369.610 640.470 ;
        RECT 370.040 640.190 370.320 640.470 ;
        RECT 370.750 640.190 371.030 640.470 ;
        RECT 371.460 640.190 371.740 640.470 ;
        RECT 372.170 640.190 372.450 640.470 ;
        RECT 372.880 640.190 373.160 640.470 ;
        RECT 373.590 640.190 373.870 640.470 ;
        RECT 374.300 640.190 374.580 640.470 ;
        RECT 375.010 640.190 375.290 640.470 ;
        RECT 375.720 640.190 376.000 640.470 ;
        RECT 376.430 640.190 376.710 640.470 ;
        RECT 369.330 639.480 369.610 639.760 ;
        RECT 370.040 639.480 370.320 639.760 ;
        RECT 370.750 639.480 371.030 639.760 ;
        RECT 371.460 639.480 371.740 639.760 ;
        RECT 372.170 639.480 372.450 639.760 ;
        RECT 372.880 639.480 373.160 639.760 ;
        RECT 373.590 639.480 373.870 639.760 ;
        RECT 374.300 639.480 374.580 639.760 ;
        RECT 375.010 639.480 375.290 639.760 ;
        RECT 375.720 639.480 376.000 639.760 ;
        RECT 376.430 639.480 376.710 639.760 ;
        RECT 369.330 638.770 369.610 639.050 ;
        RECT 370.040 638.770 370.320 639.050 ;
        RECT 370.750 638.770 371.030 639.050 ;
        RECT 371.460 638.770 371.740 639.050 ;
        RECT 372.170 638.770 372.450 639.050 ;
        RECT 372.880 638.770 373.160 639.050 ;
        RECT 373.590 638.770 373.870 639.050 ;
        RECT 374.300 638.770 374.580 639.050 ;
        RECT 375.010 638.770 375.290 639.050 ;
        RECT 375.720 638.770 376.000 639.050 ;
        RECT 376.430 638.770 376.710 639.050 ;
        RECT 369.330 638.060 369.610 638.340 ;
        RECT 370.040 638.060 370.320 638.340 ;
        RECT 370.750 638.060 371.030 638.340 ;
        RECT 371.460 638.060 371.740 638.340 ;
        RECT 372.170 638.060 372.450 638.340 ;
        RECT 372.880 638.060 373.160 638.340 ;
        RECT 373.590 638.060 373.870 638.340 ;
        RECT 374.300 638.060 374.580 638.340 ;
        RECT 375.010 638.060 375.290 638.340 ;
        RECT 375.720 638.060 376.000 638.340 ;
        RECT 376.430 638.060 376.710 638.340 ;
        RECT 369.330 637.350 369.610 637.630 ;
        RECT 370.040 637.350 370.320 637.630 ;
        RECT 370.750 637.350 371.030 637.630 ;
        RECT 371.460 637.350 371.740 637.630 ;
        RECT 372.170 637.350 372.450 637.630 ;
        RECT 372.880 637.350 373.160 637.630 ;
        RECT 373.590 637.350 373.870 637.630 ;
        RECT 374.300 637.350 374.580 637.630 ;
        RECT 375.010 637.350 375.290 637.630 ;
        RECT 375.720 637.350 376.000 637.630 ;
        RECT 376.430 637.350 376.710 637.630 ;
        RECT 369.330 636.640 369.610 636.920 ;
        RECT 370.040 636.640 370.320 636.920 ;
        RECT 370.750 636.640 371.030 636.920 ;
        RECT 371.460 636.640 371.740 636.920 ;
        RECT 372.170 636.640 372.450 636.920 ;
        RECT 372.880 636.640 373.160 636.920 ;
        RECT 373.590 636.640 373.870 636.920 ;
        RECT 374.300 636.640 374.580 636.920 ;
        RECT 375.010 636.640 375.290 636.920 ;
        RECT 375.720 636.640 376.000 636.920 ;
        RECT 376.430 636.640 376.710 636.920 ;
        RECT 369.330 635.930 369.610 636.210 ;
        RECT 370.040 635.930 370.320 636.210 ;
        RECT 370.750 635.930 371.030 636.210 ;
        RECT 371.460 635.930 371.740 636.210 ;
        RECT 372.170 635.930 372.450 636.210 ;
        RECT 372.880 635.930 373.160 636.210 ;
        RECT 373.590 635.930 373.870 636.210 ;
        RECT 374.300 635.930 374.580 636.210 ;
        RECT 375.010 635.930 375.290 636.210 ;
        RECT 375.720 635.930 376.000 636.210 ;
        RECT 376.430 635.930 376.710 636.210 ;
        RECT 369.330 635.220 369.610 635.500 ;
        RECT 370.040 635.220 370.320 635.500 ;
        RECT 370.750 635.220 371.030 635.500 ;
        RECT 371.460 635.220 371.740 635.500 ;
        RECT 372.170 635.220 372.450 635.500 ;
        RECT 372.880 635.220 373.160 635.500 ;
        RECT 373.590 635.220 373.870 635.500 ;
        RECT 374.300 635.220 374.580 635.500 ;
        RECT 375.010 635.220 375.290 635.500 ;
        RECT 375.720 635.220 376.000 635.500 ;
        RECT 376.430 635.220 376.710 635.500 ;
        RECT 369.330 634.510 369.610 634.790 ;
        RECT 370.040 634.510 370.320 634.790 ;
        RECT 370.750 634.510 371.030 634.790 ;
        RECT 371.460 634.510 371.740 634.790 ;
        RECT 372.170 634.510 372.450 634.790 ;
        RECT 372.880 634.510 373.160 634.790 ;
        RECT 373.590 634.510 373.870 634.790 ;
        RECT 374.300 634.510 374.580 634.790 ;
        RECT 375.010 634.510 375.290 634.790 ;
        RECT 375.720 634.510 376.000 634.790 ;
        RECT 376.430 634.510 376.710 634.790 ;
        RECT 369.330 633.800 369.610 634.080 ;
        RECT 370.040 633.800 370.320 634.080 ;
        RECT 370.750 633.800 371.030 634.080 ;
        RECT 371.460 633.800 371.740 634.080 ;
        RECT 372.170 633.800 372.450 634.080 ;
        RECT 372.880 633.800 373.160 634.080 ;
        RECT 373.590 633.800 373.870 634.080 ;
        RECT 374.300 633.800 374.580 634.080 ;
        RECT 375.010 633.800 375.290 634.080 ;
        RECT 375.720 633.800 376.000 634.080 ;
        RECT 376.430 633.800 376.710 634.080 ;
        RECT 369.330 633.090 369.610 633.370 ;
        RECT 370.040 633.090 370.320 633.370 ;
        RECT 370.750 633.090 371.030 633.370 ;
        RECT 371.460 633.090 371.740 633.370 ;
        RECT 372.170 633.090 372.450 633.370 ;
        RECT 372.880 633.090 373.160 633.370 ;
        RECT 373.590 633.090 373.870 633.370 ;
        RECT 374.300 633.090 374.580 633.370 ;
        RECT 375.010 633.090 375.290 633.370 ;
        RECT 375.720 633.090 376.000 633.370 ;
        RECT 376.430 633.090 376.710 633.370 ;
        RECT 369.330 632.380 369.610 632.660 ;
        RECT 370.040 632.380 370.320 632.660 ;
        RECT 370.750 632.380 371.030 632.660 ;
        RECT 371.460 632.380 371.740 632.660 ;
        RECT 372.170 632.380 372.450 632.660 ;
        RECT 372.880 632.380 373.160 632.660 ;
        RECT 373.590 632.380 373.870 632.660 ;
        RECT 374.300 632.380 374.580 632.660 ;
        RECT 375.010 632.380 375.290 632.660 ;
        RECT 375.720 632.380 376.000 632.660 ;
        RECT 376.430 632.380 376.710 632.660 ;
        RECT 369.330 631.670 369.610 631.950 ;
        RECT 370.040 631.670 370.320 631.950 ;
        RECT 370.750 631.670 371.030 631.950 ;
        RECT 371.460 631.670 371.740 631.950 ;
        RECT 372.170 631.670 372.450 631.950 ;
        RECT 372.880 631.670 373.160 631.950 ;
        RECT 373.590 631.670 373.870 631.950 ;
        RECT 374.300 631.670 374.580 631.950 ;
        RECT 375.010 631.670 375.290 631.950 ;
        RECT 375.720 631.670 376.000 631.950 ;
        RECT 376.430 631.670 376.710 631.950 ;
        RECT 369.330 497.970 369.610 498.250 ;
        RECT 370.040 497.970 370.320 498.250 ;
        RECT 370.750 497.970 371.030 498.250 ;
        RECT 371.460 497.970 371.740 498.250 ;
        RECT 372.170 497.970 372.450 498.250 ;
        RECT 372.880 497.970 373.160 498.250 ;
        RECT 373.590 497.970 373.870 498.250 ;
        RECT 374.300 497.970 374.580 498.250 ;
        RECT 375.010 497.970 375.290 498.250 ;
        RECT 375.720 497.970 376.000 498.250 ;
        RECT 376.430 497.970 376.710 498.250 ;
        RECT 369.330 497.260 369.610 497.540 ;
        RECT 370.040 497.260 370.320 497.540 ;
        RECT 370.750 497.260 371.030 497.540 ;
        RECT 371.460 497.260 371.740 497.540 ;
        RECT 372.170 497.260 372.450 497.540 ;
        RECT 372.880 497.260 373.160 497.540 ;
        RECT 373.590 497.260 373.870 497.540 ;
        RECT 374.300 497.260 374.580 497.540 ;
        RECT 375.010 497.260 375.290 497.540 ;
        RECT 375.720 497.260 376.000 497.540 ;
        RECT 376.430 497.260 376.710 497.540 ;
        RECT 369.330 496.550 369.610 496.830 ;
        RECT 370.040 496.550 370.320 496.830 ;
        RECT 370.750 496.550 371.030 496.830 ;
        RECT 371.460 496.550 371.740 496.830 ;
        RECT 372.170 496.550 372.450 496.830 ;
        RECT 372.880 496.550 373.160 496.830 ;
        RECT 373.590 496.550 373.870 496.830 ;
        RECT 374.300 496.550 374.580 496.830 ;
        RECT 375.010 496.550 375.290 496.830 ;
        RECT 375.720 496.550 376.000 496.830 ;
        RECT 376.430 496.550 376.710 496.830 ;
        RECT 369.330 495.840 369.610 496.120 ;
        RECT 370.040 495.840 370.320 496.120 ;
        RECT 370.750 495.840 371.030 496.120 ;
        RECT 371.460 495.840 371.740 496.120 ;
        RECT 372.170 495.840 372.450 496.120 ;
        RECT 372.880 495.840 373.160 496.120 ;
        RECT 373.590 495.840 373.870 496.120 ;
        RECT 374.300 495.840 374.580 496.120 ;
        RECT 375.010 495.840 375.290 496.120 ;
        RECT 375.720 495.840 376.000 496.120 ;
        RECT 376.430 495.840 376.710 496.120 ;
        RECT 369.330 495.130 369.610 495.410 ;
        RECT 370.040 495.130 370.320 495.410 ;
        RECT 370.750 495.130 371.030 495.410 ;
        RECT 371.460 495.130 371.740 495.410 ;
        RECT 372.170 495.130 372.450 495.410 ;
        RECT 372.880 495.130 373.160 495.410 ;
        RECT 373.590 495.130 373.870 495.410 ;
        RECT 374.300 495.130 374.580 495.410 ;
        RECT 375.010 495.130 375.290 495.410 ;
        RECT 375.720 495.130 376.000 495.410 ;
        RECT 376.430 495.130 376.710 495.410 ;
        RECT 369.330 494.420 369.610 494.700 ;
        RECT 370.040 494.420 370.320 494.700 ;
        RECT 370.750 494.420 371.030 494.700 ;
        RECT 371.460 494.420 371.740 494.700 ;
        RECT 372.170 494.420 372.450 494.700 ;
        RECT 372.880 494.420 373.160 494.700 ;
        RECT 373.590 494.420 373.870 494.700 ;
        RECT 374.300 494.420 374.580 494.700 ;
        RECT 375.010 494.420 375.290 494.700 ;
        RECT 375.720 494.420 376.000 494.700 ;
        RECT 376.430 494.420 376.710 494.700 ;
        RECT 369.330 493.710 369.610 493.990 ;
        RECT 370.040 493.710 370.320 493.990 ;
        RECT 370.750 493.710 371.030 493.990 ;
        RECT 371.460 493.710 371.740 493.990 ;
        RECT 372.170 493.710 372.450 493.990 ;
        RECT 372.880 493.710 373.160 493.990 ;
        RECT 373.590 493.710 373.870 493.990 ;
        RECT 374.300 493.710 374.580 493.990 ;
        RECT 375.010 493.710 375.290 493.990 ;
        RECT 375.720 493.710 376.000 493.990 ;
        RECT 376.430 493.710 376.710 493.990 ;
        RECT 369.330 493.000 369.610 493.280 ;
        RECT 370.040 493.000 370.320 493.280 ;
        RECT 370.750 493.000 371.030 493.280 ;
        RECT 371.460 493.000 371.740 493.280 ;
        RECT 372.170 493.000 372.450 493.280 ;
        RECT 372.880 493.000 373.160 493.280 ;
        RECT 373.590 493.000 373.870 493.280 ;
        RECT 374.300 493.000 374.580 493.280 ;
        RECT 375.010 493.000 375.290 493.280 ;
        RECT 375.720 493.000 376.000 493.280 ;
        RECT 376.430 493.000 376.710 493.280 ;
        RECT 369.330 492.290 369.610 492.570 ;
        RECT 370.040 492.290 370.320 492.570 ;
        RECT 370.750 492.290 371.030 492.570 ;
        RECT 371.460 492.290 371.740 492.570 ;
        RECT 372.170 492.290 372.450 492.570 ;
        RECT 372.880 492.290 373.160 492.570 ;
        RECT 373.590 492.290 373.870 492.570 ;
        RECT 374.300 492.290 374.580 492.570 ;
        RECT 375.010 492.290 375.290 492.570 ;
        RECT 375.720 492.290 376.000 492.570 ;
        RECT 376.430 492.290 376.710 492.570 ;
        RECT 369.330 491.580 369.610 491.860 ;
        RECT 370.040 491.580 370.320 491.860 ;
        RECT 370.750 491.580 371.030 491.860 ;
        RECT 371.460 491.580 371.740 491.860 ;
        RECT 372.170 491.580 372.450 491.860 ;
        RECT 372.880 491.580 373.160 491.860 ;
        RECT 373.590 491.580 373.870 491.860 ;
        RECT 374.300 491.580 374.580 491.860 ;
        RECT 375.010 491.580 375.290 491.860 ;
        RECT 375.720 491.580 376.000 491.860 ;
        RECT 376.430 491.580 376.710 491.860 ;
        RECT 369.330 490.870 369.610 491.150 ;
        RECT 370.040 490.870 370.320 491.150 ;
        RECT 370.750 490.870 371.030 491.150 ;
        RECT 371.460 490.870 371.740 491.150 ;
        RECT 372.170 490.870 372.450 491.150 ;
        RECT 372.880 490.870 373.160 491.150 ;
        RECT 373.590 490.870 373.870 491.150 ;
        RECT 374.300 490.870 374.580 491.150 ;
        RECT 375.010 490.870 375.290 491.150 ;
        RECT 375.720 490.870 376.000 491.150 ;
        RECT 376.430 490.870 376.710 491.150 ;
        RECT 369.330 490.160 369.610 490.440 ;
        RECT 370.040 490.160 370.320 490.440 ;
        RECT 370.750 490.160 371.030 490.440 ;
        RECT 371.460 490.160 371.740 490.440 ;
        RECT 372.170 490.160 372.450 490.440 ;
        RECT 372.880 490.160 373.160 490.440 ;
        RECT 373.590 490.160 373.870 490.440 ;
        RECT 374.300 490.160 374.580 490.440 ;
        RECT 375.010 490.160 375.290 490.440 ;
        RECT 375.720 490.160 376.000 490.440 ;
        RECT 376.430 490.160 376.710 490.440 ;
        RECT 369.330 489.450 369.610 489.730 ;
        RECT 370.040 489.450 370.320 489.730 ;
        RECT 370.750 489.450 371.030 489.730 ;
        RECT 371.460 489.450 371.740 489.730 ;
        RECT 372.170 489.450 372.450 489.730 ;
        RECT 372.880 489.450 373.160 489.730 ;
        RECT 373.590 489.450 373.870 489.730 ;
        RECT 374.300 489.450 374.580 489.730 ;
        RECT 375.010 489.450 375.290 489.730 ;
        RECT 375.720 489.450 376.000 489.730 ;
        RECT 376.430 489.450 376.710 489.730 ;
        RECT 369.275 485.565 369.555 485.845 ;
        RECT 369.985 485.565 370.265 485.845 ;
        RECT 370.695 485.565 370.975 485.845 ;
        RECT 371.405 485.565 371.685 485.845 ;
        RECT 372.115 485.565 372.395 485.845 ;
        RECT 372.825 485.565 373.105 485.845 ;
        RECT 373.535 485.565 373.815 485.845 ;
        RECT 374.245 485.565 374.525 485.845 ;
        RECT 374.955 485.565 375.235 485.845 ;
        RECT 375.665 485.565 375.945 485.845 ;
        RECT 376.375 485.565 376.655 485.845 ;
        RECT 369.275 484.855 369.555 485.135 ;
        RECT 369.985 484.855 370.265 485.135 ;
        RECT 370.695 484.855 370.975 485.135 ;
        RECT 371.405 484.855 371.685 485.135 ;
        RECT 372.115 484.855 372.395 485.135 ;
        RECT 372.825 484.855 373.105 485.135 ;
        RECT 373.535 484.855 373.815 485.135 ;
        RECT 374.245 484.855 374.525 485.135 ;
        RECT 374.955 484.855 375.235 485.135 ;
        RECT 375.665 484.855 375.945 485.135 ;
        RECT 376.375 484.855 376.655 485.135 ;
        RECT 369.275 484.145 369.555 484.425 ;
        RECT 369.985 484.145 370.265 484.425 ;
        RECT 370.695 484.145 370.975 484.425 ;
        RECT 371.405 484.145 371.685 484.425 ;
        RECT 372.115 484.145 372.395 484.425 ;
        RECT 372.825 484.145 373.105 484.425 ;
        RECT 373.535 484.145 373.815 484.425 ;
        RECT 374.245 484.145 374.525 484.425 ;
        RECT 374.955 484.145 375.235 484.425 ;
        RECT 375.665 484.145 375.945 484.425 ;
        RECT 376.375 484.145 376.655 484.425 ;
        RECT 369.275 483.435 369.555 483.715 ;
        RECT 369.985 483.435 370.265 483.715 ;
        RECT 370.695 483.435 370.975 483.715 ;
        RECT 371.405 483.435 371.685 483.715 ;
        RECT 372.115 483.435 372.395 483.715 ;
        RECT 372.825 483.435 373.105 483.715 ;
        RECT 373.535 483.435 373.815 483.715 ;
        RECT 374.245 483.435 374.525 483.715 ;
        RECT 374.955 483.435 375.235 483.715 ;
        RECT 375.665 483.435 375.945 483.715 ;
        RECT 376.375 483.435 376.655 483.715 ;
        RECT 369.275 482.725 369.555 483.005 ;
        RECT 369.985 482.725 370.265 483.005 ;
        RECT 370.695 482.725 370.975 483.005 ;
        RECT 371.405 482.725 371.685 483.005 ;
        RECT 372.115 482.725 372.395 483.005 ;
        RECT 372.825 482.725 373.105 483.005 ;
        RECT 373.535 482.725 373.815 483.005 ;
        RECT 374.245 482.725 374.525 483.005 ;
        RECT 374.955 482.725 375.235 483.005 ;
        RECT 375.665 482.725 375.945 483.005 ;
        RECT 376.375 482.725 376.655 483.005 ;
        RECT 369.275 482.015 369.555 482.295 ;
        RECT 369.985 482.015 370.265 482.295 ;
        RECT 370.695 482.015 370.975 482.295 ;
        RECT 371.405 482.015 371.685 482.295 ;
        RECT 372.115 482.015 372.395 482.295 ;
        RECT 372.825 482.015 373.105 482.295 ;
        RECT 373.535 482.015 373.815 482.295 ;
        RECT 374.245 482.015 374.525 482.295 ;
        RECT 374.955 482.015 375.235 482.295 ;
        RECT 375.665 482.015 375.945 482.295 ;
        RECT 376.375 482.015 376.655 482.295 ;
        RECT 369.275 481.305 369.555 481.585 ;
        RECT 369.985 481.305 370.265 481.585 ;
        RECT 370.695 481.305 370.975 481.585 ;
        RECT 371.405 481.305 371.685 481.585 ;
        RECT 372.115 481.305 372.395 481.585 ;
        RECT 372.825 481.305 373.105 481.585 ;
        RECT 373.535 481.305 373.815 481.585 ;
        RECT 374.245 481.305 374.525 481.585 ;
        RECT 374.955 481.305 375.235 481.585 ;
        RECT 375.665 481.305 375.945 481.585 ;
        RECT 376.375 481.305 376.655 481.585 ;
        RECT 369.275 480.595 369.555 480.875 ;
        RECT 369.985 480.595 370.265 480.875 ;
        RECT 370.695 480.595 370.975 480.875 ;
        RECT 371.405 480.595 371.685 480.875 ;
        RECT 372.115 480.595 372.395 480.875 ;
        RECT 372.825 480.595 373.105 480.875 ;
        RECT 373.535 480.595 373.815 480.875 ;
        RECT 374.245 480.595 374.525 480.875 ;
        RECT 374.955 480.595 375.235 480.875 ;
        RECT 375.665 480.595 375.945 480.875 ;
        RECT 376.375 480.595 376.655 480.875 ;
        RECT 369.275 479.885 369.555 480.165 ;
        RECT 369.985 479.885 370.265 480.165 ;
        RECT 370.695 479.885 370.975 480.165 ;
        RECT 371.405 479.885 371.685 480.165 ;
        RECT 372.115 479.885 372.395 480.165 ;
        RECT 372.825 479.885 373.105 480.165 ;
        RECT 373.535 479.885 373.815 480.165 ;
        RECT 374.245 479.885 374.525 480.165 ;
        RECT 374.955 479.885 375.235 480.165 ;
        RECT 375.665 479.885 375.945 480.165 ;
        RECT 376.375 479.885 376.655 480.165 ;
        RECT 369.275 479.175 369.555 479.455 ;
        RECT 369.985 479.175 370.265 479.455 ;
        RECT 370.695 479.175 370.975 479.455 ;
        RECT 371.405 479.175 371.685 479.455 ;
        RECT 372.115 479.175 372.395 479.455 ;
        RECT 372.825 479.175 373.105 479.455 ;
        RECT 373.535 479.175 373.815 479.455 ;
        RECT 374.245 479.175 374.525 479.455 ;
        RECT 374.955 479.175 375.235 479.455 ;
        RECT 375.665 479.175 375.945 479.455 ;
        RECT 376.375 479.175 376.655 479.455 ;
        RECT 369.275 478.465 369.555 478.745 ;
        RECT 369.985 478.465 370.265 478.745 ;
        RECT 370.695 478.465 370.975 478.745 ;
        RECT 371.405 478.465 371.685 478.745 ;
        RECT 372.115 478.465 372.395 478.745 ;
        RECT 372.825 478.465 373.105 478.745 ;
        RECT 373.535 478.465 373.815 478.745 ;
        RECT 374.245 478.465 374.525 478.745 ;
        RECT 374.955 478.465 375.235 478.745 ;
        RECT 375.665 478.465 375.945 478.745 ;
        RECT 376.375 478.465 376.655 478.745 ;
        RECT 369.275 477.755 369.555 478.035 ;
        RECT 369.985 477.755 370.265 478.035 ;
        RECT 370.695 477.755 370.975 478.035 ;
        RECT 371.405 477.755 371.685 478.035 ;
        RECT 372.115 477.755 372.395 478.035 ;
        RECT 372.825 477.755 373.105 478.035 ;
        RECT 373.535 477.755 373.815 478.035 ;
        RECT 374.245 477.755 374.525 478.035 ;
        RECT 374.955 477.755 375.235 478.035 ;
        RECT 375.665 477.755 375.945 478.035 ;
        RECT 376.375 477.755 376.655 478.035 ;
        RECT 369.275 477.045 369.555 477.325 ;
        RECT 369.985 477.045 370.265 477.325 ;
        RECT 370.695 477.045 370.975 477.325 ;
        RECT 371.405 477.045 371.685 477.325 ;
        RECT 372.115 477.045 372.395 477.325 ;
        RECT 372.825 477.045 373.105 477.325 ;
        RECT 373.535 477.045 373.815 477.325 ;
        RECT 374.245 477.045 374.525 477.325 ;
        RECT 374.955 477.045 375.235 477.325 ;
        RECT 375.665 477.045 375.945 477.325 ;
        RECT 376.375 477.045 376.655 477.325 ;
        RECT 369.275 476.335 369.555 476.615 ;
        RECT 369.985 476.335 370.265 476.615 ;
        RECT 370.695 476.335 370.975 476.615 ;
        RECT 371.405 476.335 371.685 476.615 ;
        RECT 372.115 476.335 372.395 476.615 ;
        RECT 372.825 476.335 373.105 476.615 ;
        RECT 373.535 476.335 373.815 476.615 ;
        RECT 374.245 476.335 374.525 476.615 ;
        RECT 374.955 476.335 375.235 476.615 ;
        RECT 375.665 476.335 375.945 476.615 ;
        RECT 376.375 476.335 376.655 476.615 ;
        RECT 369.275 473.715 369.555 473.995 ;
        RECT 369.985 473.715 370.265 473.995 ;
        RECT 370.695 473.715 370.975 473.995 ;
        RECT 371.405 473.715 371.685 473.995 ;
        RECT 372.115 473.715 372.395 473.995 ;
        RECT 372.825 473.715 373.105 473.995 ;
        RECT 373.535 473.715 373.815 473.995 ;
        RECT 374.245 473.715 374.525 473.995 ;
        RECT 374.955 473.715 375.235 473.995 ;
        RECT 375.665 473.715 375.945 473.995 ;
        RECT 376.375 473.715 376.655 473.995 ;
        RECT 369.275 473.005 369.555 473.285 ;
        RECT 369.985 473.005 370.265 473.285 ;
        RECT 370.695 473.005 370.975 473.285 ;
        RECT 371.405 473.005 371.685 473.285 ;
        RECT 372.115 473.005 372.395 473.285 ;
        RECT 372.825 473.005 373.105 473.285 ;
        RECT 373.535 473.005 373.815 473.285 ;
        RECT 374.245 473.005 374.525 473.285 ;
        RECT 374.955 473.005 375.235 473.285 ;
        RECT 375.665 473.005 375.945 473.285 ;
        RECT 376.375 473.005 376.655 473.285 ;
        RECT 369.275 472.295 369.555 472.575 ;
        RECT 369.985 472.295 370.265 472.575 ;
        RECT 370.695 472.295 370.975 472.575 ;
        RECT 371.405 472.295 371.685 472.575 ;
        RECT 372.115 472.295 372.395 472.575 ;
        RECT 372.825 472.295 373.105 472.575 ;
        RECT 373.535 472.295 373.815 472.575 ;
        RECT 374.245 472.295 374.525 472.575 ;
        RECT 374.955 472.295 375.235 472.575 ;
        RECT 375.665 472.295 375.945 472.575 ;
        RECT 376.375 472.295 376.655 472.575 ;
        RECT 369.275 471.585 369.555 471.865 ;
        RECT 369.985 471.585 370.265 471.865 ;
        RECT 370.695 471.585 370.975 471.865 ;
        RECT 371.405 471.585 371.685 471.865 ;
        RECT 372.115 471.585 372.395 471.865 ;
        RECT 372.825 471.585 373.105 471.865 ;
        RECT 373.535 471.585 373.815 471.865 ;
        RECT 374.245 471.585 374.525 471.865 ;
        RECT 374.955 471.585 375.235 471.865 ;
        RECT 375.665 471.585 375.945 471.865 ;
        RECT 376.375 471.585 376.655 471.865 ;
        RECT 369.275 470.875 369.555 471.155 ;
        RECT 369.985 470.875 370.265 471.155 ;
        RECT 370.695 470.875 370.975 471.155 ;
        RECT 371.405 470.875 371.685 471.155 ;
        RECT 372.115 470.875 372.395 471.155 ;
        RECT 372.825 470.875 373.105 471.155 ;
        RECT 373.535 470.875 373.815 471.155 ;
        RECT 374.245 470.875 374.525 471.155 ;
        RECT 374.955 470.875 375.235 471.155 ;
        RECT 375.665 470.875 375.945 471.155 ;
        RECT 376.375 470.875 376.655 471.155 ;
        RECT 369.275 470.165 369.555 470.445 ;
        RECT 369.985 470.165 370.265 470.445 ;
        RECT 370.695 470.165 370.975 470.445 ;
        RECT 371.405 470.165 371.685 470.445 ;
        RECT 372.115 470.165 372.395 470.445 ;
        RECT 372.825 470.165 373.105 470.445 ;
        RECT 373.535 470.165 373.815 470.445 ;
        RECT 374.245 470.165 374.525 470.445 ;
        RECT 374.955 470.165 375.235 470.445 ;
        RECT 375.665 470.165 375.945 470.445 ;
        RECT 376.375 470.165 376.655 470.445 ;
        RECT 369.275 469.455 369.555 469.735 ;
        RECT 369.985 469.455 370.265 469.735 ;
        RECT 370.695 469.455 370.975 469.735 ;
        RECT 371.405 469.455 371.685 469.735 ;
        RECT 372.115 469.455 372.395 469.735 ;
        RECT 372.825 469.455 373.105 469.735 ;
        RECT 373.535 469.455 373.815 469.735 ;
        RECT 374.245 469.455 374.525 469.735 ;
        RECT 374.955 469.455 375.235 469.735 ;
        RECT 375.665 469.455 375.945 469.735 ;
        RECT 376.375 469.455 376.655 469.735 ;
        RECT 369.275 468.745 369.555 469.025 ;
        RECT 369.985 468.745 370.265 469.025 ;
        RECT 370.695 468.745 370.975 469.025 ;
        RECT 371.405 468.745 371.685 469.025 ;
        RECT 372.115 468.745 372.395 469.025 ;
        RECT 372.825 468.745 373.105 469.025 ;
        RECT 373.535 468.745 373.815 469.025 ;
        RECT 374.245 468.745 374.525 469.025 ;
        RECT 374.955 468.745 375.235 469.025 ;
        RECT 375.665 468.745 375.945 469.025 ;
        RECT 376.375 468.745 376.655 469.025 ;
        RECT 369.275 468.035 369.555 468.315 ;
        RECT 369.985 468.035 370.265 468.315 ;
        RECT 370.695 468.035 370.975 468.315 ;
        RECT 371.405 468.035 371.685 468.315 ;
        RECT 372.115 468.035 372.395 468.315 ;
        RECT 372.825 468.035 373.105 468.315 ;
        RECT 373.535 468.035 373.815 468.315 ;
        RECT 374.245 468.035 374.525 468.315 ;
        RECT 374.955 468.035 375.235 468.315 ;
        RECT 375.665 468.035 375.945 468.315 ;
        RECT 376.375 468.035 376.655 468.315 ;
        RECT 369.275 467.325 369.555 467.605 ;
        RECT 369.985 467.325 370.265 467.605 ;
        RECT 370.695 467.325 370.975 467.605 ;
        RECT 371.405 467.325 371.685 467.605 ;
        RECT 372.115 467.325 372.395 467.605 ;
        RECT 372.825 467.325 373.105 467.605 ;
        RECT 373.535 467.325 373.815 467.605 ;
        RECT 374.245 467.325 374.525 467.605 ;
        RECT 374.955 467.325 375.235 467.605 ;
        RECT 375.665 467.325 375.945 467.605 ;
        RECT 376.375 467.325 376.655 467.605 ;
        RECT 369.275 466.615 369.555 466.895 ;
        RECT 369.985 466.615 370.265 466.895 ;
        RECT 370.695 466.615 370.975 466.895 ;
        RECT 371.405 466.615 371.685 466.895 ;
        RECT 372.115 466.615 372.395 466.895 ;
        RECT 372.825 466.615 373.105 466.895 ;
        RECT 373.535 466.615 373.815 466.895 ;
        RECT 374.245 466.615 374.525 466.895 ;
        RECT 374.955 466.615 375.235 466.895 ;
        RECT 375.665 466.615 375.945 466.895 ;
        RECT 376.375 466.615 376.655 466.895 ;
        RECT 369.275 465.905 369.555 466.185 ;
        RECT 369.985 465.905 370.265 466.185 ;
        RECT 370.695 465.905 370.975 466.185 ;
        RECT 371.405 465.905 371.685 466.185 ;
        RECT 372.115 465.905 372.395 466.185 ;
        RECT 372.825 465.905 373.105 466.185 ;
        RECT 373.535 465.905 373.815 466.185 ;
        RECT 374.245 465.905 374.525 466.185 ;
        RECT 374.955 465.905 375.235 466.185 ;
        RECT 375.665 465.905 375.945 466.185 ;
        RECT 376.375 465.905 376.655 466.185 ;
        RECT 369.275 465.195 369.555 465.475 ;
        RECT 369.985 465.195 370.265 465.475 ;
        RECT 370.695 465.195 370.975 465.475 ;
        RECT 371.405 465.195 371.685 465.475 ;
        RECT 372.115 465.195 372.395 465.475 ;
        RECT 372.825 465.195 373.105 465.475 ;
        RECT 373.535 465.195 373.815 465.475 ;
        RECT 374.245 465.195 374.525 465.475 ;
        RECT 374.955 465.195 375.235 465.475 ;
        RECT 375.665 465.195 375.945 465.475 ;
        RECT 376.375 465.195 376.655 465.475 ;
        RECT 369.275 464.485 369.555 464.765 ;
        RECT 369.985 464.485 370.265 464.765 ;
        RECT 370.695 464.485 370.975 464.765 ;
        RECT 371.405 464.485 371.685 464.765 ;
        RECT 372.115 464.485 372.395 464.765 ;
        RECT 372.825 464.485 373.105 464.765 ;
        RECT 373.535 464.485 373.815 464.765 ;
        RECT 374.245 464.485 374.525 464.765 ;
        RECT 374.955 464.485 375.235 464.765 ;
        RECT 375.665 464.485 375.945 464.765 ;
        RECT 376.375 464.485 376.655 464.765 ;
        RECT 369.275 460.185 369.555 460.465 ;
        RECT 369.985 460.185 370.265 460.465 ;
        RECT 370.695 460.185 370.975 460.465 ;
        RECT 371.405 460.185 371.685 460.465 ;
        RECT 372.115 460.185 372.395 460.465 ;
        RECT 372.825 460.185 373.105 460.465 ;
        RECT 373.535 460.185 373.815 460.465 ;
        RECT 374.245 460.185 374.525 460.465 ;
        RECT 374.955 460.185 375.235 460.465 ;
        RECT 375.665 460.185 375.945 460.465 ;
        RECT 376.375 460.185 376.655 460.465 ;
        RECT 369.275 459.475 369.555 459.755 ;
        RECT 369.985 459.475 370.265 459.755 ;
        RECT 370.695 459.475 370.975 459.755 ;
        RECT 371.405 459.475 371.685 459.755 ;
        RECT 372.115 459.475 372.395 459.755 ;
        RECT 372.825 459.475 373.105 459.755 ;
        RECT 373.535 459.475 373.815 459.755 ;
        RECT 374.245 459.475 374.525 459.755 ;
        RECT 374.955 459.475 375.235 459.755 ;
        RECT 375.665 459.475 375.945 459.755 ;
        RECT 376.375 459.475 376.655 459.755 ;
        RECT 369.275 458.765 369.555 459.045 ;
        RECT 369.985 458.765 370.265 459.045 ;
        RECT 370.695 458.765 370.975 459.045 ;
        RECT 371.405 458.765 371.685 459.045 ;
        RECT 372.115 458.765 372.395 459.045 ;
        RECT 372.825 458.765 373.105 459.045 ;
        RECT 373.535 458.765 373.815 459.045 ;
        RECT 374.245 458.765 374.525 459.045 ;
        RECT 374.955 458.765 375.235 459.045 ;
        RECT 375.665 458.765 375.945 459.045 ;
        RECT 376.375 458.765 376.655 459.045 ;
        RECT 369.275 458.055 369.555 458.335 ;
        RECT 369.985 458.055 370.265 458.335 ;
        RECT 370.695 458.055 370.975 458.335 ;
        RECT 371.405 458.055 371.685 458.335 ;
        RECT 372.115 458.055 372.395 458.335 ;
        RECT 372.825 458.055 373.105 458.335 ;
        RECT 373.535 458.055 373.815 458.335 ;
        RECT 374.245 458.055 374.525 458.335 ;
        RECT 374.955 458.055 375.235 458.335 ;
        RECT 375.665 458.055 375.945 458.335 ;
        RECT 376.375 458.055 376.655 458.335 ;
        RECT 369.275 457.345 369.555 457.625 ;
        RECT 369.985 457.345 370.265 457.625 ;
        RECT 370.695 457.345 370.975 457.625 ;
        RECT 371.405 457.345 371.685 457.625 ;
        RECT 372.115 457.345 372.395 457.625 ;
        RECT 372.825 457.345 373.105 457.625 ;
        RECT 373.535 457.345 373.815 457.625 ;
        RECT 374.245 457.345 374.525 457.625 ;
        RECT 374.955 457.345 375.235 457.625 ;
        RECT 375.665 457.345 375.945 457.625 ;
        RECT 376.375 457.345 376.655 457.625 ;
        RECT 369.275 456.635 369.555 456.915 ;
        RECT 369.985 456.635 370.265 456.915 ;
        RECT 370.695 456.635 370.975 456.915 ;
        RECT 371.405 456.635 371.685 456.915 ;
        RECT 372.115 456.635 372.395 456.915 ;
        RECT 372.825 456.635 373.105 456.915 ;
        RECT 373.535 456.635 373.815 456.915 ;
        RECT 374.245 456.635 374.525 456.915 ;
        RECT 374.955 456.635 375.235 456.915 ;
        RECT 375.665 456.635 375.945 456.915 ;
        RECT 376.375 456.635 376.655 456.915 ;
        RECT 369.275 455.925 369.555 456.205 ;
        RECT 369.985 455.925 370.265 456.205 ;
        RECT 370.695 455.925 370.975 456.205 ;
        RECT 371.405 455.925 371.685 456.205 ;
        RECT 372.115 455.925 372.395 456.205 ;
        RECT 372.825 455.925 373.105 456.205 ;
        RECT 373.535 455.925 373.815 456.205 ;
        RECT 374.245 455.925 374.525 456.205 ;
        RECT 374.955 455.925 375.235 456.205 ;
        RECT 375.665 455.925 375.945 456.205 ;
        RECT 376.375 455.925 376.655 456.205 ;
        RECT 369.275 455.215 369.555 455.495 ;
        RECT 369.985 455.215 370.265 455.495 ;
        RECT 370.695 455.215 370.975 455.495 ;
        RECT 371.405 455.215 371.685 455.495 ;
        RECT 372.115 455.215 372.395 455.495 ;
        RECT 372.825 455.215 373.105 455.495 ;
        RECT 373.535 455.215 373.815 455.495 ;
        RECT 374.245 455.215 374.525 455.495 ;
        RECT 374.955 455.215 375.235 455.495 ;
        RECT 375.665 455.215 375.945 455.495 ;
        RECT 376.375 455.215 376.655 455.495 ;
        RECT 369.275 454.505 369.555 454.785 ;
        RECT 369.985 454.505 370.265 454.785 ;
        RECT 370.695 454.505 370.975 454.785 ;
        RECT 371.405 454.505 371.685 454.785 ;
        RECT 372.115 454.505 372.395 454.785 ;
        RECT 372.825 454.505 373.105 454.785 ;
        RECT 373.535 454.505 373.815 454.785 ;
        RECT 374.245 454.505 374.525 454.785 ;
        RECT 374.955 454.505 375.235 454.785 ;
        RECT 375.665 454.505 375.945 454.785 ;
        RECT 376.375 454.505 376.655 454.785 ;
        RECT 369.275 453.795 369.555 454.075 ;
        RECT 369.985 453.795 370.265 454.075 ;
        RECT 370.695 453.795 370.975 454.075 ;
        RECT 371.405 453.795 371.685 454.075 ;
        RECT 372.115 453.795 372.395 454.075 ;
        RECT 372.825 453.795 373.105 454.075 ;
        RECT 373.535 453.795 373.815 454.075 ;
        RECT 374.245 453.795 374.525 454.075 ;
        RECT 374.955 453.795 375.235 454.075 ;
        RECT 375.665 453.795 375.945 454.075 ;
        RECT 376.375 453.795 376.655 454.075 ;
        RECT 369.275 453.085 369.555 453.365 ;
        RECT 369.985 453.085 370.265 453.365 ;
        RECT 370.695 453.085 370.975 453.365 ;
        RECT 371.405 453.085 371.685 453.365 ;
        RECT 372.115 453.085 372.395 453.365 ;
        RECT 372.825 453.085 373.105 453.365 ;
        RECT 373.535 453.085 373.815 453.365 ;
        RECT 374.245 453.085 374.525 453.365 ;
        RECT 374.955 453.085 375.235 453.365 ;
        RECT 375.665 453.085 375.945 453.365 ;
        RECT 376.375 453.085 376.655 453.365 ;
        RECT 369.275 452.375 369.555 452.655 ;
        RECT 369.985 452.375 370.265 452.655 ;
        RECT 370.695 452.375 370.975 452.655 ;
        RECT 371.405 452.375 371.685 452.655 ;
        RECT 372.115 452.375 372.395 452.655 ;
        RECT 372.825 452.375 373.105 452.655 ;
        RECT 373.535 452.375 373.815 452.655 ;
        RECT 374.245 452.375 374.525 452.655 ;
        RECT 374.955 452.375 375.235 452.655 ;
        RECT 375.665 452.375 375.945 452.655 ;
        RECT 376.375 452.375 376.655 452.655 ;
        RECT 369.275 451.665 369.555 451.945 ;
        RECT 369.985 451.665 370.265 451.945 ;
        RECT 370.695 451.665 370.975 451.945 ;
        RECT 371.405 451.665 371.685 451.945 ;
        RECT 372.115 451.665 372.395 451.945 ;
        RECT 372.825 451.665 373.105 451.945 ;
        RECT 373.535 451.665 373.815 451.945 ;
        RECT 374.245 451.665 374.525 451.945 ;
        RECT 374.955 451.665 375.235 451.945 ;
        RECT 375.665 451.665 375.945 451.945 ;
        RECT 376.375 451.665 376.655 451.945 ;
        RECT 369.275 450.955 369.555 451.235 ;
        RECT 369.985 450.955 370.265 451.235 ;
        RECT 370.695 450.955 370.975 451.235 ;
        RECT 371.405 450.955 371.685 451.235 ;
        RECT 372.115 450.955 372.395 451.235 ;
        RECT 372.825 450.955 373.105 451.235 ;
        RECT 373.535 450.955 373.815 451.235 ;
        RECT 374.245 450.955 374.525 451.235 ;
        RECT 374.955 450.955 375.235 451.235 ;
        RECT 375.665 450.955 375.945 451.235 ;
        RECT 376.375 450.955 376.655 451.235 ;
        RECT 369.275 448.335 369.555 448.615 ;
        RECT 369.985 448.335 370.265 448.615 ;
        RECT 370.695 448.335 370.975 448.615 ;
        RECT 371.405 448.335 371.685 448.615 ;
        RECT 372.115 448.335 372.395 448.615 ;
        RECT 372.825 448.335 373.105 448.615 ;
        RECT 373.535 448.335 373.815 448.615 ;
        RECT 374.245 448.335 374.525 448.615 ;
        RECT 374.955 448.335 375.235 448.615 ;
        RECT 375.665 448.335 375.945 448.615 ;
        RECT 376.375 448.335 376.655 448.615 ;
        RECT 369.275 447.625 369.555 447.905 ;
        RECT 369.985 447.625 370.265 447.905 ;
        RECT 370.695 447.625 370.975 447.905 ;
        RECT 371.405 447.625 371.685 447.905 ;
        RECT 372.115 447.625 372.395 447.905 ;
        RECT 372.825 447.625 373.105 447.905 ;
        RECT 373.535 447.625 373.815 447.905 ;
        RECT 374.245 447.625 374.525 447.905 ;
        RECT 374.955 447.625 375.235 447.905 ;
        RECT 375.665 447.625 375.945 447.905 ;
        RECT 376.375 447.625 376.655 447.905 ;
        RECT 369.275 446.915 369.555 447.195 ;
        RECT 369.985 446.915 370.265 447.195 ;
        RECT 370.695 446.915 370.975 447.195 ;
        RECT 371.405 446.915 371.685 447.195 ;
        RECT 372.115 446.915 372.395 447.195 ;
        RECT 372.825 446.915 373.105 447.195 ;
        RECT 373.535 446.915 373.815 447.195 ;
        RECT 374.245 446.915 374.525 447.195 ;
        RECT 374.955 446.915 375.235 447.195 ;
        RECT 375.665 446.915 375.945 447.195 ;
        RECT 376.375 446.915 376.655 447.195 ;
        RECT 369.275 446.205 369.555 446.485 ;
        RECT 369.985 446.205 370.265 446.485 ;
        RECT 370.695 446.205 370.975 446.485 ;
        RECT 371.405 446.205 371.685 446.485 ;
        RECT 372.115 446.205 372.395 446.485 ;
        RECT 372.825 446.205 373.105 446.485 ;
        RECT 373.535 446.205 373.815 446.485 ;
        RECT 374.245 446.205 374.525 446.485 ;
        RECT 374.955 446.205 375.235 446.485 ;
        RECT 375.665 446.205 375.945 446.485 ;
        RECT 376.375 446.205 376.655 446.485 ;
        RECT 369.275 445.495 369.555 445.775 ;
        RECT 369.985 445.495 370.265 445.775 ;
        RECT 370.695 445.495 370.975 445.775 ;
        RECT 371.405 445.495 371.685 445.775 ;
        RECT 372.115 445.495 372.395 445.775 ;
        RECT 372.825 445.495 373.105 445.775 ;
        RECT 373.535 445.495 373.815 445.775 ;
        RECT 374.245 445.495 374.525 445.775 ;
        RECT 374.955 445.495 375.235 445.775 ;
        RECT 375.665 445.495 375.945 445.775 ;
        RECT 376.375 445.495 376.655 445.775 ;
        RECT 369.275 444.785 369.555 445.065 ;
        RECT 369.985 444.785 370.265 445.065 ;
        RECT 370.695 444.785 370.975 445.065 ;
        RECT 371.405 444.785 371.685 445.065 ;
        RECT 372.115 444.785 372.395 445.065 ;
        RECT 372.825 444.785 373.105 445.065 ;
        RECT 373.535 444.785 373.815 445.065 ;
        RECT 374.245 444.785 374.525 445.065 ;
        RECT 374.955 444.785 375.235 445.065 ;
        RECT 375.665 444.785 375.945 445.065 ;
        RECT 376.375 444.785 376.655 445.065 ;
        RECT 369.275 444.075 369.555 444.355 ;
        RECT 369.985 444.075 370.265 444.355 ;
        RECT 370.695 444.075 370.975 444.355 ;
        RECT 371.405 444.075 371.685 444.355 ;
        RECT 372.115 444.075 372.395 444.355 ;
        RECT 372.825 444.075 373.105 444.355 ;
        RECT 373.535 444.075 373.815 444.355 ;
        RECT 374.245 444.075 374.525 444.355 ;
        RECT 374.955 444.075 375.235 444.355 ;
        RECT 375.665 444.075 375.945 444.355 ;
        RECT 376.375 444.075 376.655 444.355 ;
        RECT 369.275 443.365 369.555 443.645 ;
        RECT 369.985 443.365 370.265 443.645 ;
        RECT 370.695 443.365 370.975 443.645 ;
        RECT 371.405 443.365 371.685 443.645 ;
        RECT 372.115 443.365 372.395 443.645 ;
        RECT 372.825 443.365 373.105 443.645 ;
        RECT 373.535 443.365 373.815 443.645 ;
        RECT 374.245 443.365 374.525 443.645 ;
        RECT 374.955 443.365 375.235 443.645 ;
        RECT 375.665 443.365 375.945 443.645 ;
        RECT 376.375 443.365 376.655 443.645 ;
        RECT 369.275 442.655 369.555 442.935 ;
        RECT 369.985 442.655 370.265 442.935 ;
        RECT 370.695 442.655 370.975 442.935 ;
        RECT 371.405 442.655 371.685 442.935 ;
        RECT 372.115 442.655 372.395 442.935 ;
        RECT 372.825 442.655 373.105 442.935 ;
        RECT 373.535 442.655 373.815 442.935 ;
        RECT 374.245 442.655 374.525 442.935 ;
        RECT 374.955 442.655 375.235 442.935 ;
        RECT 375.665 442.655 375.945 442.935 ;
        RECT 376.375 442.655 376.655 442.935 ;
        RECT 369.275 441.945 369.555 442.225 ;
        RECT 369.985 441.945 370.265 442.225 ;
        RECT 370.695 441.945 370.975 442.225 ;
        RECT 371.405 441.945 371.685 442.225 ;
        RECT 372.115 441.945 372.395 442.225 ;
        RECT 372.825 441.945 373.105 442.225 ;
        RECT 373.535 441.945 373.815 442.225 ;
        RECT 374.245 441.945 374.525 442.225 ;
        RECT 374.955 441.945 375.235 442.225 ;
        RECT 375.665 441.945 375.945 442.225 ;
        RECT 376.375 441.945 376.655 442.225 ;
        RECT 369.275 441.235 369.555 441.515 ;
        RECT 369.985 441.235 370.265 441.515 ;
        RECT 370.695 441.235 370.975 441.515 ;
        RECT 371.405 441.235 371.685 441.515 ;
        RECT 372.115 441.235 372.395 441.515 ;
        RECT 372.825 441.235 373.105 441.515 ;
        RECT 373.535 441.235 373.815 441.515 ;
        RECT 374.245 441.235 374.525 441.515 ;
        RECT 374.955 441.235 375.235 441.515 ;
        RECT 375.665 441.235 375.945 441.515 ;
        RECT 376.375 441.235 376.655 441.515 ;
        RECT 369.275 440.525 369.555 440.805 ;
        RECT 369.985 440.525 370.265 440.805 ;
        RECT 370.695 440.525 370.975 440.805 ;
        RECT 371.405 440.525 371.685 440.805 ;
        RECT 372.115 440.525 372.395 440.805 ;
        RECT 372.825 440.525 373.105 440.805 ;
        RECT 373.535 440.525 373.815 440.805 ;
        RECT 374.245 440.525 374.525 440.805 ;
        RECT 374.955 440.525 375.235 440.805 ;
        RECT 375.665 440.525 375.945 440.805 ;
        RECT 376.375 440.525 376.655 440.805 ;
        RECT 369.275 439.815 369.555 440.095 ;
        RECT 369.985 439.815 370.265 440.095 ;
        RECT 370.695 439.815 370.975 440.095 ;
        RECT 371.405 439.815 371.685 440.095 ;
        RECT 372.115 439.815 372.395 440.095 ;
        RECT 372.825 439.815 373.105 440.095 ;
        RECT 373.535 439.815 373.815 440.095 ;
        RECT 374.245 439.815 374.525 440.095 ;
        RECT 374.955 439.815 375.235 440.095 ;
        RECT 375.665 439.815 375.945 440.095 ;
        RECT 376.375 439.815 376.655 440.095 ;
        RECT 369.275 439.105 369.555 439.385 ;
        RECT 369.985 439.105 370.265 439.385 ;
        RECT 370.695 439.105 370.975 439.385 ;
        RECT 371.405 439.105 371.685 439.385 ;
        RECT 372.115 439.105 372.395 439.385 ;
        RECT 372.825 439.105 373.105 439.385 ;
        RECT 373.535 439.105 373.815 439.385 ;
        RECT 374.245 439.105 374.525 439.385 ;
        RECT 374.955 439.105 375.235 439.385 ;
        RECT 375.665 439.105 375.945 439.385 ;
        RECT 376.375 439.105 376.655 439.385 ;
        RECT 369.330 435.190 369.610 435.470 ;
        RECT 370.040 435.190 370.320 435.470 ;
        RECT 370.750 435.190 371.030 435.470 ;
        RECT 371.460 435.190 371.740 435.470 ;
        RECT 372.170 435.190 372.450 435.470 ;
        RECT 372.880 435.190 373.160 435.470 ;
        RECT 373.590 435.190 373.870 435.470 ;
        RECT 374.300 435.190 374.580 435.470 ;
        RECT 375.010 435.190 375.290 435.470 ;
        RECT 375.720 435.190 376.000 435.470 ;
        RECT 376.430 435.190 376.710 435.470 ;
        RECT 369.330 434.480 369.610 434.760 ;
        RECT 370.040 434.480 370.320 434.760 ;
        RECT 370.750 434.480 371.030 434.760 ;
        RECT 371.460 434.480 371.740 434.760 ;
        RECT 372.170 434.480 372.450 434.760 ;
        RECT 372.880 434.480 373.160 434.760 ;
        RECT 373.590 434.480 373.870 434.760 ;
        RECT 374.300 434.480 374.580 434.760 ;
        RECT 375.010 434.480 375.290 434.760 ;
        RECT 375.720 434.480 376.000 434.760 ;
        RECT 376.430 434.480 376.710 434.760 ;
        RECT 369.330 433.770 369.610 434.050 ;
        RECT 370.040 433.770 370.320 434.050 ;
        RECT 370.750 433.770 371.030 434.050 ;
        RECT 371.460 433.770 371.740 434.050 ;
        RECT 372.170 433.770 372.450 434.050 ;
        RECT 372.880 433.770 373.160 434.050 ;
        RECT 373.590 433.770 373.870 434.050 ;
        RECT 374.300 433.770 374.580 434.050 ;
        RECT 375.010 433.770 375.290 434.050 ;
        RECT 375.720 433.770 376.000 434.050 ;
        RECT 376.430 433.770 376.710 434.050 ;
        RECT 369.330 433.060 369.610 433.340 ;
        RECT 370.040 433.060 370.320 433.340 ;
        RECT 370.750 433.060 371.030 433.340 ;
        RECT 371.460 433.060 371.740 433.340 ;
        RECT 372.170 433.060 372.450 433.340 ;
        RECT 372.880 433.060 373.160 433.340 ;
        RECT 373.590 433.060 373.870 433.340 ;
        RECT 374.300 433.060 374.580 433.340 ;
        RECT 375.010 433.060 375.290 433.340 ;
        RECT 375.720 433.060 376.000 433.340 ;
        RECT 376.430 433.060 376.710 433.340 ;
        RECT 369.330 432.350 369.610 432.630 ;
        RECT 370.040 432.350 370.320 432.630 ;
        RECT 370.750 432.350 371.030 432.630 ;
        RECT 371.460 432.350 371.740 432.630 ;
        RECT 372.170 432.350 372.450 432.630 ;
        RECT 372.880 432.350 373.160 432.630 ;
        RECT 373.590 432.350 373.870 432.630 ;
        RECT 374.300 432.350 374.580 432.630 ;
        RECT 375.010 432.350 375.290 432.630 ;
        RECT 375.720 432.350 376.000 432.630 ;
        RECT 376.430 432.350 376.710 432.630 ;
        RECT 369.330 431.640 369.610 431.920 ;
        RECT 370.040 431.640 370.320 431.920 ;
        RECT 370.750 431.640 371.030 431.920 ;
        RECT 371.460 431.640 371.740 431.920 ;
        RECT 372.170 431.640 372.450 431.920 ;
        RECT 372.880 431.640 373.160 431.920 ;
        RECT 373.590 431.640 373.870 431.920 ;
        RECT 374.300 431.640 374.580 431.920 ;
        RECT 375.010 431.640 375.290 431.920 ;
        RECT 375.720 431.640 376.000 431.920 ;
        RECT 376.430 431.640 376.710 431.920 ;
        RECT 369.330 430.930 369.610 431.210 ;
        RECT 370.040 430.930 370.320 431.210 ;
        RECT 370.750 430.930 371.030 431.210 ;
        RECT 371.460 430.930 371.740 431.210 ;
        RECT 372.170 430.930 372.450 431.210 ;
        RECT 372.880 430.930 373.160 431.210 ;
        RECT 373.590 430.930 373.870 431.210 ;
        RECT 374.300 430.930 374.580 431.210 ;
        RECT 375.010 430.930 375.290 431.210 ;
        RECT 375.720 430.930 376.000 431.210 ;
        RECT 376.430 430.930 376.710 431.210 ;
        RECT 369.330 430.220 369.610 430.500 ;
        RECT 370.040 430.220 370.320 430.500 ;
        RECT 370.750 430.220 371.030 430.500 ;
        RECT 371.460 430.220 371.740 430.500 ;
        RECT 372.170 430.220 372.450 430.500 ;
        RECT 372.880 430.220 373.160 430.500 ;
        RECT 373.590 430.220 373.870 430.500 ;
        RECT 374.300 430.220 374.580 430.500 ;
        RECT 375.010 430.220 375.290 430.500 ;
        RECT 375.720 430.220 376.000 430.500 ;
        RECT 376.430 430.220 376.710 430.500 ;
        RECT 369.330 429.510 369.610 429.790 ;
        RECT 370.040 429.510 370.320 429.790 ;
        RECT 370.750 429.510 371.030 429.790 ;
        RECT 371.460 429.510 371.740 429.790 ;
        RECT 372.170 429.510 372.450 429.790 ;
        RECT 372.880 429.510 373.160 429.790 ;
        RECT 373.590 429.510 373.870 429.790 ;
        RECT 374.300 429.510 374.580 429.790 ;
        RECT 375.010 429.510 375.290 429.790 ;
        RECT 375.720 429.510 376.000 429.790 ;
        RECT 376.430 429.510 376.710 429.790 ;
        RECT 369.330 428.800 369.610 429.080 ;
        RECT 370.040 428.800 370.320 429.080 ;
        RECT 370.750 428.800 371.030 429.080 ;
        RECT 371.460 428.800 371.740 429.080 ;
        RECT 372.170 428.800 372.450 429.080 ;
        RECT 372.880 428.800 373.160 429.080 ;
        RECT 373.590 428.800 373.870 429.080 ;
        RECT 374.300 428.800 374.580 429.080 ;
        RECT 375.010 428.800 375.290 429.080 ;
        RECT 375.720 428.800 376.000 429.080 ;
        RECT 376.430 428.800 376.710 429.080 ;
        RECT 369.330 428.090 369.610 428.370 ;
        RECT 370.040 428.090 370.320 428.370 ;
        RECT 370.750 428.090 371.030 428.370 ;
        RECT 371.460 428.090 371.740 428.370 ;
        RECT 372.170 428.090 372.450 428.370 ;
        RECT 372.880 428.090 373.160 428.370 ;
        RECT 373.590 428.090 373.870 428.370 ;
        RECT 374.300 428.090 374.580 428.370 ;
        RECT 375.010 428.090 375.290 428.370 ;
        RECT 375.720 428.090 376.000 428.370 ;
        RECT 376.430 428.090 376.710 428.370 ;
        RECT 369.330 427.380 369.610 427.660 ;
        RECT 370.040 427.380 370.320 427.660 ;
        RECT 370.750 427.380 371.030 427.660 ;
        RECT 371.460 427.380 371.740 427.660 ;
        RECT 372.170 427.380 372.450 427.660 ;
        RECT 372.880 427.380 373.160 427.660 ;
        RECT 373.590 427.380 373.870 427.660 ;
        RECT 374.300 427.380 374.580 427.660 ;
        RECT 375.010 427.380 375.290 427.660 ;
        RECT 375.720 427.380 376.000 427.660 ;
        RECT 376.430 427.380 376.710 427.660 ;
        RECT 369.330 426.670 369.610 426.950 ;
        RECT 370.040 426.670 370.320 426.950 ;
        RECT 370.750 426.670 371.030 426.950 ;
        RECT 371.460 426.670 371.740 426.950 ;
        RECT 372.170 426.670 372.450 426.950 ;
        RECT 372.880 426.670 373.160 426.950 ;
        RECT 373.590 426.670 373.870 426.950 ;
        RECT 374.300 426.670 374.580 426.950 ;
        RECT 375.010 426.670 375.290 426.950 ;
        RECT 375.720 426.670 376.000 426.950 ;
        RECT 376.430 426.670 376.710 426.950 ;
        RECT 3276.360 372.440 3282.100 380.440 ;
        RECT 3288.760 372.440 3299.010 380.440 ;
        RECT 3300.610 372.440 3310.860 380.440 ;
        RECT 3314.140 372.440 3324.390 380.440 ;
        RECT 3325.990 372.440 3336.240 380.440 ;
        RECT 3339.140 372.440 3348.640 380.440 ;
        RECT 526.360 360.440 535.860 370.440 ;
        RECT 544.740 360.440 549.010 370.440 ;
        RECT 550.610 360.440 560.860 370.440 ;
        RECT 564.140 360.440 574.390 370.440 ;
        RECT 575.990 360.440 586.240 370.440 ;
        RECT 589.140 360.440 598.640 370.440 ;
        RECT 1351.360 360.440 1360.860 370.440 ;
        RECT 1363.760 360.440 1374.010 370.440 ;
        RECT 1375.610 360.440 1385.860 370.440 ;
        RECT 1389.140 360.440 1399.390 370.440 ;
        RECT 1400.990 360.440 1411.240 370.440 ;
        RECT 1414.140 360.440 1420.080 370.440 ;
        RECT 3001.360 360.440 3010.860 370.440 ;
        RECT 3013.760 360.440 3020.200 370.440 ;
        RECT 3025.610 360.440 3035.860 370.440 ;
        RECT 3039.140 360.440 3049.390 370.440 ;
        RECT 3050.990 360.440 3061.240 370.440 ;
        RECT 3064.140 360.440 3073.640 370.440 ;
      LAYER Via4 ;
        RECT 1896.705 4708.095 1896.985 4708.375 ;
        RECT 1897.415 4708.095 1897.695 4708.375 ;
        RECT 1898.125 4708.095 1898.405 4708.375 ;
        RECT 1898.835 4708.095 1899.115 4708.375 ;
        RECT 1899.545 4708.095 1899.825 4708.375 ;
        RECT 1896.705 4707.385 1896.985 4707.665 ;
        RECT 1897.415 4707.385 1897.695 4707.665 ;
        RECT 1898.125 4707.385 1898.405 4707.665 ;
        RECT 1898.835 4707.385 1899.115 4707.665 ;
        RECT 1899.545 4707.385 1899.825 4707.665 ;
        RECT 1896.705 4706.675 1896.985 4706.955 ;
        RECT 1897.415 4706.675 1897.695 4706.955 ;
        RECT 1898.125 4706.675 1898.405 4706.955 ;
        RECT 1898.835 4706.675 1899.115 4706.955 ;
        RECT 1899.545 4706.675 1899.825 4706.955 ;
        RECT 1896.705 4705.965 1896.985 4706.245 ;
        RECT 1897.415 4705.965 1897.695 4706.245 ;
        RECT 1898.125 4705.965 1898.405 4706.245 ;
        RECT 1898.835 4705.965 1899.115 4706.245 ;
        RECT 1899.545 4705.965 1899.825 4706.245 ;
        RECT 1896.705 4705.255 1896.985 4705.535 ;
        RECT 1897.415 4705.255 1897.695 4705.535 ;
        RECT 1898.125 4705.255 1898.405 4705.535 ;
        RECT 1898.835 4705.255 1899.115 4705.535 ;
        RECT 1899.545 4705.255 1899.825 4705.535 ;
        RECT 1896.705 4704.545 1896.985 4704.825 ;
        RECT 1897.415 4704.545 1897.695 4704.825 ;
        RECT 1898.125 4704.545 1898.405 4704.825 ;
        RECT 1898.835 4704.545 1899.115 4704.825 ;
        RECT 1899.545 4704.545 1899.825 4704.825 ;
        RECT 1896.705 4703.835 1896.985 4704.115 ;
        RECT 1897.415 4703.835 1897.695 4704.115 ;
        RECT 1898.125 4703.835 1898.405 4704.115 ;
        RECT 1898.835 4703.835 1899.115 4704.115 ;
        RECT 1899.545 4703.835 1899.825 4704.115 ;
        RECT 1896.705 4703.125 1896.985 4703.405 ;
        RECT 1897.415 4703.125 1897.695 4703.405 ;
        RECT 1898.125 4703.125 1898.405 4703.405 ;
        RECT 1898.835 4703.125 1899.115 4703.405 ;
        RECT 1899.545 4703.125 1899.825 4703.405 ;
        RECT 1896.705 4702.415 1896.985 4702.695 ;
        RECT 1897.415 4702.415 1897.695 4702.695 ;
        RECT 1898.125 4702.415 1898.405 4702.695 ;
        RECT 1898.835 4702.415 1899.115 4702.695 ;
        RECT 1899.545 4702.415 1899.825 4702.695 ;
        RECT 1896.705 4701.705 1896.985 4701.985 ;
        RECT 1897.415 4701.705 1897.695 4701.985 ;
        RECT 1898.125 4701.705 1898.405 4701.985 ;
        RECT 1898.835 4701.705 1899.115 4701.985 ;
        RECT 1899.545 4701.705 1899.825 4701.985 ;
        RECT 1896.705 4700.995 1896.985 4701.275 ;
        RECT 1897.415 4700.995 1897.695 4701.275 ;
        RECT 1898.125 4700.995 1898.405 4701.275 ;
        RECT 1898.835 4700.995 1899.115 4701.275 ;
        RECT 1899.545 4700.995 1899.825 4701.275 ;
        RECT 1896.705 4700.285 1896.985 4700.565 ;
        RECT 1897.415 4700.285 1897.695 4700.565 ;
        RECT 1898.125 4700.285 1898.405 4700.565 ;
        RECT 1898.835 4700.285 1899.115 4700.565 ;
        RECT 1899.545 4700.285 1899.825 4700.565 ;
        RECT 1896.705 4699.575 1896.985 4699.855 ;
        RECT 1897.415 4699.575 1897.695 4699.855 ;
        RECT 1898.125 4699.575 1898.405 4699.855 ;
        RECT 1898.835 4699.575 1899.115 4699.855 ;
        RECT 1899.545 4699.575 1899.825 4699.855 ;
        RECT 1896.705 4698.865 1896.985 4699.145 ;
        RECT 1897.415 4698.865 1897.695 4699.145 ;
        RECT 1898.125 4698.865 1898.405 4699.145 ;
        RECT 1898.835 4698.865 1899.115 4699.145 ;
        RECT 1899.545 4698.865 1899.825 4699.145 ;
        RECT 1909.145 4708.095 1909.425 4708.375 ;
        RECT 1909.855 4708.095 1910.135 4708.375 ;
        RECT 1910.565 4708.095 1910.845 4708.375 ;
        RECT 1911.275 4708.095 1911.555 4708.375 ;
        RECT 1911.985 4708.095 1912.265 4708.375 ;
        RECT 1912.695 4708.095 1912.975 4708.375 ;
        RECT 1913.405 4708.095 1913.685 4708.375 ;
        RECT 1914.115 4708.095 1914.395 4708.375 ;
        RECT 1914.825 4708.095 1915.105 4708.375 ;
        RECT 1915.535 4708.095 1915.815 4708.375 ;
        RECT 1916.245 4708.095 1916.525 4708.375 ;
        RECT 1916.955 4708.095 1917.235 4708.375 ;
        RECT 1917.665 4708.095 1917.945 4708.375 ;
        RECT 1918.375 4708.095 1918.655 4708.375 ;
        RECT 1909.145 4707.385 1909.425 4707.665 ;
        RECT 1909.855 4707.385 1910.135 4707.665 ;
        RECT 1910.565 4707.385 1910.845 4707.665 ;
        RECT 1911.275 4707.385 1911.555 4707.665 ;
        RECT 1911.985 4707.385 1912.265 4707.665 ;
        RECT 1912.695 4707.385 1912.975 4707.665 ;
        RECT 1913.405 4707.385 1913.685 4707.665 ;
        RECT 1914.115 4707.385 1914.395 4707.665 ;
        RECT 1914.825 4707.385 1915.105 4707.665 ;
        RECT 1915.535 4707.385 1915.815 4707.665 ;
        RECT 1916.245 4707.385 1916.525 4707.665 ;
        RECT 1916.955 4707.385 1917.235 4707.665 ;
        RECT 1917.665 4707.385 1917.945 4707.665 ;
        RECT 1918.375 4707.385 1918.655 4707.665 ;
        RECT 1909.145 4706.675 1909.425 4706.955 ;
        RECT 1909.855 4706.675 1910.135 4706.955 ;
        RECT 1910.565 4706.675 1910.845 4706.955 ;
        RECT 1911.275 4706.675 1911.555 4706.955 ;
        RECT 1911.985 4706.675 1912.265 4706.955 ;
        RECT 1912.695 4706.675 1912.975 4706.955 ;
        RECT 1913.405 4706.675 1913.685 4706.955 ;
        RECT 1914.115 4706.675 1914.395 4706.955 ;
        RECT 1914.825 4706.675 1915.105 4706.955 ;
        RECT 1915.535 4706.675 1915.815 4706.955 ;
        RECT 1916.245 4706.675 1916.525 4706.955 ;
        RECT 1916.955 4706.675 1917.235 4706.955 ;
        RECT 1917.665 4706.675 1917.945 4706.955 ;
        RECT 1918.375 4706.675 1918.655 4706.955 ;
        RECT 1909.145 4705.965 1909.425 4706.245 ;
        RECT 1909.855 4705.965 1910.135 4706.245 ;
        RECT 1910.565 4705.965 1910.845 4706.245 ;
        RECT 1911.275 4705.965 1911.555 4706.245 ;
        RECT 1911.985 4705.965 1912.265 4706.245 ;
        RECT 1912.695 4705.965 1912.975 4706.245 ;
        RECT 1913.405 4705.965 1913.685 4706.245 ;
        RECT 1914.115 4705.965 1914.395 4706.245 ;
        RECT 1914.825 4705.965 1915.105 4706.245 ;
        RECT 1915.535 4705.965 1915.815 4706.245 ;
        RECT 1916.245 4705.965 1916.525 4706.245 ;
        RECT 1916.955 4705.965 1917.235 4706.245 ;
        RECT 1917.665 4705.965 1917.945 4706.245 ;
        RECT 1918.375 4705.965 1918.655 4706.245 ;
        RECT 1909.145 4705.255 1909.425 4705.535 ;
        RECT 1909.855 4705.255 1910.135 4705.535 ;
        RECT 1910.565 4705.255 1910.845 4705.535 ;
        RECT 1911.275 4705.255 1911.555 4705.535 ;
        RECT 1911.985 4705.255 1912.265 4705.535 ;
        RECT 1912.695 4705.255 1912.975 4705.535 ;
        RECT 1913.405 4705.255 1913.685 4705.535 ;
        RECT 1914.115 4705.255 1914.395 4705.535 ;
        RECT 1914.825 4705.255 1915.105 4705.535 ;
        RECT 1915.535 4705.255 1915.815 4705.535 ;
        RECT 1916.245 4705.255 1916.525 4705.535 ;
        RECT 1916.955 4705.255 1917.235 4705.535 ;
        RECT 1917.665 4705.255 1917.945 4705.535 ;
        RECT 1918.375 4705.255 1918.655 4705.535 ;
        RECT 1909.145 4704.545 1909.425 4704.825 ;
        RECT 1909.855 4704.545 1910.135 4704.825 ;
        RECT 1910.565 4704.545 1910.845 4704.825 ;
        RECT 1911.275 4704.545 1911.555 4704.825 ;
        RECT 1911.985 4704.545 1912.265 4704.825 ;
        RECT 1912.695 4704.545 1912.975 4704.825 ;
        RECT 1913.405 4704.545 1913.685 4704.825 ;
        RECT 1914.115 4704.545 1914.395 4704.825 ;
        RECT 1914.825 4704.545 1915.105 4704.825 ;
        RECT 1915.535 4704.545 1915.815 4704.825 ;
        RECT 1916.245 4704.545 1916.525 4704.825 ;
        RECT 1916.955 4704.545 1917.235 4704.825 ;
        RECT 1917.665 4704.545 1917.945 4704.825 ;
        RECT 1918.375 4704.545 1918.655 4704.825 ;
        RECT 1909.145 4703.835 1909.425 4704.115 ;
        RECT 1909.855 4703.835 1910.135 4704.115 ;
        RECT 1910.565 4703.835 1910.845 4704.115 ;
        RECT 1911.275 4703.835 1911.555 4704.115 ;
        RECT 1911.985 4703.835 1912.265 4704.115 ;
        RECT 1912.695 4703.835 1912.975 4704.115 ;
        RECT 1913.405 4703.835 1913.685 4704.115 ;
        RECT 1914.115 4703.835 1914.395 4704.115 ;
        RECT 1914.825 4703.835 1915.105 4704.115 ;
        RECT 1915.535 4703.835 1915.815 4704.115 ;
        RECT 1916.245 4703.835 1916.525 4704.115 ;
        RECT 1916.955 4703.835 1917.235 4704.115 ;
        RECT 1917.665 4703.835 1917.945 4704.115 ;
        RECT 1918.375 4703.835 1918.655 4704.115 ;
        RECT 1909.145 4703.125 1909.425 4703.405 ;
        RECT 1909.855 4703.125 1910.135 4703.405 ;
        RECT 1910.565 4703.125 1910.845 4703.405 ;
        RECT 1911.275 4703.125 1911.555 4703.405 ;
        RECT 1911.985 4703.125 1912.265 4703.405 ;
        RECT 1912.695 4703.125 1912.975 4703.405 ;
        RECT 1913.405 4703.125 1913.685 4703.405 ;
        RECT 1914.115 4703.125 1914.395 4703.405 ;
        RECT 1914.825 4703.125 1915.105 4703.405 ;
        RECT 1915.535 4703.125 1915.815 4703.405 ;
        RECT 1916.245 4703.125 1916.525 4703.405 ;
        RECT 1916.955 4703.125 1917.235 4703.405 ;
        RECT 1917.665 4703.125 1917.945 4703.405 ;
        RECT 1918.375 4703.125 1918.655 4703.405 ;
        RECT 1909.145 4702.415 1909.425 4702.695 ;
        RECT 1909.855 4702.415 1910.135 4702.695 ;
        RECT 1910.565 4702.415 1910.845 4702.695 ;
        RECT 1911.275 4702.415 1911.555 4702.695 ;
        RECT 1911.985 4702.415 1912.265 4702.695 ;
        RECT 1912.695 4702.415 1912.975 4702.695 ;
        RECT 1913.405 4702.415 1913.685 4702.695 ;
        RECT 1914.115 4702.415 1914.395 4702.695 ;
        RECT 1914.825 4702.415 1915.105 4702.695 ;
        RECT 1915.535 4702.415 1915.815 4702.695 ;
        RECT 1916.245 4702.415 1916.525 4702.695 ;
        RECT 1916.955 4702.415 1917.235 4702.695 ;
        RECT 1917.665 4702.415 1917.945 4702.695 ;
        RECT 1918.375 4702.415 1918.655 4702.695 ;
        RECT 1909.145 4701.705 1909.425 4701.985 ;
        RECT 1909.855 4701.705 1910.135 4701.985 ;
        RECT 1910.565 4701.705 1910.845 4701.985 ;
        RECT 1911.275 4701.705 1911.555 4701.985 ;
        RECT 1911.985 4701.705 1912.265 4701.985 ;
        RECT 1912.695 4701.705 1912.975 4701.985 ;
        RECT 1913.405 4701.705 1913.685 4701.985 ;
        RECT 1914.115 4701.705 1914.395 4701.985 ;
        RECT 1914.825 4701.705 1915.105 4701.985 ;
        RECT 1915.535 4701.705 1915.815 4701.985 ;
        RECT 1916.245 4701.705 1916.525 4701.985 ;
        RECT 1916.955 4701.705 1917.235 4701.985 ;
        RECT 1917.665 4701.705 1917.945 4701.985 ;
        RECT 1918.375 4701.705 1918.655 4701.985 ;
        RECT 1909.145 4700.995 1909.425 4701.275 ;
        RECT 1909.855 4700.995 1910.135 4701.275 ;
        RECT 1910.565 4700.995 1910.845 4701.275 ;
        RECT 1911.275 4700.995 1911.555 4701.275 ;
        RECT 1911.985 4700.995 1912.265 4701.275 ;
        RECT 1912.695 4700.995 1912.975 4701.275 ;
        RECT 1913.405 4700.995 1913.685 4701.275 ;
        RECT 1914.115 4700.995 1914.395 4701.275 ;
        RECT 1914.825 4700.995 1915.105 4701.275 ;
        RECT 1915.535 4700.995 1915.815 4701.275 ;
        RECT 1916.245 4700.995 1916.525 4701.275 ;
        RECT 1916.955 4700.995 1917.235 4701.275 ;
        RECT 1917.665 4700.995 1917.945 4701.275 ;
        RECT 1918.375 4700.995 1918.655 4701.275 ;
        RECT 1909.145 4700.285 1909.425 4700.565 ;
        RECT 1909.855 4700.285 1910.135 4700.565 ;
        RECT 1910.565 4700.285 1910.845 4700.565 ;
        RECT 1911.275 4700.285 1911.555 4700.565 ;
        RECT 1911.985 4700.285 1912.265 4700.565 ;
        RECT 1912.695 4700.285 1912.975 4700.565 ;
        RECT 1913.405 4700.285 1913.685 4700.565 ;
        RECT 1914.115 4700.285 1914.395 4700.565 ;
        RECT 1914.825 4700.285 1915.105 4700.565 ;
        RECT 1915.535 4700.285 1915.815 4700.565 ;
        RECT 1916.245 4700.285 1916.525 4700.565 ;
        RECT 1916.955 4700.285 1917.235 4700.565 ;
        RECT 1917.665 4700.285 1917.945 4700.565 ;
        RECT 1918.375 4700.285 1918.655 4700.565 ;
        RECT 1909.145 4699.575 1909.425 4699.855 ;
        RECT 1909.855 4699.575 1910.135 4699.855 ;
        RECT 1910.565 4699.575 1910.845 4699.855 ;
        RECT 1911.275 4699.575 1911.555 4699.855 ;
        RECT 1911.985 4699.575 1912.265 4699.855 ;
        RECT 1912.695 4699.575 1912.975 4699.855 ;
        RECT 1913.405 4699.575 1913.685 4699.855 ;
        RECT 1914.115 4699.575 1914.395 4699.855 ;
        RECT 1914.825 4699.575 1915.105 4699.855 ;
        RECT 1915.535 4699.575 1915.815 4699.855 ;
        RECT 1916.245 4699.575 1916.525 4699.855 ;
        RECT 1916.955 4699.575 1917.235 4699.855 ;
        RECT 1917.665 4699.575 1917.945 4699.855 ;
        RECT 1918.375 4699.575 1918.655 4699.855 ;
        RECT 1909.145 4698.865 1909.425 4699.145 ;
        RECT 1909.855 4698.865 1910.135 4699.145 ;
        RECT 1910.565 4698.865 1910.845 4699.145 ;
        RECT 1911.275 4698.865 1911.555 4699.145 ;
        RECT 1911.985 4698.865 1912.265 4699.145 ;
        RECT 1912.695 4698.865 1912.975 4699.145 ;
        RECT 1913.405 4698.865 1913.685 4699.145 ;
        RECT 1914.115 4698.865 1914.395 4699.145 ;
        RECT 1914.825 4698.865 1915.105 4699.145 ;
        RECT 1915.535 4698.865 1915.815 4699.145 ;
        RECT 1916.245 4698.865 1916.525 4699.145 ;
        RECT 1916.955 4698.865 1917.235 4699.145 ;
        RECT 1917.665 4698.865 1917.945 4699.145 ;
        RECT 1918.375 4698.865 1918.655 4699.145 ;
        RECT 1920.995 4708.095 1921.275 4708.375 ;
        RECT 1921.705 4708.095 1921.985 4708.375 ;
        RECT 1922.415 4708.095 1922.695 4708.375 ;
        RECT 1926.675 4708.095 1926.955 4708.375 ;
        RECT 1927.385 4708.095 1927.665 4708.375 ;
        RECT 1928.095 4708.095 1928.375 4708.375 ;
        RECT 1928.805 4708.095 1929.085 4708.375 ;
        RECT 1929.515 4708.095 1929.795 4708.375 ;
        RECT 1930.225 4708.095 1930.505 4708.375 ;
        RECT 1920.995 4707.385 1921.275 4707.665 ;
        RECT 1921.705 4707.385 1921.985 4707.665 ;
        RECT 1922.415 4707.385 1922.695 4707.665 ;
        RECT 1926.675 4707.385 1926.955 4707.665 ;
        RECT 1927.385 4707.385 1927.665 4707.665 ;
        RECT 1928.095 4707.385 1928.375 4707.665 ;
        RECT 1928.805 4707.385 1929.085 4707.665 ;
        RECT 1929.515 4707.385 1929.795 4707.665 ;
        RECT 1930.225 4707.385 1930.505 4707.665 ;
        RECT 1920.995 4706.675 1921.275 4706.955 ;
        RECT 1921.705 4706.675 1921.985 4706.955 ;
        RECT 1922.415 4706.675 1922.695 4706.955 ;
        RECT 1926.675 4706.675 1926.955 4706.955 ;
        RECT 1927.385 4706.675 1927.665 4706.955 ;
        RECT 1928.095 4706.675 1928.375 4706.955 ;
        RECT 1928.805 4706.675 1929.085 4706.955 ;
        RECT 1929.515 4706.675 1929.795 4706.955 ;
        RECT 1930.225 4706.675 1930.505 4706.955 ;
        RECT 1920.995 4705.965 1921.275 4706.245 ;
        RECT 1921.705 4705.965 1921.985 4706.245 ;
        RECT 1922.415 4705.965 1922.695 4706.245 ;
        RECT 1926.675 4705.965 1926.955 4706.245 ;
        RECT 1927.385 4705.965 1927.665 4706.245 ;
        RECT 1928.095 4705.965 1928.375 4706.245 ;
        RECT 1928.805 4705.965 1929.085 4706.245 ;
        RECT 1929.515 4705.965 1929.795 4706.245 ;
        RECT 1930.225 4705.965 1930.505 4706.245 ;
        RECT 1920.995 4705.255 1921.275 4705.535 ;
        RECT 1921.705 4705.255 1921.985 4705.535 ;
        RECT 1922.415 4705.255 1922.695 4705.535 ;
        RECT 1926.675 4705.255 1926.955 4705.535 ;
        RECT 1927.385 4705.255 1927.665 4705.535 ;
        RECT 1928.095 4705.255 1928.375 4705.535 ;
        RECT 1928.805 4705.255 1929.085 4705.535 ;
        RECT 1929.515 4705.255 1929.795 4705.535 ;
        RECT 1930.225 4705.255 1930.505 4705.535 ;
        RECT 1920.995 4704.545 1921.275 4704.825 ;
        RECT 1921.705 4704.545 1921.985 4704.825 ;
        RECT 1922.415 4704.545 1922.695 4704.825 ;
        RECT 1926.675 4704.545 1926.955 4704.825 ;
        RECT 1927.385 4704.545 1927.665 4704.825 ;
        RECT 1928.095 4704.545 1928.375 4704.825 ;
        RECT 1928.805 4704.545 1929.085 4704.825 ;
        RECT 1929.515 4704.545 1929.795 4704.825 ;
        RECT 1930.225 4704.545 1930.505 4704.825 ;
        RECT 1920.995 4703.835 1921.275 4704.115 ;
        RECT 1921.705 4703.835 1921.985 4704.115 ;
        RECT 1922.415 4703.835 1922.695 4704.115 ;
        RECT 1926.675 4703.835 1926.955 4704.115 ;
        RECT 1927.385 4703.835 1927.665 4704.115 ;
        RECT 1928.095 4703.835 1928.375 4704.115 ;
        RECT 1928.805 4703.835 1929.085 4704.115 ;
        RECT 1929.515 4703.835 1929.795 4704.115 ;
        RECT 1930.225 4703.835 1930.505 4704.115 ;
        RECT 1920.995 4703.125 1921.275 4703.405 ;
        RECT 1921.705 4703.125 1921.985 4703.405 ;
        RECT 1922.415 4703.125 1922.695 4703.405 ;
        RECT 1926.675 4703.125 1926.955 4703.405 ;
        RECT 1927.385 4703.125 1927.665 4703.405 ;
        RECT 1928.095 4703.125 1928.375 4703.405 ;
        RECT 1928.805 4703.125 1929.085 4703.405 ;
        RECT 1929.515 4703.125 1929.795 4703.405 ;
        RECT 1930.225 4703.125 1930.505 4703.405 ;
        RECT 1920.995 4702.415 1921.275 4702.695 ;
        RECT 1921.705 4702.415 1921.985 4702.695 ;
        RECT 1922.415 4702.415 1922.695 4702.695 ;
        RECT 1926.675 4702.415 1926.955 4702.695 ;
        RECT 1927.385 4702.415 1927.665 4702.695 ;
        RECT 1928.095 4702.415 1928.375 4702.695 ;
        RECT 1928.805 4702.415 1929.085 4702.695 ;
        RECT 1929.515 4702.415 1929.795 4702.695 ;
        RECT 1930.225 4702.415 1930.505 4702.695 ;
        RECT 1920.995 4701.705 1921.275 4701.985 ;
        RECT 1921.705 4701.705 1921.985 4701.985 ;
        RECT 1922.415 4701.705 1922.695 4701.985 ;
        RECT 1926.675 4701.705 1926.955 4701.985 ;
        RECT 1927.385 4701.705 1927.665 4701.985 ;
        RECT 1928.095 4701.705 1928.375 4701.985 ;
        RECT 1928.805 4701.705 1929.085 4701.985 ;
        RECT 1929.515 4701.705 1929.795 4701.985 ;
        RECT 1930.225 4701.705 1930.505 4701.985 ;
        RECT 1920.995 4700.995 1921.275 4701.275 ;
        RECT 1921.705 4700.995 1921.985 4701.275 ;
        RECT 1922.415 4700.995 1922.695 4701.275 ;
        RECT 1926.675 4700.995 1926.955 4701.275 ;
        RECT 1927.385 4700.995 1927.665 4701.275 ;
        RECT 1928.095 4700.995 1928.375 4701.275 ;
        RECT 1928.805 4700.995 1929.085 4701.275 ;
        RECT 1929.515 4700.995 1929.795 4701.275 ;
        RECT 1930.225 4700.995 1930.505 4701.275 ;
        RECT 1920.995 4700.285 1921.275 4700.565 ;
        RECT 1921.705 4700.285 1921.985 4700.565 ;
        RECT 1922.415 4700.285 1922.695 4700.565 ;
        RECT 1926.675 4700.285 1926.955 4700.565 ;
        RECT 1927.385 4700.285 1927.665 4700.565 ;
        RECT 1928.095 4700.285 1928.375 4700.565 ;
        RECT 1928.805 4700.285 1929.085 4700.565 ;
        RECT 1929.515 4700.285 1929.795 4700.565 ;
        RECT 1930.225 4700.285 1930.505 4700.565 ;
        RECT 1920.995 4699.575 1921.275 4699.855 ;
        RECT 1921.705 4699.575 1921.985 4699.855 ;
        RECT 1922.415 4699.575 1922.695 4699.855 ;
        RECT 1926.675 4699.575 1926.955 4699.855 ;
        RECT 1927.385 4699.575 1927.665 4699.855 ;
        RECT 1928.095 4699.575 1928.375 4699.855 ;
        RECT 1928.805 4699.575 1929.085 4699.855 ;
        RECT 1929.515 4699.575 1929.795 4699.855 ;
        RECT 1930.225 4699.575 1930.505 4699.855 ;
        RECT 1920.995 4698.865 1921.275 4699.145 ;
        RECT 1921.705 4698.865 1921.985 4699.145 ;
        RECT 1922.415 4698.865 1922.695 4699.145 ;
        RECT 1926.675 4698.865 1926.955 4699.145 ;
        RECT 1927.385 4698.865 1927.665 4699.145 ;
        RECT 1928.095 4698.865 1928.375 4699.145 ;
        RECT 1928.805 4698.865 1929.085 4699.145 ;
        RECT 1929.515 4698.865 1929.795 4699.145 ;
        RECT 1930.225 4698.865 1930.505 4699.145 ;
        RECT 1934.525 4708.095 1934.805 4708.375 ;
        RECT 1935.235 4708.095 1935.515 4708.375 ;
        RECT 1935.945 4708.095 1936.225 4708.375 ;
        RECT 1936.655 4708.095 1936.935 4708.375 ;
        RECT 1937.365 4708.095 1937.645 4708.375 ;
        RECT 1938.075 4708.095 1938.355 4708.375 ;
        RECT 1938.785 4708.095 1939.065 4708.375 ;
        RECT 1939.495 4708.095 1939.775 4708.375 ;
        RECT 1940.205 4708.095 1940.485 4708.375 ;
        RECT 1940.915 4708.095 1941.195 4708.375 ;
        RECT 1941.625 4708.095 1941.905 4708.375 ;
        RECT 1942.335 4708.095 1942.615 4708.375 ;
        RECT 1943.045 4708.095 1943.325 4708.375 ;
        RECT 1943.755 4708.095 1944.035 4708.375 ;
        RECT 1934.525 4707.385 1934.805 4707.665 ;
        RECT 1935.235 4707.385 1935.515 4707.665 ;
        RECT 1935.945 4707.385 1936.225 4707.665 ;
        RECT 1936.655 4707.385 1936.935 4707.665 ;
        RECT 1937.365 4707.385 1937.645 4707.665 ;
        RECT 1938.075 4707.385 1938.355 4707.665 ;
        RECT 1938.785 4707.385 1939.065 4707.665 ;
        RECT 1939.495 4707.385 1939.775 4707.665 ;
        RECT 1940.205 4707.385 1940.485 4707.665 ;
        RECT 1940.915 4707.385 1941.195 4707.665 ;
        RECT 1941.625 4707.385 1941.905 4707.665 ;
        RECT 1942.335 4707.385 1942.615 4707.665 ;
        RECT 1943.045 4707.385 1943.325 4707.665 ;
        RECT 1943.755 4707.385 1944.035 4707.665 ;
        RECT 1934.525 4706.675 1934.805 4706.955 ;
        RECT 1935.235 4706.675 1935.515 4706.955 ;
        RECT 1935.945 4706.675 1936.225 4706.955 ;
        RECT 1936.655 4706.675 1936.935 4706.955 ;
        RECT 1937.365 4706.675 1937.645 4706.955 ;
        RECT 1938.075 4706.675 1938.355 4706.955 ;
        RECT 1938.785 4706.675 1939.065 4706.955 ;
        RECT 1939.495 4706.675 1939.775 4706.955 ;
        RECT 1940.205 4706.675 1940.485 4706.955 ;
        RECT 1940.915 4706.675 1941.195 4706.955 ;
        RECT 1941.625 4706.675 1941.905 4706.955 ;
        RECT 1942.335 4706.675 1942.615 4706.955 ;
        RECT 1943.045 4706.675 1943.325 4706.955 ;
        RECT 1943.755 4706.675 1944.035 4706.955 ;
        RECT 1934.525 4705.965 1934.805 4706.245 ;
        RECT 1935.235 4705.965 1935.515 4706.245 ;
        RECT 1935.945 4705.965 1936.225 4706.245 ;
        RECT 1936.655 4705.965 1936.935 4706.245 ;
        RECT 1937.365 4705.965 1937.645 4706.245 ;
        RECT 1938.075 4705.965 1938.355 4706.245 ;
        RECT 1938.785 4705.965 1939.065 4706.245 ;
        RECT 1939.495 4705.965 1939.775 4706.245 ;
        RECT 1940.205 4705.965 1940.485 4706.245 ;
        RECT 1940.915 4705.965 1941.195 4706.245 ;
        RECT 1941.625 4705.965 1941.905 4706.245 ;
        RECT 1942.335 4705.965 1942.615 4706.245 ;
        RECT 1943.045 4705.965 1943.325 4706.245 ;
        RECT 1943.755 4705.965 1944.035 4706.245 ;
        RECT 1934.525 4705.255 1934.805 4705.535 ;
        RECT 1935.235 4705.255 1935.515 4705.535 ;
        RECT 1935.945 4705.255 1936.225 4705.535 ;
        RECT 1936.655 4705.255 1936.935 4705.535 ;
        RECT 1937.365 4705.255 1937.645 4705.535 ;
        RECT 1938.075 4705.255 1938.355 4705.535 ;
        RECT 1938.785 4705.255 1939.065 4705.535 ;
        RECT 1939.495 4705.255 1939.775 4705.535 ;
        RECT 1940.205 4705.255 1940.485 4705.535 ;
        RECT 1940.915 4705.255 1941.195 4705.535 ;
        RECT 1941.625 4705.255 1941.905 4705.535 ;
        RECT 1942.335 4705.255 1942.615 4705.535 ;
        RECT 1943.045 4705.255 1943.325 4705.535 ;
        RECT 1943.755 4705.255 1944.035 4705.535 ;
        RECT 1934.525 4704.545 1934.805 4704.825 ;
        RECT 1935.235 4704.545 1935.515 4704.825 ;
        RECT 1935.945 4704.545 1936.225 4704.825 ;
        RECT 1936.655 4704.545 1936.935 4704.825 ;
        RECT 1937.365 4704.545 1937.645 4704.825 ;
        RECT 1938.075 4704.545 1938.355 4704.825 ;
        RECT 1938.785 4704.545 1939.065 4704.825 ;
        RECT 1939.495 4704.545 1939.775 4704.825 ;
        RECT 1940.205 4704.545 1940.485 4704.825 ;
        RECT 1940.915 4704.545 1941.195 4704.825 ;
        RECT 1941.625 4704.545 1941.905 4704.825 ;
        RECT 1942.335 4704.545 1942.615 4704.825 ;
        RECT 1943.045 4704.545 1943.325 4704.825 ;
        RECT 1943.755 4704.545 1944.035 4704.825 ;
        RECT 1934.525 4703.835 1934.805 4704.115 ;
        RECT 1935.235 4703.835 1935.515 4704.115 ;
        RECT 1935.945 4703.835 1936.225 4704.115 ;
        RECT 1936.655 4703.835 1936.935 4704.115 ;
        RECT 1937.365 4703.835 1937.645 4704.115 ;
        RECT 1938.075 4703.835 1938.355 4704.115 ;
        RECT 1938.785 4703.835 1939.065 4704.115 ;
        RECT 1939.495 4703.835 1939.775 4704.115 ;
        RECT 1940.205 4703.835 1940.485 4704.115 ;
        RECT 1940.915 4703.835 1941.195 4704.115 ;
        RECT 1941.625 4703.835 1941.905 4704.115 ;
        RECT 1942.335 4703.835 1942.615 4704.115 ;
        RECT 1943.045 4703.835 1943.325 4704.115 ;
        RECT 1943.755 4703.835 1944.035 4704.115 ;
        RECT 1934.525 4703.125 1934.805 4703.405 ;
        RECT 1935.235 4703.125 1935.515 4703.405 ;
        RECT 1935.945 4703.125 1936.225 4703.405 ;
        RECT 1936.655 4703.125 1936.935 4703.405 ;
        RECT 1937.365 4703.125 1937.645 4703.405 ;
        RECT 1938.075 4703.125 1938.355 4703.405 ;
        RECT 1938.785 4703.125 1939.065 4703.405 ;
        RECT 1939.495 4703.125 1939.775 4703.405 ;
        RECT 1940.205 4703.125 1940.485 4703.405 ;
        RECT 1940.915 4703.125 1941.195 4703.405 ;
        RECT 1941.625 4703.125 1941.905 4703.405 ;
        RECT 1942.335 4703.125 1942.615 4703.405 ;
        RECT 1943.045 4703.125 1943.325 4703.405 ;
        RECT 1943.755 4703.125 1944.035 4703.405 ;
        RECT 1934.525 4702.415 1934.805 4702.695 ;
        RECT 1935.235 4702.415 1935.515 4702.695 ;
        RECT 1935.945 4702.415 1936.225 4702.695 ;
        RECT 1936.655 4702.415 1936.935 4702.695 ;
        RECT 1937.365 4702.415 1937.645 4702.695 ;
        RECT 1938.075 4702.415 1938.355 4702.695 ;
        RECT 1938.785 4702.415 1939.065 4702.695 ;
        RECT 1939.495 4702.415 1939.775 4702.695 ;
        RECT 1940.205 4702.415 1940.485 4702.695 ;
        RECT 1940.915 4702.415 1941.195 4702.695 ;
        RECT 1941.625 4702.415 1941.905 4702.695 ;
        RECT 1942.335 4702.415 1942.615 4702.695 ;
        RECT 1943.045 4702.415 1943.325 4702.695 ;
        RECT 1943.755 4702.415 1944.035 4702.695 ;
        RECT 1934.525 4701.705 1934.805 4701.985 ;
        RECT 1935.235 4701.705 1935.515 4701.985 ;
        RECT 1935.945 4701.705 1936.225 4701.985 ;
        RECT 1936.655 4701.705 1936.935 4701.985 ;
        RECT 1937.365 4701.705 1937.645 4701.985 ;
        RECT 1938.075 4701.705 1938.355 4701.985 ;
        RECT 1938.785 4701.705 1939.065 4701.985 ;
        RECT 1939.495 4701.705 1939.775 4701.985 ;
        RECT 1940.205 4701.705 1940.485 4701.985 ;
        RECT 1940.915 4701.705 1941.195 4701.985 ;
        RECT 1941.625 4701.705 1941.905 4701.985 ;
        RECT 1942.335 4701.705 1942.615 4701.985 ;
        RECT 1943.045 4701.705 1943.325 4701.985 ;
        RECT 1943.755 4701.705 1944.035 4701.985 ;
        RECT 1934.525 4700.995 1934.805 4701.275 ;
        RECT 1935.235 4700.995 1935.515 4701.275 ;
        RECT 1935.945 4700.995 1936.225 4701.275 ;
        RECT 1936.655 4700.995 1936.935 4701.275 ;
        RECT 1937.365 4700.995 1937.645 4701.275 ;
        RECT 1938.075 4700.995 1938.355 4701.275 ;
        RECT 1938.785 4700.995 1939.065 4701.275 ;
        RECT 1939.495 4700.995 1939.775 4701.275 ;
        RECT 1940.205 4700.995 1940.485 4701.275 ;
        RECT 1940.915 4700.995 1941.195 4701.275 ;
        RECT 1941.625 4700.995 1941.905 4701.275 ;
        RECT 1942.335 4700.995 1942.615 4701.275 ;
        RECT 1943.045 4700.995 1943.325 4701.275 ;
        RECT 1943.755 4700.995 1944.035 4701.275 ;
        RECT 1934.525 4700.285 1934.805 4700.565 ;
        RECT 1935.235 4700.285 1935.515 4700.565 ;
        RECT 1935.945 4700.285 1936.225 4700.565 ;
        RECT 1936.655 4700.285 1936.935 4700.565 ;
        RECT 1937.365 4700.285 1937.645 4700.565 ;
        RECT 1938.075 4700.285 1938.355 4700.565 ;
        RECT 1938.785 4700.285 1939.065 4700.565 ;
        RECT 1939.495 4700.285 1939.775 4700.565 ;
        RECT 1940.205 4700.285 1940.485 4700.565 ;
        RECT 1940.915 4700.285 1941.195 4700.565 ;
        RECT 1941.625 4700.285 1941.905 4700.565 ;
        RECT 1942.335 4700.285 1942.615 4700.565 ;
        RECT 1943.045 4700.285 1943.325 4700.565 ;
        RECT 1943.755 4700.285 1944.035 4700.565 ;
        RECT 1934.525 4699.575 1934.805 4699.855 ;
        RECT 1935.235 4699.575 1935.515 4699.855 ;
        RECT 1935.945 4699.575 1936.225 4699.855 ;
        RECT 1936.655 4699.575 1936.935 4699.855 ;
        RECT 1937.365 4699.575 1937.645 4699.855 ;
        RECT 1938.075 4699.575 1938.355 4699.855 ;
        RECT 1938.785 4699.575 1939.065 4699.855 ;
        RECT 1939.495 4699.575 1939.775 4699.855 ;
        RECT 1940.205 4699.575 1940.485 4699.855 ;
        RECT 1940.915 4699.575 1941.195 4699.855 ;
        RECT 1941.625 4699.575 1941.905 4699.855 ;
        RECT 1942.335 4699.575 1942.615 4699.855 ;
        RECT 1943.045 4699.575 1943.325 4699.855 ;
        RECT 1943.755 4699.575 1944.035 4699.855 ;
        RECT 1934.525 4698.865 1934.805 4699.145 ;
        RECT 1935.235 4698.865 1935.515 4699.145 ;
        RECT 1935.945 4698.865 1936.225 4699.145 ;
        RECT 1936.655 4698.865 1936.935 4699.145 ;
        RECT 1937.365 4698.865 1937.645 4699.145 ;
        RECT 1938.075 4698.865 1938.355 4699.145 ;
        RECT 1938.785 4698.865 1939.065 4699.145 ;
        RECT 1939.495 4698.865 1939.775 4699.145 ;
        RECT 1940.205 4698.865 1940.485 4699.145 ;
        RECT 1940.915 4698.865 1941.195 4699.145 ;
        RECT 1941.625 4698.865 1941.905 4699.145 ;
        RECT 1942.335 4698.865 1942.615 4699.145 ;
        RECT 1943.045 4698.865 1943.325 4699.145 ;
        RECT 1943.755 4698.865 1944.035 4699.145 ;
        RECT 1946.375 4708.095 1946.655 4708.375 ;
        RECT 1947.085 4708.095 1947.365 4708.375 ;
        RECT 1947.795 4708.095 1948.075 4708.375 ;
        RECT 1948.505 4708.095 1948.785 4708.375 ;
        RECT 1949.215 4708.095 1949.495 4708.375 ;
        RECT 1949.925 4708.095 1950.205 4708.375 ;
        RECT 1950.635 4708.095 1950.915 4708.375 ;
        RECT 1951.345 4708.095 1951.625 4708.375 ;
        RECT 1952.055 4708.095 1952.335 4708.375 ;
        RECT 1952.765 4708.095 1953.045 4708.375 ;
        RECT 1953.475 4708.095 1953.755 4708.375 ;
        RECT 1954.185 4708.095 1954.465 4708.375 ;
        RECT 1954.895 4708.095 1955.175 4708.375 ;
        RECT 1955.605 4708.095 1955.885 4708.375 ;
        RECT 1946.375 4707.385 1946.655 4707.665 ;
        RECT 1947.085 4707.385 1947.365 4707.665 ;
        RECT 1947.795 4707.385 1948.075 4707.665 ;
        RECT 1948.505 4707.385 1948.785 4707.665 ;
        RECT 1949.215 4707.385 1949.495 4707.665 ;
        RECT 1949.925 4707.385 1950.205 4707.665 ;
        RECT 1950.635 4707.385 1950.915 4707.665 ;
        RECT 1951.345 4707.385 1951.625 4707.665 ;
        RECT 1952.055 4707.385 1952.335 4707.665 ;
        RECT 1952.765 4707.385 1953.045 4707.665 ;
        RECT 1953.475 4707.385 1953.755 4707.665 ;
        RECT 1954.185 4707.385 1954.465 4707.665 ;
        RECT 1954.895 4707.385 1955.175 4707.665 ;
        RECT 1955.605 4707.385 1955.885 4707.665 ;
        RECT 1946.375 4706.675 1946.655 4706.955 ;
        RECT 1947.085 4706.675 1947.365 4706.955 ;
        RECT 1947.795 4706.675 1948.075 4706.955 ;
        RECT 1948.505 4706.675 1948.785 4706.955 ;
        RECT 1949.215 4706.675 1949.495 4706.955 ;
        RECT 1949.925 4706.675 1950.205 4706.955 ;
        RECT 1950.635 4706.675 1950.915 4706.955 ;
        RECT 1951.345 4706.675 1951.625 4706.955 ;
        RECT 1952.055 4706.675 1952.335 4706.955 ;
        RECT 1952.765 4706.675 1953.045 4706.955 ;
        RECT 1953.475 4706.675 1953.755 4706.955 ;
        RECT 1954.185 4706.675 1954.465 4706.955 ;
        RECT 1954.895 4706.675 1955.175 4706.955 ;
        RECT 1955.605 4706.675 1955.885 4706.955 ;
        RECT 1946.375 4705.965 1946.655 4706.245 ;
        RECT 1947.085 4705.965 1947.365 4706.245 ;
        RECT 1947.795 4705.965 1948.075 4706.245 ;
        RECT 1948.505 4705.965 1948.785 4706.245 ;
        RECT 1949.215 4705.965 1949.495 4706.245 ;
        RECT 1949.925 4705.965 1950.205 4706.245 ;
        RECT 1950.635 4705.965 1950.915 4706.245 ;
        RECT 1951.345 4705.965 1951.625 4706.245 ;
        RECT 1952.055 4705.965 1952.335 4706.245 ;
        RECT 1952.765 4705.965 1953.045 4706.245 ;
        RECT 1953.475 4705.965 1953.755 4706.245 ;
        RECT 1954.185 4705.965 1954.465 4706.245 ;
        RECT 1954.895 4705.965 1955.175 4706.245 ;
        RECT 1955.605 4705.965 1955.885 4706.245 ;
        RECT 1946.375 4705.255 1946.655 4705.535 ;
        RECT 1947.085 4705.255 1947.365 4705.535 ;
        RECT 1947.795 4705.255 1948.075 4705.535 ;
        RECT 1948.505 4705.255 1948.785 4705.535 ;
        RECT 1949.215 4705.255 1949.495 4705.535 ;
        RECT 1949.925 4705.255 1950.205 4705.535 ;
        RECT 1950.635 4705.255 1950.915 4705.535 ;
        RECT 1951.345 4705.255 1951.625 4705.535 ;
        RECT 1952.055 4705.255 1952.335 4705.535 ;
        RECT 1952.765 4705.255 1953.045 4705.535 ;
        RECT 1953.475 4705.255 1953.755 4705.535 ;
        RECT 1954.185 4705.255 1954.465 4705.535 ;
        RECT 1954.895 4705.255 1955.175 4705.535 ;
        RECT 1955.605 4705.255 1955.885 4705.535 ;
        RECT 1946.375 4704.545 1946.655 4704.825 ;
        RECT 1947.085 4704.545 1947.365 4704.825 ;
        RECT 1947.795 4704.545 1948.075 4704.825 ;
        RECT 1948.505 4704.545 1948.785 4704.825 ;
        RECT 1949.215 4704.545 1949.495 4704.825 ;
        RECT 1949.925 4704.545 1950.205 4704.825 ;
        RECT 1950.635 4704.545 1950.915 4704.825 ;
        RECT 1951.345 4704.545 1951.625 4704.825 ;
        RECT 1952.055 4704.545 1952.335 4704.825 ;
        RECT 1952.765 4704.545 1953.045 4704.825 ;
        RECT 1953.475 4704.545 1953.755 4704.825 ;
        RECT 1954.185 4704.545 1954.465 4704.825 ;
        RECT 1954.895 4704.545 1955.175 4704.825 ;
        RECT 1955.605 4704.545 1955.885 4704.825 ;
        RECT 1946.375 4703.835 1946.655 4704.115 ;
        RECT 1947.085 4703.835 1947.365 4704.115 ;
        RECT 1947.795 4703.835 1948.075 4704.115 ;
        RECT 1948.505 4703.835 1948.785 4704.115 ;
        RECT 1949.215 4703.835 1949.495 4704.115 ;
        RECT 1949.925 4703.835 1950.205 4704.115 ;
        RECT 1950.635 4703.835 1950.915 4704.115 ;
        RECT 1951.345 4703.835 1951.625 4704.115 ;
        RECT 1952.055 4703.835 1952.335 4704.115 ;
        RECT 1952.765 4703.835 1953.045 4704.115 ;
        RECT 1953.475 4703.835 1953.755 4704.115 ;
        RECT 1954.185 4703.835 1954.465 4704.115 ;
        RECT 1954.895 4703.835 1955.175 4704.115 ;
        RECT 1955.605 4703.835 1955.885 4704.115 ;
        RECT 1946.375 4703.125 1946.655 4703.405 ;
        RECT 1947.085 4703.125 1947.365 4703.405 ;
        RECT 1947.795 4703.125 1948.075 4703.405 ;
        RECT 1948.505 4703.125 1948.785 4703.405 ;
        RECT 1949.215 4703.125 1949.495 4703.405 ;
        RECT 1949.925 4703.125 1950.205 4703.405 ;
        RECT 1950.635 4703.125 1950.915 4703.405 ;
        RECT 1951.345 4703.125 1951.625 4703.405 ;
        RECT 1952.055 4703.125 1952.335 4703.405 ;
        RECT 1952.765 4703.125 1953.045 4703.405 ;
        RECT 1953.475 4703.125 1953.755 4703.405 ;
        RECT 1954.185 4703.125 1954.465 4703.405 ;
        RECT 1954.895 4703.125 1955.175 4703.405 ;
        RECT 1955.605 4703.125 1955.885 4703.405 ;
        RECT 1946.375 4702.415 1946.655 4702.695 ;
        RECT 1947.085 4702.415 1947.365 4702.695 ;
        RECT 1947.795 4702.415 1948.075 4702.695 ;
        RECT 1948.505 4702.415 1948.785 4702.695 ;
        RECT 1949.215 4702.415 1949.495 4702.695 ;
        RECT 1949.925 4702.415 1950.205 4702.695 ;
        RECT 1950.635 4702.415 1950.915 4702.695 ;
        RECT 1951.345 4702.415 1951.625 4702.695 ;
        RECT 1952.055 4702.415 1952.335 4702.695 ;
        RECT 1952.765 4702.415 1953.045 4702.695 ;
        RECT 1953.475 4702.415 1953.755 4702.695 ;
        RECT 1954.185 4702.415 1954.465 4702.695 ;
        RECT 1954.895 4702.415 1955.175 4702.695 ;
        RECT 1955.605 4702.415 1955.885 4702.695 ;
        RECT 1946.375 4701.705 1946.655 4701.985 ;
        RECT 1947.085 4701.705 1947.365 4701.985 ;
        RECT 1947.795 4701.705 1948.075 4701.985 ;
        RECT 1948.505 4701.705 1948.785 4701.985 ;
        RECT 1949.215 4701.705 1949.495 4701.985 ;
        RECT 1949.925 4701.705 1950.205 4701.985 ;
        RECT 1950.635 4701.705 1950.915 4701.985 ;
        RECT 1951.345 4701.705 1951.625 4701.985 ;
        RECT 1952.055 4701.705 1952.335 4701.985 ;
        RECT 1952.765 4701.705 1953.045 4701.985 ;
        RECT 1953.475 4701.705 1953.755 4701.985 ;
        RECT 1954.185 4701.705 1954.465 4701.985 ;
        RECT 1954.895 4701.705 1955.175 4701.985 ;
        RECT 1955.605 4701.705 1955.885 4701.985 ;
        RECT 1946.375 4700.995 1946.655 4701.275 ;
        RECT 1947.085 4700.995 1947.365 4701.275 ;
        RECT 1947.795 4700.995 1948.075 4701.275 ;
        RECT 1948.505 4700.995 1948.785 4701.275 ;
        RECT 1949.215 4700.995 1949.495 4701.275 ;
        RECT 1949.925 4700.995 1950.205 4701.275 ;
        RECT 1950.635 4700.995 1950.915 4701.275 ;
        RECT 1951.345 4700.995 1951.625 4701.275 ;
        RECT 1952.055 4700.995 1952.335 4701.275 ;
        RECT 1952.765 4700.995 1953.045 4701.275 ;
        RECT 1953.475 4700.995 1953.755 4701.275 ;
        RECT 1954.185 4700.995 1954.465 4701.275 ;
        RECT 1954.895 4700.995 1955.175 4701.275 ;
        RECT 1955.605 4700.995 1955.885 4701.275 ;
        RECT 1946.375 4700.285 1946.655 4700.565 ;
        RECT 1947.085 4700.285 1947.365 4700.565 ;
        RECT 1947.795 4700.285 1948.075 4700.565 ;
        RECT 1948.505 4700.285 1948.785 4700.565 ;
        RECT 1949.215 4700.285 1949.495 4700.565 ;
        RECT 1949.925 4700.285 1950.205 4700.565 ;
        RECT 1950.635 4700.285 1950.915 4700.565 ;
        RECT 1951.345 4700.285 1951.625 4700.565 ;
        RECT 1952.055 4700.285 1952.335 4700.565 ;
        RECT 1952.765 4700.285 1953.045 4700.565 ;
        RECT 1953.475 4700.285 1953.755 4700.565 ;
        RECT 1954.185 4700.285 1954.465 4700.565 ;
        RECT 1954.895 4700.285 1955.175 4700.565 ;
        RECT 1955.605 4700.285 1955.885 4700.565 ;
        RECT 1946.375 4699.575 1946.655 4699.855 ;
        RECT 1947.085 4699.575 1947.365 4699.855 ;
        RECT 1947.795 4699.575 1948.075 4699.855 ;
        RECT 1948.505 4699.575 1948.785 4699.855 ;
        RECT 1949.215 4699.575 1949.495 4699.855 ;
        RECT 1949.925 4699.575 1950.205 4699.855 ;
        RECT 1950.635 4699.575 1950.915 4699.855 ;
        RECT 1951.345 4699.575 1951.625 4699.855 ;
        RECT 1952.055 4699.575 1952.335 4699.855 ;
        RECT 1952.765 4699.575 1953.045 4699.855 ;
        RECT 1953.475 4699.575 1953.755 4699.855 ;
        RECT 1954.185 4699.575 1954.465 4699.855 ;
        RECT 1954.895 4699.575 1955.175 4699.855 ;
        RECT 1955.605 4699.575 1955.885 4699.855 ;
        RECT 1946.375 4698.865 1946.655 4699.145 ;
        RECT 1947.085 4698.865 1947.365 4699.145 ;
        RECT 1947.795 4698.865 1948.075 4699.145 ;
        RECT 1948.505 4698.865 1948.785 4699.145 ;
        RECT 1949.215 4698.865 1949.495 4699.145 ;
        RECT 1949.925 4698.865 1950.205 4699.145 ;
        RECT 1950.635 4698.865 1950.915 4699.145 ;
        RECT 1951.345 4698.865 1951.625 4699.145 ;
        RECT 1952.055 4698.865 1952.335 4699.145 ;
        RECT 1952.765 4698.865 1953.045 4699.145 ;
        RECT 1953.475 4698.865 1953.755 4699.145 ;
        RECT 1954.185 4698.865 1954.465 4699.145 ;
        RECT 1954.895 4698.865 1955.175 4699.145 ;
        RECT 1955.605 4698.865 1955.885 4699.145 ;
        RECT 1959.485 4708.095 1959.765 4708.375 ;
        RECT 1960.195 4708.095 1960.475 4708.375 ;
        RECT 1960.905 4708.095 1961.185 4708.375 ;
        RECT 1961.615 4708.095 1961.895 4708.375 ;
        RECT 1962.325 4708.095 1962.605 4708.375 ;
        RECT 1963.035 4708.095 1963.315 4708.375 ;
        RECT 1963.745 4708.095 1964.025 4708.375 ;
        RECT 1964.455 4708.095 1964.735 4708.375 ;
        RECT 1965.165 4708.095 1965.445 4708.375 ;
        RECT 1965.875 4708.095 1966.155 4708.375 ;
        RECT 1966.585 4708.095 1966.865 4708.375 ;
        RECT 1967.295 4708.095 1967.575 4708.375 ;
        RECT 1968.005 4708.095 1968.285 4708.375 ;
        RECT 1959.485 4707.385 1959.765 4707.665 ;
        RECT 1960.195 4707.385 1960.475 4707.665 ;
        RECT 1960.905 4707.385 1961.185 4707.665 ;
        RECT 1961.615 4707.385 1961.895 4707.665 ;
        RECT 1962.325 4707.385 1962.605 4707.665 ;
        RECT 1963.035 4707.385 1963.315 4707.665 ;
        RECT 1963.745 4707.385 1964.025 4707.665 ;
        RECT 1964.455 4707.385 1964.735 4707.665 ;
        RECT 1965.165 4707.385 1965.445 4707.665 ;
        RECT 1965.875 4707.385 1966.155 4707.665 ;
        RECT 1966.585 4707.385 1966.865 4707.665 ;
        RECT 1967.295 4707.385 1967.575 4707.665 ;
        RECT 1968.005 4707.385 1968.285 4707.665 ;
        RECT 1959.485 4706.675 1959.765 4706.955 ;
        RECT 1960.195 4706.675 1960.475 4706.955 ;
        RECT 1960.905 4706.675 1961.185 4706.955 ;
        RECT 1961.615 4706.675 1961.895 4706.955 ;
        RECT 1962.325 4706.675 1962.605 4706.955 ;
        RECT 1963.035 4706.675 1963.315 4706.955 ;
        RECT 1963.745 4706.675 1964.025 4706.955 ;
        RECT 1964.455 4706.675 1964.735 4706.955 ;
        RECT 1965.165 4706.675 1965.445 4706.955 ;
        RECT 1965.875 4706.675 1966.155 4706.955 ;
        RECT 1966.585 4706.675 1966.865 4706.955 ;
        RECT 1967.295 4706.675 1967.575 4706.955 ;
        RECT 1968.005 4706.675 1968.285 4706.955 ;
        RECT 1959.485 4705.965 1959.765 4706.245 ;
        RECT 1960.195 4705.965 1960.475 4706.245 ;
        RECT 1960.905 4705.965 1961.185 4706.245 ;
        RECT 1961.615 4705.965 1961.895 4706.245 ;
        RECT 1962.325 4705.965 1962.605 4706.245 ;
        RECT 1963.035 4705.965 1963.315 4706.245 ;
        RECT 1963.745 4705.965 1964.025 4706.245 ;
        RECT 1964.455 4705.965 1964.735 4706.245 ;
        RECT 1965.165 4705.965 1965.445 4706.245 ;
        RECT 1965.875 4705.965 1966.155 4706.245 ;
        RECT 1966.585 4705.965 1966.865 4706.245 ;
        RECT 1967.295 4705.965 1967.575 4706.245 ;
        RECT 1968.005 4705.965 1968.285 4706.245 ;
        RECT 1959.485 4705.255 1959.765 4705.535 ;
        RECT 1960.195 4705.255 1960.475 4705.535 ;
        RECT 1960.905 4705.255 1961.185 4705.535 ;
        RECT 1961.615 4705.255 1961.895 4705.535 ;
        RECT 1962.325 4705.255 1962.605 4705.535 ;
        RECT 1963.035 4705.255 1963.315 4705.535 ;
        RECT 1963.745 4705.255 1964.025 4705.535 ;
        RECT 1964.455 4705.255 1964.735 4705.535 ;
        RECT 1965.165 4705.255 1965.445 4705.535 ;
        RECT 1965.875 4705.255 1966.155 4705.535 ;
        RECT 1966.585 4705.255 1966.865 4705.535 ;
        RECT 1967.295 4705.255 1967.575 4705.535 ;
        RECT 1968.005 4705.255 1968.285 4705.535 ;
        RECT 1959.485 4704.545 1959.765 4704.825 ;
        RECT 1960.195 4704.545 1960.475 4704.825 ;
        RECT 1960.905 4704.545 1961.185 4704.825 ;
        RECT 1961.615 4704.545 1961.895 4704.825 ;
        RECT 1962.325 4704.545 1962.605 4704.825 ;
        RECT 1963.035 4704.545 1963.315 4704.825 ;
        RECT 1963.745 4704.545 1964.025 4704.825 ;
        RECT 1964.455 4704.545 1964.735 4704.825 ;
        RECT 1965.165 4704.545 1965.445 4704.825 ;
        RECT 1965.875 4704.545 1966.155 4704.825 ;
        RECT 1966.585 4704.545 1966.865 4704.825 ;
        RECT 1967.295 4704.545 1967.575 4704.825 ;
        RECT 1968.005 4704.545 1968.285 4704.825 ;
        RECT 1959.485 4703.835 1959.765 4704.115 ;
        RECT 1960.195 4703.835 1960.475 4704.115 ;
        RECT 1960.905 4703.835 1961.185 4704.115 ;
        RECT 1961.615 4703.835 1961.895 4704.115 ;
        RECT 1962.325 4703.835 1962.605 4704.115 ;
        RECT 1963.035 4703.835 1963.315 4704.115 ;
        RECT 1963.745 4703.835 1964.025 4704.115 ;
        RECT 1964.455 4703.835 1964.735 4704.115 ;
        RECT 1965.165 4703.835 1965.445 4704.115 ;
        RECT 1965.875 4703.835 1966.155 4704.115 ;
        RECT 1966.585 4703.835 1966.865 4704.115 ;
        RECT 1967.295 4703.835 1967.575 4704.115 ;
        RECT 1968.005 4703.835 1968.285 4704.115 ;
        RECT 1959.485 4703.125 1959.765 4703.405 ;
        RECT 1960.195 4703.125 1960.475 4703.405 ;
        RECT 1960.905 4703.125 1961.185 4703.405 ;
        RECT 1961.615 4703.125 1961.895 4703.405 ;
        RECT 1962.325 4703.125 1962.605 4703.405 ;
        RECT 1963.035 4703.125 1963.315 4703.405 ;
        RECT 1963.745 4703.125 1964.025 4703.405 ;
        RECT 1964.455 4703.125 1964.735 4703.405 ;
        RECT 1965.165 4703.125 1965.445 4703.405 ;
        RECT 1965.875 4703.125 1966.155 4703.405 ;
        RECT 1966.585 4703.125 1966.865 4703.405 ;
        RECT 1967.295 4703.125 1967.575 4703.405 ;
        RECT 1968.005 4703.125 1968.285 4703.405 ;
        RECT 1959.485 4702.415 1959.765 4702.695 ;
        RECT 1960.195 4702.415 1960.475 4702.695 ;
        RECT 1960.905 4702.415 1961.185 4702.695 ;
        RECT 1961.615 4702.415 1961.895 4702.695 ;
        RECT 1962.325 4702.415 1962.605 4702.695 ;
        RECT 1963.035 4702.415 1963.315 4702.695 ;
        RECT 1963.745 4702.415 1964.025 4702.695 ;
        RECT 1964.455 4702.415 1964.735 4702.695 ;
        RECT 1965.165 4702.415 1965.445 4702.695 ;
        RECT 1965.875 4702.415 1966.155 4702.695 ;
        RECT 1966.585 4702.415 1966.865 4702.695 ;
        RECT 1967.295 4702.415 1967.575 4702.695 ;
        RECT 1968.005 4702.415 1968.285 4702.695 ;
        RECT 1959.485 4701.705 1959.765 4701.985 ;
        RECT 1960.195 4701.705 1960.475 4701.985 ;
        RECT 1960.905 4701.705 1961.185 4701.985 ;
        RECT 1961.615 4701.705 1961.895 4701.985 ;
        RECT 1962.325 4701.705 1962.605 4701.985 ;
        RECT 1963.035 4701.705 1963.315 4701.985 ;
        RECT 1963.745 4701.705 1964.025 4701.985 ;
        RECT 1964.455 4701.705 1964.735 4701.985 ;
        RECT 1965.165 4701.705 1965.445 4701.985 ;
        RECT 1965.875 4701.705 1966.155 4701.985 ;
        RECT 1966.585 4701.705 1966.865 4701.985 ;
        RECT 1967.295 4701.705 1967.575 4701.985 ;
        RECT 1968.005 4701.705 1968.285 4701.985 ;
        RECT 1959.485 4700.995 1959.765 4701.275 ;
        RECT 1960.195 4700.995 1960.475 4701.275 ;
        RECT 1960.905 4700.995 1961.185 4701.275 ;
        RECT 1961.615 4700.995 1961.895 4701.275 ;
        RECT 1962.325 4700.995 1962.605 4701.275 ;
        RECT 1963.035 4700.995 1963.315 4701.275 ;
        RECT 1963.745 4700.995 1964.025 4701.275 ;
        RECT 1964.455 4700.995 1964.735 4701.275 ;
        RECT 1965.165 4700.995 1965.445 4701.275 ;
        RECT 1965.875 4700.995 1966.155 4701.275 ;
        RECT 1966.585 4700.995 1966.865 4701.275 ;
        RECT 1967.295 4700.995 1967.575 4701.275 ;
        RECT 1968.005 4700.995 1968.285 4701.275 ;
        RECT 1959.485 4700.285 1959.765 4700.565 ;
        RECT 1960.195 4700.285 1960.475 4700.565 ;
        RECT 1960.905 4700.285 1961.185 4700.565 ;
        RECT 1961.615 4700.285 1961.895 4700.565 ;
        RECT 1962.325 4700.285 1962.605 4700.565 ;
        RECT 1963.035 4700.285 1963.315 4700.565 ;
        RECT 1963.745 4700.285 1964.025 4700.565 ;
        RECT 1964.455 4700.285 1964.735 4700.565 ;
        RECT 1965.165 4700.285 1965.445 4700.565 ;
        RECT 1965.875 4700.285 1966.155 4700.565 ;
        RECT 1966.585 4700.285 1966.865 4700.565 ;
        RECT 1967.295 4700.285 1967.575 4700.565 ;
        RECT 1968.005 4700.285 1968.285 4700.565 ;
        RECT 1959.485 4699.575 1959.765 4699.855 ;
        RECT 1960.195 4699.575 1960.475 4699.855 ;
        RECT 1960.905 4699.575 1961.185 4699.855 ;
        RECT 1961.615 4699.575 1961.895 4699.855 ;
        RECT 1962.325 4699.575 1962.605 4699.855 ;
        RECT 1963.035 4699.575 1963.315 4699.855 ;
        RECT 1963.745 4699.575 1964.025 4699.855 ;
        RECT 1964.455 4699.575 1964.735 4699.855 ;
        RECT 1965.165 4699.575 1965.445 4699.855 ;
        RECT 1965.875 4699.575 1966.155 4699.855 ;
        RECT 1966.585 4699.575 1966.865 4699.855 ;
        RECT 1967.295 4699.575 1967.575 4699.855 ;
        RECT 1968.005 4699.575 1968.285 4699.855 ;
        RECT 1959.485 4698.865 1959.765 4699.145 ;
        RECT 1960.195 4698.865 1960.475 4699.145 ;
        RECT 1960.905 4698.865 1961.185 4699.145 ;
        RECT 1961.615 4698.865 1961.895 4699.145 ;
        RECT 1962.325 4698.865 1962.605 4699.145 ;
        RECT 1963.035 4698.865 1963.315 4699.145 ;
        RECT 1963.745 4698.865 1964.025 4699.145 ;
        RECT 1964.455 4698.865 1964.735 4699.145 ;
        RECT 1965.165 4698.865 1965.445 4699.145 ;
        RECT 1965.875 4698.865 1966.155 4699.145 ;
        RECT 1966.585 4698.865 1966.865 4699.145 ;
        RECT 1967.295 4698.865 1967.575 4699.145 ;
        RECT 1968.005 4698.865 1968.285 4699.145 ;
        RECT 2996.705 4708.095 2996.985 4708.375 ;
        RECT 2997.415 4708.095 2997.695 4708.375 ;
        RECT 2998.125 4708.095 2998.405 4708.375 ;
        RECT 2998.835 4708.095 2999.115 4708.375 ;
        RECT 2999.545 4708.095 2999.825 4708.375 ;
        RECT 3000.255 4708.095 3000.535 4708.375 ;
        RECT 3000.965 4708.095 3001.245 4708.375 ;
        RECT 3001.675 4708.095 3001.955 4708.375 ;
        RECT 3002.385 4708.095 3002.665 4708.375 ;
        RECT 3003.095 4708.095 3003.375 4708.375 ;
        RECT 3003.805 4708.095 3004.085 4708.375 ;
        RECT 3004.515 4708.095 3004.795 4708.375 ;
        RECT 3005.225 4708.095 3005.505 4708.375 ;
        RECT 2996.705 4707.385 2996.985 4707.665 ;
        RECT 2997.415 4707.385 2997.695 4707.665 ;
        RECT 2998.125 4707.385 2998.405 4707.665 ;
        RECT 2998.835 4707.385 2999.115 4707.665 ;
        RECT 2999.545 4707.385 2999.825 4707.665 ;
        RECT 3000.255 4707.385 3000.535 4707.665 ;
        RECT 3000.965 4707.385 3001.245 4707.665 ;
        RECT 3001.675 4707.385 3001.955 4707.665 ;
        RECT 3002.385 4707.385 3002.665 4707.665 ;
        RECT 3003.095 4707.385 3003.375 4707.665 ;
        RECT 3003.805 4707.385 3004.085 4707.665 ;
        RECT 3004.515 4707.385 3004.795 4707.665 ;
        RECT 3005.225 4707.385 3005.505 4707.665 ;
        RECT 2996.705 4706.675 2996.985 4706.955 ;
        RECT 2997.415 4706.675 2997.695 4706.955 ;
        RECT 2998.125 4706.675 2998.405 4706.955 ;
        RECT 2998.835 4706.675 2999.115 4706.955 ;
        RECT 2999.545 4706.675 2999.825 4706.955 ;
        RECT 3000.255 4706.675 3000.535 4706.955 ;
        RECT 3000.965 4706.675 3001.245 4706.955 ;
        RECT 3001.675 4706.675 3001.955 4706.955 ;
        RECT 3002.385 4706.675 3002.665 4706.955 ;
        RECT 3003.095 4706.675 3003.375 4706.955 ;
        RECT 3003.805 4706.675 3004.085 4706.955 ;
        RECT 3004.515 4706.675 3004.795 4706.955 ;
        RECT 3005.225 4706.675 3005.505 4706.955 ;
        RECT 2996.705 4705.965 2996.985 4706.245 ;
        RECT 2997.415 4705.965 2997.695 4706.245 ;
        RECT 2998.125 4705.965 2998.405 4706.245 ;
        RECT 2998.835 4705.965 2999.115 4706.245 ;
        RECT 2999.545 4705.965 2999.825 4706.245 ;
        RECT 3000.255 4705.965 3000.535 4706.245 ;
        RECT 3000.965 4705.965 3001.245 4706.245 ;
        RECT 3001.675 4705.965 3001.955 4706.245 ;
        RECT 3002.385 4705.965 3002.665 4706.245 ;
        RECT 3003.095 4705.965 3003.375 4706.245 ;
        RECT 3003.805 4705.965 3004.085 4706.245 ;
        RECT 3004.515 4705.965 3004.795 4706.245 ;
        RECT 3005.225 4705.965 3005.505 4706.245 ;
        RECT 2996.705 4705.255 2996.985 4705.535 ;
        RECT 2997.415 4705.255 2997.695 4705.535 ;
        RECT 2998.125 4705.255 2998.405 4705.535 ;
        RECT 2998.835 4705.255 2999.115 4705.535 ;
        RECT 2999.545 4705.255 2999.825 4705.535 ;
        RECT 3000.255 4705.255 3000.535 4705.535 ;
        RECT 3000.965 4705.255 3001.245 4705.535 ;
        RECT 3001.675 4705.255 3001.955 4705.535 ;
        RECT 3002.385 4705.255 3002.665 4705.535 ;
        RECT 3003.095 4705.255 3003.375 4705.535 ;
        RECT 3003.805 4705.255 3004.085 4705.535 ;
        RECT 3004.515 4705.255 3004.795 4705.535 ;
        RECT 3005.225 4705.255 3005.505 4705.535 ;
        RECT 2996.705 4704.545 2996.985 4704.825 ;
        RECT 2997.415 4704.545 2997.695 4704.825 ;
        RECT 2998.125 4704.545 2998.405 4704.825 ;
        RECT 2998.835 4704.545 2999.115 4704.825 ;
        RECT 2999.545 4704.545 2999.825 4704.825 ;
        RECT 3000.255 4704.545 3000.535 4704.825 ;
        RECT 3000.965 4704.545 3001.245 4704.825 ;
        RECT 3001.675 4704.545 3001.955 4704.825 ;
        RECT 3002.385 4704.545 3002.665 4704.825 ;
        RECT 3003.095 4704.545 3003.375 4704.825 ;
        RECT 3003.805 4704.545 3004.085 4704.825 ;
        RECT 3004.515 4704.545 3004.795 4704.825 ;
        RECT 3005.225 4704.545 3005.505 4704.825 ;
        RECT 2996.705 4703.835 2996.985 4704.115 ;
        RECT 2997.415 4703.835 2997.695 4704.115 ;
        RECT 2998.125 4703.835 2998.405 4704.115 ;
        RECT 2998.835 4703.835 2999.115 4704.115 ;
        RECT 2999.545 4703.835 2999.825 4704.115 ;
        RECT 3000.255 4703.835 3000.535 4704.115 ;
        RECT 3000.965 4703.835 3001.245 4704.115 ;
        RECT 3001.675 4703.835 3001.955 4704.115 ;
        RECT 3002.385 4703.835 3002.665 4704.115 ;
        RECT 3003.095 4703.835 3003.375 4704.115 ;
        RECT 3003.805 4703.835 3004.085 4704.115 ;
        RECT 3004.515 4703.835 3004.795 4704.115 ;
        RECT 3005.225 4703.835 3005.505 4704.115 ;
        RECT 2996.705 4703.125 2996.985 4703.405 ;
        RECT 2997.415 4703.125 2997.695 4703.405 ;
        RECT 2998.125 4703.125 2998.405 4703.405 ;
        RECT 2998.835 4703.125 2999.115 4703.405 ;
        RECT 2999.545 4703.125 2999.825 4703.405 ;
        RECT 3000.255 4703.125 3000.535 4703.405 ;
        RECT 3000.965 4703.125 3001.245 4703.405 ;
        RECT 3001.675 4703.125 3001.955 4703.405 ;
        RECT 3002.385 4703.125 3002.665 4703.405 ;
        RECT 3003.095 4703.125 3003.375 4703.405 ;
        RECT 3003.805 4703.125 3004.085 4703.405 ;
        RECT 3004.515 4703.125 3004.795 4703.405 ;
        RECT 3005.225 4703.125 3005.505 4703.405 ;
        RECT 2996.705 4702.415 2996.985 4702.695 ;
        RECT 2997.415 4702.415 2997.695 4702.695 ;
        RECT 2998.125 4702.415 2998.405 4702.695 ;
        RECT 2998.835 4702.415 2999.115 4702.695 ;
        RECT 2999.545 4702.415 2999.825 4702.695 ;
        RECT 3000.255 4702.415 3000.535 4702.695 ;
        RECT 3000.965 4702.415 3001.245 4702.695 ;
        RECT 3001.675 4702.415 3001.955 4702.695 ;
        RECT 3002.385 4702.415 3002.665 4702.695 ;
        RECT 3003.095 4702.415 3003.375 4702.695 ;
        RECT 3003.805 4702.415 3004.085 4702.695 ;
        RECT 3004.515 4702.415 3004.795 4702.695 ;
        RECT 3005.225 4702.415 3005.505 4702.695 ;
        RECT 2996.705 4701.705 2996.985 4701.985 ;
        RECT 2997.415 4701.705 2997.695 4701.985 ;
        RECT 2998.125 4701.705 2998.405 4701.985 ;
        RECT 2998.835 4701.705 2999.115 4701.985 ;
        RECT 2999.545 4701.705 2999.825 4701.985 ;
        RECT 3000.255 4701.705 3000.535 4701.985 ;
        RECT 3000.965 4701.705 3001.245 4701.985 ;
        RECT 3001.675 4701.705 3001.955 4701.985 ;
        RECT 3002.385 4701.705 3002.665 4701.985 ;
        RECT 3003.095 4701.705 3003.375 4701.985 ;
        RECT 3003.805 4701.705 3004.085 4701.985 ;
        RECT 3004.515 4701.705 3004.795 4701.985 ;
        RECT 3005.225 4701.705 3005.505 4701.985 ;
        RECT 2996.705 4700.995 2996.985 4701.275 ;
        RECT 2997.415 4700.995 2997.695 4701.275 ;
        RECT 2998.125 4700.995 2998.405 4701.275 ;
        RECT 2998.835 4700.995 2999.115 4701.275 ;
        RECT 2999.545 4700.995 2999.825 4701.275 ;
        RECT 3000.255 4700.995 3000.535 4701.275 ;
        RECT 3000.965 4700.995 3001.245 4701.275 ;
        RECT 3001.675 4700.995 3001.955 4701.275 ;
        RECT 3002.385 4700.995 3002.665 4701.275 ;
        RECT 3003.095 4700.995 3003.375 4701.275 ;
        RECT 3003.805 4700.995 3004.085 4701.275 ;
        RECT 3004.515 4700.995 3004.795 4701.275 ;
        RECT 3005.225 4700.995 3005.505 4701.275 ;
        RECT 2996.705 4700.285 2996.985 4700.565 ;
        RECT 2997.415 4700.285 2997.695 4700.565 ;
        RECT 2998.125 4700.285 2998.405 4700.565 ;
        RECT 2998.835 4700.285 2999.115 4700.565 ;
        RECT 2999.545 4700.285 2999.825 4700.565 ;
        RECT 3000.255 4700.285 3000.535 4700.565 ;
        RECT 3000.965 4700.285 3001.245 4700.565 ;
        RECT 3001.675 4700.285 3001.955 4700.565 ;
        RECT 3002.385 4700.285 3002.665 4700.565 ;
        RECT 3003.095 4700.285 3003.375 4700.565 ;
        RECT 3003.805 4700.285 3004.085 4700.565 ;
        RECT 3004.515 4700.285 3004.795 4700.565 ;
        RECT 3005.225 4700.285 3005.505 4700.565 ;
        RECT 2996.705 4699.575 2996.985 4699.855 ;
        RECT 2997.415 4699.575 2997.695 4699.855 ;
        RECT 2998.125 4699.575 2998.405 4699.855 ;
        RECT 2998.835 4699.575 2999.115 4699.855 ;
        RECT 2999.545 4699.575 2999.825 4699.855 ;
        RECT 3000.255 4699.575 3000.535 4699.855 ;
        RECT 3000.965 4699.575 3001.245 4699.855 ;
        RECT 3001.675 4699.575 3001.955 4699.855 ;
        RECT 3002.385 4699.575 3002.665 4699.855 ;
        RECT 3003.095 4699.575 3003.375 4699.855 ;
        RECT 3003.805 4699.575 3004.085 4699.855 ;
        RECT 3004.515 4699.575 3004.795 4699.855 ;
        RECT 3005.225 4699.575 3005.505 4699.855 ;
        RECT 2996.705 4698.865 2996.985 4699.145 ;
        RECT 2997.415 4698.865 2997.695 4699.145 ;
        RECT 2998.125 4698.865 2998.405 4699.145 ;
        RECT 2998.835 4698.865 2999.115 4699.145 ;
        RECT 2999.545 4698.865 2999.825 4699.145 ;
        RECT 3000.255 4698.865 3000.535 4699.145 ;
        RECT 3000.965 4698.865 3001.245 4699.145 ;
        RECT 3001.675 4698.865 3001.955 4699.145 ;
        RECT 3002.385 4698.865 3002.665 4699.145 ;
        RECT 3003.095 4698.865 3003.375 4699.145 ;
        RECT 3003.805 4698.865 3004.085 4699.145 ;
        RECT 3004.515 4698.865 3004.795 4699.145 ;
        RECT 3005.225 4698.865 3005.505 4699.145 ;
        RECT 3009.145 4708.095 3009.425 4708.375 ;
        RECT 3009.855 4708.095 3010.135 4708.375 ;
        RECT 3010.565 4708.095 3010.845 4708.375 ;
        RECT 3011.275 4708.095 3011.555 4708.375 ;
        RECT 3011.985 4708.095 3012.265 4708.375 ;
        RECT 3012.695 4708.095 3012.975 4708.375 ;
        RECT 3013.405 4708.095 3013.685 4708.375 ;
        RECT 3014.115 4708.095 3014.395 4708.375 ;
        RECT 3014.825 4708.095 3015.105 4708.375 ;
        RECT 3015.535 4708.095 3015.815 4708.375 ;
        RECT 3016.245 4708.095 3016.525 4708.375 ;
        RECT 3016.955 4708.095 3017.235 4708.375 ;
        RECT 3017.665 4708.095 3017.945 4708.375 ;
        RECT 3018.375 4708.095 3018.655 4708.375 ;
        RECT 3009.145 4707.385 3009.425 4707.665 ;
        RECT 3009.855 4707.385 3010.135 4707.665 ;
        RECT 3010.565 4707.385 3010.845 4707.665 ;
        RECT 3011.275 4707.385 3011.555 4707.665 ;
        RECT 3011.985 4707.385 3012.265 4707.665 ;
        RECT 3012.695 4707.385 3012.975 4707.665 ;
        RECT 3013.405 4707.385 3013.685 4707.665 ;
        RECT 3014.115 4707.385 3014.395 4707.665 ;
        RECT 3014.825 4707.385 3015.105 4707.665 ;
        RECT 3015.535 4707.385 3015.815 4707.665 ;
        RECT 3016.245 4707.385 3016.525 4707.665 ;
        RECT 3016.955 4707.385 3017.235 4707.665 ;
        RECT 3017.665 4707.385 3017.945 4707.665 ;
        RECT 3018.375 4707.385 3018.655 4707.665 ;
        RECT 3009.145 4706.675 3009.425 4706.955 ;
        RECT 3009.855 4706.675 3010.135 4706.955 ;
        RECT 3010.565 4706.675 3010.845 4706.955 ;
        RECT 3011.275 4706.675 3011.555 4706.955 ;
        RECT 3011.985 4706.675 3012.265 4706.955 ;
        RECT 3012.695 4706.675 3012.975 4706.955 ;
        RECT 3013.405 4706.675 3013.685 4706.955 ;
        RECT 3014.115 4706.675 3014.395 4706.955 ;
        RECT 3014.825 4706.675 3015.105 4706.955 ;
        RECT 3015.535 4706.675 3015.815 4706.955 ;
        RECT 3016.245 4706.675 3016.525 4706.955 ;
        RECT 3016.955 4706.675 3017.235 4706.955 ;
        RECT 3017.665 4706.675 3017.945 4706.955 ;
        RECT 3018.375 4706.675 3018.655 4706.955 ;
        RECT 3009.145 4705.965 3009.425 4706.245 ;
        RECT 3009.855 4705.965 3010.135 4706.245 ;
        RECT 3010.565 4705.965 3010.845 4706.245 ;
        RECT 3011.275 4705.965 3011.555 4706.245 ;
        RECT 3011.985 4705.965 3012.265 4706.245 ;
        RECT 3012.695 4705.965 3012.975 4706.245 ;
        RECT 3013.405 4705.965 3013.685 4706.245 ;
        RECT 3014.115 4705.965 3014.395 4706.245 ;
        RECT 3014.825 4705.965 3015.105 4706.245 ;
        RECT 3015.535 4705.965 3015.815 4706.245 ;
        RECT 3016.245 4705.965 3016.525 4706.245 ;
        RECT 3016.955 4705.965 3017.235 4706.245 ;
        RECT 3017.665 4705.965 3017.945 4706.245 ;
        RECT 3018.375 4705.965 3018.655 4706.245 ;
        RECT 3009.145 4705.255 3009.425 4705.535 ;
        RECT 3009.855 4705.255 3010.135 4705.535 ;
        RECT 3010.565 4705.255 3010.845 4705.535 ;
        RECT 3011.275 4705.255 3011.555 4705.535 ;
        RECT 3011.985 4705.255 3012.265 4705.535 ;
        RECT 3012.695 4705.255 3012.975 4705.535 ;
        RECT 3013.405 4705.255 3013.685 4705.535 ;
        RECT 3014.115 4705.255 3014.395 4705.535 ;
        RECT 3014.825 4705.255 3015.105 4705.535 ;
        RECT 3015.535 4705.255 3015.815 4705.535 ;
        RECT 3016.245 4705.255 3016.525 4705.535 ;
        RECT 3016.955 4705.255 3017.235 4705.535 ;
        RECT 3017.665 4705.255 3017.945 4705.535 ;
        RECT 3018.375 4705.255 3018.655 4705.535 ;
        RECT 3009.145 4704.545 3009.425 4704.825 ;
        RECT 3009.855 4704.545 3010.135 4704.825 ;
        RECT 3010.565 4704.545 3010.845 4704.825 ;
        RECT 3011.275 4704.545 3011.555 4704.825 ;
        RECT 3011.985 4704.545 3012.265 4704.825 ;
        RECT 3012.695 4704.545 3012.975 4704.825 ;
        RECT 3013.405 4704.545 3013.685 4704.825 ;
        RECT 3014.115 4704.545 3014.395 4704.825 ;
        RECT 3014.825 4704.545 3015.105 4704.825 ;
        RECT 3015.535 4704.545 3015.815 4704.825 ;
        RECT 3016.245 4704.545 3016.525 4704.825 ;
        RECT 3016.955 4704.545 3017.235 4704.825 ;
        RECT 3017.665 4704.545 3017.945 4704.825 ;
        RECT 3018.375 4704.545 3018.655 4704.825 ;
        RECT 3009.145 4703.835 3009.425 4704.115 ;
        RECT 3009.855 4703.835 3010.135 4704.115 ;
        RECT 3010.565 4703.835 3010.845 4704.115 ;
        RECT 3011.275 4703.835 3011.555 4704.115 ;
        RECT 3011.985 4703.835 3012.265 4704.115 ;
        RECT 3012.695 4703.835 3012.975 4704.115 ;
        RECT 3013.405 4703.835 3013.685 4704.115 ;
        RECT 3014.115 4703.835 3014.395 4704.115 ;
        RECT 3014.825 4703.835 3015.105 4704.115 ;
        RECT 3015.535 4703.835 3015.815 4704.115 ;
        RECT 3016.245 4703.835 3016.525 4704.115 ;
        RECT 3016.955 4703.835 3017.235 4704.115 ;
        RECT 3017.665 4703.835 3017.945 4704.115 ;
        RECT 3018.375 4703.835 3018.655 4704.115 ;
        RECT 3009.145 4703.125 3009.425 4703.405 ;
        RECT 3009.855 4703.125 3010.135 4703.405 ;
        RECT 3010.565 4703.125 3010.845 4703.405 ;
        RECT 3011.275 4703.125 3011.555 4703.405 ;
        RECT 3011.985 4703.125 3012.265 4703.405 ;
        RECT 3012.695 4703.125 3012.975 4703.405 ;
        RECT 3013.405 4703.125 3013.685 4703.405 ;
        RECT 3014.115 4703.125 3014.395 4703.405 ;
        RECT 3014.825 4703.125 3015.105 4703.405 ;
        RECT 3015.535 4703.125 3015.815 4703.405 ;
        RECT 3016.245 4703.125 3016.525 4703.405 ;
        RECT 3016.955 4703.125 3017.235 4703.405 ;
        RECT 3017.665 4703.125 3017.945 4703.405 ;
        RECT 3018.375 4703.125 3018.655 4703.405 ;
        RECT 3009.145 4702.415 3009.425 4702.695 ;
        RECT 3009.855 4702.415 3010.135 4702.695 ;
        RECT 3010.565 4702.415 3010.845 4702.695 ;
        RECT 3011.275 4702.415 3011.555 4702.695 ;
        RECT 3011.985 4702.415 3012.265 4702.695 ;
        RECT 3012.695 4702.415 3012.975 4702.695 ;
        RECT 3013.405 4702.415 3013.685 4702.695 ;
        RECT 3014.115 4702.415 3014.395 4702.695 ;
        RECT 3014.825 4702.415 3015.105 4702.695 ;
        RECT 3015.535 4702.415 3015.815 4702.695 ;
        RECT 3016.245 4702.415 3016.525 4702.695 ;
        RECT 3016.955 4702.415 3017.235 4702.695 ;
        RECT 3017.665 4702.415 3017.945 4702.695 ;
        RECT 3018.375 4702.415 3018.655 4702.695 ;
        RECT 3009.145 4701.705 3009.425 4701.985 ;
        RECT 3009.855 4701.705 3010.135 4701.985 ;
        RECT 3010.565 4701.705 3010.845 4701.985 ;
        RECT 3011.275 4701.705 3011.555 4701.985 ;
        RECT 3011.985 4701.705 3012.265 4701.985 ;
        RECT 3012.695 4701.705 3012.975 4701.985 ;
        RECT 3013.405 4701.705 3013.685 4701.985 ;
        RECT 3014.115 4701.705 3014.395 4701.985 ;
        RECT 3014.825 4701.705 3015.105 4701.985 ;
        RECT 3015.535 4701.705 3015.815 4701.985 ;
        RECT 3016.245 4701.705 3016.525 4701.985 ;
        RECT 3016.955 4701.705 3017.235 4701.985 ;
        RECT 3017.665 4701.705 3017.945 4701.985 ;
        RECT 3018.375 4701.705 3018.655 4701.985 ;
        RECT 3009.145 4700.995 3009.425 4701.275 ;
        RECT 3009.855 4700.995 3010.135 4701.275 ;
        RECT 3010.565 4700.995 3010.845 4701.275 ;
        RECT 3011.275 4700.995 3011.555 4701.275 ;
        RECT 3011.985 4700.995 3012.265 4701.275 ;
        RECT 3012.695 4700.995 3012.975 4701.275 ;
        RECT 3013.405 4700.995 3013.685 4701.275 ;
        RECT 3014.115 4700.995 3014.395 4701.275 ;
        RECT 3014.825 4700.995 3015.105 4701.275 ;
        RECT 3015.535 4700.995 3015.815 4701.275 ;
        RECT 3016.245 4700.995 3016.525 4701.275 ;
        RECT 3016.955 4700.995 3017.235 4701.275 ;
        RECT 3017.665 4700.995 3017.945 4701.275 ;
        RECT 3018.375 4700.995 3018.655 4701.275 ;
        RECT 3009.145 4700.285 3009.425 4700.565 ;
        RECT 3009.855 4700.285 3010.135 4700.565 ;
        RECT 3010.565 4700.285 3010.845 4700.565 ;
        RECT 3011.275 4700.285 3011.555 4700.565 ;
        RECT 3011.985 4700.285 3012.265 4700.565 ;
        RECT 3012.695 4700.285 3012.975 4700.565 ;
        RECT 3013.405 4700.285 3013.685 4700.565 ;
        RECT 3014.115 4700.285 3014.395 4700.565 ;
        RECT 3014.825 4700.285 3015.105 4700.565 ;
        RECT 3015.535 4700.285 3015.815 4700.565 ;
        RECT 3016.245 4700.285 3016.525 4700.565 ;
        RECT 3016.955 4700.285 3017.235 4700.565 ;
        RECT 3017.665 4700.285 3017.945 4700.565 ;
        RECT 3018.375 4700.285 3018.655 4700.565 ;
        RECT 3009.145 4699.575 3009.425 4699.855 ;
        RECT 3009.855 4699.575 3010.135 4699.855 ;
        RECT 3010.565 4699.575 3010.845 4699.855 ;
        RECT 3011.275 4699.575 3011.555 4699.855 ;
        RECT 3011.985 4699.575 3012.265 4699.855 ;
        RECT 3012.695 4699.575 3012.975 4699.855 ;
        RECT 3013.405 4699.575 3013.685 4699.855 ;
        RECT 3014.115 4699.575 3014.395 4699.855 ;
        RECT 3014.825 4699.575 3015.105 4699.855 ;
        RECT 3015.535 4699.575 3015.815 4699.855 ;
        RECT 3016.245 4699.575 3016.525 4699.855 ;
        RECT 3016.955 4699.575 3017.235 4699.855 ;
        RECT 3017.665 4699.575 3017.945 4699.855 ;
        RECT 3018.375 4699.575 3018.655 4699.855 ;
        RECT 3009.145 4698.865 3009.425 4699.145 ;
        RECT 3009.855 4698.865 3010.135 4699.145 ;
        RECT 3010.565 4698.865 3010.845 4699.145 ;
        RECT 3011.275 4698.865 3011.555 4699.145 ;
        RECT 3011.985 4698.865 3012.265 4699.145 ;
        RECT 3012.695 4698.865 3012.975 4699.145 ;
        RECT 3013.405 4698.865 3013.685 4699.145 ;
        RECT 3014.115 4698.865 3014.395 4699.145 ;
        RECT 3014.825 4698.865 3015.105 4699.145 ;
        RECT 3015.535 4698.865 3015.815 4699.145 ;
        RECT 3016.245 4698.865 3016.525 4699.145 ;
        RECT 3016.955 4698.865 3017.235 4699.145 ;
        RECT 3017.665 4698.865 3017.945 4699.145 ;
        RECT 3018.375 4698.865 3018.655 4699.145 ;
        RECT 3025.255 4708.095 3025.535 4708.375 ;
        RECT 3025.965 4708.095 3026.245 4708.375 ;
        RECT 3026.675 4708.095 3026.955 4708.375 ;
        RECT 3027.385 4708.095 3027.665 4708.375 ;
        RECT 3028.095 4708.095 3028.375 4708.375 ;
        RECT 3028.805 4708.095 3029.085 4708.375 ;
        RECT 3029.515 4708.095 3029.795 4708.375 ;
        RECT 3030.225 4708.095 3030.505 4708.375 ;
        RECT 3025.255 4707.385 3025.535 4707.665 ;
        RECT 3025.965 4707.385 3026.245 4707.665 ;
        RECT 3026.675 4707.385 3026.955 4707.665 ;
        RECT 3027.385 4707.385 3027.665 4707.665 ;
        RECT 3028.095 4707.385 3028.375 4707.665 ;
        RECT 3028.805 4707.385 3029.085 4707.665 ;
        RECT 3029.515 4707.385 3029.795 4707.665 ;
        RECT 3030.225 4707.385 3030.505 4707.665 ;
        RECT 3025.255 4706.675 3025.535 4706.955 ;
        RECT 3025.965 4706.675 3026.245 4706.955 ;
        RECT 3026.675 4706.675 3026.955 4706.955 ;
        RECT 3027.385 4706.675 3027.665 4706.955 ;
        RECT 3028.095 4706.675 3028.375 4706.955 ;
        RECT 3028.805 4706.675 3029.085 4706.955 ;
        RECT 3029.515 4706.675 3029.795 4706.955 ;
        RECT 3030.225 4706.675 3030.505 4706.955 ;
        RECT 3025.255 4705.965 3025.535 4706.245 ;
        RECT 3025.965 4705.965 3026.245 4706.245 ;
        RECT 3026.675 4705.965 3026.955 4706.245 ;
        RECT 3027.385 4705.965 3027.665 4706.245 ;
        RECT 3028.095 4705.965 3028.375 4706.245 ;
        RECT 3028.805 4705.965 3029.085 4706.245 ;
        RECT 3029.515 4705.965 3029.795 4706.245 ;
        RECT 3030.225 4705.965 3030.505 4706.245 ;
        RECT 3025.255 4705.255 3025.535 4705.535 ;
        RECT 3025.965 4705.255 3026.245 4705.535 ;
        RECT 3026.675 4705.255 3026.955 4705.535 ;
        RECT 3027.385 4705.255 3027.665 4705.535 ;
        RECT 3028.095 4705.255 3028.375 4705.535 ;
        RECT 3028.805 4705.255 3029.085 4705.535 ;
        RECT 3029.515 4705.255 3029.795 4705.535 ;
        RECT 3030.225 4705.255 3030.505 4705.535 ;
        RECT 3025.255 4704.545 3025.535 4704.825 ;
        RECT 3025.965 4704.545 3026.245 4704.825 ;
        RECT 3026.675 4704.545 3026.955 4704.825 ;
        RECT 3027.385 4704.545 3027.665 4704.825 ;
        RECT 3028.095 4704.545 3028.375 4704.825 ;
        RECT 3028.805 4704.545 3029.085 4704.825 ;
        RECT 3029.515 4704.545 3029.795 4704.825 ;
        RECT 3030.225 4704.545 3030.505 4704.825 ;
        RECT 3025.255 4703.835 3025.535 4704.115 ;
        RECT 3025.965 4703.835 3026.245 4704.115 ;
        RECT 3026.675 4703.835 3026.955 4704.115 ;
        RECT 3027.385 4703.835 3027.665 4704.115 ;
        RECT 3028.095 4703.835 3028.375 4704.115 ;
        RECT 3028.805 4703.835 3029.085 4704.115 ;
        RECT 3029.515 4703.835 3029.795 4704.115 ;
        RECT 3030.225 4703.835 3030.505 4704.115 ;
        RECT 3025.255 4703.125 3025.535 4703.405 ;
        RECT 3025.965 4703.125 3026.245 4703.405 ;
        RECT 3026.675 4703.125 3026.955 4703.405 ;
        RECT 3027.385 4703.125 3027.665 4703.405 ;
        RECT 3028.095 4703.125 3028.375 4703.405 ;
        RECT 3028.805 4703.125 3029.085 4703.405 ;
        RECT 3029.515 4703.125 3029.795 4703.405 ;
        RECT 3030.225 4703.125 3030.505 4703.405 ;
        RECT 3025.255 4702.415 3025.535 4702.695 ;
        RECT 3025.965 4702.415 3026.245 4702.695 ;
        RECT 3026.675 4702.415 3026.955 4702.695 ;
        RECT 3027.385 4702.415 3027.665 4702.695 ;
        RECT 3028.095 4702.415 3028.375 4702.695 ;
        RECT 3028.805 4702.415 3029.085 4702.695 ;
        RECT 3029.515 4702.415 3029.795 4702.695 ;
        RECT 3030.225 4702.415 3030.505 4702.695 ;
        RECT 3025.255 4701.705 3025.535 4701.985 ;
        RECT 3025.965 4701.705 3026.245 4701.985 ;
        RECT 3026.675 4701.705 3026.955 4701.985 ;
        RECT 3027.385 4701.705 3027.665 4701.985 ;
        RECT 3028.095 4701.705 3028.375 4701.985 ;
        RECT 3028.805 4701.705 3029.085 4701.985 ;
        RECT 3029.515 4701.705 3029.795 4701.985 ;
        RECT 3030.225 4701.705 3030.505 4701.985 ;
        RECT 3025.255 4700.995 3025.535 4701.275 ;
        RECT 3025.965 4700.995 3026.245 4701.275 ;
        RECT 3026.675 4700.995 3026.955 4701.275 ;
        RECT 3027.385 4700.995 3027.665 4701.275 ;
        RECT 3028.095 4700.995 3028.375 4701.275 ;
        RECT 3028.805 4700.995 3029.085 4701.275 ;
        RECT 3029.515 4700.995 3029.795 4701.275 ;
        RECT 3030.225 4700.995 3030.505 4701.275 ;
        RECT 3025.255 4700.285 3025.535 4700.565 ;
        RECT 3025.965 4700.285 3026.245 4700.565 ;
        RECT 3026.675 4700.285 3026.955 4700.565 ;
        RECT 3027.385 4700.285 3027.665 4700.565 ;
        RECT 3028.095 4700.285 3028.375 4700.565 ;
        RECT 3028.805 4700.285 3029.085 4700.565 ;
        RECT 3029.515 4700.285 3029.795 4700.565 ;
        RECT 3030.225 4700.285 3030.505 4700.565 ;
        RECT 3025.255 4699.575 3025.535 4699.855 ;
        RECT 3025.965 4699.575 3026.245 4699.855 ;
        RECT 3026.675 4699.575 3026.955 4699.855 ;
        RECT 3027.385 4699.575 3027.665 4699.855 ;
        RECT 3028.095 4699.575 3028.375 4699.855 ;
        RECT 3028.805 4699.575 3029.085 4699.855 ;
        RECT 3029.515 4699.575 3029.795 4699.855 ;
        RECT 3030.225 4699.575 3030.505 4699.855 ;
        RECT 3025.255 4698.865 3025.535 4699.145 ;
        RECT 3025.965 4698.865 3026.245 4699.145 ;
        RECT 3026.675 4698.865 3026.955 4699.145 ;
        RECT 3027.385 4698.865 3027.665 4699.145 ;
        RECT 3028.095 4698.865 3028.375 4699.145 ;
        RECT 3028.805 4698.865 3029.085 4699.145 ;
        RECT 3029.515 4698.865 3029.795 4699.145 ;
        RECT 3030.225 4698.865 3030.505 4699.145 ;
        RECT 3034.525 4708.095 3034.805 4708.375 ;
        RECT 3035.235 4708.095 3035.515 4708.375 ;
        RECT 3035.945 4708.095 3036.225 4708.375 ;
        RECT 3036.655 4708.095 3036.935 4708.375 ;
        RECT 3037.365 4708.095 3037.645 4708.375 ;
        RECT 3038.075 4708.095 3038.355 4708.375 ;
        RECT 3038.785 4708.095 3039.065 4708.375 ;
        RECT 3039.495 4708.095 3039.775 4708.375 ;
        RECT 3040.205 4708.095 3040.485 4708.375 ;
        RECT 3040.915 4708.095 3041.195 4708.375 ;
        RECT 3041.625 4708.095 3041.905 4708.375 ;
        RECT 3042.335 4708.095 3042.615 4708.375 ;
        RECT 3034.525 4707.385 3034.805 4707.665 ;
        RECT 3035.235 4707.385 3035.515 4707.665 ;
        RECT 3035.945 4707.385 3036.225 4707.665 ;
        RECT 3036.655 4707.385 3036.935 4707.665 ;
        RECT 3037.365 4707.385 3037.645 4707.665 ;
        RECT 3038.075 4707.385 3038.355 4707.665 ;
        RECT 3038.785 4707.385 3039.065 4707.665 ;
        RECT 3039.495 4707.385 3039.775 4707.665 ;
        RECT 3040.205 4707.385 3040.485 4707.665 ;
        RECT 3040.915 4707.385 3041.195 4707.665 ;
        RECT 3041.625 4707.385 3041.905 4707.665 ;
        RECT 3042.335 4707.385 3042.615 4707.665 ;
        RECT 3034.525 4706.675 3034.805 4706.955 ;
        RECT 3035.235 4706.675 3035.515 4706.955 ;
        RECT 3035.945 4706.675 3036.225 4706.955 ;
        RECT 3036.655 4706.675 3036.935 4706.955 ;
        RECT 3037.365 4706.675 3037.645 4706.955 ;
        RECT 3038.075 4706.675 3038.355 4706.955 ;
        RECT 3038.785 4706.675 3039.065 4706.955 ;
        RECT 3039.495 4706.675 3039.775 4706.955 ;
        RECT 3040.205 4706.675 3040.485 4706.955 ;
        RECT 3040.915 4706.675 3041.195 4706.955 ;
        RECT 3041.625 4706.675 3041.905 4706.955 ;
        RECT 3042.335 4706.675 3042.615 4706.955 ;
        RECT 3034.525 4705.965 3034.805 4706.245 ;
        RECT 3035.235 4705.965 3035.515 4706.245 ;
        RECT 3035.945 4705.965 3036.225 4706.245 ;
        RECT 3036.655 4705.965 3036.935 4706.245 ;
        RECT 3037.365 4705.965 3037.645 4706.245 ;
        RECT 3038.075 4705.965 3038.355 4706.245 ;
        RECT 3038.785 4705.965 3039.065 4706.245 ;
        RECT 3039.495 4705.965 3039.775 4706.245 ;
        RECT 3040.205 4705.965 3040.485 4706.245 ;
        RECT 3040.915 4705.965 3041.195 4706.245 ;
        RECT 3041.625 4705.965 3041.905 4706.245 ;
        RECT 3042.335 4705.965 3042.615 4706.245 ;
        RECT 3034.525 4705.255 3034.805 4705.535 ;
        RECT 3035.235 4705.255 3035.515 4705.535 ;
        RECT 3035.945 4705.255 3036.225 4705.535 ;
        RECT 3036.655 4705.255 3036.935 4705.535 ;
        RECT 3037.365 4705.255 3037.645 4705.535 ;
        RECT 3038.075 4705.255 3038.355 4705.535 ;
        RECT 3038.785 4705.255 3039.065 4705.535 ;
        RECT 3039.495 4705.255 3039.775 4705.535 ;
        RECT 3040.205 4705.255 3040.485 4705.535 ;
        RECT 3040.915 4705.255 3041.195 4705.535 ;
        RECT 3041.625 4705.255 3041.905 4705.535 ;
        RECT 3042.335 4705.255 3042.615 4705.535 ;
        RECT 3034.525 4704.545 3034.805 4704.825 ;
        RECT 3035.235 4704.545 3035.515 4704.825 ;
        RECT 3035.945 4704.545 3036.225 4704.825 ;
        RECT 3036.655 4704.545 3036.935 4704.825 ;
        RECT 3037.365 4704.545 3037.645 4704.825 ;
        RECT 3038.075 4704.545 3038.355 4704.825 ;
        RECT 3038.785 4704.545 3039.065 4704.825 ;
        RECT 3039.495 4704.545 3039.775 4704.825 ;
        RECT 3040.205 4704.545 3040.485 4704.825 ;
        RECT 3040.915 4704.545 3041.195 4704.825 ;
        RECT 3041.625 4704.545 3041.905 4704.825 ;
        RECT 3042.335 4704.545 3042.615 4704.825 ;
        RECT 3034.525 4703.835 3034.805 4704.115 ;
        RECT 3035.235 4703.835 3035.515 4704.115 ;
        RECT 3035.945 4703.835 3036.225 4704.115 ;
        RECT 3036.655 4703.835 3036.935 4704.115 ;
        RECT 3037.365 4703.835 3037.645 4704.115 ;
        RECT 3038.075 4703.835 3038.355 4704.115 ;
        RECT 3038.785 4703.835 3039.065 4704.115 ;
        RECT 3039.495 4703.835 3039.775 4704.115 ;
        RECT 3040.205 4703.835 3040.485 4704.115 ;
        RECT 3040.915 4703.835 3041.195 4704.115 ;
        RECT 3041.625 4703.835 3041.905 4704.115 ;
        RECT 3042.335 4703.835 3042.615 4704.115 ;
        RECT 3034.525 4703.125 3034.805 4703.405 ;
        RECT 3035.235 4703.125 3035.515 4703.405 ;
        RECT 3035.945 4703.125 3036.225 4703.405 ;
        RECT 3036.655 4703.125 3036.935 4703.405 ;
        RECT 3037.365 4703.125 3037.645 4703.405 ;
        RECT 3038.075 4703.125 3038.355 4703.405 ;
        RECT 3038.785 4703.125 3039.065 4703.405 ;
        RECT 3039.495 4703.125 3039.775 4703.405 ;
        RECT 3040.205 4703.125 3040.485 4703.405 ;
        RECT 3040.915 4703.125 3041.195 4703.405 ;
        RECT 3041.625 4703.125 3041.905 4703.405 ;
        RECT 3042.335 4703.125 3042.615 4703.405 ;
        RECT 3034.525 4702.415 3034.805 4702.695 ;
        RECT 3035.235 4702.415 3035.515 4702.695 ;
        RECT 3035.945 4702.415 3036.225 4702.695 ;
        RECT 3036.655 4702.415 3036.935 4702.695 ;
        RECT 3037.365 4702.415 3037.645 4702.695 ;
        RECT 3038.075 4702.415 3038.355 4702.695 ;
        RECT 3038.785 4702.415 3039.065 4702.695 ;
        RECT 3039.495 4702.415 3039.775 4702.695 ;
        RECT 3040.205 4702.415 3040.485 4702.695 ;
        RECT 3040.915 4702.415 3041.195 4702.695 ;
        RECT 3041.625 4702.415 3041.905 4702.695 ;
        RECT 3042.335 4702.415 3042.615 4702.695 ;
        RECT 3034.525 4701.705 3034.805 4701.985 ;
        RECT 3035.235 4701.705 3035.515 4701.985 ;
        RECT 3035.945 4701.705 3036.225 4701.985 ;
        RECT 3036.655 4701.705 3036.935 4701.985 ;
        RECT 3037.365 4701.705 3037.645 4701.985 ;
        RECT 3038.075 4701.705 3038.355 4701.985 ;
        RECT 3038.785 4701.705 3039.065 4701.985 ;
        RECT 3039.495 4701.705 3039.775 4701.985 ;
        RECT 3040.205 4701.705 3040.485 4701.985 ;
        RECT 3040.915 4701.705 3041.195 4701.985 ;
        RECT 3041.625 4701.705 3041.905 4701.985 ;
        RECT 3042.335 4701.705 3042.615 4701.985 ;
        RECT 3034.525 4700.995 3034.805 4701.275 ;
        RECT 3035.235 4700.995 3035.515 4701.275 ;
        RECT 3035.945 4700.995 3036.225 4701.275 ;
        RECT 3036.655 4700.995 3036.935 4701.275 ;
        RECT 3037.365 4700.995 3037.645 4701.275 ;
        RECT 3038.075 4700.995 3038.355 4701.275 ;
        RECT 3038.785 4700.995 3039.065 4701.275 ;
        RECT 3039.495 4700.995 3039.775 4701.275 ;
        RECT 3040.205 4700.995 3040.485 4701.275 ;
        RECT 3040.915 4700.995 3041.195 4701.275 ;
        RECT 3041.625 4700.995 3041.905 4701.275 ;
        RECT 3042.335 4700.995 3042.615 4701.275 ;
        RECT 3034.525 4700.285 3034.805 4700.565 ;
        RECT 3035.235 4700.285 3035.515 4700.565 ;
        RECT 3035.945 4700.285 3036.225 4700.565 ;
        RECT 3036.655 4700.285 3036.935 4700.565 ;
        RECT 3037.365 4700.285 3037.645 4700.565 ;
        RECT 3038.075 4700.285 3038.355 4700.565 ;
        RECT 3038.785 4700.285 3039.065 4700.565 ;
        RECT 3039.495 4700.285 3039.775 4700.565 ;
        RECT 3040.205 4700.285 3040.485 4700.565 ;
        RECT 3040.915 4700.285 3041.195 4700.565 ;
        RECT 3041.625 4700.285 3041.905 4700.565 ;
        RECT 3042.335 4700.285 3042.615 4700.565 ;
        RECT 3034.525 4699.575 3034.805 4699.855 ;
        RECT 3035.235 4699.575 3035.515 4699.855 ;
        RECT 3035.945 4699.575 3036.225 4699.855 ;
        RECT 3036.655 4699.575 3036.935 4699.855 ;
        RECT 3037.365 4699.575 3037.645 4699.855 ;
        RECT 3038.075 4699.575 3038.355 4699.855 ;
        RECT 3038.785 4699.575 3039.065 4699.855 ;
        RECT 3039.495 4699.575 3039.775 4699.855 ;
        RECT 3040.205 4699.575 3040.485 4699.855 ;
        RECT 3040.915 4699.575 3041.195 4699.855 ;
        RECT 3041.625 4699.575 3041.905 4699.855 ;
        RECT 3042.335 4699.575 3042.615 4699.855 ;
        RECT 3034.525 4698.865 3034.805 4699.145 ;
        RECT 3035.235 4698.865 3035.515 4699.145 ;
        RECT 3035.945 4698.865 3036.225 4699.145 ;
        RECT 3036.655 4698.865 3036.935 4699.145 ;
        RECT 3037.365 4698.865 3037.645 4699.145 ;
        RECT 3038.075 4698.865 3038.355 4699.145 ;
        RECT 3038.785 4698.865 3039.065 4699.145 ;
        RECT 3039.495 4698.865 3039.775 4699.145 ;
        RECT 3040.205 4698.865 3040.485 4699.145 ;
        RECT 3040.915 4698.865 3041.195 4699.145 ;
        RECT 3041.625 4698.865 3041.905 4699.145 ;
        RECT 3042.335 4698.865 3042.615 4699.145 ;
        RECT 3046.375 4708.095 3046.655 4708.375 ;
        RECT 3047.085 4708.095 3047.365 4708.375 ;
        RECT 3047.795 4708.095 3048.075 4708.375 ;
        RECT 3048.505 4708.095 3048.785 4708.375 ;
        RECT 3049.215 4708.095 3049.495 4708.375 ;
        RECT 3049.925 4708.095 3050.205 4708.375 ;
        RECT 3050.635 4708.095 3050.915 4708.375 ;
        RECT 3051.345 4708.095 3051.625 4708.375 ;
        RECT 3052.055 4708.095 3052.335 4708.375 ;
        RECT 3052.765 4708.095 3053.045 4708.375 ;
        RECT 3053.475 4708.095 3053.755 4708.375 ;
        RECT 3054.185 4708.095 3054.465 4708.375 ;
        RECT 3054.895 4708.095 3055.175 4708.375 ;
        RECT 3055.605 4708.095 3055.885 4708.375 ;
        RECT 3046.375 4707.385 3046.655 4707.665 ;
        RECT 3047.085 4707.385 3047.365 4707.665 ;
        RECT 3047.795 4707.385 3048.075 4707.665 ;
        RECT 3048.505 4707.385 3048.785 4707.665 ;
        RECT 3049.215 4707.385 3049.495 4707.665 ;
        RECT 3049.925 4707.385 3050.205 4707.665 ;
        RECT 3050.635 4707.385 3050.915 4707.665 ;
        RECT 3051.345 4707.385 3051.625 4707.665 ;
        RECT 3052.055 4707.385 3052.335 4707.665 ;
        RECT 3052.765 4707.385 3053.045 4707.665 ;
        RECT 3053.475 4707.385 3053.755 4707.665 ;
        RECT 3054.185 4707.385 3054.465 4707.665 ;
        RECT 3054.895 4707.385 3055.175 4707.665 ;
        RECT 3055.605 4707.385 3055.885 4707.665 ;
        RECT 3046.375 4706.675 3046.655 4706.955 ;
        RECT 3047.085 4706.675 3047.365 4706.955 ;
        RECT 3047.795 4706.675 3048.075 4706.955 ;
        RECT 3048.505 4706.675 3048.785 4706.955 ;
        RECT 3049.215 4706.675 3049.495 4706.955 ;
        RECT 3049.925 4706.675 3050.205 4706.955 ;
        RECT 3050.635 4706.675 3050.915 4706.955 ;
        RECT 3051.345 4706.675 3051.625 4706.955 ;
        RECT 3052.055 4706.675 3052.335 4706.955 ;
        RECT 3052.765 4706.675 3053.045 4706.955 ;
        RECT 3053.475 4706.675 3053.755 4706.955 ;
        RECT 3054.185 4706.675 3054.465 4706.955 ;
        RECT 3054.895 4706.675 3055.175 4706.955 ;
        RECT 3055.605 4706.675 3055.885 4706.955 ;
        RECT 3046.375 4705.965 3046.655 4706.245 ;
        RECT 3047.085 4705.965 3047.365 4706.245 ;
        RECT 3047.795 4705.965 3048.075 4706.245 ;
        RECT 3048.505 4705.965 3048.785 4706.245 ;
        RECT 3049.215 4705.965 3049.495 4706.245 ;
        RECT 3049.925 4705.965 3050.205 4706.245 ;
        RECT 3050.635 4705.965 3050.915 4706.245 ;
        RECT 3051.345 4705.965 3051.625 4706.245 ;
        RECT 3052.055 4705.965 3052.335 4706.245 ;
        RECT 3052.765 4705.965 3053.045 4706.245 ;
        RECT 3053.475 4705.965 3053.755 4706.245 ;
        RECT 3054.185 4705.965 3054.465 4706.245 ;
        RECT 3054.895 4705.965 3055.175 4706.245 ;
        RECT 3055.605 4705.965 3055.885 4706.245 ;
        RECT 3046.375 4705.255 3046.655 4705.535 ;
        RECT 3047.085 4705.255 3047.365 4705.535 ;
        RECT 3047.795 4705.255 3048.075 4705.535 ;
        RECT 3048.505 4705.255 3048.785 4705.535 ;
        RECT 3049.215 4705.255 3049.495 4705.535 ;
        RECT 3049.925 4705.255 3050.205 4705.535 ;
        RECT 3050.635 4705.255 3050.915 4705.535 ;
        RECT 3051.345 4705.255 3051.625 4705.535 ;
        RECT 3052.055 4705.255 3052.335 4705.535 ;
        RECT 3052.765 4705.255 3053.045 4705.535 ;
        RECT 3053.475 4705.255 3053.755 4705.535 ;
        RECT 3054.185 4705.255 3054.465 4705.535 ;
        RECT 3054.895 4705.255 3055.175 4705.535 ;
        RECT 3055.605 4705.255 3055.885 4705.535 ;
        RECT 3046.375 4704.545 3046.655 4704.825 ;
        RECT 3047.085 4704.545 3047.365 4704.825 ;
        RECT 3047.795 4704.545 3048.075 4704.825 ;
        RECT 3048.505 4704.545 3048.785 4704.825 ;
        RECT 3049.215 4704.545 3049.495 4704.825 ;
        RECT 3049.925 4704.545 3050.205 4704.825 ;
        RECT 3050.635 4704.545 3050.915 4704.825 ;
        RECT 3051.345 4704.545 3051.625 4704.825 ;
        RECT 3052.055 4704.545 3052.335 4704.825 ;
        RECT 3052.765 4704.545 3053.045 4704.825 ;
        RECT 3053.475 4704.545 3053.755 4704.825 ;
        RECT 3054.185 4704.545 3054.465 4704.825 ;
        RECT 3054.895 4704.545 3055.175 4704.825 ;
        RECT 3055.605 4704.545 3055.885 4704.825 ;
        RECT 3046.375 4703.835 3046.655 4704.115 ;
        RECT 3047.085 4703.835 3047.365 4704.115 ;
        RECT 3047.795 4703.835 3048.075 4704.115 ;
        RECT 3048.505 4703.835 3048.785 4704.115 ;
        RECT 3049.215 4703.835 3049.495 4704.115 ;
        RECT 3049.925 4703.835 3050.205 4704.115 ;
        RECT 3050.635 4703.835 3050.915 4704.115 ;
        RECT 3051.345 4703.835 3051.625 4704.115 ;
        RECT 3052.055 4703.835 3052.335 4704.115 ;
        RECT 3052.765 4703.835 3053.045 4704.115 ;
        RECT 3053.475 4703.835 3053.755 4704.115 ;
        RECT 3054.185 4703.835 3054.465 4704.115 ;
        RECT 3054.895 4703.835 3055.175 4704.115 ;
        RECT 3055.605 4703.835 3055.885 4704.115 ;
        RECT 3046.375 4703.125 3046.655 4703.405 ;
        RECT 3047.085 4703.125 3047.365 4703.405 ;
        RECT 3047.795 4703.125 3048.075 4703.405 ;
        RECT 3048.505 4703.125 3048.785 4703.405 ;
        RECT 3049.215 4703.125 3049.495 4703.405 ;
        RECT 3049.925 4703.125 3050.205 4703.405 ;
        RECT 3050.635 4703.125 3050.915 4703.405 ;
        RECT 3051.345 4703.125 3051.625 4703.405 ;
        RECT 3052.055 4703.125 3052.335 4703.405 ;
        RECT 3052.765 4703.125 3053.045 4703.405 ;
        RECT 3053.475 4703.125 3053.755 4703.405 ;
        RECT 3054.185 4703.125 3054.465 4703.405 ;
        RECT 3054.895 4703.125 3055.175 4703.405 ;
        RECT 3055.605 4703.125 3055.885 4703.405 ;
        RECT 3046.375 4702.415 3046.655 4702.695 ;
        RECT 3047.085 4702.415 3047.365 4702.695 ;
        RECT 3047.795 4702.415 3048.075 4702.695 ;
        RECT 3048.505 4702.415 3048.785 4702.695 ;
        RECT 3049.215 4702.415 3049.495 4702.695 ;
        RECT 3049.925 4702.415 3050.205 4702.695 ;
        RECT 3050.635 4702.415 3050.915 4702.695 ;
        RECT 3051.345 4702.415 3051.625 4702.695 ;
        RECT 3052.055 4702.415 3052.335 4702.695 ;
        RECT 3052.765 4702.415 3053.045 4702.695 ;
        RECT 3053.475 4702.415 3053.755 4702.695 ;
        RECT 3054.185 4702.415 3054.465 4702.695 ;
        RECT 3054.895 4702.415 3055.175 4702.695 ;
        RECT 3055.605 4702.415 3055.885 4702.695 ;
        RECT 3046.375 4701.705 3046.655 4701.985 ;
        RECT 3047.085 4701.705 3047.365 4701.985 ;
        RECT 3047.795 4701.705 3048.075 4701.985 ;
        RECT 3048.505 4701.705 3048.785 4701.985 ;
        RECT 3049.215 4701.705 3049.495 4701.985 ;
        RECT 3049.925 4701.705 3050.205 4701.985 ;
        RECT 3050.635 4701.705 3050.915 4701.985 ;
        RECT 3051.345 4701.705 3051.625 4701.985 ;
        RECT 3052.055 4701.705 3052.335 4701.985 ;
        RECT 3052.765 4701.705 3053.045 4701.985 ;
        RECT 3053.475 4701.705 3053.755 4701.985 ;
        RECT 3054.185 4701.705 3054.465 4701.985 ;
        RECT 3054.895 4701.705 3055.175 4701.985 ;
        RECT 3055.605 4701.705 3055.885 4701.985 ;
        RECT 3046.375 4700.995 3046.655 4701.275 ;
        RECT 3047.085 4700.995 3047.365 4701.275 ;
        RECT 3047.795 4700.995 3048.075 4701.275 ;
        RECT 3048.505 4700.995 3048.785 4701.275 ;
        RECT 3049.215 4700.995 3049.495 4701.275 ;
        RECT 3049.925 4700.995 3050.205 4701.275 ;
        RECT 3050.635 4700.995 3050.915 4701.275 ;
        RECT 3051.345 4700.995 3051.625 4701.275 ;
        RECT 3052.055 4700.995 3052.335 4701.275 ;
        RECT 3052.765 4700.995 3053.045 4701.275 ;
        RECT 3053.475 4700.995 3053.755 4701.275 ;
        RECT 3054.185 4700.995 3054.465 4701.275 ;
        RECT 3054.895 4700.995 3055.175 4701.275 ;
        RECT 3055.605 4700.995 3055.885 4701.275 ;
        RECT 3046.375 4700.285 3046.655 4700.565 ;
        RECT 3047.085 4700.285 3047.365 4700.565 ;
        RECT 3047.795 4700.285 3048.075 4700.565 ;
        RECT 3048.505 4700.285 3048.785 4700.565 ;
        RECT 3049.215 4700.285 3049.495 4700.565 ;
        RECT 3049.925 4700.285 3050.205 4700.565 ;
        RECT 3050.635 4700.285 3050.915 4700.565 ;
        RECT 3051.345 4700.285 3051.625 4700.565 ;
        RECT 3052.055 4700.285 3052.335 4700.565 ;
        RECT 3052.765 4700.285 3053.045 4700.565 ;
        RECT 3053.475 4700.285 3053.755 4700.565 ;
        RECT 3054.185 4700.285 3054.465 4700.565 ;
        RECT 3054.895 4700.285 3055.175 4700.565 ;
        RECT 3055.605 4700.285 3055.885 4700.565 ;
        RECT 3046.375 4699.575 3046.655 4699.855 ;
        RECT 3047.085 4699.575 3047.365 4699.855 ;
        RECT 3047.795 4699.575 3048.075 4699.855 ;
        RECT 3048.505 4699.575 3048.785 4699.855 ;
        RECT 3049.215 4699.575 3049.495 4699.855 ;
        RECT 3049.925 4699.575 3050.205 4699.855 ;
        RECT 3050.635 4699.575 3050.915 4699.855 ;
        RECT 3051.345 4699.575 3051.625 4699.855 ;
        RECT 3052.055 4699.575 3052.335 4699.855 ;
        RECT 3052.765 4699.575 3053.045 4699.855 ;
        RECT 3053.475 4699.575 3053.755 4699.855 ;
        RECT 3054.185 4699.575 3054.465 4699.855 ;
        RECT 3054.895 4699.575 3055.175 4699.855 ;
        RECT 3055.605 4699.575 3055.885 4699.855 ;
        RECT 3046.375 4698.865 3046.655 4699.145 ;
        RECT 3047.085 4698.865 3047.365 4699.145 ;
        RECT 3047.795 4698.865 3048.075 4699.145 ;
        RECT 3048.505 4698.865 3048.785 4699.145 ;
        RECT 3049.215 4698.865 3049.495 4699.145 ;
        RECT 3049.925 4698.865 3050.205 4699.145 ;
        RECT 3050.635 4698.865 3050.915 4699.145 ;
        RECT 3051.345 4698.865 3051.625 4699.145 ;
        RECT 3052.055 4698.865 3052.335 4699.145 ;
        RECT 3052.765 4698.865 3053.045 4699.145 ;
        RECT 3053.475 4698.865 3053.755 4699.145 ;
        RECT 3054.185 4698.865 3054.465 4699.145 ;
        RECT 3054.895 4698.865 3055.175 4699.145 ;
        RECT 3055.605 4698.865 3055.885 4699.145 ;
        RECT 3059.485 4708.095 3059.765 4708.375 ;
        RECT 3060.195 4708.095 3060.475 4708.375 ;
        RECT 3060.905 4708.095 3061.185 4708.375 ;
        RECT 3061.615 4708.095 3061.895 4708.375 ;
        RECT 3062.325 4708.095 3062.605 4708.375 ;
        RECT 3063.035 4708.095 3063.315 4708.375 ;
        RECT 3063.745 4708.095 3064.025 4708.375 ;
        RECT 3064.455 4708.095 3064.735 4708.375 ;
        RECT 3065.165 4708.095 3065.445 4708.375 ;
        RECT 3065.875 4708.095 3066.155 4708.375 ;
        RECT 3066.585 4708.095 3066.865 4708.375 ;
        RECT 3067.295 4708.095 3067.575 4708.375 ;
        RECT 3068.005 4708.095 3068.285 4708.375 ;
        RECT 3059.485 4707.385 3059.765 4707.665 ;
        RECT 3060.195 4707.385 3060.475 4707.665 ;
        RECT 3060.905 4707.385 3061.185 4707.665 ;
        RECT 3061.615 4707.385 3061.895 4707.665 ;
        RECT 3062.325 4707.385 3062.605 4707.665 ;
        RECT 3063.035 4707.385 3063.315 4707.665 ;
        RECT 3063.745 4707.385 3064.025 4707.665 ;
        RECT 3064.455 4707.385 3064.735 4707.665 ;
        RECT 3065.165 4707.385 3065.445 4707.665 ;
        RECT 3065.875 4707.385 3066.155 4707.665 ;
        RECT 3066.585 4707.385 3066.865 4707.665 ;
        RECT 3067.295 4707.385 3067.575 4707.665 ;
        RECT 3068.005 4707.385 3068.285 4707.665 ;
        RECT 3059.485 4706.675 3059.765 4706.955 ;
        RECT 3060.195 4706.675 3060.475 4706.955 ;
        RECT 3060.905 4706.675 3061.185 4706.955 ;
        RECT 3061.615 4706.675 3061.895 4706.955 ;
        RECT 3062.325 4706.675 3062.605 4706.955 ;
        RECT 3063.035 4706.675 3063.315 4706.955 ;
        RECT 3063.745 4706.675 3064.025 4706.955 ;
        RECT 3064.455 4706.675 3064.735 4706.955 ;
        RECT 3065.165 4706.675 3065.445 4706.955 ;
        RECT 3065.875 4706.675 3066.155 4706.955 ;
        RECT 3066.585 4706.675 3066.865 4706.955 ;
        RECT 3067.295 4706.675 3067.575 4706.955 ;
        RECT 3068.005 4706.675 3068.285 4706.955 ;
        RECT 3059.485 4705.965 3059.765 4706.245 ;
        RECT 3060.195 4705.965 3060.475 4706.245 ;
        RECT 3060.905 4705.965 3061.185 4706.245 ;
        RECT 3061.615 4705.965 3061.895 4706.245 ;
        RECT 3062.325 4705.965 3062.605 4706.245 ;
        RECT 3063.035 4705.965 3063.315 4706.245 ;
        RECT 3063.745 4705.965 3064.025 4706.245 ;
        RECT 3064.455 4705.965 3064.735 4706.245 ;
        RECT 3065.165 4705.965 3065.445 4706.245 ;
        RECT 3065.875 4705.965 3066.155 4706.245 ;
        RECT 3066.585 4705.965 3066.865 4706.245 ;
        RECT 3067.295 4705.965 3067.575 4706.245 ;
        RECT 3068.005 4705.965 3068.285 4706.245 ;
        RECT 3059.485 4705.255 3059.765 4705.535 ;
        RECT 3060.195 4705.255 3060.475 4705.535 ;
        RECT 3060.905 4705.255 3061.185 4705.535 ;
        RECT 3061.615 4705.255 3061.895 4705.535 ;
        RECT 3062.325 4705.255 3062.605 4705.535 ;
        RECT 3063.035 4705.255 3063.315 4705.535 ;
        RECT 3063.745 4705.255 3064.025 4705.535 ;
        RECT 3064.455 4705.255 3064.735 4705.535 ;
        RECT 3065.165 4705.255 3065.445 4705.535 ;
        RECT 3065.875 4705.255 3066.155 4705.535 ;
        RECT 3066.585 4705.255 3066.865 4705.535 ;
        RECT 3067.295 4705.255 3067.575 4705.535 ;
        RECT 3068.005 4705.255 3068.285 4705.535 ;
        RECT 3059.485 4704.545 3059.765 4704.825 ;
        RECT 3060.195 4704.545 3060.475 4704.825 ;
        RECT 3060.905 4704.545 3061.185 4704.825 ;
        RECT 3061.615 4704.545 3061.895 4704.825 ;
        RECT 3062.325 4704.545 3062.605 4704.825 ;
        RECT 3063.035 4704.545 3063.315 4704.825 ;
        RECT 3063.745 4704.545 3064.025 4704.825 ;
        RECT 3064.455 4704.545 3064.735 4704.825 ;
        RECT 3065.165 4704.545 3065.445 4704.825 ;
        RECT 3065.875 4704.545 3066.155 4704.825 ;
        RECT 3066.585 4704.545 3066.865 4704.825 ;
        RECT 3067.295 4704.545 3067.575 4704.825 ;
        RECT 3068.005 4704.545 3068.285 4704.825 ;
        RECT 3059.485 4703.835 3059.765 4704.115 ;
        RECT 3060.195 4703.835 3060.475 4704.115 ;
        RECT 3060.905 4703.835 3061.185 4704.115 ;
        RECT 3061.615 4703.835 3061.895 4704.115 ;
        RECT 3062.325 4703.835 3062.605 4704.115 ;
        RECT 3063.035 4703.835 3063.315 4704.115 ;
        RECT 3063.745 4703.835 3064.025 4704.115 ;
        RECT 3064.455 4703.835 3064.735 4704.115 ;
        RECT 3065.165 4703.835 3065.445 4704.115 ;
        RECT 3065.875 4703.835 3066.155 4704.115 ;
        RECT 3066.585 4703.835 3066.865 4704.115 ;
        RECT 3067.295 4703.835 3067.575 4704.115 ;
        RECT 3068.005 4703.835 3068.285 4704.115 ;
        RECT 3059.485 4703.125 3059.765 4703.405 ;
        RECT 3060.195 4703.125 3060.475 4703.405 ;
        RECT 3060.905 4703.125 3061.185 4703.405 ;
        RECT 3061.615 4703.125 3061.895 4703.405 ;
        RECT 3062.325 4703.125 3062.605 4703.405 ;
        RECT 3063.035 4703.125 3063.315 4703.405 ;
        RECT 3063.745 4703.125 3064.025 4703.405 ;
        RECT 3064.455 4703.125 3064.735 4703.405 ;
        RECT 3065.165 4703.125 3065.445 4703.405 ;
        RECT 3065.875 4703.125 3066.155 4703.405 ;
        RECT 3066.585 4703.125 3066.865 4703.405 ;
        RECT 3067.295 4703.125 3067.575 4703.405 ;
        RECT 3068.005 4703.125 3068.285 4703.405 ;
        RECT 3059.485 4702.415 3059.765 4702.695 ;
        RECT 3060.195 4702.415 3060.475 4702.695 ;
        RECT 3060.905 4702.415 3061.185 4702.695 ;
        RECT 3061.615 4702.415 3061.895 4702.695 ;
        RECT 3062.325 4702.415 3062.605 4702.695 ;
        RECT 3063.035 4702.415 3063.315 4702.695 ;
        RECT 3063.745 4702.415 3064.025 4702.695 ;
        RECT 3064.455 4702.415 3064.735 4702.695 ;
        RECT 3065.165 4702.415 3065.445 4702.695 ;
        RECT 3065.875 4702.415 3066.155 4702.695 ;
        RECT 3066.585 4702.415 3066.865 4702.695 ;
        RECT 3067.295 4702.415 3067.575 4702.695 ;
        RECT 3068.005 4702.415 3068.285 4702.695 ;
        RECT 3059.485 4701.705 3059.765 4701.985 ;
        RECT 3060.195 4701.705 3060.475 4701.985 ;
        RECT 3060.905 4701.705 3061.185 4701.985 ;
        RECT 3061.615 4701.705 3061.895 4701.985 ;
        RECT 3062.325 4701.705 3062.605 4701.985 ;
        RECT 3063.035 4701.705 3063.315 4701.985 ;
        RECT 3063.745 4701.705 3064.025 4701.985 ;
        RECT 3064.455 4701.705 3064.735 4701.985 ;
        RECT 3065.165 4701.705 3065.445 4701.985 ;
        RECT 3065.875 4701.705 3066.155 4701.985 ;
        RECT 3066.585 4701.705 3066.865 4701.985 ;
        RECT 3067.295 4701.705 3067.575 4701.985 ;
        RECT 3068.005 4701.705 3068.285 4701.985 ;
        RECT 3059.485 4700.995 3059.765 4701.275 ;
        RECT 3060.195 4700.995 3060.475 4701.275 ;
        RECT 3060.905 4700.995 3061.185 4701.275 ;
        RECT 3061.615 4700.995 3061.895 4701.275 ;
        RECT 3062.325 4700.995 3062.605 4701.275 ;
        RECT 3063.035 4700.995 3063.315 4701.275 ;
        RECT 3063.745 4700.995 3064.025 4701.275 ;
        RECT 3064.455 4700.995 3064.735 4701.275 ;
        RECT 3065.165 4700.995 3065.445 4701.275 ;
        RECT 3065.875 4700.995 3066.155 4701.275 ;
        RECT 3066.585 4700.995 3066.865 4701.275 ;
        RECT 3067.295 4700.995 3067.575 4701.275 ;
        RECT 3068.005 4700.995 3068.285 4701.275 ;
        RECT 3059.485 4700.285 3059.765 4700.565 ;
        RECT 3060.195 4700.285 3060.475 4700.565 ;
        RECT 3060.905 4700.285 3061.185 4700.565 ;
        RECT 3061.615 4700.285 3061.895 4700.565 ;
        RECT 3062.325 4700.285 3062.605 4700.565 ;
        RECT 3063.035 4700.285 3063.315 4700.565 ;
        RECT 3063.745 4700.285 3064.025 4700.565 ;
        RECT 3064.455 4700.285 3064.735 4700.565 ;
        RECT 3065.165 4700.285 3065.445 4700.565 ;
        RECT 3065.875 4700.285 3066.155 4700.565 ;
        RECT 3066.585 4700.285 3066.865 4700.565 ;
        RECT 3067.295 4700.285 3067.575 4700.565 ;
        RECT 3068.005 4700.285 3068.285 4700.565 ;
        RECT 3059.485 4699.575 3059.765 4699.855 ;
        RECT 3060.195 4699.575 3060.475 4699.855 ;
        RECT 3060.905 4699.575 3061.185 4699.855 ;
        RECT 3061.615 4699.575 3061.895 4699.855 ;
        RECT 3062.325 4699.575 3062.605 4699.855 ;
        RECT 3063.035 4699.575 3063.315 4699.855 ;
        RECT 3063.745 4699.575 3064.025 4699.855 ;
        RECT 3064.455 4699.575 3064.735 4699.855 ;
        RECT 3065.165 4699.575 3065.445 4699.855 ;
        RECT 3065.875 4699.575 3066.155 4699.855 ;
        RECT 3066.585 4699.575 3066.865 4699.855 ;
        RECT 3067.295 4699.575 3067.575 4699.855 ;
        RECT 3068.005 4699.575 3068.285 4699.855 ;
        RECT 3059.485 4698.865 3059.765 4699.145 ;
        RECT 3060.195 4698.865 3060.475 4699.145 ;
        RECT 3060.905 4698.865 3061.185 4699.145 ;
        RECT 3061.615 4698.865 3061.895 4699.145 ;
        RECT 3062.325 4698.865 3062.605 4699.145 ;
        RECT 3063.035 4698.865 3063.315 4699.145 ;
        RECT 3063.745 4698.865 3064.025 4699.145 ;
        RECT 3064.455 4698.865 3064.735 4699.145 ;
        RECT 3065.165 4698.865 3065.445 4699.145 ;
        RECT 3065.875 4698.865 3066.155 4699.145 ;
        RECT 3066.585 4698.865 3066.865 4699.145 ;
        RECT 3067.295 4698.865 3067.575 4699.145 ;
        RECT 3068.005 4698.865 3068.285 4699.145 ;
        RECT 3276.715 379.895 3276.995 380.175 ;
        RECT 3277.425 379.895 3277.705 380.175 ;
        RECT 3278.135 379.895 3278.415 380.175 ;
        RECT 3278.845 379.895 3279.125 380.175 ;
        RECT 3279.555 379.895 3279.835 380.175 ;
        RECT 3280.265 379.895 3280.545 380.175 ;
        RECT 3280.975 379.895 3281.255 380.175 ;
        RECT 3281.685 379.895 3281.965 380.175 ;
        RECT 3276.715 379.185 3276.995 379.465 ;
        RECT 3277.425 379.185 3277.705 379.465 ;
        RECT 3278.135 379.185 3278.415 379.465 ;
        RECT 3278.845 379.185 3279.125 379.465 ;
        RECT 3279.555 379.185 3279.835 379.465 ;
        RECT 3280.265 379.185 3280.545 379.465 ;
        RECT 3280.975 379.185 3281.255 379.465 ;
        RECT 3281.685 379.185 3281.965 379.465 ;
        RECT 3276.715 378.475 3276.995 378.755 ;
        RECT 3277.425 378.475 3277.705 378.755 ;
        RECT 3278.135 378.475 3278.415 378.755 ;
        RECT 3278.845 378.475 3279.125 378.755 ;
        RECT 3279.555 378.475 3279.835 378.755 ;
        RECT 3280.265 378.475 3280.545 378.755 ;
        RECT 3280.975 378.475 3281.255 378.755 ;
        RECT 3281.685 378.475 3281.965 378.755 ;
        RECT 3276.715 377.765 3276.995 378.045 ;
        RECT 3277.425 377.765 3277.705 378.045 ;
        RECT 3278.135 377.765 3278.415 378.045 ;
        RECT 3278.845 377.765 3279.125 378.045 ;
        RECT 3279.555 377.765 3279.835 378.045 ;
        RECT 3280.265 377.765 3280.545 378.045 ;
        RECT 3280.975 377.765 3281.255 378.045 ;
        RECT 3281.685 377.765 3281.965 378.045 ;
        RECT 3276.715 377.055 3276.995 377.335 ;
        RECT 3277.425 377.055 3277.705 377.335 ;
        RECT 3278.135 377.055 3278.415 377.335 ;
        RECT 3278.845 377.055 3279.125 377.335 ;
        RECT 3279.555 377.055 3279.835 377.335 ;
        RECT 3280.265 377.055 3280.545 377.335 ;
        RECT 3280.975 377.055 3281.255 377.335 ;
        RECT 3281.685 377.055 3281.965 377.335 ;
        RECT 3276.715 376.345 3276.995 376.625 ;
        RECT 3277.425 376.345 3277.705 376.625 ;
        RECT 3278.135 376.345 3278.415 376.625 ;
        RECT 3278.845 376.345 3279.125 376.625 ;
        RECT 3279.555 376.345 3279.835 376.625 ;
        RECT 3280.265 376.345 3280.545 376.625 ;
        RECT 3280.975 376.345 3281.255 376.625 ;
        RECT 3281.685 376.345 3281.965 376.625 ;
        RECT 3276.715 375.635 3276.995 375.915 ;
        RECT 3277.425 375.635 3277.705 375.915 ;
        RECT 3278.135 375.635 3278.415 375.915 ;
        RECT 3278.845 375.635 3279.125 375.915 ;
        RECT 3279.555 375.635 3279.835 375.915 ;
        RECT 3280.265 375.635 3280.545 375.915 ;
        RECT 3280.975 375.635 3281.255 375.915 ;
        RECT 3281.685 375.635 3281.965 375.915 ;
        RECT 3276.715 374.925 3276.995 375.205 ;
        RECT 3277.425 374.925 3277.705 375.205 ;
        RECT 3278.135 374.925 3278.415 375.205 ;
        RECT 3278.845 374.925 3279.125 375.205 ;
        RECT 3279.555 374.925 3279.835 375.205 ;
        RECT 3280.265 374.925 3280.545 375.205 ;
        RECT 3280.975 374.925 3281.255 375.205 ;
        RECT 3281.685 374.925 3281.965 375.205 ;
        RECT 3276.715 374.215 3276.995 374.495 ;
        RECT 3277.425 374.215 3277.705 374.495 ;
        RECT 3278.135 374.215 3278.415 374.495 ;
        RECT 3278.845 374.215 3279.125 374.495 ;
        RECT 3279.555 374.215 3279.835 374.495 ;
        RECT 3280.265 374.215 3280.545 374.495 ;
        RECT 3280.975 374.215 3281.255 374.495 ;
        RECT 3281.685 374.215 3281.965 374.495 ;
        RECT 3276.715 373.505 3276.995 373.785 ;
        RECT 3277.425 373.505 3277.705 373.785 ;
        RECT 3278.135 373.505 3278.415 373.785 ;
        RECT 3278.845 373.505 3279.125 373.785 ;
        RECT 3279.555 373.505 3279.835 373.785 ;
        RECT 3280.265 373.505 3280.545 373.785 ;
        RECT 3280.975 373.505 3281.255 373.785 ;
        RECT 3281.685 373.505 3281.965 373.785 ;
        RECT 3276.715 372.795 3276.995 373.075 ;
        RECT 3277.425 372.795 3277.705 373.075 ;
        RECT 3278.135 372.795 3278.415 373.075 ;
        RECT 3278.845 372.795 3279.125 373.075 ;
        RECT 3279.555 372.795 3279.835 373.075 ;
        RECT 3280.265 372.795 3280.545 373.075 ;
        RECT 3280.975 372.795 3281.255 373.075 ;
        RECT 3281.685 372.795 3281.965 373.075 ;
        RECT 3289.115 379.895 3289.395 380.175 ;
        RECT 3289.825 379.895 3290.105 380.175 ;
        RECT 3290.535 379.895 3290.815 380.175 ;
        RECT 3291.245 379.895 3291.525 380.175 ;
        RECT 3291.955 379.895 3292.235 380.175 ;
        RECT 3292.665 379.895 3292.945 380.175 ;
        RECT 3293.375 379.895 3293.655 380.175 ;
        RECT 3294.085 379.895 3294.365 380.175 ;
        RECT 3294.795 379.895 3295.075 380.175 ;
        RECT 3295.505 379.895 3295.785 380.175 ;
        RECT 3296.215 379.895 3296.495 380.175 ;
        RECT 3296.925 379.895 3297.205 380.175 ;
        RECT 3297.635 379.895 3297.915 380.175 ;
        RECT 3298.345 379.895 3298.625 380.175 ;
        RECT 3289.115 379.185 3289.395 379.465 ;
        RECT 3289.825 379.185 3290.105 379.465 ;
        RECT 3290.535 379.185 3290.815 379.465 ;
        RECT 3291.245 379.185 3291.525 379.465 ;
        RECT 3291.955 379.185 3292.235 379.465 ;
        RECT 3292.665 379.185 3292.945 379.465 ;
        RECT 3293.375 379.185 3293.655 379.465 ;
        RECT 3294.085 379.185 3294.365 379.465 ;
        RECT 3294.795 379.185 3295.075 379.465 ;
        RECT 3295.505 379.185 3295.785 379.465 ;
        RECT 3296.215 379.185 3296.495 379.465 ;
        RECT 3296.925 379.185 3297.205 379.465 ;
        RECT 3297.635 379.185 3297.915 379.465 ;
        RECT 3298.345 379.185 3298.625 379.465 ;
        RECT 3289.115 378.475 3289.395 378.755 ;
        RECT 3289.825 378.475 3290.105 378.755 ;
        RECT 3290.535 378.475 3290.815 378.755 ;
        RECT 3291.245 378.475 3291.525 378.755 ;
        RECT 3291.955 378.475 3292.235 378.755 ;
        RECT 3292.665 378.475 3292.945 378.755 ;
        RECT 3293.375 378.475 3293.655 378.755 ;
        RECT 3294.085 378.475 3294.365 378.755 ;
        RECT 3294.795 378.475 3295.075 378.755 ;
        RECT 3295.505 378.475 3295.785 378.755 ;
        RECT 3296.215 378.475 3296.495 378.755 ;
        RECT 3296.925 378.475 3297.205 378.755 ;
        RECT 3297.635 378.475 3297.915 378.755 ;
        RECT 3298.345 378.475 3298.625 378.755 ;
        RECT 3289.115 377.765 3289.395 378.045 ;
        RECT 3289.825 377.765 3290.105 378.045 ;
        RECT 3290.535 377.765 3290.815 378.045 ;
        RECT 3291.245 377.765 3291.525 378.045 ;
        RECT 3291.955 377.765 3292.235 378.045 ;
        RECT 3292.665 377.765 3292.945 378.045 ;
        RECT 3293.375 377.765 3293.655 378.045 ;
        RECT 3294.085 377.765 3294.365 378.045 ;
        RECT 3294.795 377.765 3295.075 378.045 ;
        RECT 3295.505 377.765 3295.785 378.045 ;
        RECT 3296.215 377.765 3296.495 378.045 ;
        RECT 3296.925 377.765 3297.205 378.045 ;
        RECT 3297.635 377.765 3297.915 378.045 ;
        RECT 3298.345 377.765 3298.625 378.045 ;
        RECT 3289.115 377.055 3289.395 377.335 ;
        RECT 3289.825 377.055 3290.105 377.335 ;
        RECT 3290.535 377.055 3290.815 377.335 ;
        RECT 3291.245 377.055 3291.525 377.335 ;
        RECT 3291.955 377.055 3292.235 377.335 ;
        RECT 3292.665 377.055 3292.945 377.335 ;
        RECT 3293.375 377.055 3293.655 377.335 ;
        RECT 3294.085 377.055 3294.365 377.335 ;
        RECT 3294.795 377.055 3295.075 377.335 ;
        RECT 3295.505 377.055 3295.785 377.335 ;
        RECT 3296.215 377.055 3296.495 377.335 ;
        RECT 3296.925 377.055 3297.205 377.335 ;
        RECT 3297.635 377.055 3297.915 377.335 ;
        RECT 3298.345 377.055 3298.625 377.335 ;
        RECT 3289.115 376.345 3289.395 376.625 ;
        RECT 3289.825 376.345 3290.105 376.625 ;
        RECT 3290.535 376.345 3290.815 376.625 ;
        RECT 3291.245 376.345 3291.525 376.625 ;
        RECT 3291.955 376.345 3292.235 376.625 ;
        RECT 3292.665 376.345 3292.945 376.625 ;
        RECT 3293.375 376.345 3293.655 376.625 ;
        RECT 3294.085 376.345 3294.365 376.625 ;
        RECT 3294.795 376.345 3295.075 376.625 ;
        RECT 3295.505 376.345 3295.785 376.625 ;
        RECT 3296.215 376.345 3296.495 376.625 ;
        RECT 3296.925 376.345 3297.205 376.625 ;
        RECT 3297.635 376.345 3297.915 376.625 ;
        RECT 3298.345 376.345 3298.625 376.625 ;
        RECT 3289.115 375.635 3289.395 375.915 ;
        RECT 3289.825 375.635 3290.105 375.915 ;
        RECT 3290.535 375.635 3290.815 375.915 ;
        RECT 3291.245 375.635 3291.525 375.915 ;
        RECT 3291.955 375.635 3292.235 375.915 ;
        RECT 3292.665 375.635 3292.945 375.915 ;
        RECT 3293.375 375.635 3293.655 375.915 ;
        RECT 3294.085 375.635 3294.365 375.915 ;
        RECT 3294.795 375.635 3295.075 375.915 ;
        RECT 3295.505 375.635 3295.785 375.915 ;
        RECT 3296.215 375.635 3296.495 375.915 ;
        RECT 3296.925 375.635 3297.205 375.915 ;
        RECT 3297.635 375.635 3297.915 375.915 ;
        RECT 3298.345 375.635 3298.625 375.915 ;
        RECT 3289.115 374.925 3289.395 375.205 ;
        RECT 3289.825 374.925 3290.105 375.205 ;
        RECT 3290.535 374.925 3290.815 375.205 ;
        RECT 3291.245 374.925 3291.525 375.205 ;
        RECT 3291.955 374.925 3292.235 375.205 ;
        RECT 3292.665 374.925 3292.945 375.205 ;
        RECT 3293.375 374.925 3293.655 375.205 ;
        RECT 3294.085 374.925 3294.365 375.205 ;
        RECT 3294.795 374.925 3295.075 375.205 ;
        RECT 3295.505 374.925 3295.785 375.205 ;
        RECT 3296.215 374.925 3296.495 375.205 ;
        RECT 3296.925 374.925 3297.205 375.205 ;
        RECT 3297.635 374.925 3297.915 375.205 ;
        RECT 3298.345 374.925 3298.625 375.205 ;
        RECT 3289.115 374.215 3289.395 374.495 ;
        RECT 3289.825 374.215 3290.105 374.495 ;
        RECT 3290.535 374.215 3290.815 374.495 ;
        RECT 3291.245 374.215 3291.525 374.495 ;
        RECT 3291.955 374.215 3292.235 374.495 ;
        RECT 3292.665 374.215 3292.945 374.495 ;
        RECT 3293.375 374.215 3293.655 374.495 ;
        RECT 3294.085 374.215 3294.365 374.495 ;
        RECT 3294.795 374.215 3295.075 374.495 ;
        RECT 3295.505 374.215 3295.785 374.495 ;
        RECT 3296.215 374.215 3296.495 374.495 ;
        RECT 3296.925 374.215 3297.205 374.495 ;
        RECT 3297.635 374.215 3297.915 374.495 ;
        RECT 3298.345 374.215 3298.625 374.495 ;
        RECT 3289.115 373.505 3289.395 373.785 ;
        RECT 3289.825 373.505 3290.105 373.785 ;
        RECT 3290.535 373.505 3290.815 373.785 ;
        RECT 3291.245 373.505 3291.525 373.785 ;
        RECT 3291.955 373.505 3292.235 373.785 ;
        RECT 3292.665 373.505 3292.945 373.785 ;
        RECT 3293.375 373.505 3293.655 373.785 ;
        RECT 3294.085 373.505 3294.365 373.785 ;
        RECT 3294.795 373.505 3295.075 373.785 ;
        RECT 3295.505 373.505 3295.785 373.785 ;
        RECT 3296.215 373.505 3296.495 373.785 ;
        RECT 3296.925 373.505 3297.205 373.785 ;
        RECT 3297.635 373.505 3297.915 373.785 ;
        RECT 3298.345 373.505 3298.625 373.785 ;
        RECT 3289.115 372.795 3289.395 373.075 ;
        RECT 3289.825 372.795 3290.105 373.075 ;
        RECT 3290.535 372.795 3290.815 373.075 ;
        RECT 3291.245 372.795 3291.525 373.075 ;
        RECT 3291.955 372.795 3292.235 373.075 ;
        RECT 3292.665 372.795 3292.945 373.075 ;
        RECT 3293.375 372.795 3293.655 373.075 ;
        RECT 3294.085 372.795 3294.365 373.075 ;
        RECT 3294.795 372.795 3295.075 373.075 ;
        RECT 3295.505 372.795 3295.785 373.075 ;
        RECT 3296.215 372.795 3296.495 373.075 ;
        RECT 3296.925 372.795 3297.205 373.075 ;
        RECT 3297.635 372.795 3297.915 373.075 ;
        RECT 3298.345 372.795 3298.625 373.075 ;
        RECT 3300.965 379.895 3301.245 380.175 ;
        RECT 3301.675 379.895 3301.955 380.175 ;
        RECT 3302.385 379.895 3302.665 380.175 ;
        RECT 3303.095 379.895 3303.375 380.175 ;
        RECT 3303.805 379.895 3304.085 380.175 ;
        RECT 3304.515 379.895 3304.795 380.175 ;
        RECT 3305.225 379.895 3305.505 380.175 ;
        RECT 3305.935 379.895 3306.215 380.175 ;
        RECT 3306.645 379.895 3306.925 380.175 ;
        RECT 3307.355 379.895 3307.635 380.175 ;
        RECT 3308.065 379.895 3308.345 380.175 ;
        RECT 3308.775 379.895 3309.055 380.175 ;
        RECT 3309.485 379.895 3309.765 380.175 ;
        RECT 3310.195 379.895 3310.475 380.175 ;
        RECT 3300.965 379.185 3301.245 379.465 ;
        RECT 3301.675 379.185 3301.955 379.465 ;
        RECT 3302.385 379.185 3302.665 379.465 ;
        RECT 3303.095 379.185 3303.375 379.465 ;
        RECT 3303.805 379.185 3304.085 379.465 ;
        RECT 3304.515 379.185 3304.795 379.465 ;
        RECT 3305.225 379.185 3305.505 379.465 ;
        RECT 3305.935 379.185 3306.215 379.465 ;
        RECT 3306.645 379.185 3306.925 379.465 ;
        RECT 3307.355 379.185 3307.635 379.465 ;
        RECT 3308.065 379.185 3308.345 379.465 ;
        RECT 3308.775 379.185 3309.055 379.465 ;
        RECT 3309.485 379.185 3309.765 379.465 ;
        RECT 3310.195 379.185 3310.475 379.465 ;
        RECT 3300.965 378.475 3301.245 378.755 ;
        RECT 3301.675 378.475 3301.955 378.755 ;
        RECT 3302.385 378.475 3302.665 378.755 ;
        RECT 3303.095 378.475 3303.375 378.755 ;
        RECT 3303.805 378.475 3304.085 378.755 ;
        RECT 3304.515 378.475 3304.795 378.755 ;
        RECT 3305.225 378.475 3305.505 378.755 ;
        RECT 3305.935 378.475 3306.215 378.755 ;
        RECT 3306.645 378.475 3306.925 378.755 ;
        RECT 3307.355 378.475 3307.635 378.755 ;
        RECT 3308.065 378.475 3308.345 378.755 ;
        RECT 3308.775 378.475 3309.055 378.755 ;
        RECT 3309.485 378.475 3309.765 378.755 ;
        RECT 3310.195 378.475 3310.475 378.755 ;
        RECT 3300.965 377.765 3301.245 378.045 ;
        RECT 3301.675 377.765 3301.955 378.045 ;
        RECT 3302.385 377.765 3302.665 378.045 ;
        RECT 3303.095 377.765 3303.375 378.045 ;
        RECT 3303.805 377.765 3304.085 378.045 ;
        RECT 3304.515 377.765 3304.795 378.045 ;
        RECT 3305.225 377.765 3305.505 378.045 ;
        RECT 3305.935 377.765 3306.215 378.045 ;
        RECT 3306.645 377.765 3306.925 378.045 ;
        RECT 3307.355 377.765 3307.635 378.045 ;
        RECT 3308.065 377.765 3308.345 378.045 ;
        RECT 3308.775 377.765 3309.055 378.045 ;
        RECT 3309.485 377.765 3309.765 378.045 ;
        RECT 3310.195 377.765 3310.475 378.045 ;
        RECT 3300.965 377.055 3301.245 377.335 ;
        RECT 3301.675 377.055 3301.955 377.335 ;
        RECT 3302.385 377.055 3302.665 377.335 ;
        RECT 3303.095 377.055 3303.375 377.335 ;
        RECT 3303.805 377.055 3304.085 377.335 ;
        RECT 3304.515 377.055 3304.795 377.335 ;
        RECT 3305.225 377.055 3305.505 377.335 ;
        RECT 3305.935 377.055 3306.215 377.335 ;
        RECT 3306.645 377.055 3306.925 377.335 ;
        RECT 3307.355 377.055 3307.635 377.335 ;
        RECT 3308.065 377.055 3308.345 377.335 ;
        RECT 3308.775 377.055 3309.055 377.335 ;
        RECT 3309.485 377.055 3309.765 377.335 ;
        RECT 3310.195 377.055 3310.475 377.335 ;
        RECT 3300.965 376.345 3301.245 376.625 ;
        RECT 3301.675 376.345 3301.955 376.625 ;
        RECT 3302.385 376.345 3302.665 376.625 ;
        RECT 3303.095 376.345 3303.375 376.625 ;
        RECT 3303.805 376.345 3304.085 376.625 ;
        RECT 3304.515 376.345 3304.795 376.625 ;
        RECT 3305.225 376.345 3305.505 376.625 ;
        RECT 3305.935 376.345 3306.215 376.625 ;
        RECT 3306.645 376.345 3306.925 376.625 ;
        RECT 3307.355 376.345 3307.635 376.625 ;
        RECT 3308.065 376.345 3308.345 376.625 ;
        RECT 3308.775 376.345 3309.055 376.625 ;
        RECT 3309.485 376.345 3309.765 376.625 ;
        RECT 3310.195 376.345 3310.475 376.625 ;
        RECT 3300.965 375.635 3301.245 375.915 ;
        RECT 3301.675 375.635 3301.955 375.915 ;
        RECT 3302.385 375.635 3302.665 375.915 ;
        RECT 3303.095 375.635 3303.375 375.915 ;
        RECT 3303.805 375.635 3304.085 375.915 ;
        RECT 3304.515 375.635 3304.795 375.915 ;
        RECT 3305.225 375.635 3305.505 375.915 ;
        RECT 3305.935 375.635 3306.215 375.915 ;
        RECT 3306.645 375.635 3306.925 375.915 ;
        RECT 3307.355 375.635 3307.635 375.915 ;
        RECT 3308.065 375.635 3308.345 375.915 ;
        RECT 3308.775 375.635 3309.055 375.915 ;
        RECT 3309.485 375.635 3309.765 375.915 ;
        RECT 3310.195 375.635 3310.475 375.915 ;
        RECT 3300.965 374.925 3301.245 375.205 ;
        RECT 3301.675 374.925 3301.955 375.205 ;
        RECT 3302.385 374.925 3302.665 375.205 ;
        RECT 3303.095 374.925 3303.375 375.205 ;
        RECT 3303.805 374.925 3304.085 375.205 ;
        RECT 3304.515 374.925 3304.795 375.205 ;
        RECT 3305.225 374.925 3305.505 375.205 ;
        RECT 3305.935 374.925 3306.215 375.205 ;
        RECT 3306.645 374.925 3306.925 375.205 ;
        RECT 3307.355 374.925 3307.635 375.205 ;
        RECT 3308.065 374.925 3308.345 375.205 ;
        RECT 3308.775 374.925 3309.055 375.205 ;
        RECT 3309.485 374.925 3309.765 375.205 ;
        RECT 3310.195 374.925 3310.475 375.205 ;
        RECT 3300.965 374.215 3301.245 374.495 ;
        RECT 3301.675 374.215 3301.955 374.495 ;
        RECT 3302.385 374.215 3302.665 374.495 ;
        RECT 3303.095 374.215 3303.375 374.495 ;
        RECT 3303.805 374.215 3304.085 374.495 ;
        RECT 3304.515 374.215 3304.795 374.495 ;
        RECT 3305.225 374.215 3305.505 374.495 ;
        RECT 3305.935 374.215 3306.215 374.495 ;
        RECT 3306.645 374.215 3306.925 374.495 ;
        RECT 3307.355 374.215 3307.635 374.495 ;
        RECT 3308.065 374.215 3308.345 374.495 ;
        RECT 3308.775 374.215 3309.055 374.495 ;
        RECT 3309.485 374.215 3309.765 374.495 ;
        RECT 3310.195 374.215 3310.475 374.495 ;
        RECT 3300.965 373.505 3301.245 373.785 ;
        RECT 3301.675 373.505 3301.955 373.785 ;
        RECT 3302.385 373.505 3302.665 373.785 ;
        RECT 3303.095 373.505 3303.375 373.785 ;
        RECT 3303.805 373.505 3304.085 373.785 ;
        RECT 3304.515 373.505 3304.795 373.785 ;
        RECT 3305.225 373.505 3305.505 373.785 ;
        RECT 3305.935 373.505 3306.215 373.785 ;
        RECT 3306.645 373.505 3306.925 373.785 ;
        RECT 3307.355 373.505 3307.635 373.785 ;
        RECT 3308.065 373.505 3308.345 373.785 ;
        RECT 3308.775 373.505 3309.055 373.785 ;
        RECT 3309.485 373.505 3309.765 373.785 ;
        RECT 3310.195 373.505 3310.475 373.785 ;
        RECT 3300.965 372.795 3301.245 373.075 ;
        RECT 3301.675 372.795 3301.955 373.075 ;
        RECT 3302.385 372.795 3302.665 373.075 ;
        RECT 3303.095 372.795 3303.375 373.075 ;
        RECT 3303.805 372.795 3304.085 373.075 ;
        RECT 3304.515 372.795 3304.795 373.075 ;
        RECT 3305.225 372.795 3305.505 373.075 ;
        RECT 3305.935 372.795 3306.215 373.075 ;
        RECT 3306.645 372.795 3306.925 373.075 ;
        RECT 3307.355 372.795 3307.635 373.075 ;
        RECT 3308.065 372.795 3308.345 373.075 ;
        RECT 3308.775 372.795 3309.055 373.075 ;
        RECT 3309.485 372.795 3309.765 373.075 ;
        RECT 3310.195 372.795 3310.475 373.075 ;
        RECT 3314.495 379.895 3314.775 380.175 ;
        RECT 3315.205 379.895 3315.485 380.175 ;
        RECT 3315.915 379.895 3316.195 380.175 ;
        RECT 3316.625 379.895 3316.905 380.175 ;
        RECT 3317.335 379.895 3317.615 380.175 ;
        RECT 3318.045 379.895 3318.325 380.175 ;
        RECT 3318.755 379.895 3319.035 380.175 ;
        RECT 3319.465 379.895 3319.745 380.175 ;
        RECT 3320.175 379.895 3320.455 380.175 ;
        RECT 3320.885 379.895 3321.165 380.175 ;
        RECT 3321.595 379.895 3321.875 380.175 ;
        RECT 3322.305 379.895 3322.585 380.175 ;
        RECT 3323.015 379.895 3323.295 380.175 ;
        RECT 3323.725 379.895 3324.005 380.175 ;
        RECT 3314.495 379.185 3314.775 379.465 ;
        RECT 3315.205 379.185 3315.485 379.465 ;
        RECT 3315.915 379.185 3316.195 379.465 ;
        RECT 3316.625 379.185 3316.905 379.465 ;
        RECT 3317.335 379.185 3317.615 379.465 ;
        RECT 3318.045 379.185 3318.325 379.465 ;
        RECT 3318.755 379.185 3319.035 379.465 ;
        RECT 3319.465 379.185 3319.745 379.465 ;
        RECT 3320.175 379.185 3320.455 379.465 ;
        RECT 3320.885 379.185 3321.165 379.465 ;
        RECT 3321.595 379.185 3321.875 379.465 ;
        RECT 3322.305 379.185 3322.585 379.465 ;
        RECT 3323.015 379.185 3323.295 379.465 ;
        RECT 3323.725 379.185 3324.005 379.465 ;
        RECT 3314.495 378.475 3314.775 378.755 ;
        RECT 3315.205 378.475 3315.485 378.755 ;
        RECT 3315.915 378.475 3316.195 378.755 ;
        RECT 3316.625 378.475 3316.905 378.755 ;
        RECT 3317.335 378.475 3317.615 378.755 ;
        RECT 3318.045 378.475 3318.325 378.755 ;
        RECT 3318.755 378.475 3319.035 378.755 ;
        RECT 3319.465 378.475 3319.745 378.755 ;
        RECT 3320.175 378.475 3320.455 378.755 ;
        RECT 3320.885 378.475 3321.165 378.755 ;
        RECT 3321.595 378.475 3321.875 378.755 ;
        RECT 3322.305 378.475 3322.585 378.755 ;
        RECT 3323.015 378.475 3323.295 378.755 ;
        RECT 3323.725 378.475 3324.005 378.755 ;
        RECT 3314.495 377.765 3314.775 378.045 ;
        RECT 3315.205 377.765 3315.485 378.045 ;
        RECT 3315.915 377.765 3316.195 378.045 ;
        RECT 3316.625 377.765 3316.905 378.045 ;
        RECT 3317.335 377.765 3317.615 378.045 ;
        RECT 3318.045 377.765 3318.325 378.045 ;
        RECT 3318.755 377.765 3319.035 378.045 ;
        RECT 3319.465 377.765 3319.745 378.045 ;
        RECT 3320.175 377.765 3320.455 378.045 ;
        RECT 3320.885 377.765 3321.165 378.045 ;
        RECT 3321.595 377.765 3321.875 378.045 ;
        RECT 3322.305 377.765 3322.585 378.045 ;
        RECT 3323.015 377.765 3323.295 378.045 ;
        RECT 3323.725 377.765 3324.005 378.045 ;
        RECT 3314.495 377.055 3314.775 377.335 ;
        RECT 3315.205 377.055 3315.485 377.335 ;
        RECT 3315.915 377.055 3316.195 377.335 ;
        RECT 3316.625 377.055 3316.905 377.335 ;
        RECT 3317.335 377.055 3317.615 377.335 ;
        RECT 3318.045 377.055 3318.325 377.335 ;
        RECT 3318.755 377.055 3319.035 377.335 ;
        RECT 3319.465 377.055 3319.745 377.335 ;
        RECT 3320.175 377.055 3320.455 377.335 ;
        RECT 3320.885 377.055 3321.165 377.335 ;
        RECT 3321.595 377.055 3321.875 377.335 ;
        RECT 3322.305 377.055 3322.585 377.335 ;
        RECT 3323.015 377.055 3323.295 377.335 ;
        RECT 3323.725 377.055 3324.005 377.335 ;
        RECT 3314.495 376.345 3314.775 376.625 ;
        RECT 3315.205 376.345 3315.485 376.625 ;
        RECT 3315.915 376.345 3316.195 376.625 ;
        RECT 3316.625 376.345 3316.905 376.625 ;
        RECT 3317.335 376.345 3317.615 376.625 ;
        RECT 3318.045 376.345 3318.325 376.625 ;
        RECT 3318.755 376.345 3319.035 376.625 ;
        RECT 3319.465 376.345 3319.745 376.625 ;
        RECT 3320.175 376.345 3320.455 376.625 ;
        RECT 3320.885 376.345 3321.165 376.625 ;
        RECT 3321.595 376.345 3321.875 376.625 ;
        RECT 3322.305 376.345 3322.585 376.625 ;
        RECT 3323.015 376.345 3323.295 376.625 ;
        RECT 3323.725 376.345 3324.005 376.625 ;
        RECT 3314.495 375.635 3314.775 375.915 ;
        RECT 3315.205 375.635 3315.485 375.915 ;
        RECT 3315.915 375.635 3316.195 375.915 ;
        RECT 3316.625 375.635 3316.905 375.915 ;
        RECT 3317.335 375.635 3317.615 375.915 ;
        RECT 3318.045 375.635 3318.325 375.915 ;
        RECT 3318.755 375.635 3319.035 375.915 ;
        RECT 3319.465 375.635 3319.745 375.915 ;
        RECT 3320.175 375.635 3320.455 375.915 ;
        RECT 3320.885 375.635 3321.165 375.915 ;
        RECT 3321.595 375.635 3321.875 375.915 ;
        RECT 3322.305 375.635 3322.585 375.915 ;
        RECT 3323.015 375.635 3323.295 375.915 ;
        RECT 3323.725 375.635 3324.005 375.915 ;
        RECT 3314.495 374.925 3314.775 375.205 ;
        RECT 3315.205 374.925 3315.485 375.205 ;
        RECT 3315.915 374.925 3316.195 375.205 ;
        RECT 3316.625 374.925 3316.905 375.205 ;
        RECT 3317.335 374.925 3317.615 375.205 ;
        RECT 3318.045 374.925 3318.325 375.205 ;
        RECT 3318.755 374.925 3319.035 375.205 ;
        RECT 3319.465 374.925 3319.745 375.205 ;
        RECT 3320.175 374.925 3320.455 375.205 ;
        RECT 3320.885 374.925 3321.165 375.205 ;
        RECT 3321.595 374.925 3321.875 375.205 ;
        RECT 3322.305 374.925 3322.585 375.205 ;
        RECT 3323.015 374.925 3323.295 375.205 ;
        RECT 3323.725 374.925 3324.005 375.205 ;
        RECT 3314.495 374.215 3314.775 374.495 ;
        RECT 3315.205 374.215 3315.485 374.495 ;
        RECT 3315.915 374.215 3316.195 374.495 ;
        RECT 3316.625 374.215 3316.905 374.495 ;
        RECT 3317.335 374.215 3317.615 374.495 ;
        RECT 3318.045 374.215 3318.325 374.495 ;
        RECT 3318.755 374.215 3319.035 374.495 ;
        RECT 3319.465 374.215 3319.745 374.495 ;
        RECT 3320.175 374.215 3320.455 374.495 ;
        RECT 3320.885 374.215 3321.165 374.495 ;
        RECT 3321.595 374.215 3321.875 374.495 ;
        RECT 3322.305 374.215 3322.585 374.495 ;
        RECT 3323.015 374.215 3323.295 374.495 ;
        RECT 3323.725 374.215 3324.005 374.495 ;
        RECT 3314.495 373.505 3314.775 373.785 ;
        RECT 3315.205 373.505 3315.485 373.785 ;
        RECT 3315.915 373.505 3316.195 373.785 ;
        RECT 3316.625 373.505 3316.905 373.785 ;
        RECT 3317.335 373.505 3317.615 373.785 ;
        RECT 3318.045 373.505 3318.325 373.785 ;
        RECT 3318.755 373.505 3319.035 373.785 ;
        RECT 3319.465 373.505 3319.745 373.785 ;
        RECT 3320.175 373.505 3320.455 373.785 ;
        RECT 3320.885 373.505 3321.165 373.785 ;
        RECT 3321.595 373.505 3321.875 373.785 ;
        RECT 3322.305 373.505 3322.585 373.785 ;
        RECT 3323.015 373.505 3323.295 373.785 ;
        RECT 3323.725 373.505 3324.005 373.785 ;
        RECT 3314.495 372.795 3314.775 373.075 ;
        RECT 3315.205 372.795 3315.485 373.075 ;
        RECT 3315.915 372.795 3316.195 373.075 ;
        RECT 3316.625 372.795 3316.905 373.075 ;
        RECT 3317.335 372.795 3317.615 373.075 ;
        RECT 3318.045 372.795 3318.325 373.075 ;
        RECT 3318.755 372.795 3319.035 373.075 ;
        RECT 3319.465 372.795 3319.745 373.075 ;
        RECT 3320.175 372.795 3320.455 373.075 ;
        RECT 3320.885 372.795 3321.165 373.075 ;
        RECT 3321.595 372.795 3321.875 373.075 ;
        RECT 3322.305 372.795 3322.585 373.075 ;
        RECT 3323.015 372.795 3323.295 373.075 ;
        RECT 3323.725 372.795 3324.005 373.075 ;
        RECT 3326.345 379.895 3326.625 380.175 ;
        RECT 3327.055 379.895 3327.335 380.175 ;
        RECT 3327.765 379.895 3328.045 380.175 ;
        RECT 3328.475 379.895 3328.755 380.175 ;
        RECT 3329.185 379.895 3329.465 380.175 ;
        RECT 3329.895 379.895 3330.175 380.175 ;
        RECT 3330.605 379.895 3330.885 380.175 ;
        RECT 3331.315 379.895 3331.595 380.175 ;
        RECT 3332.025 379.895 3332.305 380.175 ;
        RECT 3332.735 379.895 3333.015 380.175 ;
        RECT 3333.445 379.895 3333.725 380.175 ;
        RECT 3334.155 379.895 3334.435 380.175 ;
        RECT 3334.865 379.895 3335.145 380.175 ;
        RECT 3335.575 379.895 3335.855 380.175 ;
        RECT 3326.345 379.185 3326.625 379.465 ;
        RECT 3327.055 379.185 3327.335 379.465 ;
        RECT 3327.765 379.185 3328.045 379.465 ;
        RECT 3328.475 379.185 3328.755 379.465 ;
        RECT 3329.185 379.185 3329.465 379.465 ;
        RECT 3329.895 379.185 3330.175 379.465 ;
        RECT 3330.605 379.185 3330.885 379.465 ;
        RECT 3331.315 379.185 3331.595 379.465 ;
        RECT 3332.025 379.185 3332.305 379.465 ;
        RECT 3332.735 379.185 3333.015 379.465 ;
        RECT 3333.445 379.185 3333.725 379.465 ;
        RECT 3334.155 379.185 3334.435 379.465 ;
        RECT 3334.865 379.185 3335.145 379.465 ;
        RECT 3335.575 379.185 3335.855 379.465 ;
        RECT 3326.345 378.475 3326.625 378.755 ;
        RECT 3327.055 378.475 3327.335 378.755 ;
        RECT 3327.765 378.475 3328.045 378.755 ;
        RECT 3328.475 378.475 3328.755 378.755 ;
        RECT 3329.185 378.475 3329.465 378.755 ;
        RECT 3329.895 378.475 3330.175 378.755 ;
        RECT 3330.605 378.475 3330.885 378.755 ;
        RECT 3331.315 378.475 3331.595 378.755 ;
        RECT 3332.025 378.475 3332.305 378.755 ;
        RECT 3332.735 378.475 3333.015 378.755 ;
        RECT 3333.445 378.475 3333.725 378.755 ;
        RECT 3334.155 378.475 3334.435 378.755 ;
        RECT 3334.865 378.475 3335.145 378.755 ;
        RECT 3335.575 378.475 3335.855 378.755 ;
        RECT 3326.345 377.765 3326.625 378.045 ;
        RECT 3327.055 377.765 3327.335 378.045 ;
        RECT 3327.765 377.765 3328.045 378.045 ;
        RECT 3328.475 377.765 3328.755 378.045 ;
        RECT 3329.185 377.765 3329.465 378.045 ;
        RECT 3329.895 377.765 3330.175 378.045 ;
        RECT 3330.605 377.765 3330.885 378.045 ;
        RECT 3331.315 377.765 3331.595 378.045 ;
        RECT 3332.025 377.765 3332.305 378.045 ;
        RECT 3332.735 377.765 3333.015 378.045 ;
        RECT 3333.445 377.765 3333.725 378.045 ;
        RECT 3334.155 377.765 3334.435 378.045 ;
        RECT 3334.865 377.765 3335.145 378.045 ;
        RECT 3335.575 377.765 3335.855 378.045 ;
        RECT 3326.345 377.055 3326.625 377.335 ;
        RECT 3327.055 377.055 3327.335 377.335 ;
        RECT 3327.765 377.055 3328.045 377.335 ;
        RECT 3328.475 377.055 3328.755 377.335 ;
        RECT 3329.185 377.055 3329.465 377.335 ;
        RECT 3329.895 377.055 3330.175 377.335 ;
        RECT 3330.605 377.055 3330.885 377.335 ;
        RECT 3331.315 377.055 3331.595 377.335 ;
        RECT 3332.025 377.055 3332.305 377.335 ;
        RECT 3332.735 377.055 3333.015 377.335 ;
        RECT 3333.445 377.055 3333.725 377.335 ;
        RECT 3334.155 377.055 3334.435 377.335 ;
        RECT 3334.865 377.055 3335.145 377.335 ;
        RECT 3335.575 377.055 3335.855 377.335 ;
        RECT 3326.345 376.345 3326.625 376.625 ;
        RECT 3327.055 376.345 3327.335 376.625 ;
        RECT 3327.765 376.345 3328.045 376.625 ;
        RECT 3328.475 376.345 3328.755 376.625 ;
        RECT 3329.185 376.345 3329.465 376.625 ;
        RECT 3329.895 376.345 3330.175 376.625 ;
        RECT 3330.605 376.345 3330.885 376.625 ;
        RECT 3331.315 376.345 3331.595 376.625 ;
        RECT 3332.025 376.345 3332.305 376.625 ;
        RECT 3332.735 376.345 3333.015 376.625 ;
        RECT 3333.445 376.345 3333.725 376.625 ;
        RECT 3334.155 376.345 3334.435 376.625 ;
        RECT 3334.865 376.345 3335.145 376.625 ;
        RECT 3335.575 376.345 3335.855 376.625 ;
        RECT 3326.345 375.635 3326.625 375.915 ;
        RECT 3327.055 375.635 3327.335 375.915 ;
        RECT 3327.765 375.635 3328.045 375.915 ;
        RECT 3328.475 375.635 3328.755 375.915 ;
        RECT 3329.185 375.635 3329.465 375.915 ;
        RECT 3329.895 375.635 3330.175 375.915 ;
        RECT 3330.605 375.635 3330.885 375.915 ;
        RECT 3331.315 375.635 3331.595 375.915 ;
        RECT 3332.025 375.635 3332.305 375.915 ;
        RECT 3332.735 375.635 3333.015 375.915 ;
        RECT 3333.445 375.635 3333.725 375.915 ;
        RECT 3334.155 375.635 3334.435 375.915 ;
        RECT 3334.865 375.635 3335.145 375.915 ;
        RECT 3335.575 375.635 3335.855 375.915 ;
        RECT 3326.345 374.925 3326.625 375.205 ;
        RECT 3327.055 374.925 3327.335 375.205 ;
        RECT 3327.765 374.925 3328.045 375.205 ;
        RECT 3328.475 374.925 3328.755 375.205 ;
        RECT 3329.185 374.925 3329.465 375.205 ;
        RECT 3329.895 374.925 3330.175 375.205 ;
        RECT 3330.605 374.925 3330.885 375.205 ;
        RECT 3331.315 374.925 3331.595 375.205 ;
        RECT 3332.025 374.925 3332.305 375.205 ;
        RECT 3332.735 374.925 3333.015 375.205 ;
        RECT 3333.445 374.925 3333.725 375.205 ;
        RECT 3334.155 374.925 3334.435 375.205 ;
        RECT 3334.865 374.925 3335.145 375.205 ;
        RECT 3335.575 374.925 3335.855 375.205 ;
        RECT 3326.345 374.215 3326.625 374.495 ;
        RECT 3327.055 374.215 3327.335 374.495 ;
        RECT 3327.765 374.215 3328.045 374.495 ;
        RECT 3328.475 374.215 3328.755 374.495 ;
        RECT 3329.185 374.215 3329.465 374.495 ;
        RECT 3329.895 374.215 3330.175 374.495 ;
        RECT 3330.605 374.215 3330.885 374.495 ;
        RECT 3331.315 374.215 3331.595 374.495 ;
        RECT 3332.025 374.215 3332.305 374.495 ;
        RECT 3332.735 374.215 3333.015 374.495 ;
        RECT 3333.445 374.215 3333.725 374.495 ;
        RECT 3334.155 374.215 3334.435 374.495 ;
        RECT 3334.865 374.215 3335.145 374.495 ;
        RECT 3335.575 374.215 3335.855 374.495 ;
        RECT 3326.345 373.505 3326.625 373.785 ;
        RECT 3327.055 373.505 3327.335 373.785 ;
        RECT 3327.765 373.505 3328.045 373.785 ;
        RECT 3328.475 373.505 3328.755 373.785 ;
        RECT 3329.185 373.505 3329.465 373.785 ;
        RECT 3329.895 373.505 3330.175 373.785 ;
        RECT 3330.605 373.505 3330.885 373.785 ;
        RECT 3331.315 373.505 3331.595 373.785 ;
        RECT 3332.025 373.505 3332.305 373.785 ;
        RECT 3332.735 373.505 3333.015 373.785 ;
        RECT 3333.445 373.505 3333.725 373.785 ;
        RECT 3334.155 373.505 3334.435 373.785 ;
        RECT 3334.865 373.505 3335.145 373.785 ;
        RECT 3335.575 373.505 3335.855 373.785 ;
        RECT 3326.345 372.795 3326.625 373.075 ;
        RECT 3327.055 372.795 3327.335 373.075 ;
        RECT 3327.765 372.795 3328.045 373.075 ;
        RECT 3328.475 372.795 3328.755 373.075 ;
        RECT 3329.185 372.795 3329.465 373.075 ;
        RECT 3329.895 372.795 3330.175 373.075 ;
        RECT 3330.605 372.795 3330.885 373.075 ;
        RECT 3331.315 372.795 3331.595 373.075 ;
        RECT 3332.025 372.795 3332.305 373.075 ;
        RECT 3332.735 372.795 3333.015 373.075 ;
        RECT 3333.445 372.795 3333.725 373.075 ;
        RECT 3334.155 372.795 3334.435 373.075 ;
        RECT 3334.865 372.795 3335.145 373.075 ;
        RECT 3335.575 372.795 3335.855 373.075 ;
        RECT 3339.495 379.895 3339.775 380.175 ;
        RECT 3340.205 379.895 3340.485 380.175 ;
        RECT 3344.465 379.895 3344.745 380.175 ;
        RECT 3345.175 379.895 3345.455 380.175 ;
        RECT 3345.885 379.895 3346.165 380.175 ;
        RECT 3346.595 379.895 3346.875 380.175 ;
        RECT 3347.305 379.895 3347.585 380.175 ;
        RECT 3348.015 379.895 3348.295 380.175 ;
        RECT 3339.495 379.185 3339.775 379.465 ;
        RECT 3340.205 379.185 3340.485 379.465 ;
        RECT 3344.465 379.185 3344.745 379.465 ;
        RECT 3345.175 379.185 3345.455 379.465 ;
        RECT 3345.885 379.185 3346.165 379.465 ;
        RECT 3346.595 379.185 3346.875 379.465 ;
        RECT 3347.305 379.185 3347.585 379.465 ;
        RECT 3348.015 379.185 3348.295 379.465 ;
        RECT 3339.495 378.475 3339.775 378.755 ;
        RECT 3340.205 378.475 3340.485 378.755 ;
        RECT 3344.465 378.475 3344.745 378.755 ;
        RECT 3345.175 378.475 3345.455 378.755 ;
        RECT 3345.885 378.475 3346.165 378.755 ;
        RECT 3346.595 378.475 3346.875 378.755 ;
        RECT 3347.305 378.475 3347.585 378.755 ;
        RECT 3348.015 378.475 3348.295 378.755 ;
        RECT 3339.495 377.765 3339.775 378.045 ;
        RECT 3340.205 377.765 3340.485 378.045 ;
        RECT 3344.465 377.765 3344.745 378.045 ;
        RECT 3345.175 377.765 3345.455 378.045 ;
        RECT 3345.885 377.765 3346.165 378.045 ;
        RECT 3346.595 377.765 3346.875 378.045 ;
        RECT 3347.305 377.765 3347.585 378.045 ;
        RECT 3348.015 377.765 3348.295 378.045 ;
        RECT 3339.495 377.055 3339.775 377.335 ;
        RECT 3340.205 377.055 3340.485 377.335 ;
        RECT 3344.465 377.055 3344.745 377.335 ;
        RECT 3345.175 377.055 3345.455 377.335 ;
        RECT 3345.885 377.055 3346.165 377.335 ;
        RECT 3346.595 377.055 3346.875 377.335 ;
        RECT 3347.305 377.055 3347.585 377.335 ;
        RECT 3348.015 377.055 3348.295 377.335 ;
        RECT 3339.495 376.345 3339.775 376.625 ;
        RECT 3340.205 376.345 3340.485 376.625 ;
        RECT 3344.465 376.345 3344.745 376.625 ;
        RECT 3345.175 376.345 3345.455 376.625 ;
        RECT 3345.885 376.345 3346.165 376.625 ;
        RECT 3346.595 376.345 3346.875 376.625 ;
        RECT 3347.305 376.345 3347.585 376.625 ;
        RECT 3348.015 376.345 3348.295 376.625 ;
        RECT 3339.495 375.635 3339.775 375.915 ;
        RECT 3340.205 375.635 3340.485 375.915 ;
        RECT 3344.465 375.635 3344.745 375.915 ;
        RECT 3345.175 375.635 3345.455 375.915 ;
        RECT 3345.885 375.635 3346.165 375.915 ;
        RECT 3346.595 375.635 3346.875 375.915 ;
        RECT 3347.305 375.635 3347.585 375.915 ;
        RECT 3348.015 375.635 3348.295 375.915 ;
        RECT 3339.495 374.925 3339.775 375.205 ;
        RECT 3340.205 374.925 3340.485 375.205 ;
        RECT 3344.465 374.925 3344.745 375.205 ;
        RECT 3345.175 374.925 3345.455 375.205 ;
        RECT 3345.885 374.925 3346.165 375.205 ;
        RECT 3346.595 374.925 3346.875 375.205 ;
        RECT 3347.305 374.925 3347.585 375.205 ;
        RECT 3348.015 374.925 3348.295 375.205 ;
        RECT 3339.495 374.215 3339.775 374.495 ;
        RECT 3340.205 374.215 3340.485 374.495 ;
        RECT 3344.465 374.215 3344.745 374.495 ;
        RECT 3345.175 374.215 3345.455 374.495 ;
        RECT 3345.885 374.215 3346.165 374.495 ;
        RECT 3346.595 374.215 3346.875 374.495 ;
        RECT 3347.305 374.215 3347.585 374.495 ;
        RECT 3348.015 374.215 3348.295 374.495 ;
        RECT 3339.495 373.505 3339.775 373.785 ;
        RECT 3340.205 373.505 3340.485 373.785 ;
        RECT 3344.465 373.505 3344.745 373.785 ;
        RECT 3345.175 373.505 3345.455 373.785 ;
        RECT 3345.885 373.505 3346.165 373.785 ;
        RECT 3346.595 373.505 3346.875 373.785 ;
        RECT 3347.305 373.505 3347.585 373.785 ;
        RECT 3348.015 373.505 3348.295 373.785 ;
        RECT 3339.495 372.795 3339.775 373.075 ;
        RECT 3340.205 372.795 3340.485 373.075 ;
        RECT 3344.465 372.795 3344.745 373.075 ;
        RECT 3345.175 372.795 3345.455 373.075 ;
        RECT 3345.885 372.795 3346.165 373.075 ;
        RECT 3346.595 372.795 3346.875 373.075 ;
        RECT 3347.305 372.795 3347.585 373.075 ;
        RECT 3348.015 372.795 3348.295 373.075 ;
        RECT 526.715 369.895 526.995 370.175 ;
        RECT 527.425 369.895 527.705 370.175 ;
        RECT 528.135 369.895 528.415 370.175 ;
        RECT 528.845 369.895 529.125 370.175 ;
        RECT 529.555 369.895 529.835 370.175 ;
        RECT 530.265 369.895 530.545 370.175 ;
        RECT 530.975 369.895 531.255 370.175 ;
        RECT 531.685 369.895 531.965 370.175 ;
        RECT 532.395 369.895 532.675 370.175 ;
        RECT 533.105 369.895 533.385 370.175 ;
        RECT 533.815 369.895 534.095 370.175 ;
        RECT 534.525 369.895 534.805 370.175 ;
        RECT 535.235 369.895 535.515 370.175 ;
        RECT 526.715 369.185 526.995 369.465 ;
        RECT 527.425 369.185 527.705 369.465 ;
        RECT 528.135 369.185 528.415 369.465 ;
        RECT 528.845 369.185 529.125 369.465 ;
        RECT 529.555 369.185 529.835 369.465 ;
        RECT 530.265 369.185 530.545 369.465 ;
        RECT 530.975 369.185 531.255 369.465 ;
        RECT 531.685 369.185 531.965 369.465 ;
        RECT 532.395 369.185 532.675 369.465 ;
        RECT 533.105 369.185 533.385 369.465 ;
        RECT 533.815 369.185 534.095 369.465 ;
        RECT 534.525 369.185 534.805 369.465 ;
        RECT 535.235 369.185 535.515 369.465 ;
        RECT 526.715 368.475 526.995 368.755 ;
        RECT 527.425 368.475 527.705 368.755 ;
        RECT 528.135 368.475 528.415 368.755 ;
        RECT 528.845 368.475 529.125 368.755 ;
        RECT 529.555 368.475 529.835 368.755 ;
        RECT 530.265 368.475 530.545 368.755 ;
        RECT 530.975 368.475 531.255 368.755 ;
        RECT 531.685 368.475 531.965 368.755 ;
        RECT 532.395 368.475 532.675 368.755 ;
        RECT 533.105 368.475 533.385 368.755 ;
        RECT 533.815 368.475 534.095 368.755 ;
        RECT 534.525 368.475 534.805 368.755 ;
        RECT 535.235 368.475 535.515 368.755 ;
        RECT 526.715 367.765 526.995 368.045 ;
        RECT 527.425 367.765 527.705 368.045 ;
        RECT 528.135 367.765 528.415 368.045 ;
        RECT 528.845 367.765 529.125 368.045 ;
        RECT 529.555 367.765 529.835 368.045 ;
        RECT 530.265 367.765 530.545 368.045 ;
        RECT 530.975 367.765 531.255 368.045 ;
        RECT 531.685 367.765 531.965 368.045 ;
        RECT 532.395 367.765 532.675 368.045 ;
        RECT 533.105 367.765 533.385 368.045 ;
        RECT 533.815 367.765 534.095 368.045 ;
        RECT 534.525 367.765 534.805 368.045 ;
        RECT 535.235 367.765 535.515 368.045 ;
        RECT 526.715 367.055 526.995 367.335 ;
        RECT 527.425 367.055 527.705 367.335 ;
        RECT 528.135 367.055 528.415 367.335 ;
        RECT 528.845 367.055 529.125 367.335 ;
        RECT 529.555 367.055 529.835 367.335 ;
        RECT 530.265 367.055 530.545 367.335 ;
        RECT 530.975 367.055 531.255 367.335 ;
        RECT 531.685 367.055 531.965 367.335 ;
        RECT 532.395 367.055 532.675 367.335 ;
        RECT 533.105 367.055 533.385 367.335 ;
        RECT 533.815 367.055 534.095 367.335 ;
        RECT 534.525 367.055 534.805 367.335 ;
        RECT 535.235 367.055 535.515 367.335 ;
        RECT 526.715 366.345 526.995 366.625 ;
        RECT 527.425 366.345 527.705 366.625 ;
        RECT 528.135 366.345 528.415 366.625 ;
        RECT 528.845 366.345 529.125 366.625 ;
        RECT 529.555 366.345 529.835 366.625 ;
        RECT 530.265 366.345 530.545 366.625 ;
        RECT 530.975 366.345 531.255 366.625 ;
        RECT 531.685 366.345 531.965 366.625 ;
        RECT 532.395 366.345 532.675 366.625 ;
        RECT 533.105 366.345 533.385 366.625 ;
        RECT 533.815 366.345 534.095 366.625 ;
        RECT 534.525 366.345 534.805 366.625 ;
        RECT 535.235 366.345 535.515 366.625 ;
        RECT 526.715 365.635 526.995 365.915 ;
        RECT 527.425 365.635 527.705 365.915 ;
        RECT 528.135 365.635 528.415 365.915 ;
        RECT 528.845 365.635 529.125 365.915 ;
        RECT 529.555 365.635 529.835 365.915 ;
        RECT 530.265 365.635 530.545 365.915 ;
        RECT 530.975 365.635 531.255 365.915 ;
        RECT 531.685 365.635 531.965 365.915 ;
        RECT 532.395 365.635 532.675 365.915 ;
        RECT 533.105 365.635 533.385 365.915 ;
        RECT 533.815 365.635 534.095 365.915 ;
        RECT 534.525 365.635 534.805 365.915 ;
        RECT 535.235 365.635 535.515 365.915 ;
        RECT 526.715 364.925 526.995 365.205 ;
        RECT 527.425 364.925 527.705 365.205 ;
        RECT 528.135 364.925 528.415 365.205 ;
        RECT 528.845 364.925 529.125 365.205 ;
        RECT 529.555 364.925 529.835 365.205 ;
        RECT 530.265 364.925 530.545 365.205 ;
        RECT 530.975 364.925 531.255 365.205 ;
        RECT 531.685 364.925 531.965 365.205 ;
        RECT 532.395 364.925 532.675 365.205 ;
        RECT 533.105 364.925 533.385 365.205 ;
        RECT 533.815 364.925 534.095 365.205 ;
        RECT 534.525 364.925 534.805 365.205 ;
        RECT 535.235 364.925 535.515 365.205 ;
        RECT 526.715 364.215 526.995 364.495 ;
        RECT 527.425 364.215 527.705 364.495 ;
        RECT 528.135 364.215 528.415 364.495 ;
        RECT 528.845 364.215 529.125 364.495 ;
        RECT 529.555 364.215 529.835 364.495 ;
        RECT 530.265 364.215 530.545 364.495 ;
        RECT 530.975 364.215 531.255 364.495 ;
        RECT 531.685 364.215 531.965 364.495 ;
        RECT 532.395 364.215 532.675 364.495 ;
        RECT 533.105 364.215 533.385 364.495 ;
        RECT 533.815 364.215 534.095 364.495 ;
        RECT 534.525 364.215 534.805 364.495 ;
        RECT 535.235 364.215 535.515 364.495 ;
        RECT 526.715 363.505 526.995 363.785 ;
        RECT 527.425 363.505 527.705 363.785 ;
        RECT 528.135 363.505 528.415 363.785 ;
        RECT 528.845 363.505 529.125 363.785 ;
        RECT 529.555 363.505 529.835 363.785 ;
        RECT 530.265 363.505 530.545 363.785 ;
        RECT 530.975 363.505 531.255 363.785 ;
        RECT 531.685 363.505 531.965 363.785 ;
        RECT 532.395 363.505 532.675 363.785 ;
        RECT 533.105 363.505 533.385 363.785 ;
        RECT 533.815 363.505 534.095 363.785 ;
        RECT 534.525 363.505 534.805 363.785 ;
        RECT 535.235 363.505 535.515 363.785 ;
        RECT 526.715 362.795 526.995 363.075 ;
        RECT 527.425 362.795 527.705 363.075 ;
        RECT 528.135 362.795 528.415 363.075 ;
        RECT 528.845 362.795 529.125 363.075 ;
        RECT 529.555 362.795 529.835 363.075 ;
        RECT 530.265 362.795 530.545 363.075 ;
        RECT 530.975 362.795 531.255 363.075 ;
        RECT 531.685 362.795 531.965 363.075 ;
        RECT 532.395 362.795 532.675 363.075 ;
        RECT 533.105 362.795 533.385 363.075 ;
        RECT 533.815 362.795 534.095 363.075 ;
        RECT 534.525 362.795 534.805 363.075 ;
        RECT 535.235 362.795 535.515 363.075 ;
        RECT 526.715 362.085 526.995 362.365 ;
        RECT 527.425 362.085 527.705 362.365 ;
        RECT 528.135 362.085 528.415 362.365 ;
        RECT 528.845 362.085 529.125 362.365 ;
        RECT 529.555 362.085 529.835 362.365 ;
        RECT 530.265 362.085 530.545 362.365 ;
        RECT 530.975 362.085 531.255 362.365 ;
        RECT 531.685 362.085 531.965 362.365 ;
        RECT 532.395 362.085 532.675 362.365 ;
        RECT 533.105 362.085 533.385 362.365 ;
        RECT 533.815 362.085 534.095 362.365 ;
        RECT 534.525 362.085 534.805 362.365 ;
        RECT 535.235 362.085 535.515 362.365 ;
        RECT 526.715 361.375 526.995 361.655 ;
        RECT 527.425 361.375 527.705 361.655 ;
        RECT 528.135 361.375 528.415 361.655 ;
        RECT 528.845 361.375 529.125 361.655 ;
        RECT 529.555 361.375 529.835 361.655 ;
        RECT 530.265 361.375 530.545 361.655 ;
        RECT 530.975 361.375 531.255 361.655 ;
        RECT 531.685 361.375 531.965 361.655 ;
        RECT 532.395 361.375 532.675 361.655 ;
        RECT 533.105 361.375 533.385 361.655 ;
        RECT 533.815 361.375 534.095 361.655 ;
        RECT 534.525 361.375 534.805 361.655 ;
        RECT 535.235 361.375 535.515 361.655 ;
        RECT 526.715 360.665 526.995 360.945 ;
        RECT 527.425 360.665 527.705 360.945 ;
        RECT 528.135 360.665 528.415 360.945 ;
        RECT 528.845 360.665 529.125 360.945 ;
        RECT 529.555 360.665 529.835 360.945 ;
        RECT 530.265 360.665 530.545 360.945 ;
        RECT 530.975 360.665 531.255 360.945 ;
        RECT 531.685 360.665 531.965 360.945 ;
        RECT 532.395 360.665 532.675 360.945 ;
        RECT 533.105 360.665 533.385 360.945 ;
        RECT 533.815 360.665 534.095 360.945 ;
        RECT 534.525 360.665 534.805 360.945 ;
        RECT 535.235 360.665 535.515 360.945 ;
        RECT 544.975 369.895 545.255 370.175 ;
        RECT 545.685 369.895 545.965 370.175 ;
        RECT 546.395 369.895 546.675 370.175 ;
        RECT 547.105 369.895 547.385 370.175 ;
        RECT 547.815 369.895 548.095 370.175 ;
        RECT 548.525 369.895 548.805 370.175 ;
        RECT 544.975 369.185 545.255 369.465 ;
        RECT 545.685 369.185 545.965 369.465 ;
        RECT 546.395 369.185 546.675 369.465 ;
        RECT 547.105 369.185 547.385 369.465 ;
        RECT 547.815 369.185 548.095 369.465 ;
        RECT 548.525 369.185 548.805 369.465 ;
        RECT 544.975 368.475 545.255 368.755 ;
        RECT 545.685 368.475 545.965 368.755 ;
        RECT 546.395 368.475 546.675 368.755 ;
        RECT 547.105 368.475 547.385 368.755 ;
        RECT 547.815 368.475 548.095 368.755 ;
        RECT 548.525 368.475 548.805 368.755 ;
        RECT 544.975 367.765 545.255 368.045 ;
        RECT 545.685 367.765 545.965 368.045 ;
        RECT 546.395 367.765 546.675 368.045 ;
        RECT 547.105 367.765 547.385 368.045 ;
        RECT 547.815 367.765 548.095 368.045 ;
        RECT 548.525 367.765 548.805 368.045 ;
        RECT 544.975 367.055 545.255 367.335 ;
        RECT 545.685 367.055 545.965 367.335 ;
        RECT 546.395 367.055 546.675 367.335 ;
        RECT 547.105 367.055 547.385 367.335 ;
        RECT 547.815 367.055 548.095 367.335 ;
        RECT 548.525 367.055 548.805 367.335 ;
        RECT 544.975 366.345 545.255 366.625 ;
        RECT 545.685 366.345 545.965 366.625 ;
        RECT 546.395 366.345 546.675 366.625 ;
        RECT 547.105 366.345 547.385 366.625 ;
        RECT 547.815 366.345 548.095 366.625 ;
        RECT 548.525 366.345 548.805 366.625 ;
        RECT 544.975 365.635 545.255 365.915 ;
        RECT 545.685 365.635 545.965 365.915 ;
        RECT 546.395 365.635 546.675 365.915 ;
        RECT 547.105 365.635 547.385 365.915 ;
        RECT 547.815 365.635 548.095 365.915 ;
        RECT 548.525 365.635 548.805 365.915 ;
        RECT 544.975 364.925 545.255 365.205 ;
        RECT 545.685 364.925 545.965 365.205 ;
        RECT 546.395 364.925 546.675 365.205 ;
        RECT 547.105 364.925 547.385 365.205 ;
        RECT 547.815 364.925 548.095 365.205 ;
        RECT 548.525 364.925 548.805 365.205 ;
        RECT 544.975 364.215 545.255 364.495 ;
        RECT 545.685 364.215 545.965 364.495 ;
        RECT 546.395 364.215 546.675 364.495 ;
        RECT 547.105 364.215 547.385 364.495 ;
        RECT 547.815 364.215 548.095 364.495 ;
        RECT 548.525 364.215 548.805 364.495 ;
        RECT 544.975 363.505 545.255 363.785 ;
        RECT 545.685 363.505 545.965 363.785 ;
        RECT 546.395 363.505 546.675 363.785 ;
        RECT 547.105 363.505 547.385 363.785 ;
        RECT 547.815 363.505 548.095 363.785 ;
        RECT 548.525 363.505 548.805 363.785 ;
        RECT 544.975 362.795 545.255 363.075 ;
        RECT 545.685 362.795 545.965 363.075 ;
        RECT 546.395 362.795 546.675 363.075 ;
        RECT 547.105 362.795 547.385 363.075 ;
        RECT 547.815 362.795 548.095 363.075 ;
        RECT 548.525 362.795 548.805 363.075 ;
        RECT 544.975 362.085 545.255 362.365 ;
        RECT 545.685 362.085 545.965 362.365 ;
        RECT 546.395 362.085 546.675 362.365 ;
        RECT 547.105 362.085 547.385 362.365 ;
        RECT 547.815 362.085 548.095 362.365 ;
        RECT 548.525 362.085 548.805 362.365 ;
        RECT 544.975 361.375 545.255 361.655 ;
        RECT 545.685 361.375 545.965 361.655 ;
        RECT 546.395 361.375 546.675 361.655 ;
        RECT 547.105 361.375 547.385 361.655 ;
        RECT 547.815 361.375 548.095 361.655 ;
        RECT 548.525 361.375 548.805 361.655 ;
        RECT 544.975 360.665 545.255 360.945 ;
        RECT 545.685 360.665 545.965 360.945 ;
        RECT 546.395 360.665 546.675 360.945 ;
        RECT 547.105 360.665 547.385 360.945 ;
        RECT 547.815 360.665 548.095 360.945 ;
        RECT 548.525 360.665 548.805 360.945 ;
        RECT 550.965 369.895 551.245 370.175 ;
        RECT 551.675 369.895 551.955 370.175 ;
        RECT 552.385 369.895 552.665 370.175 ;
        RECT 553.095 369.895 553.375 370.175 ;
        RECT 553.805 369.895 554.085 370.175 ;
        RECT 554.515 369.895 554.795 370.175 ;
        RECT 555.225 369.895 555.505 370.175 ;
        RECT 555.935 369.895 556.215 370.175 ;
        RECT 556.645 369.895 556.925 370.175 ;
        RECT 557.355 369.895 557.635 370.175 ;
        RECT 558.065 369.895 558.345 370.175 ;
        RECT 558.775 369.895 559.055 370.175 ;
        RECT 559.485 369.895 559.765 370.175 ;
        RECT 560.195 369.895 560.475 370.175 ;
        RECT 550.965 369.185 551.245 369.465 ;
        RECT 551.675 369.185 551.955 369.465 ;
        RECT 552.385 369.185 552.665 369.465 ;
        RECT 553.095 369.185 553.375 369.465 ;
        RECT 553.805 369.185 554.085 369.465 ;
        RECT 554.515 369.185 554.795 369.465 ;
        RECT 555.225 369.185 555.505 369.465 ;
        RECT 555.935 369.185 556.215 369.465 ;
        RECT 556.645 369.185 556.925 369.465 ;
        RECT 557.355 369.185 557.635 369.465 ;
        RECT 558.065 369.185 558.345 369.465 ;
        RECT 558.775 369.185 559.055 369.465 ;
        RECT 559.485 369.185 559.765 369.465 ;
        RECT 560.195 369.185 560.475 369.465 ;
        RECT 550.965 368.475 551.245 368.755 ;
        RECT 551.675 368.475 551.955 368.755 ;
        RECT 552.385 368.475 552.665 368.755 ;
        RECT 553.095 368.475 553.375 368.755 ;
        RECT 553.805 368.475 554.085 368.755 ;
        RECT 554.515 368.475 554.795 368.755 ;
        RECT 555.225 368.475 555.505 368.755 ;
        RECT 555.935 368.475 556.215 368.755 ;
        RECT 556.645 368.475 556.925 368.755 ;
        RECT 557.355 368.475 557.635 368.755 ;
        RECT 558.065 368.475 558.345 368.755 ;
        RECT 558.775 368.475 559.055 368.755 ;
        RECT 559.485 368.475 559.765 368.755 ;
        RECT 560.195 368.475 560.475 368.755 ;
        RECT 550.965 367.765 551.245 368.045 ;
        RECT 551.675 367.765 551.955 368.045 ;
        RECT 552.385 367.765 552.665 368.045 ;
        RECT 553.095 367.765 553.375 368.045 ;
        RECT 553.805 367.765 554.085 368.045 ;
        RECT 554.515 367.765 554.795 368.045 ;
        RECT 555.225 367.765 555.505 368.045 ;
        RECT 555.935 367.765 556.215 368.045 ;
        RECT 556.645 367.765 556.925 368.045 ;
        RECT 557.355 367.765 557.635 368.045 ;
        RECT 558.065 367.765 558.345 368.045 ;
        RECT 558.775 367.765 559.055 368.045 ;
        RECT 559.485 367.765 559.765 368.045 ;
        RECT 560.195 367.765 560.475 368.045 ;
        RECT 550.965 367.055 551.245 367.335 ;
        RECT 551.675 367.055 551.955 367.335 ;
        RECT 552.385 367.055 552.665 367.335 ;
        RECT 553.095 367.055 553.375 367.335 ;
        RECT 553.805 367.055 554.085 367.335 ;
        RECT 554.515 367.055 554.795 367.335 ;
        RECT 555.225 367.055 555.505 367.335 ;
        RECT 555.935 367.055 556.215 367.335 ;
        RECT 556.645 367.055 556.925 367.335 ;
        RECT 557.355 367.055 557.635 367.335 ;
        RECT 558.065 367.055 558.345 367.335 ;
        RECT 558.775 367.055 559.055 367.335 ;
        RECT 559.485 367.055 559.765 367.335 ;
        RECT 560.195 367.055 560.475 367.335 ;
        RECT 550.965 366.345 551.245 366.625 ;
        RECT 551.675 366.345 551.955 366.625 ;
        RECT 552.385 366.345 552.665 366.625 ;
        RECT 553.095 366.345 553.375 366.625 ;
        RECT 553.805 366.345 554.085 366.625 ;
        RECT 554.515 366.345 554.795 366.625 ;
        RECT 555.225 366.345 555.505 366.625 ;
        RECT 555.935 366.345 556.215 366.625 ;
        RECT 556.645 366.345 556.925 366.625 ;
        RECT 557.355 366.345 557.635 366.625 ;
        RECT 558.065 366.345 558.345 366.625 ;
        RECT 558.775 366.345 559.055 366.625 ;
        RECT 559.485 366.345 559.765 366.625 ;
        RECT 560.195 366.345 560.475 366.625 ;
        RECT 550.965 365.635 551.245 365.915 ;
        RECT 551.675 365.635 551.955 365.915 ;
        RECT 552.385 365.635 552.665 365.915 ;
        RECT 553.095 365.635 553.375 365.915 ;
        RECT 553.805 365.635 554.085 365.915 ;
        RECT 554.515 365.635 554.795 365.915 ;
        RECT 555.225 365.635 555.505 365.915 ;
        RECT 555.935 365.635 556.215 365.915 ;
        RECT 556.645 365.635 556.925 365.915 ;
        RECT 557.355 365.635 557.635 365.915 ;
        RECT 558.065 365.635 558.345 365.915 ;
        RECT 558.775 365.635 559.055 365.915 ;
        RECT 559.485 365.635 559.765 365.915 ;
        RECT 560.195 365.635 560.475 365.915 ;
        RECT 550.965 364.925 551.245 365.205 ;
        RECT 551.675 364.925 551.955 365.205 ;
        RECT 552.385 364.925 552.665 365.205 ;
        RECT 553.095 364.925 553.375 365.205 ;
        RECT 553.805 364.925 554.085 365.205 ;
        RECT 554.515 364.925 554.795 365.205 ;
        RECT 555.225 364.925 555.505 365.205 ;
        RECT 555.935 364.925 556.215 365.205 ;
        RECT 556.645 364.925 556.925 365.205 ;
        RECT 557.355 364.925 557.635 365.205 ;
        RECT 558.065 364.925 558.345 365.205 ;
        RECT 558.775 364.925 559.055 365.205 ;
        RECT 559.485 364.925 559.765 365.205 ;
        RECT 560.195 364.925 560.475 365.205 ;
        RECT 550.965 364.215 551.245 364.495 ;
        RECT 551.675 364.215 551.955 364.495 ;
        RECT 552.385 364.215 552.665 364.495 ;
        RECT 553.095 364.215 553.375 364.495 ;
        RECT 553.805 364.215 554.085 364.495 ;
        RECT 554.515 364.215 554.795 364.495 ;
        RECT 555.225 364.215 555.505 364.495 ;
        RECT 555.935 364.215 556.215 364.495 ;
        RECT 556.645 364.215 556.925 364.495 ;
        RECT 557.355 364.215 557.635 364.495 ;
        RECT 558.065 364.215 558.345 364.495 ;
        RECT 558.775 364.215 559.055 364.495 ;
        RECT 559.485 364.215 559.765 364.495 ;
        RECT 560.195 364.215 560.475 364.495 ;
        RECT 550.965 363.505 551.245 363.785 ;
        RECT 551.675 363.505 551.955 363.785 ;
        RECT 552.385 363.505 552.665 363.785 ;
        RECT 553.095 363.505 553.375 363.785 ;
        RECT 553.805 363.505 554.085 363.785 ;
        RECT 554.515 363.505 554.795 363.785 ;
        RECT 555.225 363.505 555.505 363.785 ;
        RECT 555.935 363.505 556.215 363.785 ;
        RECT 556.645 363.505 556.925 363.785 ;
        RECT 557.355 363.505 557.635 363.785 ;
        RECT 558.065 363.505 558.345 363.785 ;
        RECT 558.775 363.505 559.055 363.785 ;
        RECT 559.485 363.505 559.765 363.785 ;
        RECT 560.195 363.505 560.475 363.785 ;
        RECT 550.965 362.795 551.245 363.075 ;
        RECT 551.675 362.795 551.955 363.075 ;
        RECT 552.385 362.795 552.665 363.075 ;
        RECT 553.095 362.795 553.375 363.075 ;
        RECT 553.805 362.795 554.085 363.075 ;
        RECT 554.515 362.795 554.795 363.075 ;
        RECT 555.225 362.795 555.505 363.075 ;
        RECT 555.935 362.795 556.215 363.075 ;
        RECT 556.645 362.795 556.925 363.075 ;
        RECT 557.355 362.795 557.635 363.075 ;
        RECT 558.065 362.795 558.345 363.075 ;
        RECT 558.775 362.795 559.055 363.075 ;
        RECT 559.485 362.795 559.765 363.075 ;
        RECT 560.195 362.795 560.475 363.075 ;
        RECT 550.965 362.085 551.245 362.365 ;
        RECT 551.675 362.085 551.955 362.365 ;
        RECT 552.385 362.085 552.665 362.365 ;
        RECT 553.095 362.085 553.375 362.365 ;
        RECT 553.805 362.085 554.085 362.365 ;
        RECT 554.515 362.085 554.795 362.365 ;
        RECT 555.225 362.085 555.505 362.365 ;
        RECT 555.935 362.085 556.215 362.365 ;
        RECT 556.645 362.085 556.925 362.365 ;
        RECT 557.355 362.085 557.635 362.365 ;
        RECT 558.065 362.085 558.345 362.365 ;
        RECT 558.775 362.085 559.055 362.365 ;
        RECT 559.485 362.085 559.765 362.365 ;
        RECT 560.195 362.085 560.475 362.365 ;
        RECT 550.965 361.375 551.245 361.655 ;
        RECT 551.675 361.375 551.955 361.655 ;
        RECT 552.385 361.375 552.665 361.655 ;
        RECT 553.095 361.375 553.375 361.655 ;
        RECT 553.805 361.375 554.085 361.655 ;
        RECT 554.515 361.375 554.795 361.655 ;
        RECT 555.225 361.375 555.505 361.655 ;
        RECT 555.935 361.375 556.215 361.655 ;
        RECT 556.645 361.375 556.925 361.655 ;
        RECT 557.355 361.375 557.635 361.655 ;
        RECT 558.065 361.375 558.345 361.655 ;
        RECT 558.775 361.375 559.055 361.655 ;
        RECT 559.485 361.375 559.765 361.655 ;
        RECT 560.195 361.375 560.475 361.655 ;
        RECT 550.965 360.665 551.245 360.945 ;
        RECT 551.675 360.665 551.955 360.945 ;
        RECT 552.385 360.665 552.665 360.945 ;
        RECT 553.095 360.665 553.375 360.945 ;
        RECT 553.805 360.665 554.085 360.945 ;
        RECT 554.515 360.665 554.795 360.945 ;
        RECT 555.225 360.665 555.505 360.945 ;
        RECT 555.935 360.665 556.215 360.945 ;
        RECT 556.645 360.665 556.925 360.945 ;
        RECT 557.355 360.665 557.635 360.945 ;
        RECT 558.065 360.665 558.345 360.945 ;
        RECT 558.775 360.665 559.055 360.945 ;
        RECT 559.485 360.665 559.765 360.945 ;
        RECT 560.195 360.665 560.475 360.945 ;
        RECT 566.625 369.895 566.905 370.175 ;
        RECT 567.335 369.895 567.615 370.175 ;
        RECT 568.045 369.895 568.325 370.175 ;
        RECT 568.755 369.895 569.035 370.175 ;
        RECT 569.465 369.895 569.745 370.175 ;
        RECT 570.175 369.895 570.455 370.175 ;
        RECT 570.885 369.895 571.165 370.175 ;
        RECT 571.595 369.895 571.875 370.175 ;
        RECT 572.305 369.895 572.585 370.175 ;
        RECT 573.015 369.895 573.295 370.175 ;
        RECT 573.725 369.895 574.005 370.175 ;
        RECT 566.625 369.185 566.905 369.465 ;
        RECT 567.335 369.185 567.615 369.465 ;
        RECT 568.045 369.185 568.325 369.465 ;
        RECT 568.755 369.185 569.035 369.465 ;
        RECT 569.465 369.185 569.745 369.465 ;
        RECT 570.175 369.185 570.455 369.465 ;
        RECT 570.885 369.185 571.165 369.465 ;
        RECT 571.595 369.185 571.875 369.465 ;
        RECT 572.305 369.185 572.585 369.465 ;
        RECT 573.015 369.185 573.295 369.465 ;
        RECT 573.725 369.185 574.005 369.465 ;
        RECT 566.625 368.475 566.905 368.755 ;
        RECT 567.335 368.475 567.615 368.755 ;
        RECT 568.045 368.475 568.325 368.755 ;
        RECT 568.755 368.475 569.035 368.755 ;
        RECT 569.465 368.475 569.745 368.755 ;
        RECT 570.175 368.475 570.455 368.755 ;
        RECT 570.885 368.475 571.165 368.755 ;
        RECT 571.595 368.475 571.875 368.755 ;
        RECT 572.305 368.475 572.585 368.755 ;
        RECT 573.015 368.475 573.295 368.755 ;
        RECT 573.725 368.475 574.005 368.755 ;
        RECT 566.625 367.765 566.905 368.045 ;
        RECT 567.335 367.765 567.615 368.045 ;
        RECT 568.045 367.765 568.325 368.045 ;
        RECT 568.755 367.765 569.035 368.045 ;
        RECT 569.465 367.765 569.745 368.045 ;
        RECT 570.175 367.765 570.455 368.045 ;
        RECT 570.885 367.765 571.165 368.045 ;
        RECT 571.595 367.765 571.875 368.045 ;
        RECT 572.305 367.765 572.585 368.045 ;
        RECT 573.015 367.765 573.295 368.045 ;
        RECT 573.725 367.765 574.005 368.045 ;
        RECT 566.625 367.055 566.905 367.335 ;
        RECT 567.335 367.055 567.615 367.335 ;
        RECT 568.045 367.055 568.325 367.335 ;
        RECT 568.755 367.055 569.035 367.335 ;
        RECT 569.465 367.055 569.745 367.335 ;
        RECT 570.175 367.055 570.455 367.335 ;
        RECT 570.885 367.055 571.165 367.335 ;
        RECT 571.595 367.055 571.875 367.335 ;
        RECT 572.305 367.055 572.585 367.335 ;
        RECT 573.015 367.055 573.295 367.335 ;
        RECT 573.725 367.055 574.005 367.335 ;
        RECT 566.625 366.345 566.905 366.625 ;
        RECT 567.335 366.345 567.615 366.625 ;
        RECT 568.045 366.345 568.325 366.625 ;
        RECT 568.755 366.345 569.035 366.625 ;
        RECT 569.465 366.345 569.745 366.625 ;
        RECT 570.175 366.345 570.455 366.625 ;
        RECT 570.885 366.345 571.165 366.625 ;
        RECT 571.595 366.345 571.875 366.625 ;
        RECT 572.305 366.345 572.585 366.625 ;
        RECT 573.015 366.345 573.295 366.625 ;
        RECT 573.725 366.345 574.005 366.625 ;
        RECT 566.625 365.635 566.905 365.915 ;
        RECT 567.335 365.635 567.615 365.915 ;
        RECT 568.045 365.635 568.325 365.915 ;
        RECT 568.755 365.635 569.035 365.915 ;
        RECT 569.465 365.635 569.745 365.915 ;
        RECT 570.175 365.635 570.455 365.915 ;
        RECT 570.885 365.635 571.165 365.915 ;
        RECT 571.595 365.635 571.875 365.915 ;
        RECT 572.305 365.635 572.585 365.915 ;
        RECT 573.015 365.635 573.295 365.915 ;
        RECT 573.725 365.635 574.005 365.915 ;
        RECT 566.625 364.925 566.905 365.205 ;
        RECT 567.335 364.925 567.615 365.205 ;
        RECT 568.045 364.925 568.325 365.205 ;
        RECT 568.755 364.925 569.035 365.205 ;
        RECT 569.465 364.925 569.745 365.205 ;
        RECT 570.175 364.925 570.455 365.205 ;
        RECT 570.885 364.925 571.165 365.205 ;
        RECT 571.595 364.925 571.875 365.205 ;
        RECT 572.305 364.925 572.585 365.205 ;
        RECT 573.015 364.925 573.295 365.205 ;
        RECT 573.725 364.925 574.005 365.205 ;
        RECT 566.625 364.215 566.905 364.495 ;
        RECT 567.335 364.215 567.615 364.495 ;
        RECT 568.045 364.215 568.325 364.495 ;
        RECT 568.755 364.215 569.035 364.495 ;
        RECT 569.465 364.215 569.745 364.495 ;
        RECT 570.175 364.215 570.455 364.495 ;
        RECT 570.885 364.215 571.165 364.495 ;
        RECT 571.595 364.215 571.875 364.495 ;
        RECT 572.305 364.215 572.585 364.495 ;
        RECT 573.015 364.215 573.295 364.495 ;
        RECT 573.725 364.215 574.005 364.495 ;
        RECT 566.625 363.505 566.905 363.785 ;
        RECT 567.335 363.505 567.615 363.785 ;
        RECT 568.045 363.505 568.325 363.785 ;
        RECT 568.755 363.505 569.035 363.785 ;
        RECT 569.465 363.505 569.745 363.785 ;
        RECT 570.175 363.505 570.455 363.785 ;
        RECT 570.885 363.505 571.165 363.785 ;
        RECT 571.595 363.505 571.875 363.785 ;
        RECT 572.305 363.505 572.585 363.785 ;
        RECT 573.015 363.505 573.295 363.785 ;
        RECT 573.725 363.505 574.005 363.785 ;
        RECT 566.625 362.795 566.905 363.075 ;
        RECT 567.335 362.795 567.615 363.075 ;
        RECT 568.045 362.795 568.325 363.075 ;
        RECT 568.755 362.795 569.035 363.075 ;
        RECT 569.465 362.795 569.745 363.075 ;
        RECT 570.175 362.795 570.455 363.075 ;
        RECT 570.885 362.795 571.165 363.075 ;
        RECT 571.595 362.795 571.875 363.075 ;
        RECT 572.305 362.795 572.585 363.075 ;
        RECT 573.015 362.795 573.295 363.075 ;
        RECT 573.725 362.795 574.005 363.075 ;
        RECT 566.625 362.085 566.905 362.365 ;
        RECT 567.335 362.085 567.615 362.365 ;
        RECT 568.045 362.085 568.325 362.365 ;
        RECT 568.755 362.085 569.035 362.365 ;
        RECT 569.465 362.085 569.745 362.365 ;
        RECT 570.175 362.085 570.455 362.365 ;
        RECT 570.885 362.085 571.165 362.365 ;
        RECT 571.595 362.085 571.875 362.365 ;
        RECT 572.305 362.085 572.585 362.365 ;
        RECT 573.015 362.085 573.295 362.365 ;
        RECT 573.725 362.085 574.005 362.365 ;
        RECT 566.625 361.375 566.905 361.655 ;
        RECT 567.335 361.375 567.615 361.655 ;
        RECT 568.045 361.375 568.325 361.655 ;
        RECT 568.755 361.375 569.035 361.655 ;
        RECT 569.465 361.375 569.745 361.655 ;
        RECT 570.175 361.375 570.455 361.655 ;
        RECT 570.885 361.375 571.165 361.655 ;
        RECT 571.595 361.375 571.875 361.655 ;
        RECT 572.305 361.375 572.585 361.655 ;
        RECT 573.015 361.375 573.295 361.655 ;
        RECT 573.725 361.375 574.005 361.655 ;
        RECT 566.625 360.665 566.905 360.945 ;
        RECT 567.335 360.665 567.615 360.945 ;
        RECT 568.045 360.665 568.325 360.945 ;
        RECT 568.755 360.665 569.035 360.945 ;
        RECT 569.465 360.665 569.745 360.945 ;
        RECT 570.175 360.665 570.455 360.945 ;
        RECT 570.885 360.665 571.165 360.945 ;
        RECT 571.595 360.665 571.875 360.945 ;
        RECT 572.305 360.665 572.585 360.945 ;
        RECT 573.015 360.665 573.295 360.945 ;
        RECT 573.725 360.665 574.005 360.945 ;
        RECT 576.345 369.895 576.625 370.175 ;
        RECT 577.055 369.895 577.335 370.175 ;
        RECT 577.765 369.895 578.045 370.175 ;
        RECT 578.475 369.895 578.755 370.175 ;
        RECT 579.185 369.895 579.465 370.175 ;
        RECT 579.895 369.895 580.175 370.175 ;
        RECT 580.605 369.895 580.885 370.175 ;
        RECT 581.315 369.895 581.595 370.175 ;
        RECT 582.025 369.895 582.305 370.175 ;
        RECT 582.735 369.895 583.015 370.175 ;
        RECT 583.445 369.895 583.725 370.175 ;
        RECT 584.155 369.895 584.435 370.175 ;
        RECT 584.865 369.895 585.145 370.175 ;
        RECT 585.575 369.895 585.855 370.175 ;
        RECT 576.345 369.185 576.625 369.465 ;
        RECT 577.055 369.185 577.335 369.465 ;
        RECT 577.765 369.185 578.045 369.465 ;
        RECT 578.475 369.185 578.755 369.465 ;
        RECT 579.185 369.185 579.465 369.465 ;
        RECT 579.895 369.185 580.175 369.465 ;
        RECT 580.605 369.185 580.885 369.465 ;
        RECT 581.315 369.185 581.595 369.465 ;
        RECT 582.025 369.185 582.305 369.465 ;
        RECT 582.735 369.185 583.015 369.465 ;
        RECT 583.445 369.185 583.725 369.465 ;
        RECT 584.155 369.185 584.435 369.465 ;
        RECT 584.865 369.185 585.145 369.465 ;
        RECT 585.575 369.185 585.855 369.465 ;
        RECT 576.345 368.475 576.625 368.755 ;
        RECT 577.055 368.475 577.335 368.755 ;
        RECT 577.765 368.475 578.045 368.755 ;
        RECT 578.475 368.475 578.755 368.755 ;
        RECT 579.185 368.475 579.465 368.755 ;
        RECT 579.895 368.475 580.175 368.755 ;
        RECT 580.605 368.475 580.885 368.755 ;
        RECT 581.315 368.475 581.595 368.755 ;
        RECT 582.025 368.475 582.305 368.755 ;
        RECT 582.735 368.475 583.015 368.755 ;
        RECT 583.445 368.475 583.725 368.755 ;
        RECT 584.155 368.475 584.435 368.755 ;
        RECT 584.865 368.475 585.145 368.755 ;
        RECT 585.575 368.475 585.855 368.755 ;
        RECT 576.345 367.765 576.625 368.045 ;
        RECT 577.055 367.765 577.335 368.045 ;
        RECT 577.765 367.765 578.045 368.045 ;
        RECT 578.475 367.765 578.755 368.045 ;
        RECT 579.185 367.765 579.465 368.045 ;
        RECT 579.895 367.765 580.175 368.045 ;
        RECT 580.605 367.765 580.885 368.045 ;
        RECT 581.315 367.765 581.595 368.045 ;
        RECT 582.025 367.765 582.305 368.045 ;
        RECT 582.735 367.765 583.015 368.045 ;
        RECT 583.445 367.765 583.725 368.045 ;
        RECT 584.155 367.765 584.435 368.045 ;
        RECT 584.865 367.765 585.145 368.045 ;
        RECT 585.575 367.765 585.855 368.045 ;
        RECT 576.345 367.055 576.625 367.335 ;
        RECT 577.055 367.055 577.335 367.335 ;
        RECT 577.765 367.055 578.045 367.335 ;
        RECT 578.475 367.055 578.755 367.335 ;
        RECT 579.185 367.055 579.465 367.335 ;
        RECT 579.895 367.055 580.175 367.335 ;
        RECT 580.605 367.055 580.885 367.335 ;
        RECT 581.315 367.055 581.595 367.335 ;
        RECT 582.025 367.055 582.305 367.335 ;
        RECT 582.735 367.055 583.015 367.335 ;
        RECT 583.445 367.055 583.725 367.335 ;
        RECT 584.155 367.055 584.435 367.335 ;
        RECT 584.865 367.055 585.145 367.335 ;
        RECT 585.575 367.055 585.855 367.335 ;
        RECT 576.345 366.345 576.625 366.625 ;
        RECT 577.055 366.345 577.335 366.625 ;
        RECT 577.765 366.345 578.045 366.625 ;
        RECT 578.475 366.345 578.755 366.625 ;
        RECT 579.185 366.345 579.465 366.625 ;
        RECT 579.895 366.345 580.175 366.625 ;
        RECT 580.605 366.345 580.885 366.625 ;
        RECT 581.315 366.345 581.595 366.625 ;
        RECT 582.025 366.345 582.305 366.625 ;
        RECT 582.735 366.345 583.015 366.625 ;
        RECT 583.445 366.345 583.725 366.625 ;
        RECT 584.155 366.345 584.435 366.625 ;
        RECT 584.865 366.345 585.145 366.625 ;
        RECT 585.575 366.345 585.855 366.625 ;
        RECT 576.345 365.635 576.625 365.915 ;
        RECT 577.055 365.635 577.335 365.915 ;
        RECT 577.765 365.635 578.045 365.915 ;
        RECT 578.475 365.635 578.755 365.915 ;
        RECT 579.185 365.635 579.465 365.915 ;
        RECT 579.895 365.635 580.175 365.915 ;
        RECT 580.605 365.635 580.885 365.915 ;
        RECT 581.315 365.635 581.595 365.915 ;
        RECT 582.025 365.635 582.305 365.915 ;
        RECT 582.735 365.635 583.015 365.915 ;
        RECT 583.445 365.635 583.725 365.915 ;
        RECT 584.155 365.635 584.435 365.915 ;
        RECT 584.865 365.635 585.145 365.915 ;
        RECT 585.575 365.635 585.855 365.915 ;
        RECT 576.345 364.925 576.625 365.205 ;
        RECT 577.055 364.925 577.335 365.205 ;
        RECT 577.765 364.925 578.045 365.205 ;
        RECT 578.475 364.925 578.755 365.205 ;
        RECT 579.185 364.925 579.465 365.205 ;
        RECT 579.895 364.925 580.175 365.205 ;
        RECT 580.605 364.925 580.885 365.205 ;
        RECT 581.315 364.925 581.595 365.205 ;
        RECT 582.025 364.925 582.305 365.205 ;
        RECT 582.735 364.925 583.015 365.205 ;
        RECT 583.445 364.925 583.725 365.205 ;
        RECT 584.155 364.925 584.435 365.205 ;
        RECT 584.865 364.925 585.145 365.205 ;
        RECT 585.575 364.925 585.855 365.205 ;
        RECT 576.345 364.215 576.625 364.495 ;
        RECT 577.055 364.215 577.335 364.495 ;
        RECT 577.765 364.215 578.045 364.495 ;
        RECT 578.475 364.215 578.755 364.495 ;
        RECT 579.185 364.215 579.465 364.495 ;
        RECT 579.895 364.215 580.175 364.495 ;
        RECT 580.605 364.215 580.885 364.495 ;
        RECT 581.315 364.215 581.595 364.495 ;
        RECT 582.025 364.215 582.305 364.495 ;
        RECT 582.735 364.215 583.015 364.495 ;
        RECT 583.445 364.215 583.725 364.495 ;
        RECT 584.155 364.215 584.435 364.495 ;
        RECT 584.865 364.215 585.145 364.495 ;
        RECT 585.575 364.215 585.855 364.495 ;
        RECT 576.345 363.505 576.625 363.785 ;
        RECT 577.055 363.505 577.335 363.785 ;
        RECT 577.765 363.505 578.045 363.785 ;
        RECT 578.475 363.505 578.755 363.785 ;
        RECT 579.185 363.505 579.465 363.785 ;
        RECT 579.895 363.505 580.175 363.785 ;
        RECT 580.605 363.505 580.885 363.785 ;
        RECT 581.315 363.505 581.595 363.785 ;
        RECT 582.025 363.505 582.305 363.785 ;
        RECT 582.735 363.505 583.015 363.785 ;
        RECT 583.445 363.505 583.725 363.785 ;
        RECT 584.155 363.505 584.435 363.785 ;
        RECT 584.865 363.505 585.145 363.785 ;
        RECT 585.575 363.505 585.855 363.785 ;
        RECT 576.345 362.795 576.625 363.075 ;
        RECT 577.055 362.795 577.335 363.075 ;
        RECT 577.765 362.795 578.045 363.075 ;
        RECT 578.475 362.795 578.755 363.075 ;
        RECT 579.185 362.795 579.465 363.075 ;
        RECT 579.895 362.795 580.175 363.075 ;
        RECT 580.605 362.795 580.885 363.075 ;
        RECT 581.315 362.795 581.595 363.075 ;
        RECT 582.025 362.795 582.305 363.075 ;
        RECT 582.735 362.795 583.015 363.075 ;
        RECT 583.445 362.795 583.725 363.075 ;
        RECT 584.155 362.795 584.435 363.075 ;
        RECT 584.865 362.795 585.145 363.075 ;
        RECT 585.575 362.795 585.855 363.075 ;
        RECT 576.345 362.085 576.625 362.365 ;
        RECT 577.055 362.085 577.335 362.365 ;
        RECT 577.765 362.085 578.045 362.365 ;
        RECT 578.475 362.085 578.755 362.365 ;
        RECT 579.185 362.085 579.465 362.365 ;
        RECT 579.895 362.085 580.175 362.365 ;
        RECT 580.605 362.085 580.885 362.365 ;
        RECT 581.315 362.085 581.595 362.365 ;
        RECT 582.025 362.085 582.305 362.365 ;
        RECT 582.735 362.085 583.015 362.365 ;
        RECT 583.445 362.085 583.725 362.365 ;
        RECT 584.155 362.085 584.435 362.365 ;
        RECT 584.865 362.085 585.145 362.365 ;
        RECT 585.575 362.085 585.855 362.365 ;
        RECT 576.345 361.375 576.625 361.655 ;
        RECT 577.055 361.375 577.335 361.655 ;
        RECT 577.765 361.375 578.045 361.655 ;
        RECT 578.475 361.375 578.755 361.655 ;
        RECT 579.185 361.375 579.465 361.655 ;
        RECT 579.895 361.375 580.175 361.655 ;
        RECT 580.605 361.375 580.885 361.655 ;
        RECT 581.315 361.375 581.595 361.655 ;
        RECT 582.025 361.375 582.305 361.655 ;
        RECT 582.735 361.375 583.015 361.655 ;
        RECT 583.445 361.375 583.725 361.655 ;
        RECT 584.155 361.375 584.435 361.655 ;
        RECT 584.865 361.375 585.145 361.655 ;
        RECT 585.575 361.375 585.855 361.655 ;
        RECT 576.345 360.665 576.625 360.945 ;
        RECT 577.055 360.665 577.335 360.945 ;
        RECT 577.765 360.665 578.045 360.945 ;
        RECT 578.475 360.665 578.755 360.945 ;
        RECT 579.185 360.665 579.465 360.945 ;
        RECT 579.895 360.665 580.175 360.945 ;
        RECT 580.605 360.665 580.885 360.945 ;
        RECT 581.315 360.665 581.595 360.945 ;
        RECT 582.025 360.665 582.305 360.945 ;
        RECT 582.735 360.665 583.015 360.945 ;
        RECT 583.445 360.665 583.725 360.945 ;
        RECT 584.155 360.665 584.435 360.945 ;
        RECT 584.865 360.665 585.145 360.945 ;
        RECT 585.575 360.665 585.855 360.945 ;
        RECT 589.495 369.895 589.775 370.175 ;
        RECT 590.205 369.895 590.485 370.175 ;
        RECT 590.915 369.895 591.195 370.175 ;
        RECT 591.625 369.895 591.905 370.175 ;
        RECT 592.335 369.895 592.615 370.175 ;
        RECT 593.045 369.895 593.325 370.175 ;
        RECT 593.755 369.895 594.035 370.175 ;
        RECT 594.465 369.895 594.745 370.175 ;
        RECT 595.175 369.895 595.455 370.175 ;
        RECT 595.885 369.895 596.165 370.175 ;
        RECT 596.595 369.895 596.875 370.175 ;
        RECT 597.305 369.895 597.585 370.175 ;
        RECT 598.015 369.895 598.295 370.175 ;
        RECT 589.495 369.185 589.775 369.465 ;
        RECT 590.205 369.185 590.485 369.465 ;
        RECT 590.915 369.185 591.195 369.465 ;
        RECT 591.625 369.185 591.905 369.465 ;
        RECT 592.335 369.185 592.615 369.465 ;
        RECT 593.045 369.185 593.325 369.465 ;
        RECT 593.755 369.185 594.035 369.465 ;
        RECT 594.465 369.185 594.745 369.465 ;
        RECT 595.175 369.185 595.455 369.465 ;
        RECT 595.885 369.185 596.165 369.465 ;
        RECT 596.595 369.185 596.875 369.465 ;
        RECT 597.305 369.185 597.585 369.465 ;
        RECT 598.015 369.185 598.295 369.465 ;
        RECT 589.495 368.475 589.775 368.755 ;
        RECT 590.205 368.475 590.485 368.755 ;
        RECT 590.915 368.475 591.195 368.755 ;
        RECT 591.625 368.475 591.905 368.755 ;
        RECT 592.335 368.475 592.615 368.755 ;
        RECT 593.045 368.475 593.325 368.755 ;
        RECT 593.755 368.475 594.035 368.755 ;
        RECT 594.465 368.475 594.745 368.755 ;
        RECT 595.175 368.475 595.455 368.755 ;
        RECT 595.885 368.475 596.165 368.755 ;
        RECT 596.595 368.475 596.875 368.755 ;
        RECT 597.305 368.475 597.585 368.755 ;
        RECT 598.015 368.475 598.295 368.755 ;
        RECT 589.495 367.765 589.775 368.045 ;
        RECT 590.205 367.765 590.485 368.045 ;
        RECT 590.915 367.765 591.195 368.045 ;
        RECT 591.625 367.765 591.905 368.045 ;
        RECT 592.335 367.765 592.615 368.045 ;
        RECT 593.045 367.765 593.325 368.045 ;
        RECT 593.755 367.765 594.035 368.045 ;
        RECT 594.465 367.765 594.745 368.045 ;
        RECT 595.175 367.765 595.455 368.045 ;
        RECT 595.885 367.765 596.165 368.045 ;
        RECT 596.595 367.765 596.875 368.045 ;
        RECT 597.305 367.765 597.585 368.045 ;
        RECT 598.015 367.765 598.295 368.045 ;
        RECT 589.495 367.055 589.775 367.335 ;
        RECT 590.205 367.055 590.485 367.335 ;
        RECT 590.915 367.055 591.195 367.335 ;
        RECT 591.625 367.055 591.905 367.335 ;
        RECT 592.335 367.055 592.615 367.335 ;
        RECT 593.045 367.055 593.325 367.335 ;
        RECT 593.755 367.055 594.035 367.335 ;
        RECT 594.465 367.055 594.745 367.335 ;
        RECT 595.175 367.055 595.455 367.335 ;
        RECT 595.885 367.055 596.165 367.335 ;
        RECT 596.595 367.055 596.875 367.335 ;
        RECT 597.305 367.055 597.585 367.335 ;
        RECT 598.015 367.055 598.295 367.335 ;
        RECT 589.495 366.345 589.775 366.625 ;
        RECT 590.205 366.345 590.485 366.625 ;
        RECT 590.915 366.345 591.195 366.625 ;
        RECT 591.625 366.345 591.905 366.625 ;
        RECT 592.335 366.345 592.615 366.625 ;
        RECT 593.045 366.345 593.325 366.625 ;
        RECT 593.755 366.345 594.035 366.625 ;
        RECT 594.465 366.345 594.745 366.625 ;
        RECT 595.175 366.345 595.455 366.625 ;
        RECT 595.885 366.345 596.165 366.625 ;
        RECT 596.595 366.345 596.875 366.625 ;
        RECT 597.305 366.345 597.585 366.625 ;
        RECT 598.015 366.345 598.295 366.625 ;
        RECT 589.495 365.635 589.775 365.915 ;
        RECT 590.205 365.635 590.485 365.915 ;
        RECT 590.915 365.635 591.195 365.915 ;
        RECT 591.625 365.635 591.905 365.915 ;
        RECT 592.335 365.635 592.615 365.915 ;
        RECT 593.045 365.635 593.325 365.915 ;
        RECT 593.755 365.635 594.035 365.915 ;
        RECT 594.465 365.635 594.745 365.915 ;
        RECT 595.175 365.635 595.455 365.915 ;
        RECT 595.885 365.635 596.165 365.915 ;
        RECT 596.595 365.635 596.875 365.915 ;
        RECT 597.305 365.635 597.585 365.915 ;
        RECT 598.015 365.635 598.295 365.915 ;
        RECT 589.495 364.925 589.775 365.205 ;
        RECT 590.205 364.925 590.485 365.205 ;
        RECT 590.915 364.925 591.195 365.205 ;
        RECT 591.625 364.925 591.905 365.205 ;
        RECT 592.335 364.925 592.615 365.205 ;
        RECT 593.045 364.925 593.325 365.205 ;
        RECT 593.755 364.925 594.035 365.205 ;
        RECT 594.465 364.925 594.745 365.205 ;
        RECT 595.175 364.925 595.455 365.205 ;
        RECT 595.885 364.925 596.165 365.205 ;
        RECT 596.595 364.925 596.875 365.205 ;
        RECT 597.305 364.925 597.585 365.205 ;
        RECT 598.015 364.925 598.295 365.205 ;
        RECT 589.495 364.215 589.775 364.495 ;
        RECT 590.205 364.215 590.485 364.495 ;
        RECT 590.915 364.215 591.195 364.495 ;
        RECT 591.625 364.215 591.905 364.495 ;
        RECT 592.335 364.215 592.615 364.495 ;
        RECT 593.045 364.215 593.325 364.495 ;
        RECT 593.755 364.215 594.035 364.495 ;
        RECT 594.465 364.215 594.745 364.495 ;
        RECT 595.175 364.215 595.455 364.495 ;
        RECT 595.885 364.215 596.165 364.495 ;
        RECT 596.595 364.215 596.875 364.495 ;
        RECT 597.305 364.215 597.585 364.495 ;
        RECT 598.015 364.215 598.295 364.495 ;
        RECT 589.495 363.505 589.775 363.785 ;
        RECT 590.205 363.505 590.485 363.785 ;
        RECT 590.915 363.505 591.195 363.785 ;
        RECT 591.625 363.505 591.905 363.785 ;
        RECT 592.335 363.505 592.615 363.785 ;
        RECT 593.045 363.505 593.325 363.785 ;
        RECT 593.755 363.505 594.035 363.785 ;
        RECT 594.465 363.505 594.745 363.785 ;
        RECT 595.175 363.505 595.455 363.785 ;
        RECT 595.885 363.505 596.165 363.785 ;
        RECT 596.595 363.505 596.875 363.785 ;
        RECT 597.305 363.505 597.585 363.785 ;
        RECT 598.015 363.505 598.295 363.785 ;
        RECT 589.495 362.795 589.775 363.075 ;
        RECT 590.205 362.795 590.485 363.075 ;
        RECT 590.915 362.795 591.195 363.075 ;
        RECT 591.625 362.795 591.905 363.075 ;
        RECT 592.335 362.795 592.615 363.075 ;
        RECT 593.045 362.795 593.325 363.075 ;
        RECT 593.755 362.795 594.035 363.075 ;
        RECT 594.465 362.795 594.745 363.075 ;
        RECT 595.175 362.795 595.455 363.075 ;
        RECT 595.885 362.795 596.165 363.075 ;
        RECT 596.595 362.795 596.875 363.075 ;
        RECT 597.305 362.795 597.585 363.075 ;
        RECT 598.015 362.795 598.295 363.075 ;
        RECT 589.495 362.085 589.775 362.365 ;
        RECT 590.205 362.085 590.485 362.365 ;
        RECT 590.915 362.085 591.195 362.365 ;
        RECT 591.625 362.085 591.905 362.365 ;
        RECT 592.335 362.085 592.615 362.365 ;
        RECT 593.045 362.085 593.325 362.365 ;
        RECT 593.755 362.085 594.035 362.365 ;
        RECT 594.465 362.085 594.745 362.365 ;
        RECT 595.175 362.085 595.455 362.365 ;
        RECT 595.885 362.085 596.165 362.365 ;
        RECT 596.595 362.085 596.875 362.365 ;
        RECT 597.305 362.085 597.585 362.365 ;
        RECT 598.015 362.085 598.295 362.365 ;
        RECT 589.495 361.375 589.775 361.655 ;
        RECT 590.205 361.375 590.485 361.655 ;
        RECT 590.915 361.375 591.195 361.655 ;
        RECT 591.625 361.375 591.905 361.655 ;
        RECT 592.335 361.375 592.615 361.655 ;
        RECT 593.045 361.375 593.325 361.655 ;
        RECT 593.755 361.375 594.035 361.655 ;
        RECT 594.465 361.375 594.745 361.655 ;
        RECT 595.175 361.375 595.455 361.655 ;
        RECT 595.885 361.375 596.165 361.655 ;
        RECT 596.595 361.375 596.875 361.655 ;
        RECT 597.305 361.375 597.585 361.655 ;
        RECT 598.015 361.375 598.295 361.655 ;
        RECT 589.495 360.665 589.775 360.945 ;
        RECT 590.205 360.665 590.485 360.945 ;
        RECT 590.915 360.665 591.195 360.945 ;
        RECT 591.625 360.665 591.905 360.945 ;
        RECT 592.335 360.665 592.615 360.945 ;
        RECT 593.045 360.665 593.325 360.945 ;
        RECT 593.755 360.665 594.035 360.945 ;
        RECT 594.465 360.665 594.745 360.945 ;
        RECT 595.175 360.665 595.455 360.945 ;
        RECT 595.885 360.665 596.165 360.945 ;
        RECT 596.595 360.665 596.875 360.945 ;
        RECT 597.305 360.665 597.585 360.945 ;
        RECT 598.015 360.665 598.295 360.945 ;
        RECT 1351.715 369.895 1351.995 370.175 ;
        RECT 1352.425 369.895 1352.705 370.175 ;
        RECT 1353.135 369.895 1353.415 370.175 ;
        RECT 1353.845 369.895 1354.125 370.175 ;
        RECT 1354.555 369.895 1354.835 370.175 ;
        RECT 1355.265 369.895 1355.545 370.175 ;
        RECT 1355.975 369.895 1356.255 370.175 ;
        RECT 1356.685 369.895 1356.965 370.175 ;
        RECT 1357.395 369.895 1357.675 370.175 ;
        RECT 1358.105 369.895 1358.385 370.175 ;
        RECT 1358.815 369.895 1359.095 370.175 ;
        RECT 1359.525 369.895 1359.805 370.175 ;
        RECT 1360.235 369.895 1360.515 370.175 ;
        RECT 1351.715 369.185 1351.995 369.465 ;
        RECT 1352.425 369.185 1352.705 369.465 ;
        RECT 1353.135 369.185 1353.415 369.465 ;
        RECT 1353.845 369.185 1354.125 369.465 ;
        RECT 1354.555 369.185 1354.835 369.465 ;
        RECT 1355.265 369.185 1355.545 369.465 ;
        RECT 1355.975 369.185 1356.255 369.465 ;
        RECT 1356.685 369.185 1356.965 369.465 ;
        RECT 1357.395 369.185 1357.675 369.465 ;
        RECT 1358.105 369.185 1358.385 369.465 ;
        RECT 1358.815 369.185 1359.095 369.465 ;
        RECT 1359.525 369.185 1359.805 369.465 ;
        RECT 1360.235 369.185 1360.515 369.465 ;
        RECT 1351.715 368.475 1351.995 368.755 ;
        RECT 1352.425 368.475 1352.705 368.755 ;
        RECT 1353.135 368.475 1353.415 368.755 ;
        RECT 1353.845 368.475 1354.125 368.755 ;
        RECT 1354.555 368.475 1354.835 368.755 ;
        RECT 1355.265 368.475 1355.545 368.755 ;
        RECT 1355.975 368.475 1356.255 368.755 ;
        RECT 1356.685 368.475 1356.965 368.755 ;
        RECT 1357.395 368.475 1357.675 368.755 ;
        RECT 1358.105 368.475 1358.385 368.755 ;
        RECT 1358.815 368.475 1359.095 368.755 ;
        RECT 1359.525 368.475 1359.805 368.755 ;
        RECT 1360.235 368.475 1360.515 368.755 ;
        RECT 1351.715 367.765 1351.995 368.045 ;
        RECT 1352.425 367.765 1352.705 368.045 ;
        RECT 1353.135 367.765 1353.415 368.045 ;
        RECT 1353.845 367.765 1354.125 368.045 ;
        RECT 1354.555 367.765 1354.835 368.045 ;
        RECT 1355.265 367.765 1355.545 368.045 ;
        RECT 1355.975 367.765 1356.255 368.045 ;
        RECT 1356.685 367.765 1356.965 368.045 ;
        RECT 1357.395 367.765 1357.675 368.045 ;
        RECT 1358.105 367.765 1358.385 368.045 ;
        RECT 1358.815 367.765 1359.095 368.045 ;
        RECT 1359.525 367.765 1359.805 368.045 ;
        RECT 1360.235 367.765 1360.515 368.045 ;
        RECT 1351.715 367.055 1351.995 367.335 ;
        RECT 1352.425 367.055 1352.705 367.335 ;
        RECT 1353.135 367.055 1353.415 367.335 ;
        RECT 1353.845 367.055 1354.125 367.335 ;
        RECT 1354.555 367.055 1354.835 367.335 ;
        RECT 1355.265 367.055 1355.545 367.335 ;
        RECT 1355.975 367.055 1356.255 367.335 ;
        RECT 1356.685 367.055 1356.965 367.335 ;
        RECT 1357.395 367.055 1357.675 367.335 ;
        RECT 1358.105 367.055 1358.385 367.335 ;
        RECT 1358.815 367.055 1359.095 367.335 ;
        RECT 1359.525 367.055 1359.805 367.335 ;
        RECT 1360.235 367.055 1360.515 367.335 ;
        RECT 1351.715 366.345 1351.995 366.625 ;
        RECT 1352.425 366.345 1352.705 366.625 ;
        RECT 1353.135 366.345 1353.415 366.625 ;
        RECT 1353.845 366.345 1354.125 366.625 ;
        RECT 1354.555 366.345 1354.835 366.625 ;
        RECT 1355.265 366.345 1355.545 366.625 ;
        RECT 1355.975 366.345 1356.255 366.625 ;
        RECT 1356.685 366.345 1356.965 366.625 ;
        RECT 1357.395 366.345 1357.675 366.625 ;
        RECT 1358.105 366.345 1358.385 366.625 ;
        RECT 1358.815 366.345 1359.095 366.625 ;
        RECT 1359.525 366.345 1359.805 366.625 ;
        RECT 1360.235 366.345 1360.515 366.625 ;
        RECT 1351.715 365.635 1351.995 365.915 ;
        RECT 1352.425 365.635 1352.705 365.915 ;
        RECT 1353.135 365.635 1353.415 365.915 ;
        RECT 1353.845 365.635 1354.125 365.915 ;
        RECT 1354.555 365.635 1354.835 365.915 ;
        RECT 1355.265 365.635 1355.545 365.915 ;
        RECT 1355.975 365.635 1356.255 365.915 ;
        RECT 1356.685 365.635 1356.965 365.915 ;
        RECT 1357.395 365.635 1357.675 365.915 ;
        RECT 1358.105 365.635 1358.385 365.915 ;
        RECT 1358.815 365.635 1359.095 365.915 ;
        RECT 1359.525 365.635 1359.805 365.915 ;
        RECT 1360.235 365.635 1360.515 365.915 ;
        RECT 1351.715 364.925 1351.995 365.205 ;
        RECT 1352.425 364.925 1352.705 365.205 ;
        RECT 1353.135 364.925 1353.415 365.205 ;
        RECT 1353.845 364.925 1354.125 365.205 ;
        RECT 1354.555 364.925 1354.835 365.205 ;
        RECT 1355.265 364.925 1355.545 365.205 ;
        RECT 1355.975 364.925 1356.255 365.205 ;
        RECT 1356.685 364.925 1356.965 365.205 ;
        RECT 1357.395 364.925 1357.675 365.205 ;
        RECT 1358.105 364.925 1358.385 365.205 ;
        RECT 1358.815 364.925 1359.095 365.205 ;
        RECT 1359.525 364.925 1359.805 365.205 ;
        RECT 1360.235 364.925 1360.515 365.205 ;
        RECT 1351.715 364.215 1351.995 364.495 ;
        RECT 1352.425 364.215 1352.705 364.495 ;
        RECT 1353.135 364.215 1353.415 364.495 ;
        RECT 1353.845 364.215 1354.125 364.495 ;
        RECT 1354.555 364.215 1354.835 364.495 ;
        RECT 1355.265 364.215 1355.545 364.495 ;
        RECT 1355.975 364.215 1356.255 364.495 ;
        RECT 1356.685 364.215 1356.965 364.495 ;
        RECT 1357.395 364.215 1357.675 364.495 ;
        RECT 1358.105 364.215 1358.385 364.495 ;
        RECT 1358.815 364.215 1359.095 364.495 ;
        RECT 1359.525 364.215 1359.805 364.495 ;
        RECT 1360.235 364.215 1360.515 364.495 ;
        RECT 1351.715 363.505 1351.995 363.785 ;
        RECT 1352.425 363.505 1352.705 363.785 ;
        RECT 1353.135 363.505 1353.415 363.785 ;
        RECT 1353.845 363.505 1354.125 363.785 ;
        RECT 1354.555 363.505 1354.835 363.785 ;
        RECT 1355.265 363.505 1355.545 363.785 ;
        RECT 1355.975 363.505 1356.255 363.785 ;
        RECT 1356.685 363.505 1356.965 363.785 ;
        RECT 1357.395 363.505 1357.675 363.785 ;
        RECT 1358.105 363.505 1358.385 363.785 ;
        RECT 1358.815 363.505 1359.095 363.785 ;
        RECT 1359.525 363.505 1359.805 363.785 ;
        RECT 1360.235 363.505 1360.515 363.785 ;
        RECT 1351.715 362.795 1351.995 363.075 ;
        RECT 1352.425 362.795 1352.705 363.075 ;
        RECT 1353.135 362.795 1353.415 363.075 ;
        RECT 1353.845 362.795 1354.125 363.075 ;
        RECT 1354.555 362.795 1354.835 363.075 ;
        RECT 1355.265 362.795 1355.545 363.075 ;
        RECT 1355.975 362.795 1356.255 363.075 ;
        RECT 1356.685 362.795 1356.965 363.075 ;
        RECT 1357.395 362.795 1357.675 363.075 ;
        RECT 1358.105 362.795 1358.385 363.075 ;
        RECT 1358.815 362.795 1359.095 363.075 ;
        RECT 1359.525 362.795 1359.805 363.075 ;
        RECT 1360.235 362.795 1360.515 363.075 ;
        RECT 1351.715 362.085 1351.995 362.365 ;
        RECT 1352.425 362.085 1352.705 362.365 ;
        RECT 1353.135 362.085 1353.415 362.365 ;
        RECT 1353.845 362.085 1354.125 362.365 ;
        RECT 1354.555 362.085 1354.835 362.365 ;
        RECT 1355.265 362.085 1355.545 362.365 ;
        RECT 1355.975 362.085 1356.255 362.365 ;
        RECT 1356.685 362.085 1356.965 362.365 ;
        RECT 1357.395 362.085 1357.675 362.365 ;
        RECT 1358.105 362.085 1358.385 362.365 ;
        RECT 1358.815 362.085 1359.095 362.365 ;
        RECT 1359.525 362.085 1359.805 362.365 ;
        RECT 1360.235 362.085 1360.515 362.365 ;
        RECT 1351.715 361.375 1351.995 361.655 ;
        RECT 1352.425 361.375 1352.705 361.655 ;
        RECT 1353.135 361.375 1353.415 361.655 ;
        RECT 1353.845 361.375 1354.125 361.655 ;
        RECT 1354.555 361.375 1354.835 361.655 ;
        RECT 1355.265 361.375 1355.545 361.655 ;
        RECT 1355.975 361.375 1356.255 361.655 ;
        RECT 1356.685 361.375 1356.965 361.655 ;
        RECT 1357.395 361.375 1357.675 361.655 ;
        RECT 1358.105 361.375 1358.385 361.655 ;
        RECT 1358.815 361.375 1359.095 361.655 ;
        RECT 1359.525 361.375 1359.805 361.655 ;
        RECT 1360.235 361.375 1360.515 361.655 ;
        RECT 1351.715 360.665 1351.995 360.945 ;
        RECT 1352.425 360.665 1352.705 360.945 ;
        RECT 1353.135 360.665 1353.415 360.945 ;
        RECT 1353.845 360.665 1354.125 360.945 ;
        RECT 1354.555 360.665 1354.835 360.945 ;
        RECT 1355.265 360.665 1355.545 360.945 ;
        RECT 1355.975 360.665 1356.255 360.945 ;
        RECT 1356.685 360.665 1356.965 360.945 ;
        RECT 1357.395 360.665 1357.675 360.945 ;
        RECT 1358.105 360.665 1358.385 360.945 ;
        RECT 1358.815 360.665 1359.095 360.945 ;
        RECT 1359.525 360.665 1359.805 360.945 ;
        RECT 1360.235 360.665 1360.515 360.945 ;
        RECT 1366.245 369.895 1366.525 370.175 ;
        RECT 1366.955 369.895 1367.235 370.175 ;
        RECT 1367.665 369.895 1367.945 370.175 ;
        RECT 1368.375 369.895 1368.655 370.175 ;
        RECT 1369.085 369.895 1369.365 370.175 ;
        RECT 1369.795 369.895 1370.075 370.175 ;
        RECT 1370.505 369.895 1370.785 370.175 ;
        RECT 1371.215 369.895 1371.495 370.175 ;
        RECT 1371.925 369.895 1372.205 370.175 ;
        RECT 1372.635 369.895 1372.915 370.175 ;
        RECT 1373.345 369.895 1373.625 370.175 ;
        RECT 1366.245 369.185 1366.525 369.465 ;
        RECT 1366.955 369.185 1367.235 369.465 ;
        RECT 1367.665 369.185 1367.945 369.465 ;
        RECT 1368.375 369.185 1368.655 369.465 ;
        RECT 1369.085 369.185 1369.365 369.465 ;
        RECT 1369.795 369.185 1370.075 369.465 ;
        RECT 1370.505 369.185 1370.785 369.465 ;
        RECT 1371.215 369.185 1371.495 369.465 ;
        RECT 1371.925 369.185 1372.205 369.465 ;
        RECT 1372.635 369.185 1372.915 369.465 ;
        RECT 1373.345 369.185 1373.625 369.465 ;
        RECT 1366.245 368.475 1366.525 368.755 ;
        RECT 1366.955 368.475 1367.235 368.755 ;
        RECT 1367.665 368.475 1367.945 368.755 ;
        RECT 1368.375 368.475 1368.655 368.755 ;
        RECT 1369.085 368.475 1369.365 368.755 ;
        RECT 1369.795 368.475 1370.075 368.755 ;
        RECT 1370.505 368.475 1370.785 368.755 ;
        RECT 1371.215 368.475 1371.495 368.755 ;
        RECT 1371.925 368.475 1372.205 368.755 ;
        RECT 1372.635 368.475 1372.915 368.755 ;
        RECT 1373.345 368.475 1373.625 368.755 ;
        RECT 1366.245 367.765 1366.525 368.045 ;
        RECT 1366.955 367.765 1367.235 368.045 ;
        RECT 1367.665 367.765 1367.945 368.045 ;
        RECT 1368.375 367.765 1368.655 368.045 ;
        RECT 1369.085 367.765 1369.365 368.045 ;
        RECT 1369.795 367.765 1370.075 368.045 ;
        RECT 1370.505 367.765 1370.785 368.045 ;
        RECT 1371.215 367.765 1371.495 368.045 ;
        RECT 1371.925 367.765 1372.205 368.045 ;
        RECT 1372.635 367.765 1372.915 368.045 ;
        RECT 1373.345 367.765 1373.625 368.045 ;
        RECT 1366.245 367.055 1366.525 367.335 ;
        RECT 1366.955 367.055 1367.235 367.335 ;
        RECT 1367.665 367.055 1367.945 367.335 ;
        RECT 1368.375 367.055 1368.655 367.335 ;
        RECT 1369.085 367.055 1369.365 367.335 ;
        RECT 1369.795 367.055 1370.075 367.335 ;
        RECT 1370.505 367.055 1370.785 367.335 ;
        RECT 1371.215 367.055 1371.495 367.335 ;
        RECT 1371.925 367.055 1372.205 367.335 ;
        RECT 1372.635 367.055 1372.915 367.335 ;
        RECT 1373.345 367.055 1373.625 367.335 ;
        RECT 1366.245 366.345 1366.525 366.625 ;
        RECT 1366.955 366.345 1367.235 366.625 ;
        RECT 1367.665 366.345 1367.945 366.625 ;
        RECT 1368.375 366.345 1368.655 366.625 ;
        RECT 1369.085 366.345 1369.365 366.625 ;
        RECT 1369.795 366.345 1370.075 366.625 ;
        RECT 1370.505 366.345 1370.785 366.625 ;
        RECT 1371.215 366.345 1371.495 366.625 ;
        RECT 1371.925 366.345 1372.205 366.625 ;
        RECT 1372.635 366.345 1372.915 366.625 ;
        RECT 1373.345 366.345 1373.625 366.625 ;
        RECT 1366.245 365.635 1366.525 365.915 ;
        RECT 1366.955 365.635 1367.235 365.915 ;
        RECT 1367.665 365.635 1367.945 365.915 ;
        RECT 1368.375 365.635 1368.655 365.915 ;
        RECT 1369.085 365.635 1369.365 365.915 ;
        RECT 1369.795 365.635 1370.075 365.915 ;
        RECT 1370.505 365.635 1370.785 365.915 ;
        RECT 1371.215 365.635 1371.495 365.915 ;
        RECT 1371.925 365.635 1372.205 365.915 ;
        RECT 1372.635 365.635 1372.915 365.915 ;
        RECT 1373.345 365.635 1373.625 365.915 ;
        RECT 1366.245 364.925 1366.525 365.205 ;
        RECT 1366.955 364.925 1367.235 365.205 ;
        RECT 1367.665 364.925 1367.945 365.205 ;
        RECT 1368.375 364.925 1368.655 365.205 ;
        RECT 1369.085 364.925 1369.365 365.205 ;
        RECT 1369.795 364.925 1370.075 365.205 ;
        RECT 1370.505 364.925 1370.785 365.205 ;
        RECT 1371.215 364.925 1371.495 365.205 ;
        RECT 1371.925 364.925 1372.205 365.205 ;
        RECT 1372.635 364.925 1372.915 365.205 ;
        RECT 1373.345 364.925 1373.625 365.205 ;
        RECT 1366.245 364.215 1366.525 364.495 ;
        RECT 1366.955 364.215 1367.235 364.495 ;
        RECT 1367.665 364.215 1367.945 364.495 ;
        RECT 1368.375 364.215 1368.655 364.495 ;
        RECT 1369.085 364.215 1369.365 364.495 ;
        RECT 1369.795 364.215 1370.075 364.495 ;
        RECT 1370.505 364.215 1370.785 364.495 ;
        RECT 1371.215 364.215 1371.495 364.495 ;
        RECT 1371.925 364.215 1372.205 364.495 ;
        RECT 1372.635 364.215 1372.915 364.495 ;
        RECT 1373.345 364.215 1373.625 364.495 ;
        RECT 1366.245 363.505 1366.525 363.785 ;
        RECT 1366.955 363.505 1367.235 363.785 ;
        RECT 1367.665 363.505 1367.945 363.785 ;
        RECT 1368.375 363.505 1368.655 363.785 ;
        RECT 1369.085 363.505 1369.365 363.785 ;
        RECT 1369.795 363.505 1370.075 363.785 ;
        RECT 1370.505 363.505 1370.785 363.785 ;
        RECT 1371.215 363.505 1371.495 363.785 ;
        RECT 1371.925 363.505 1372.205 363.785 ;
        RECT 1372.635 363.505 1372.915 363.785 ;
        RECT 1373.345 363.505 1373.625 363.785 ;
        RECT 1366.245 362.795 1366.525 363.075 ;
        RECT 1366.955 362.795 1367.235 363.075 ;
        RECT 1367.665 362.795 1367.945 363.075 ;
        RECT 1368.375 362.795 1368.655 363.075 ;
        RECT 1369.085 362.795 1369.365 363.075 ;
        RECT 1369.795 362.795 1370.075 363.075 ;
        RECT 1370.505 362.795 1370.785 363.075 ;
        RECT 1371.215 362.795 1371.495 363.075 ;
        RECT 1371.925 362.795 1372.205 363.075 ;
        RECT 1372.635 362.795 1372.915 363.075 ;
        RECT 1373.345 362.795 1373.625 363.075 ;
        RECT 1366.245 362.085 1366.525 362.365 ;
        RECT 1366.955 362.085 1367.235 362.365 ;
        RECT 1367.665 362.085 1367.945 362.365 ;
        RECT 1368.375 362.085 1368.655 362.365 ;
        RECT 1369.085 362.085 1369.365 362.365 ;
        RECT 1369.795 362.085 1370.075 362.365 ;
        RECT 1370.505 362.085 1370.785 362.365 ;
        RECT 1371.215 362.085 1371.495 362.365 ;
        RECT 1371.925 362.085 1372.205 362.365 ;
        RECT 1372.635 362.085 1372.915 362.365 ;
        RECT 1373.345 362.085 1373.625 362.365 ;
        RECT 1366.245 361.375 1366.525 361.655 ;
        RECT 1366.955 361.375 1367.235 361.655 ;
        RECT 1367.665 361.375 1367.945 361.655 ;
        RECT 1368.375 361.375 1368.655 361.655 ;
        RECT 1369.085 361.375 1369.365 361.655 ;
        RECT 1369.795 361.375 1370.075 361.655 ;
        RECT 1370.505 361.375 1370.785 361.655 ;
        RECT 1371.215 361.375 1371.495 361.655 ;
        RECT 1371.925 361.375 1372.205 361.655 ;
        RECT 1372.635 361.375 1372.915 361.655 ;
        RECT 1373.345 361.375 1373.625 361.655 ;
        RECT 1366.245 360.665 1366.525 360.945 ;
        RECT 1366.955 360.665 1367.235 360.945 ;
        RECT 1367.665 360.665 1367.945 360.945 ;
        RECT 1368.375 360.665 1368.655 360.945 ;
        RECT 1369.085 360.665 1369.365 360.945 ;
        RECT 1369.795 360.665 1370.075 360.945 ;
        RECT 1370.505 360.665 1370.785 360.945 ;
        RECT 1371.215 360.665 1371.495 360.945 ;
        RECT 1371.925 360.665 1372.205 360.945 ;
        RECT 1372.635 360.665 1372.915 360.945 ;
        RECT 1373.345 360.665 1373.625 360.945 ;
        RECT 1375.965 369.895 1376.245 370.175 ;
        RECT 1376.675 369.895 1376.955 370.175 ;
        RECT 1377.385 369.895 1377.665 370.175 ;
        RECT 1378.095 369.895 1378.375 370.175 ;
        RECT 1378.805 369.895 1379.085 370.175 ;
        RECT 1379.515 369.895 1379.795 370.175 ;
        RECT 1380.225 369.895 1380.505 370.175 ;
        RECT 1380.935 369.895 1381.215 370.175 ;
        RECT 1381.645 369.895 1381.925 370.175 ;
        RECT 1382.355 369.895 1382.635 370.175 ;
        RECT 1383.065 369.895 1383.345 370.175 ;
        RECT 1383.775 369.895 1384.055 370.175 ;
        RECT 1384.485 369.895 1384.765 370.175 ;
        RECT 1385.195 369.895 1385.475 370.175 ;
        RECT 1375.965 369.185 1376.245 369.465 ;
        RECT 1376.675 369.185 1376.955 369.465 ;
        RECT 1377.385 369.185 1377.665 369.465 ;
        RECT 1378.095 369.185 1378.375 369.465 ;
        RECT 1378.805 369.185 1379.085 369.465 ;
        RECT 1379.515 369.185 1379.795 369.465 ;
        RECT 1380.225 369.185 1380.505 369.465 ;
        RECT 1380.935 369.185 1381.215 369.465 ;
        RECT 1381.645 369.185 1381.925 369.465 ;
        RECT 1382.355 369.185 1382.635 369.465 ;
        RECT 1383.065 369.185 1383.345 369.465 ;
        RECT 1383.775 369.185 1384.055 369.465 ;
        RECT 1384.485 369.185 1384.765 369.465 ;
        RECT 1385.195 369.185 1385.475 369.465 ;
        RECT 1375.965 368.475 1376.245 368.755 ;
        RECT 1376.675 368.475 1376.955 368.755 ;
        RECT 1377.385 368.475 1377.665 368.755 ;
        RECT 1378.095 368.475 1378.375 368.755 ;
        RECT 1378.805 368.475 1379.085 368.755 ;
        RECT 1379.515 368.475 1379.795 368.755 ;
        RECT 1380.225 368.475 1380.505 368.755 ;
        RECT 1380.935 368.475 1381.215 368.755 ;
        RECT 1381.645 368.475 1381.925 368.755 ;
        RECT 1382.355 368.475 1382.635 368.755 ;
        RECT 1383.065 368.475 1383.345 368.755 ;
        RECT 1383.775 368.475 1384.055 368.755 ;
        RECT 1384.485 368.475 1384.765 368.755 ;
        RECT 1385.195 368.475 1385.475 368.755 ;
        RECT 1375.965 367.765 1376.245 368.045 ;
        RECT 1376.675 367.765 1376.955 368.045 ;
        RECT 1377.385 367.765 1377.665 368.045 ;
        RECT 1378.095 367.765 1378.375 368.045 ;
        RECT 1378.805 367.765 1379.085 368.045 ;
        RECT 1379.515 367.765 1379.795 368.045 ;
        RECT 1380.225 367.765 1380.505 368.045 ;
        RECT 1380.935 367.765 1381.215 368.045 ;
        RECT 1381.645 367.765 1381.925 368.045 ;
        RECT 1382.355 367.765 1382.635 368.045 ;
        RECT 1383.065 367.765 1383.345 368.045 ;
        RECT 1383.775 367.765 1384.055 368.045 ;
        RECT 1384.485 367.765 1384.765 368.045 ;
        RECT 1385.195 367.765 1385.475 368.045 ;
        RECT 1375.965 367.055 1376.245 367.335 ;
        RECT 1376.675 367.055 1376.955 367.335 ;
        RECT 1377.385 367.055 1377.665 367.335 ;
        RECT 1378.095 367.055 1378.375 367.335 ;
        RECT 1378.805 367.055 1379.085 367.335 ;
        RECT 1379.515 367.055 1379.795 367.335 ;
        RECT 1380.225 367.055 1380.505 367.335 ;
        RECT 1380.935 367.055 1381.215 367.335 ;
        RECT 1381.645 367.055 1381.925 367.335 ;
        RECT 1382.355 367.055 1382.635 367.335 ;
        RECT 1383.065 367.055 1383.345 367.335 ;
        RECT 1383.775 367.055 1384.055 367.335 ;
        RECT 1384.485 367.055 1384.765 367.335 ;
        RECT 1385.195 367.055 1385.475 367.335 ;
        RECT 1375.965 366.345 1376.245 366.625 ;
        RECT 1376.675 366.345 1376.955 366.625 ;
        RECT 1377.385 366.345 1377.665 366.625 ;
        RECT 1378.095 366.345 1378.375 366.625 ;
        RECT 1378.805 366.345 1379.085 366.625 ;
        RECT 1379.515 366.345 1379.795 366.625 ;
        RECT 1380.225 366.345 1380.505 366.625 ;
        RECT 1380.935 366.345 1381.215 366.625 ;
        RECT 1381.645 366.345 1381.925 366.625 ;
        RECT 1382.355 366.345 1382.635 366.625 ;
        RECT 1383.065 366.345 1383.345 366.625 ;
        RECT 1383.775 366.345 1384.055 366.625 ;
        RECT 1384.485 366.345 1384.765 366.625 ;
        RECT 1385.195 366.345 1385.475 366.625 ;
        RECT 1375.965 365.635 1376.245 365.915 ;
        RECT 1376.675 365.635 1376.955 365.915 ;
        RECT 1377.385 365.635 1377.665 365.915 ;
        RECT 1378.095 365.635 1378.375 365.915 ;
        RECT 1378.805 365.635 1379.085 365.915 ;
        RECT 1379.515 365.635 1379.795 365.915 ;
        RECT 1380.225 365.635 1380.505 365.915 ;
        RECT 1380.935 365.635 1381.215 365.915 ;
        RECT 1381.645 365.635 1381.925 365.915 ;
        RECT 1382.355 365.635 1382.635 365.915 ;
        RECT 1383.065 365.635 1383.345 365.915 ;
        RECT 1383.775 365.635 1384.055 365.915 ;
        RECT 1384.485 365.635 1384.765 365.915 ;
        RECT 1385.195 365.635 1385.475 365.915 ;
        RECT 1375.965 364.925 1376.245 365.205 ;
        RECT 1376.675 364.925 1376.955 365.205 ;
        RECT 1377.385 364.925 1377.665 365.205 ;
        RECT 1378.095 364.925 1378.375 365.205 ;
        RECT 1378.805 364.925 1379.085 365.205 ;
        RECT 1379.515 364.925 1379.795 365.205 ;
        RECT 1380.225 364.925 1380.505 365.205 ;
        RECT 1380.935 364.925 1381.215 365.205 ;
        RECT 1381.645 364.925 1381.925 365.205 ;
        RECT 1382.355 364.925 1382.635 365.205 ;
        RECT 1383.065 364.925 1383.345 365.205 ;
        RECT 1383.775 364.925 1384.055 365.205 ;
        RECT 1384.485 364.925 1384.765 365.205 ;
        RECT 1385.195 364.925 1385.475 365.205 ;
        RECT 1375.965 364.215 1376.245 364.495 ;
        RECT 1376.675 364.215 1376.955 364.495 ;
        RECT 1377.385 364.215 1377.665 364.495 ;
        RECT 1378.095 364.215 1378.375 364.495 ;
        RECT 1378.805 364.215 1379.085 364.495 ;
        RECT 1379.515 364.215 1379.795 364.495 ;
        RECT 1380.225 364.215 1380.505 364.495 ;
        RECT 1380.935 364.215 1381.215 364.495 ;
        RECT 1381.645 364.215 1381.925 364.495 ;
        RECT 1382.355 364.215 1382.635 364.495 ;
        RECT 1383.065 364.215 1383.345 364.495 ;
        RECT 1383.775 364.215 1384.055 364.495 ;
        RECT 1384.485 364.215 1384.765 364.495 ;
        RECT 1385.195 364.215 1385.475 364.495 ;
        RECT 1375.965 363.505 1376.245 363.785 ;
        RECT 1376.675 363.505 1376.955 363.785 ;
        RECT 1377.385 363.505 1377.665 363.785 ;
        RECT 1378.095 363.505 1378.375 363.785 ;
        RECT 1378.805 363.505 1379.085 363.785 ;
        RECT 1379.515 363.505 1379.795 363.785 ;
        RECT 1380.225 363.505 1380.505 363.785 ;
        RECT 1380.935 363.505 1381.215 363.785 ;
        RECT 1381.645 363.505 1381.925 363.785 ;
        RECT 1382.355 363.505 1382.635 363.785 ;
        RECT 1383.065 363.505 1383.345 363.785 ;
        RECT 1383.775 363.505 1384.055 363.785 ;
        RECT 1384.485 363.505 1384.765 363.785 ;
        RECT 1385.195 363.505 1385.475 363.785 ;
        RECT 1375.965 362.795 1376.245 363.075 ;
        RECT 1376.675 362.795 1376.955 363.075 ;
        RECT 1377.385 362.795 1377.665 363.075 ;
        RECT 1378.095 362.795 1378.375 363.075 ;
        RECT 1378.805 362.795 1379.085 363.075 ;
        RECT 1379.515 362.795 1379.795 363.075 ;
        RECT 1380.225 362.795 1380.505 363.075 ;
        RECT 1380.935 362.795 1381.215 363.075 ;
        RECT 1381.645 362.795 1381.925 363.075 ;
        RECT 1382.355 362.795 1382.635 363.075 ;
        RECT 1383.065 362.795 1383.345 363.075 ;
        RECT 1383.775 362.795 1384.055 363.075 ;
        RECT 1384.485 362.795 1384.765 363.075 ;
        RECT 1385.195 362.795 1385.475 363.075 ;
        RECT 1375.965 362.085 1376.245 362.365 ;
        RECT 1376.675 362.085 1376.955 362.365 ;
        RECT 1377.385 362.085 1377.665 362.365 ;
        RECT 1378.095 362.085 1378.375 362.365 ;
        RECT 1378.805 362.085 1379.085 362.365 ;
        RECT 1379.515 362.085 1379.795 362.365 ;
        RECT 1380.225 362.085 1380.505 362.365 ;
        RECT 1380.935 362.085 1381.215 362.365 ;
        RECT 1381.645 362.085 1381.925 362.365 ;
        RECT 1382.355 362.085 1382.635 362.365 ;
        RECT 1383.065 362.085 1383.345 362.365 ;
        RECT 1383.775 362.085 1384.055 362.365 ;
        RECT 1384.485 362.085 1384.765 362.365 ;
        RECT 1385.195 362.085 1385.475 362.365 ;
        RECT 1375.965 361.375 1376.245 361.655 ;
        RECT 1376.675 361.375 1376.955 361.655 ;
        RECT 1377.385 361.375 1377.665 361.655 ;
        RECT 1378.095 361.375 1378.375 361.655 ;
        RECT 1378.805 361.375 1379.085 361.655 ;
        RECT 1379.515 361.375 1379.795 361.655 ;
        RECT 1380.225 361.375 1380.505 361.655 ;
        RECT 1380.935 361.375 1381.215 361.655 ;
        RECT 1381.645 361.375 1381.925 361.655 ;
        RECT 1382.355 361.375 1382.635 361.655 ;
        RECT 1383.065 361.375 1383.345 361.655 ;
        RECT 1383.775 361.375 1384.055 361.655 ;
        RECT 1384.485 361.375 1384.765 361.655 ;
        RECT 1385.195 361.375 1385.475 361.655 ;
        RECT 1375.965 360.665 1376.245 360.945 ;
        RECT 1376.675 360.665 1376.955 360.945 ;
        RECT 1377.385 360.665 1377.665 360.945 ;
        RECT 1378.095 360.665 1378.375 360.945 ;
        RECT 1378.805 360.665 1379.085 360.945 ;
        RECT 1379.515 360.665 1379.795 360.945 ;
        RECT 1380.225 360.665 1380.505 360.945 ;
        RECT 1380.935 360.665 1381.215 360.945 ;
        RECT 1381.645 360.665 1381.925 360.945 ;
        RECT 1382.355 360.665 1382.635 360.945 ;
        RECT 1383.065 360.665 1383.345 360.945 ;
        RECT 1383.775 360.665 1384.055 360.945 ;
        RECT 1384.485 360.665 1384.765 360.945 ;
        RECT 1385.195 360.665 1385.475 360.945 ;
        RECT 1389.495 369.895 1389.775 370.175 ;
        RECT 1390.205 369.895 1390.485 370.175 ;
        RECT 1390.915 369.895 1391.195 370.175 ;
        RECT 1391.625 369.895 1391.905 370.175 ;
        RECT 1392.335 369.895 1392.615 370.175 ;
        RECT 1393.045 369.895 1393.325 370.175 ;
        RECT 1393.755 369.895 1394.035 370.175 ;
        RECT 1394.465 369.895 1394.745 370.175 ;
        RECT 1395.175 369.895 1395.455 370.175 ;
        RECT 1395.885 369.895 1396.165 370.175 ;
        RECT 1396.595 369.895 1396.875 370.175 ;
        RECT 1397.305 369.895 1397.585 370.175 ;
        RECT 1398.015 369.895 1398.295 370.175 ;
        RECT 1398.725 369.895 1399.005 370.175 ;
        RECT 1389.495 369.185 1389.775 369.465 ;
        RECT 1390.205 369.185 1390.485 369.465 ;
        RECT 1390.915 369.185 1391.195 369.465 ;
        RECT 1391.625 369.185 1391.905 369.465 ;
        RECT 1392.335 369.185 1392.615 369.465 ;
        RECT 1393.045 369.185 1393.325 369.465 ;
        RECT 1393.755 369.185 1394.035 369.465 ;
        RECT 1394.465 369.185 1394.745 369.465 ;
        RECT 1395.175 369.185 1395.455 369.465 ;
        RECT 1395.885 369.185 1396.165 369.465 ;
        RECT 1396.595 369.185 1396.875 369.465 ;
        RECT 1397.305 369.185 1397.585 369.465 ;
        RECT 1398.015 369.185 1398.295 369.465 ;
        RECT 1398.725 369.185 1399.005 369.465 ;
        RECT 1389.495 368.475 1389.775 368.755 ;
        RECT 1390.205 368.475 1390.485 368.755 ;
        RECT 1390.915 368.475 1391.195 368.755 ;
        RECT 1391.625 368.475 1391.905 368.755 ;
        RECT 1392.335 368.475 1392.615 368.755 ;
        RECT 1393.045 368.475 1393.325 368.755 ;
        RECT 1393.755 368.475 1394.035 368.755 ;
        RECT 1394.465 368.475 1394.745 368.755 ;
        RECT 1395.175 368.475 1395.455 368.755 ;
        RECT 1395.885 368.475 1396.165 368.755 ;
        RECT 1396.595 368.475 1396.875 368.755 ;
        RECT 1397.305 368.475 1397.585 368.755 ;
        RECT 1398.015 368.475 1398.295 368.755 ;
        RECT 1398.725 368.475 1399.005 368.755 ;
        RECT 1389.495 367.765 1389.775 368.045 ;
        RECT 1390.205 367.765 1390.485 368.045 ;
        RECT 1390.915 367.765 1391.195 368.045 ;
        RECT 1391.625 367.765 1391.905 368.045 ;
        RECT 1392.335 367.765 1392.615 368.045 ;
        RECT 1393.045 367.765 1393.325 368.045 ;
        RECT 1393.755 367.765 1394.035 368.045 ;
        RECT 1394.465 367.765 1394.745 368.045 ;
        RECT 1395.175 367.765 1395.455 368.045 ;
        RECT 1395.885 367.765 1396.165 368.045 ;
        RECT 1396.595 367.765 1396.875 368.045 ;
        RECT 1397.305 367.765 1397.585 368.045 ;
        RECT 1398.015 367.765 1398.295 368.045 ;
        RECT 1398.725 367.765 1399.005 368.045 ;
        RECT 1389.495 367.055 1389.775 367.335 ;
        RECT 1390.205 367.055 1390.485 367.335 ;
        RECT 1390.915 367.055 1391.195 367.335 ;
        RECT 1391.625 367.055 1391.905 367.335 ;
        RECT 1392.335 367.055 1392.615 367.335 ;
        RECT 1393.045 367.055 1393.325 367.335 ;
        RECT 1393.755 367.055 1394.035 367.335 ;
        RECT 1394.465 367.055 1394.745 367.335 ;
        RECT 1395.175 367.055 1395.455 367.335 ;
        RECT 1395.885 367.055 1396.165 367.335 ;
        RECT 1396.595 367.055 1396.875 367.335 ;
        RECT 1397.305 367.055 1397.585 367.335 ;
        RECT 1398.015 367.055 1398.295 367.335 ;
        RECT 1398.725 367.055 1399.005 367.335 ;
        RECT 1389.495 366.345 1389.775 366.625 ;
        RECT 1390.205 366.345 1390.485 366.625 ;
        RECT 1390.915 366.345 1391.195 366.625 ;
        RECT 1391.625 366.345 1391.905 366.625 ;
        RECT 1392.335 366.345 1392.615 366.625 ;
        RECT 1393.045 366.345 1393.325 366.625 ;
        RECT 1393.755 366.345 1394.035 366.625 ;
        RECT 1394.465 366.345 1394.745 366.625 ;
        RECT 1395.175 366.345 1395.455 366.625 ;
        RECT 1395.885 366.345 1396.165 366.625 ;
        RECT 1396.595 366.345 1396.875 366.625 ;
        RECT 1397.305 366.345 1397.585 366.625 ;
        RECT 1398.015 366.345 1398.295 366.625 ;
        RECT 1398.725 366.345 1399.005 366.625 ;
        RECT 1389.495 365.635 1389.775 365.915 ;
        RECT 1390.205 365.635 1390.485 365.915 ;
        RECT 1390.915 365.635 1391.195 365.915 ;
        RECT 1391.625 365.635 1391.905 365.915 ;
        RECT 1392.335 365.635 1392.615 365.915 ;
        RECT 1393.045 365.635 1393.325 365.915 ;
        RECT 1393.755 365.635 1394.035 365.915 ;
        RECT 1394.465 365.635 1394.745 365.915 ;
        RECT 1395.175 365.635 1395.455 365.915 ;
        RECT 1395.885 365.635 1396.165 365.915 ;
        RECT 1396.595 365.635 1396.875 365.915 ;
        RECT 1397.305 365.635 1397.585 365.915 ;
        RECT 1398.015 365.635 1398.295 365.915 ;
        RECT 1398.725 365.635 1399.005 365.915 ;
        RECT 1389.495 364.925 1389.775 365.205 ;
        RECT 1390.205 364.925 1390.485 365.205 ;
        RECT 1390.915 364.925 1391.195 365.205 ;
        RECT 1391.625 364.925 1391.905 365.205 ;
        RECT 1392.335 364.925 1392.615 365.205 ;
        RECT 1393.045 364.925 1393.325 365.205 ;
        RECT 1393.755 364.925 1394.035 365.205 ;
        RECT 1394.465 364.925 1394.745 365.205 ;
        RECT 1395.175 364.925 1395.455 365.205 ;
        RECT 1395.885 364.925 1396.165 365.205 ;
        RECT 1396.595 364.925 1396.875 365.205 ;
        RECT 1397.305 364.925 1397.585 365.205 ;
        RECT 1398.015 364.925 1398.295 365.205 ;
        RECT 1398.725 364.925 1399.005 365.205 ;
        RECT 1389.495 364.215 1389.775 364.495 ;
        RECT 1390.205 364.215 1390.485 364.495 ;
        RECT 1390.915 364.215 1391.195 364.495 ;
        RECT 1391.625 364.215 1391.905 364.495 ;
        RECT 1392.335 364.215 1392.615 364.495 ;
        RECT 1393.045 364.215 1393.325 364.495 ;
        RECT 1393.755 364.215 1394.035 364.495 ;
        RECT 1394.465 364.215 1394.745 364.495 ;
        RECT 1395.175 364.215 1395.455 364.495 ;
        RECT 1395.885 364.215 1396.165 364.495 ;
        RECT 1396.595 364.215 1396.875 364.495 ;
        RECT 1397.305 364.215 1397.585 364.495 ;
        RECT 1398.015 364.215 1398.295 364.495 ;
        RECT 1398.725 364.215 1399.005 364.495 ;
        RECT 1389.495 363.505 1389.775 363.785 ;
        RECT 1390.205 363.505 1390.485 363.785 ;
        RECT 1390.915 363.505 1391.195 363.785 ;
        RECT 1391.625 363.505 1391.905 363.785 ;
        RECT 1392.335 363.505 1392.615 363.785 ;
        RECT 1393.045 363.505 1393.325 363.785 ;
        RECT 1393.755 363.505 1394.035 363.785 ;
        RECT 1394.465 363.505 1394.745 363.785 ;
        RECT 1395.175 363.505 1395.455 363.785 ;
        RECT 1395.885 363.505 1396.165 363.785 ;
        RECT 1396.595 363.505 1396.875 363.785 ;
        RECT 1397.305 363.505 1397.585 363.785 ;
        RECT 1398.015 363.505 1398.295 363.785 ;
        RECT 1398.725 363.505 1399.005 363.785 ;
        RECT 1389.495 362.795 1389.775 363.075 ;
        RECT 1390.205 362.795 1390.485 363.075 ;
        RECT 1390.915 362.795 1391.195 363.075 ;
        RECT 1391.625 362.795 1391.905 363.075 ;
        RECT 1392.335 362.795 1392.615 363.075 ;
        RECT 1393.045 362.795 1393.325 363.075 ;
        RECT 1393.755 362.795 1394.035 363.075 ;
        RECT 1394.465 362.795 1394.745 363.075 ;
        RECT 1395.175 362.795 1395.455 363.075 ;
        RECT 1395.885 362.795 1396.165 363.075 ;
        RECT 1396.595 362.795 1396.875 363.075 ;
        RECT 1397.305 362.795 1397.585 363.075 ;
        RECT 1398.015 362.795 1398.295 363.075 ;
        RECT 1398.725 362.795 1399.005 363.075 ;
        RECT 1389.495 362.085 1389.775 362.365 ;
        RECT 1390.205 362.085 1390.485 362.365 ;
        RECT 1390.915 362.085 1391.195 362.365 ;
        RECT 1391.625 362.085 1391.905 362.365 ;
        RECT 1392.335 362.085 1392.615 362.365 ;
        RECT 1393.045 362.085 1393.325 362.365 ;
        RECT 1393.755 362.085 1394.035 362.365 ;
        RECT 1394.465 362.085 1394.745 362.365 ;
        RECT 1395.175 362.085 1395.455 362.365 ;
        RECT 1395.885 362.085 1396.165 362.365 ;
        RECT 1396.595 362.085 1396.875 362.365 ;
        RECT 1397.305 362.085 1397.585 362.365 ;
        RECT 1398.015 362.085 1398.295 362.365 ;
        RECT 1398.725 362.085 1399.005 362.365 ;
        RECT 1389.495 361.375 1389.775 361.655 ;
        RECT 1390.205 361.375 1390.485 361.655 ;
        RECT 1390.915 361.375 1391.195 361.655 ;
        RECT 1391.625 361.375 1391.905 361.655 ;
        RECT 1392.335 361.375 1392.615 361.655 ;
        RECT 1393.045 361.375 1393.325 361.655 ;
        RECT 1393.755 361.375 1394.035 361.655 ;
        RECT 1394.465 361.375 1394.745 361.655 ;
        RECT 1395.175 361.375 1395.455 361.655 ;
        RECT 1395.885 361.375 1396.165 361.655 ;
        RECT 1396.595 361.375 1396.875 361.655 ;
        RECT 1397.305 361.375 1397.585 361.655 ;
        RECT 1398.015 361.375 1398.295 361.655 ;
        RECT 1398.725 361.375 1399.005 361.655 ;
        RECT 1389.495 360.665 1389.775 360.945 ;
        RECT 1390.205 360.665 1390.485 360.945 ;
        RECT 1390.915 360.665 1391.195 360.945 ;
        RECT 1391.625 360.665 1391.905 360.945 ;
        RECT 1392.335 360.665 1392.615 360.945 ;
        RECT 1393.045 360.665 1393.325 360.945 ;
        RECT 1393.755 360.665 1394.035 360.945 ;
        RECT 1394.465 360.665 1394.745 360.945 ;
        RECT 1395.175 360.665 1395.455 360.945 ;
        RECT 1395.885 360.665 1396.165 360.945 ;
        RECT 1396.595 360.665 1396.875 360.945 ;
        RECT 1397.305 360.665 1397.585 360.945 ;
        RECT 1398.015 360.665 1398.295 360.945 ;
        RECT 1398.725 360.665 1399.005 360.945 ;
        RECT 1401.345 369.895 1401.625 370.175 ;
        RECT 1402.055 369.895 1402.335 370.175 ;
        RECT 1402.765 369.895 1403.045 370.175 ;
        RECT 1403.475 369.895 1403.755 370.175 ;
        RECT 1404.185 369.895 1404.465 370.175 ;
        RECT 1404.895 369.895 1405.175 370.175 ;
        RECT 1405.605 369.895 1405.885 370.175 ;
        RECT 1406.315 369.895 1406.595 370.175 ;
        RECT 1407.025 369.895 1407.305 370.175 ;
        RECT 1407.735 369.895 1408.015 370.175 ;
        RECT 1408.445 369.895 1408.725 370.175 ;
        RECT 1409.155 369.895 1409.435 370.175 ;
        RECT 1409.865 369.895 1410.145 370.175 ;
        RECT 1410.575 369.895 1410.855 370.175 ;
        RECT 1401.345 369.185 1401.625 369.465 ;
        RECT 1402.055 369.185 1402.335 369.465 ;
        RECT 1402.765 369.185 1403.045 369.465 ;
        RECT 1403.475 369.185 1403.755 369.465 ;
        RECT 1404.185 369.185 1404.465 369.465 ;
        RECT 1404.895 369.185 1405.175 369.465 ;
        RECT 1405.605 369.185 1405.885 369.465 ;
        RECT 1406.315 369.185 1406.595 369.465 ;
        RECT 1407.025 369.185 1407.305 369.465 ;
        RECT 1407.735 369.185 1408.015 369.465 ;
        RECT 1408.445 369.185 1408.725 369.465 ;
        RECT 1409.155 369.185 1409.435 369.465 ;
        RECT 1409.865 369.185 1410.145 369.465 ;
        RECT 1410.575 369.185 1410.855 369.465 ;
        RECT 1401.345 368.475 1401.625 368.755 ;
        RECT 1402.055 368.475 1402.335 368.755 ;
        RECT 1402.765 368.475 1403.045 368.755 ;
        RECT 1403.475 368.475 1403.755 368.755 ;
        RECT 1404.185 368.475 1404.465 368.755 ;
        RECT 1404.895 368.475 1405.175 368.755 ;
        RECT 1405.605 368.475 1405.885 368.755 ;
        RECT 1406.315 368.475 1406.595 368.755 ;
        RECT 1407.025 368.475 1407.305 368.755 ;
        RECT 1407.735 368.475 1408.015 368.755 ;
        RECT 1408.445 368.475 1408.725 368.755 ;
        RECT 1409.155 368.475 1409.435 368.755 ;
        RECT 1409.865 368.475 1410.145 368.755 ;
        RECT 1410.575 368.475 1410.855 368.755 ;
        RECT 1401.345 367.765 1401.625 368.045 ;
        RECT 1402.055 367.765 1402.335 368.045 ;
        RECT 1402.765 367.765 1403.045 368.045 ;
        RECT 1403.475 367.765 1403.755 368.045 ;
        RECT 1404.185 367.765 1404.465 368.045 ;
        RECT 1404.895 367.765 1405.175 368.045 ;
        RECT 1405.605 367.765 1405.885 368.045 ;
        RECT 1406.315 367.765 1406.595 368.045 ;
        RECT 1407.025 367.765 1407.305 368.045 ;
        RECT 1407.735 367.765 1408.015 368.045 ;
        RECT 1408.445 367.765 1408.725 368.045 ;
        RECT 1409.155 367.765 1409.435 368.045 ;
        RECT 1409.865 367.765 1410.145 368.045 ;
        RECT 1410.575 367.765 1410.855 368.045 ;
        RECT 1401.345 367.055 1401.625 367.335 ;
        RECT 1402.055 367.055 1402.335 367.335 ;
        RECT 1402.765 367.055 1403.045 367.335 ;
        RECT 1403.475 367.055 1403.755 367.335 ;
        RECT 1404.185 367.055 1404.465 367.335 ;
        RECT 1404.895 367.055 1405.175 367.335 ;
        RECT 1405.605 367.055 1405.885 367.335 ;
        RECT 1406.315 367.055 1406.595 367.335 ;
        RECT 1407.025 367.055 1407.305 367.335 ;
        RECT 1407.735 367.055 1408.015 367.335 ;
        RECT 1408.445 367.055 1408.725 367.335 ;
        RECT 1409.155 367.055 1409.435 367.335 ;
        RECT 1409.865 367.055 1410.145 367.335 ;
        RECT 1410.575 367.055 1410.855 367.335 ;
        RECT 1401.345 366.345 1401.625 366.625 ;
        RECT 1402.055 366.345 1402.335 366.625 ;
        RECT 1402.765 366.345 1403.045 366.625 ;
        RECT 1403.475 366.345 1403.755 366.625 ;
        RECT 1404.185 366.345 1404.465 366.625 ;
        RECT 1404.895 366.345 1405.175 366.625 ;
        RECT 1405.605 366.345 1405.885 366.625 ;
        RECT 1406.315 366.345 1406.595 366.625 ;
        RECT 1407.025 366.345 1407.305 366.625 ;
        RECT 1407.735 366.345 1408.015 366.625 ;
        RECT 1408.445 366.345 1408.725 366.625 ;
        RECT 1409.155 366.345 1409.435 366.625 ;
        RECT 1409.865 366.345 1410.145 366.625 ;
        RECT 1410.575 366.345 1410.855 366.625 ;
        RECT 1401.345 365.635 1401.625 365.915 ;
        RECT 1402.055 365.635 1402.335 365.915 ;
        RECT 1402.765 365.635 1403.045 365.915 ;
        RECT 1403.475 365.635 1403.755 365.915 ;
        RECT 1404.185 365.635 1404.465 365.915 ;
        RECT 1404.895 365.635 1405.175 365.915 ;
        RECT 1405.605 365.635 1405.885 365.915 ;
        RECT 1406.315 365.635 1406.595 365.915 ;
        RECT 1407.025 365.635 1407.305 365.915 ;
        RECT 1407.735 365.635 1408.015 365.915 ;
        RECT 1408.445 365.635 1408.725 365.915 ;
        RECT 1409.155 365.635 1409.435 365.915 ;
        RECT 1409.865 365.635 1410.145 365.915 ;
        RECT 1410.575 365.635 1410.855 365.915 ;
        RECT 1401.345 364.925 1401.625 365.205 ;
        RECT 1402.055 364.925 1402.335 365.205 ;
        RECT 1402.765 364.925 1403.045 365.205 ;
        RECT 1403.475 364.925 1403.755 365.205 ;
        RECT 1404.185 364.925 1404.465 365.205 ;
        RECT 1404.895 364.925 1405.175 365.205 ;
        RECT 1405.605 364.925 1405.885 365.205 ;
        RECT 1406.315 364.925 1406.595 365.205 ;
        RECT 1407.025 364.925 1407.305 365.205 ;
        RECT 1407.735 364.925 1408.015 365.205 ;
        RECT 1408.445 364.925 1408.725 365.205 ;
        RECT 1409.155 364.925 1409.435 365.205 ;
        RECT 1409.865 364.925 1410.145 365.205 ;
        RECT 1410.575 364.925 1410.855 365.205 ;
        RECT 1401.345 364.215 1401.625 364.495 ;
        RECT 1402.055 364.215 1402.335 364.495 ;
        RECT 1402.765 364.215 1403.045 364.495 ;
        RECT 1403.475 364.215 1403.755 364.495 ;
        RECT 1404.185 364.215 1404.465 364.495 ;
        RECT 1404.895 364.215 1405.175 364.495 ;
        RECT 1405.605 364.215 1405.885 364.495 ;
        RECT 1406.315 364.215 1406.595 364.495 ;
        RECT 1407.025 364.215 1407.305 364.495 ;
        RECT 1407.735 364.215 1408.015 364.495 ;
        RECT 1408.445 364.215 1408.725 364.495 ;
        RECT 1409.155 364.215 1409.435 364.495 ;
        RECT 1409.865 364.215 1410.145 364.495 ;
        RECT 1410.575 364.215 1410.855 364.495 ;
        RECT 1401.345 363.505 1401.625 363.785 ;
        RECT 1402.055 363.505 1402.335 363.785 ;
        RECT 1402.765 363.505 1403.045 363.785 ;
        RECT 1403.475 363.505 1403.755 363.785 ;
        RECT 1404.185 363.505 1404.465 363.785 ;
        RECT 1404.895 363.505 1405.175 363.785 ;
        RECT 1405.605 363.505 1405.885 363.785 ;
        RECT 1406.315 363.505 1406.595 363.785 ;
        RECT 1407.025 363.505 1407.305 363.785 ;
        RECT 1407.735 363.505 1408.015 363.785 ;
        RECT 1408.445 363.505 1408.725 363.785 ;
        RECT 1409.155 363.505 1409.435 363.785 ;
        RECT 1409.865 363.505 1410.145 363.785 ;
        RECT 1410.575 363.505 1410.855 363.785 ;
        RECT 1401.345 362.795 1401.625 363.075 ;
        RECT 1402.055 362.795 1402.335 363.075 ;
        RECT 1402.765 362.795 1403.045 363.075 ;
        RECT 1403.475 362.795 1403.755 363.075 ;
        RECT 1404.185 362.795 1404.465 363.075 ;
        RECT 1404.895 362.795 1405.175 363.075 ;
        RECT 1405.605 362.795 1405.885 363.075 ;
        RECT 1406.315 362.795 1406.595 363.075 ;
        RECT 1407.025 362.795 1407.305 363.075 ;
        RECT 1407.735 362.795 1408.015 363.075 ;
        RECT 1408.445 362.795 1408.725 363.075 ;
        RECT 1409.155 362.795 1409.435 363.075 ;
        RECT 1409.865 362.795 1410.145 363.075 ;
        RECT 1410.575 362.795 1410.855 363.075 ;
        RECT 1401.345 362.085 1401.625 362.365 ;
        RECT 1402.055 362.085 1402.335 362.365 ;
        RECT 1402.765 362.085 1403.045 362.365 ;
        RECT 1403.475 362.085 1403.755 362.365 ;
        RECT 1404.185 362.085 1404.465 362.365 ;
        RECT 1404.895 362.085 1405.175 362.365 ;
        RECT 1405.605 362.085 1405.885 362.365 ;
        RECT 1406.315 362.085 1406.595 362.365 ;
        RECT 1407.025 362.085 1407.305 362.365 ;
        RECT 1407.735 362.085 1408.015 362.365 ;
        RECT 1408.445 362.085 1408.725 362.365 ;
        RECT 1409.155 362.085 1409.435 362.365 ;
        RECT 1409.865 362.085 1410.145 362.365 ;
        RECT 1410.575 362.085 1410.855 362.365 ;
        RECT 1401.345 361.375 1401.625 361.655 ;
        RECT 1402.055 361.375 1402.335 361.655 ;
        RECT 1402.765 361.375 1403.045 361.655 ;
        RECT 1403.475 361.375 1403.755 361.655 ;
        RECT 1404.185 361.375 1404.465 361.655 ;
        RECT 1404.895 361.375 1405.175 361.655 ;
        RECT 1405.605 361.375 1405.885 361.655 ;
        RECT 1406.315 361.375 1406.595 361.655 ;
        RECT 1407.025 361.375 1407.305 361.655 ;
        RECT 1407.735 361.375 1408.015 361.655 ;
        RECT 1408.445 361.375 1408.725 361.655 ;
        RECT 1409.155 361.375 1409.435 361.655 ;
        RECT 1409.865 361.375 1410.145 361.655 ;
        RECT 1410.575 361.375 1410.855 361.655 ;
        RECT 1401.345 360.665 1401.625 360.945 ;
        RECT 1402.055 360.665 1402.335 360.945 ;
        RECT 1402.765 360.665 1403.045 360.945 ;
        RECT 1403.475 360.665 1403.755 360.945 ;
        RECT 1404.185 360.665 1404.465 360.945 ;
        RECT 1404.895 360.665 1405.175 360.945 ;
        RECT 1405.605 360.665 1405.885 360.945 ;
        RECT 1406.315 360.665 1406.595 360.945 ;
        RECT 1407.025 360.665 1407.305 360.945 ;
        RECT 1407.735 360.665 1408.015 360.945 ;
        RECT 1408.445 360.665 1408.725 360.945 ;
        RECT 1409.155 360.665 1409.435 360.945 ;
        RECT 1409.865 360.665 1410.145 360.945 ;
        RECT 1410.575 360.665 1410.855 360.945 ;
        RECT 1414.495 369.895 1414.775 370.175 ;
        RECT 1415.205 369.895 1415.485 370.175 ;
        RECT 1415.915 369.895 1416.195 370.175 ;
        RECT 1416.625 369.895 1416.905 370.175 ;
        RECT 1417.335 369.895 1417.615 370.175 ;
        RECT 1418.045 369.895 1418.325 370.175 ;
        RECT 1418.755 369.895 1419.035 370.175 ;
        RECT 1419.465 369.895 1419.745 370.175 ;
        RECT 1414.495 369.185 1414.775 369.465 ;
        RECT 1415.205 369.185 1415.485 369.465 ;
        RECT 1415.915 369.185 1416.195 369.465 ;
        RECT 1416.625 369.185 1416.905 369.465 ;
        RECT 1417.335 369.185 1417.615 369.465 ;
        RECT 1418.045 369.185 1418.325 369.465 ;
        RECT 1418.755 369.185 1419.035 369.465 ;
        RECT 1419.465 369.185 1419.745 369.465 ;
        RECT 1414.495 368.475 1414.775 368.755 ;
        RECT 1415.205 368.475 1415.485 368.755 ;
        RECT 1415.915 368.475 1416.195 368.755 ;
        RECT 1416.625 368.475 1416.905 368.755 ;
        RECT 1417.335 368.475 1417.615 368.755 ;
        RECT 1418.045 368.475 1418.325 368.755 ;
        RECT 1418.755 368.475 1419.035 368.755 ;
        RECT 1419.465 368.475 1419.745 368.755 ;
        RECT 1414.495 367.765 1414.775 368.045 ;
        RECT 1415.205 367.765 1415.485 368.045 ;
        RECT 1415.915 367.765 1416.195 368.045 ;
        RECT 1416.625 367.765 1416.905 368.045 ;
        RECT 1417.335 367.765 1417.615 368.045 ;
        RECT 1418.045 367.765 1418.325 368.045 ;
        RECT 1418.755 367.765 1419.035 368.045 ;
        RECT 1419.465 367.765 1419.745 368.045 ;
        RECT 1414.495 367.055 1414.775 367.335 ;
        RECT 1415.205 367.055 1415.485 367.335 ;
        RECT 1415.915 367.055 1416.195 367.335 ;
        RECT 1416.625 367.055 1416.905 367.335 ;
        RECT 1417.335 367.055 1417.615 367.335 ;
        RECT 1418.045 367.055 1418.325 367.335 ;
        RECT 1418.755 367.055 1419.035 367.335 ;
        RECT 1419.465 367.055 1419.745 367.335 ;
        RECT 1414.495 366.345 1414.775 366.625 ;
        RECT 1415.205 366.345 1415.485 366.625 ;
        RECT 1415.915 366.345 1416.195 366.625 ;
        RECT 1416.625 366.345 1416.905 366.625 ;
        RECT 1417.335 366.345 1417.615 366.625 ;
        RECT 1418.045 366.345 1418.325 366.625 ;
        RECT 1418.755 366.345 1419.035 366.625 ;
        RECT 1419.465 366.345 1419.745 366.625 ;
        RECT 1414.495 365.635 1414.775 365.915 ;
        RECT 1415.205 365.635 1415.485 365.915 ;
        RECT 1415.915 365.635 1416.195 365.915 ;
        RECT 1416.625 365.635 1416.905 365.915 ;
        RECT 1417.335 365.635 1417.615 365.915 ;
        RECT 1418.045 365.635 1418.325 365.915 ;
        RECT 1418.755 365.635 1419.035 365.915 ;
        RECT 1419.465 365.635 1419.745 365.915 ;
        RECT 1414.495 364.925 1414.775 365.205 ;
        RECT 1415.205 364.925 1415.485 365.205 ;
        RECT 1415.915 364.925 1416.195 365.205 ;
        RECT 1416.625 364.925 1416.905 365.205 ;
        RECT 1417.335 364.925 1417.615 365.205 ;
        RECT 1418.045 364.925 1418.325 365.205 ;
        RECT 1418.755 364.925 1419.035 365.205 ;
        RECT 1419.465 364.925 1419.745 365.205 ;
        RECT 1414.495 364.215 1414.775 364.495 ;
        RECT 1415.205 364.215 1415.485 364.495 ;
        RECT 1415.915 364.215 1416.195 364.495 ;
        RECT 1416.625 364.215 1416.905 364.495 ;
        RECT 1417.335 364.215 1417.615 364.495 ;
        RECT 1418.045 364.215 1418.325 364.495 ;
        RECT 1418.755 364.215 1419.035 364.495 ;
        RECT 1419.465 364.215 1419.745 364.495 ;
        RECT 1414.495 363.505 1414.775 363.785 ;
        RECT 1415.205 363.505 1415.485 363.785 ;
        RECT 1415.915 363.505 1416.195 363.785 ;
        RECT 1416.625 363.505 1416.905 363.785 ;
        RECT 1417.335 363.505 1417.615 363.785 ;
        RECT 1418.045 363.505 1418.325 363.785 ;
        RECT 1418.755 363.505 1419.035 363.785 ;
        RECT 1419.465 363.505 1419.745 363.785 ;
        RECT 1414.495 362.795 1414.775 363.075 ;
        RECT 1415.205 362.795 1415.485 363.075 ;
        RECT 1415.915 362.795 1416.195 363.075 ;
        RECT 1416.625 362.795 1416.905 363.075 ;
        RECT 1417.335 362.795 1417.615 363.075 ;
        RECT 1418.045 362.795 1418.325 363.075 ;
        RECT 1418.755 362.795 1419.035 363.075 ;
        RECT 1419.465 362.795 1419.745 363.075 ;
        RECT 1414.495 362.085 1414.775 362.365 ;
        RECT 1415.205 362.085 1415.485 362.365 ;
        RECT 1415.915 362.085 1416.195 362.365 ;
        RECT 1416.625 362.085 1416.905 362.365 ;
        RECT 1417.335 362.085 1417.615 362.365 ;
        RECT 1418.045 362.085 1418.325 362.365 ;
        RECT 1418.755 362.085 1419.035 362.365 ;
        RECT 1419.465 362.085 1419.745 362.365 ;
        RECT 1414.495 361.375 1414.775 361.655 ;
        RECT 1415.205 361.375 1415.485 361.655 ;
        RECT 1415.915 361.375 1416.195 361.655 ;
        RECT 1416.625 361.375 1416.905 361.655 ;
        RECT 1417.335 361.375 1417.615 361.655 ;
        RECT 1418.045 361.375 1418.325 361.655 ;
        RECT 1418.755 361.375 1419.035 361.655 ;
        RECT 1419.465 361.375 1419.745 361.655 ;
        RECT 1414.495 360.665 1414.775 360.945 ;
        RECT 1415.205 360.665 1415.485 360.945 ;
        RECT 1415.915 360.665 1416.195 360.945 ;
        RECT 1416.625 360.665 1416.905 360.945 ;
        RECT 1417.335 360.665 1417.615 360.945 ;
        RECT 1418.045 360.665 1418.325 360.945 ;
        RECT 1418.755 360.665 1419.035 360.945 ;
        RECT 1419.465 360.665 1419.745 360.945 ;
        RECT 3001.715 369.895 3001.995 370.175 ;
        RECT 3002.425 369.895 3002.705 370.175 ;
        RECT 3003.135 369.895 3003.415 370.175 ;
        RECT 3003.845 369.895 3004.125 370.175 ;
        RECT 3004.555 369.895 3004.835 370.175 ;
        RECT 3005.265 369.895 3005.545 370.175 ;
        RECT 3005.975 369.895 3006.255 370.175 ;
        RECT 3006.685 369.895 3006.965 370.175 ;
        RECT 3007.395 369.895 3007.675 370.175 ;
        RECT 3008.105 369.895 3008.385 370.175 ;
        RECT 3008.815 369.895 3009.095 370.175 ;
        RECT 3009.525 369.895 3009.805 370.175 ;
        RECT 3010.235 369.895 3010.515 370.175 ;
        RECT 3001.715 369.185 3001.995 369.465 ;
        RECT 3002.425 369.185 3002.705 369.465 ;
        RECT 3003.135 369.185 3003.415 369.465 ;
        RECT 3003.845 369.185 3004.125 369.465 ;
        RECT 3004.555 369.185 3004.835 369.465 ;
        RECT 3005.265 369.185 3005.545 369.465 ;
        RECT 3005.975 369.185 3006.255 369.465 ;
        RECT 3006.685 369.185 3006.965 369.465 ;
        RECT 3007.395 369.185 3007.675 369.465 ;
        RECT 3008.105 369.185 3008.385 369.465 ;
        RECT 3008.815 369.185 3009.095 369.465 ;
        RECT 3009.525 369.185 3009.805 369.465 ;
        RECT 3010.235 369.185 3010.515 369.465 ;
        RECT 3001.715 368.475 3001.995 368.755 ;
        RECT 3002.425 368.475 3002.705 368.755 ;
        RECT 3003.135 368.475 3003.415 368.755 ;
        RECT 3003.845 368.475 3004.125 368.755 ;
        RECT 3004.555 368.475 3004.835 368.755 ;
        RECT 3005.265 368.475 3005.545 368.755 ;
        RECT 3005.975 368.475 3006.255 368.755 ;
        RECT 3006.685 368.475 3006.965 368.755 ;
        RECT 3007.395 368.475 3007.675 368.755 ;
        RECT 3008.105 368.475 3008.385 368.755 ;
        RECT 3008.815 368.475 3009.095 368.755 ;
        RECT 3009.525 368.475 3009.805 368.755 ;
        RECT 3010.235 368.475 3010.515 368.755 ;
        RECT 3001.715 367.765 3001.995 368.045 ;
        RECT 3002.425 367.765 3002.705 368.045 ;
        RECT 3003.135 367.765 3003.415 368.045 ;
        RECT 3003.845 367.765 3004.125 368.045 ;
        RECT 3004.555 367.765 3004.835 368.045 ;
        RECT 3005.265 367.765 3005.545 368.045 ;
        RECT 3005.975 367.765 3006.255 368.045 ;
        RECT 3006.685 367.765 3006.965 368.045 ;
        RECT 3007.395 367.765 3007.675 368.045 ;
        RECT 3008.105 367.765 3008.385 368.045 ;
        RECT 3008.815 367.765 3009.095 368.045 ;
        RECT 3009.525 367.765 3009.805 368.045 ;
        RECT 3010.235 367.765 3010.515 368.045 ;
        RECT 3001.715 367.055 3001.995 367.335 ;
        RECT 3002.425 367.055 3002.705 367.335 ;
        RECT 3003.135 367.055 3003.415 367.335 ;
        RECT 3003.845 367.055 3004.125 367.335 ;
        RECT 3004.555 367.055 3004.835 367.335 ;
        RECT 3005.265 367.055 3005.545 367.335 ;
        RECT 3005.975 367.055 3006.255 367.335 ;
        RECT 3006.685 367.055 3006.965 367.335 ;
        RECT 3007.395 367.055 3007.675 367.335 ;
        RECT 3008.105 367.055 3008.385 367.335 ;
        RECT 3008.815 367.055 3009.095 367.335 ;
        RECT 3009.525 367.055 3009.805 367.335 ;
        RECT 3010.235 367.055 3010.515 367.335 ;
        RECT 3001.715 366.345 3001.995 366.625 ;
        RECT 3002.425 366.345 3002.705 366.625 ;
        RECT 3003.135 366.345 3003.415 366.625 ;
        RECT 3003.845 366.345 3004.125 366.625 ;
        RECT 3004.555 366.345 3004.835 366.625 ;
        RECT 3005.265 366.345 3005.545 366.625 ;
        RECT 3005.975 366.345 3006.255 366.625 ;
        RECT 3006.685 366.345 3006.965 366.625 ;
        RECT 3007.395 366.345 3007.675 366.625 ;
        RECT 3008.105 366.345 3008.385 366.625 ;
        RECT 3008.815 366.345 3009.095 366.625 ;
        RECT 3009.525 366.345 3009.805 366.625 ;
        RECT 3010.235 366.345 3010.515 366.625 ;
        RECT 3001.715 365.635 3001.995 365.915 ;
        RECT 3002.425 365.635 3002.705 365.915 ;
        RECT 3003.135 365.635 3003.415 365.915 ;
        RECT 3003.845 365.635 3004.125 365.915 ;
        RECT 3004.555 365.635 3004.835 365.915 ;
        RECT 3005.265 365.635 3005.545 365.915 ;
        RECT 3005.975 365.635 3006.255 365.915 ;
        RECT 3006.685 365.635 3006.965 365.915 ;
        RECT 3007.395 365.635 3007.675 365.915 ;
        RECT 3008.105 365.635 3008.385 365.915 ;
        RECT 3008.815 365.635 3009.095 365.915 ;
        RECT 3009.525 365.635 3009.805 365.915 ;
        RECT 3010.235 365.635 3010.515 365.915 ;
        RECT 3001.715 364.925 3001.995 365.205 ;
        RECT 3002.425 364.925 3002.705 365.205 ;
        RECT 3003.135 364.925 3003.415 365.205 ;
        RECT 3003.845 364.925 3004.125 365.205 ;
        RECT 3004.555 364.925 3004.835 365.205 ;
        RECT 3005.265 364.925 3005.545 365.205 ;
        RECT 3005.975 364.925 3006.255 365.205 ;
        RECT 3006.685 364.925 3006.965 365.205 ;
        RECT 3007.395 364.925 3007.675 365.205 ;
        RECT 3008.105 364.925 3008.385 365.205 ;
        RECT 3008.815 364.925 3009.095 365.205 ;
        RECT 3009.525 364.925 3009.805 365.205 ;
        RECT 3010.235 364.925 3010.515 365.205 ;
        RECT 3001.715 364.215 3001.995 364.495 ;
        RECT 3002.425 364.215 3002.705 364.495 ;
        RECT 3003.135 364.215 3003.415 364.495 ;
        RECT 3003.845 364.215 3004.125 364.495 ;
        RECT 3004.555 364.215 3004.835 364.495 ;
        RECT 3005.265 364.215 3005.545 364.495 ;
        RECT 3005.975 364.215 3006.255 364.495 ;
        RECT 3006.685 364.215 3006.965 364.495 ;
        RECT 3007.395 364.215 3007.675 364.495 ;
        RECT 3008.105 364.215 3008.385 364.495 ;
        RECT 3008.815 364.215 3009.095 364.495 ;
        RECT 3009.525 364.215 3009.805 364.495 ;
        RECT 3010.235 364.215 3010.515 364.495 ;
        RECT 3001.715 363.505 3001.995 363.785 ;
        RECT 3002.425 363.505 3002.705 363.785 ;
        RECT 3003.135 363.505 3003.415 363.785 ;
        RECT 3003.845 363.505 3004.125 363.785 ;
        RECT 3004.555 363.505 3004.835 363.785 ;
        RECT 3005.265 363.505 3005.545 363.785 ;
        RECT 3005.975 363.505 3006.255 363.785 ;
        RECT 3006.685 363.505 3006.965 363.785 ;
        RECT 3007.395 363.505 3007.675 363.785 ;
        RECT 3008.105 363.505 3008.385 363.785 ;
        RECT 3008.815 363.505 3009.095 363.785 ;
        RECT 3009.525 363.505 3009.805 363.785 ;
        RECT 3010.235 363.505 3010.515 363.785 ;
        RECT 3001.715 362.795 3001.995 363.075 ;
        RECT 3002.425 362.795 3002.705 363.075 ;
        RECT 3003.135 362.795 3003.415 363.075 ;
        RECT 3003.845 362.795 3004.125 363.075 ;
        RECT 3004.555 362.795 3004.835 363.075 ;
        RECT 3005.265 362.795 3005.545 363.075 ;
        RECT 3005.975 362.795 3006.255 363.075 ;
        RECT 3006.685 362.795 3006.965 363.075 ;
        RECT 3007.395 362.795 3007.675 363.075 ;
        RECT 3008.105 362.795 3008.385 363.075 ;
        RECT 3008.815 362.795 3009.095 363.075 ;
        RECT 3009.525 362.795 3009.805 363.075 ;
        RECT 3010.235 362.795 3010.515 363.075 ;
        RECT 3001.715 362.085 3001.995 362.365 ;
        RECT 3002.425 362.085 3002.705 362.365 ;
        RECT 3003.135 362.085 3003.415 362.365 ;
        RECT 3003.845 362.085 3004.125 362.365 ;
        RECT 3004.555 362.085 3004.835 362.365 ;
        RECT 3005.265 362.085 3005.545 362.365 ;
        RECT 3005.975 362.085 3006.255 362.365 ;
        RECT 3006.685 362.085 3006.965 362.365 ;
        RECT 3007.395 362.085 3007.675 362.365 ;
        RECT 3008.105 362.085 3008.385 362.365 ;
        RECT 3008.815 362.085 3009.095 362.365 ;
        RECT 3009.525 362.085 3009.805 362.365 ;
        RECT 3010.235 362.085 3010.515 362.365 ;
        RECT 3001.715 361.375 3001.995 361.655 ;
        RECT 3002.425 361.375 3002.705 361.655 ;
        RECT 3003.135 361.375 3003.415 361.655 ;
        RECT 3003.845 361.375 3004.125 361.655 ;
        RECT 3004.555 361.375 3004.835 361.655 ;
        RECT 3005.265 361.375 3005.545 361.655 ;
        RECT 3005.975 361.375 3006.255 361.655 ;
        RECT 3006.685 361.375 3006.965 361.655 ;
        RECT 3007.395 361.375 3007.675 361.655 ;
        RECT 3008.105 361.375 3008.385 361.655 ;
        RECT 3008.815 361.375 3009.095 361.655 ;
        RECT 3009.525 361.375 3009.805 361.655 ;
        RECT 3010.235 361.375 3010.515 361.655 ;
        RECT 3001.715 360.665 3001.995 360.945 ;
        RECT 3002.425 360.665 3002.705 360.945 ;
        RECT 3003.135 360.665 3003.415 360.945 ;
        RECT 3003.845 360.665 3004.125 360.945 ;
        RECT 3004.555 360.665 3004.835 360.945 ;
        RECT 3005.265 360.665 3005.545 360.945 ;
        RECT 3005.975 360.665 3006.255 360.945 ;
        RECT 3006.685 360.665 3006.965 360.945 ;
        RECT 3007.395 360.665 3007.675 360.945 ;
        RECT 3008.105 360.665 3008.385 360.945 ;
        RECT 3008.815 360.665 3009.095 360.945 ;
        RECT 3009.525 360.665 3009.805 360.945 ;
        RECT 3010.235 360.665 3010.515 360.945 ;
        RECT 3014.115 369.895 3014.395 370.175 ;
        RECT 3014.825 369.895 3015.105 370.175 ;
        RECT 3015.535 369.895 3015.815 370.175 ;
        RECT 3016.245 369.895 3016.525 370.175 ;
        RECT 3016.955 369.895 3017.235 370.175 ;
        RECT 3017.665 369.895 3017.945 370.175 ;
        RECT 3018.375 369.895 3018.655 370.175 ;
        RECT 3019.085 369.895 3019.365 370.175 ;
        RECT 3019.795 369.895 3020.075 370.175 ;
        RECT 3014.115 369.185 3014.395 369.465 ;
        RECT 3014.825 369.185 3015.105 369.465 ;
        RECT 3015.535 369.185 3015.815 369.465 ;
        RECT 3016.245 369.185 3016.525 369.465 ;
        RECT 3016.955 369.185 3017.235 369.465 ;
        RECT 3017.665 369.185 3017.945 369.465 ;
        RECT 3018.375 369.185 3018.655 369.465 ;
        RECT 3019.085 369.185 3019.365 369.465 ;
        RECT 3019.795 369.185 3020.075 369.465 ;
        RECT 3014.115 368.475 3014.395 368.755 ;
        RECT 3014.825 368.475 3015.105 368.755 ;
        RECT 3015.535 368.475 3015.815 368.755 ;
        RECT 3016.245 368.475 3016.525 368.755 ;
        RECT 3016.955 368.475 3017.235 368.755 ;
        RECT 3017.665 368.475 3017.945 368.755 ;
        RECT 3018.375 368.475 3018.655 368.755 ;
        RECT 3019.085 368.475 3019.365 368.755 ;
        RECT 3019.795 368.475 3020.075 368.755 ;
        RECT 3014.115 367.765 3014.395 368.045 ;
        RECT 3014.825 367.765 3015.105 368.045 ;
        RECT 3015.535 367.765 3015.815 368.045 ;
        RECT 3016.245 367.765 3016.525 368.045 ;
        RECT 3016.955 367.765 3017.235 368.045 ;
        RECT 3017.665 367.765 3017.945 368.045 ;
        RECT 3018.375 367.765 3018.655 368.045 ;
        RECT 3019.085 367.765 3019.365 368.045 ;
        RECT 3019.795 367.765 3020.075 368.045 ;
        RECT 3014.115 367.055 3014.395 367.335 ;
        RECT 3014.825 367.055 3015.105 367.335 ;
        RECT 3015.535 367.055 3015.815 367.335 ;
        RECT 3016.245 367.055 3016.525 367.335 ;
        RECT 3016.955 367.055 3017.235 367.335 ;
        RECT 3017.665 367.055 3017.945 367.335 ;
        RECT 3018.375 367.055 3018.655 367.335 ;
        RECT 3019.085 367.055 3019.365 367.335 ;
        RECT 3019.795 367.055 3020.075 367.335 ;
        RECT 3014.115 366.345 3014.395 366.625 ;
        RECT 3014.825 366.345 3015.105 366.625 ;
        RECT 3015.535 366.345 3015.815 366.625 ;
        RECT 3016.245 366.345 3016.525 366.625 ;
        RECT 3016.955 366.345 3017.235 366.625 ;
        RECT 3017.665 366.345 3017.945 366.625 ;
        RECT 3018.375 366.345 3018.655 366.625 ;
        RECT 3019.085 366.345 3019.365 366.625 ;
        RECT 3019.795 366.345 3020.075 366.625 ;
        RECT 3014.115 365.635 3014.395 365.915 ;
        RECT 3014.825 365.635 3015.105 365.915 ;
        RECT 3015.535 365.635 3015.815 365.915 ;
        RECT 3016.245 365.635 3016.525 365.915 ;
        RECT 3016.955 365.635 3017.235 365.915 ;
        RECT 3017.665 365.635 3017.945 365.915 ;
        RECT 3018.375 365.635 3018.655 365.915 ;
        RECT 3019.085 365.635 3019.365 365.915 ;
        RECT 3019.795 365.635 3020.075 365.915 ;
        RECT 3014.115 364.925 3014.395 365.205 ;
        RECT 3014.825 364.925 3015.105 365.205 ;
        RECT 3015.535 364.925 3015.815 365.205 ;
        RECT 3016.245 364.925 3016.525 365.205 ;
        RECT 3016.955 364.925 3017.235 365.205 ;
        RECT 3017.665 364.925 3017.945 365.205 ;
        RECT 3018.375 364.925 3018.655 365.205 ;
        RECT 3019.085 364.925 3019.365 365.205 ;
        RECT 3019.795 364.925 3020.075 365.205 ;
        RECT 3014.115 364.215 3014.395 364.495 ;
        RECT 3014.825 364.215 3015.105 364.495 ;
        RECT 3015.535 364.215 3015.815 364.495 ;
        RECT 3016.245 364.215 3016.525 364.495 ;
        RECT 3016.955 364.215 3017.235 364.495 ;
        RECT 3017.665 364.215 3017.945 364.495 ;
        RECT 3018.375 364.215 3018.655 364.495 ;
        RECT 3019.085 364.215 3019.365 364.495 ;
        RECT 3019.795 364.215 3020.075 364.495 ;
        RECT 3014.115 363.505 3014.395 363.785 ;
        RECT 3014.825 363.505 3015.105 363.785 ;
        RECT 3015.535 363.505 3015.815 363.785 ;
        RECT 3016.245 363.505 3016.525 363.785 ;
        RECT 3016.955 363.505 3017.235 363.785 ;
        RECT 3017.665 363.505 3017.945 363.785 ;
        RECT 3018.375 363.505 3018.655 363.785 ;
        RECT 3019.085 363.505 3019.365 363.785 ;
        RECT 3019.795 363.505 3020.075 363.785 ;
        RECT 3014.115 362.795 3014.395 363.075 ;
        RECT 3014.825 362.795 3015.105 363.075 ;
        RECT 3015.535 362.795 3015.815 363.075 ;
        RECT 3016.245 362.795 3016.525 363.075 ;
        RECT 3016.955 362.795 3017.235 363.075 ;
        RECT 3017.665 362.795 3017.945 363.075 ;
        RECT 3018.375 362.795 3018.655 363.075 ;
        RECT 3019.085 362.795 3019.365 363.075 ;
        RECT 3019.795 362.795 3020.075 363.075 ;
        RECT 3014.115 362.085 3014.395 362.365 ;
        RECT 3014.825 362.085 3015.105 362.365 ;
        RECT 3015.535 362.085 3015.815 362.365 ;
        RECT 3016.245 362.085 3016.525 362.365 ;
        RECT 3016.955 362.085 3017.235 362.365 ;
        RECT 3017.665 362.085 3017.945 362.365 ;
        RECT 3018.375 362.085 3018.655 362.365 ;
        RECT 3019.085 362.085 3019.365 362.365 ;
        RECT 3019.795 362.085 3020.075 362.365 ;
        RECT 3014.115 361.375 3014.395 361.655 ;
        RECT 3014.825 361.375 3015.105 361.655 ;
        RECT 3015.535 361.375 3015.815 361.655 ;
        RECT 3016.245 361.375 3016.525 361.655 ;
        RECT 3016.955 361.375 3017.235 361.655 ;
        RECT 3017.665 361.375 3017.945 361.655 ;
        RECT 3018.375 361.375 3018.655 361.655 ;
        RECT 3019.085 361.375 3019.365 361.655 ;
        RECT 3019.795 361.375 3020.075 361.655 ;
        RECT 3014.115 360.665 3014.395 360.945 ;
        RECT 3014.825 360.665 3015.105 360.945 ;
        RECT 3015.535 360.665 3015.815 360.945 ;
        RECT 3016.245 360.665 3016.525 360.945 ;
        RECT 3016.955 360.665 3017.235 360.945 ;
        RECT 3017.665 360.665 3017.945 360.945 ;
        RECT 3018.375 360.665 3018.655 360.945 ;
        RECT 3019.085 360.665 3019.365 360.945 ;
        RECT 3019.795 360.665 3020.075 360.945 ;
        RECT 3025.965 369.895 3026.245 370.175 ;
        RECT 3026.675 369.895 3026.955 370.175 ;
        RECT 3027.385 369.895 3027.665 370.175 ;
        RECT 3028.095 369.895 3028.375 370.175 ;
        RECT 3028.805 369.895 3029.085 370.175 ;
        RECT 3029.515 369.895 3029.795 370.175 ;
        RECT 3030.225 369.895 3030.505 370.175 ;
        RECT 3030.935 369.895 3031.215 370.175 ;
        RECT 3031.645 369.895 3031.925 370.175 ;
        RECT 3032.355 369.895 3032.635 370.175 ;
        RECT 3033.065 369.895 3033.345 370.175 ;
        RECT 3033.775 369.895 3034.055 370.175 ;
        RECT 3034.485 369.895 3034.765 370.175 ;
        RECT 3035.195 369.895 3035.475 370.175 ;
        RECT 3025.965 369.185 3026.245 369.465 ;
        RECT 3026.675 369.185 3026.955 369.465 ;
        RECT 3027.385 369.185 3027.665 369.465 ;
        RECT 3028.095 369.185 3028.375 369.465 ;
        RECT 3028.805 369.185 3029.085 369.465 ;
        RECT 3029.515 369.185 3029.795 369.465 ;
        RECT 3030.225 369.185 3030.505 369.465 ;
        RECT 3030.935 369.185 3031.215 369.465 ;
        RECT 3031.645 369.185 3031.925 369.465 ;
        RECT 3032.355 369.185 3032.635 369.465 ;
        RECT 3033.065 369.185 3033.345 369.465 ;
        RECT 3033.775 369.185 3034.055 369.465 ;
        RECT 3034.485 369.185 3034.765 369.465 ;
        RECT 3035.195 369.185 3035.475 369.465 ;
        RECT 3025.965 368.475 3026.245 368.755 ;
        RECT 3026.675 368.475 3026.955 368.755 ;
        RECT 3027.385 368.475 3027.665 368.755 ;
        RECT 3028.095 368.475 3028.375 368.755 ;
        RECT 3028.805 368.475 3029.085 368.755 ;
        RECT 3029.515 368.475 3029.795 368.755 ;
        RECT 3030.225 368.475 3030.505 368.755 ;
        RECT 3030.935 368.475 3031.215 368.755 ;
        RECT 3031.645 368.475 3031.925 368.755 ;
        RECT 3032.355 368.475 3032.635 368.755 ;
        RECT 3033.065 368.475 3033.345 368.755 ;
        RECT 3033.775 368.475 3034.055 368.755 ;
        RECT 3034.485 368.475 3034.765 368.755 ;
        RECT 3035.195 368.475 3035.475 368.755 ;
        RECT 3025.965 367.765 3026.245 368.045 ;
        RECT 3026.675 367.765 3026.955 368.045 ;
        RECT 3027.385 367.765 3027.665 368.045 ;
        RECT 3028.095 367.765 3028.375 368.045 ;
        RECT 3028.805 367.765 3029.085 368.045 ;
        RECT 3029.515 367.765 3029.795 368.045 ;
        RECT 3030.225 367.765 3030.505 368.045 ;
        RECT 3030.935 367.765 3031.215 368.045 ;
        RECT 3031.645 367.765 3031.925 368.045 ;
        RECT 3032.355 367.765 3032.635 368.045 ;
        RECT 3033.065 367.765 3033.345 368.045 ;
        RECT 3033.775 367.765 3034.055 368.045 ;
        RECT 3034.485 367.765 3034.765 368.045 ;
        RECT 3035.195 367.765 3035.475 368.045 ;
        RECT 3025.965 367.055 3026.245 367.335 ;
        RECT 3026.675 367.055 3026.955 367.335 ;
        RECT 3027.385 367.055 3027.665 367.335 ;
        RECT 3028.095 367.055 3028.375 367.335 ;
        RECT 3028.805 367.055 3029.085 367.335 ;
        RECT 3029.515 367.055 3029.795 367.335 ;
        RECT 3030.225 367.055 3030.505 367.335 ;
        RECT 3030.935 367.055 3031.215 367.335 ;
        RECT 3031.645 367.055 3031.925 367.335 ;
        RECT 3032.355 367.055 3032.635 367.335 ;
        RECT 3033.065 367.055 3033.345 367.335 ;
        RECT 3033.775 367.055 3034.055 367.335 ;
        RECT 3034.485 367.055 3034.765 367.335 ;
        RECT 3035.195 367.055 3035.475 367.335 ;
        RECT 3025.965 366.345 3026.245 366.625 ;
        RECT 3026.675 366.345 3026.955 366.625 ;
        RECT 3027.385 366.345 3027.665 366.625 ;
        RECT 3028.095 366.345 3028.375 366.625 ;
        RECT 3028.805 366.345 3029.085 366.625 ;
        RECT 3029.515 366.345 3029.795 366.625 ;
        RECT 3030.225 366.345 3030.505 366.625 ;
        RECT 3030.935 366.345 3031.215 366.625 ;
        RECT 3031.645 366.345 3031.925 366.625 ;
        RECT 3032.355 366.345 3032.635 366.625 ;
        RECT 3033.065 366.345 3033.345 366.625 ;
        RECT 3033.775 366.345 3034.055 366.625 ;
        RECT 3034.485 366.345 3034.765 366.625 ;
        RECT 3035.195 366.345 3035.475 366.625 ;
        RECT 3025.965 365.635 3026.245 365.915 ;
        RECT 3026.675 365.635 3026.955 365.915 ;
        RECT 3027.385 365.635 3027.665 365.915 ;
        RECT 3028.095 365.635 3028.375 365.915 ;
        RECT 3028.805 365.635 3029.085 365.915 ;
        RECT 3029.515 365.635 3029.795 365.915 ;
        RECT 3030.225 365.635 3030.505 365.915 ;
        RECT 3030.935 365.635 3031.215 365.915 ;
        RECT 3031.645 365.635 3031.925 365.915 ;
        RECT 3032.355 365.635 3032.635 365.915 ;
        RECT 3033.065 365.635 3033.345 365.915 ;
        RECT 3033.775 365.635 3034.055 365.915 ;
        RECT 3034.485 365.635 3034.765 365.915 ;
        RECT 3035.195 365.635 3035.475 365.915 ;
        RECT 3025.965 364.925 3026.245 365.205 ;
        RECT 3026.675 364.925 3026.955 365.205 ;
        RECT 3027.385 364.925 3027.665 365.205 ;
        RECT 3028.095 364.925 3028.375 365.205 ;
        RECT 3028.805 364.925 3029.085 365.205 ;
        RECT 3029.515 364.925 3029.795 365.205 ;
        RECT 3030.225 364.925 3030.505 365.205 ;
        RECT 3030.935 364.925 3031.215 365.205 ;
        RECT 3031.645 364.925 3031.925 365.205 ;
        RECT 3032.355 364.925 3032.635 365.205 ;
        RECT 3033.065 364.925 3033.345 365.205 ;
        RECT 3033.775 364.925 3034.055 365.205 ;
        RECT 3034.485 364.925 3034.765 365.205 ;
        RECT 3035.195 364.925 3035.475 365.205 ;
        RECT 3025.965 364.215 3026.245 364.495 ;
        RECT 3026.675 364.215 3026.955 364.495 ;
        RECT 3027.385 364.215 3027.665 364.495 ;
        RECT 3028.095 364.215 3028.375 364.495 ;
        RECT 3028.805 364.215 3029.085 364.495 ;
        RECT 3029.515 364.215 3029.795 364.495 ;
        RECT 3030.225 364.215 3030.505 364.495 ;
        RECT 3030.935 364.215 3031.215 364.495 ;
        RECT 3031.645 364.215 3031.925 364.495 ;
        RECT 3032.355 364.215 3032.635 364.495 ;
        RECT 3033.065 364.215 3033.345 364.495 ;
        RECT 3033.775 364.215 3034.055 364.495 ;
        RECT 3034.485 364.215 3034.765 364.495 ;
        RECT 3035.195 364.215 3035.475 364.495 ;
        RECT 3025.965 363.505 3026.245 363.785 ;
        RECT 3026.675 363.505 3026.955 363.785 ;
        RECT 3027.385 363.505 3027.665 363.785 ;
        RECT 3028.095 363.505 3028.375 363.785 ;
        RECT 3028.805 363.505 3029.085 363.785 ;
        RECT 3029.515 363.505 3029.795 363.785 ;
        RECT 3030.225 363.505 3030.505 363.785 ;
        RECT 3030.935 363.505 3031.215 363.785 ;
        RECT 3031.645 363.505 3031.925 363.785 ;
        RECT 3032.355 363.505 3032.635 363.785 ;
        RECT 3033.065 363.505 3033.345 363.785 ;
        RECT 3033.775 363.505 3034.055 363.785 ;
        RECT 3034.485 363.505 3034.765 363.785 ;
        RECT 3035.195 363.505 3035.475 363.785 ;
        RECT 3025.965 362.795 3026.245 363.075 ;
        RECT 3026.675 362.795 3026.955 363.075 ;
        RECT 3027.385 362.795 3027.665 363.075 ;
        RECT 3028.095 362.795 3028.375 363.075 ;
        RECT 3028.805 362.795 3029.085 363.075 ;
        RECT 3029.515 362.795 3029.795 363.075 ;
        RECT 3030.225 362.795 3030.505 363.075 ;
        RECT 3030.935 362.795 3031.215 363.075 ;
        RECT 3031.645 362.795 3031.925 363.075 ;
        RECT 3032.355 362.795 3032.635 363.075 ;
        RECT 3033.065 362.795 3033.345 363.075 ;
        RECT 3033.775 362.795 3034.055 363.075 ;
        RECT 3034.485 362.795 3034.765 363.075 ;
        RECT 3035.195 362.795 3035.475 363.075 ;
        RECT 3025.965 362.085 3026.245 362.365 ;
        RECT 3026.675 362.085 3026.955 362.365 ;
        RECT 3027.385 362.085 3027.665 362.365 ;
        RECT 3028.095 362.085 3028.375 362.365 ;
        RECT 3028.805 362.085 3029.085 362.365 ;
        RECT 3029.515 362.085 3029.795 362.365 ;
        RECT 3030.225 362.085 3030.505 362.365 ;
        RECT 3030.935 362.085 3031.215 362.365 ;
        RECT 3031.645 362.085 3031.925 362.365 ;
        RECT 3032.355 362.085 3032.635 362.365 ;
        RECT 3033.065 362.085 3033.345 362.365 ;
        RECT 3033.775 362.085 3034.055 362.365 ;
        RECT 3034.485 362.085 3034.765 362.365 ;
        RECT 3035.195 362.085 3035.475 362.365 ;
        RECT 3025.965 361.375 3026.245 361.655 ;
        RECT 3026.675 361.375 3026.955 361.655 ;
        RECT 3027.385 361.375 3027.665 361.655 ;
        RECT 3028.095 361.375 3028.375 361.655 ;
        RECT 3028.805 361.375 3029.085 361.655 ;
        RECT 3029.515 361.375 3029.795 361.655 ;
        RECT 3030.225 361.375 3030.505 361.655 ;
        RECT 3030.935 361.375 3031.215 361.655 ;
        RECT 3031.645 361.375 3031.925 361.655 ;
        RECT 3032.355 361.375 3032.635 361.655 ;
        RECT 3033.065 361.375 3033.345 361.655 ;
        RECT 3033.775 361.375 3034.055 361.655 ;
        RECT 3034.485 361.375 3034.765 361.655 ;
        RECT 3035.195 361.375 3035.475 361.655 ;
        RECT 3025.965 360.665 3026.245 360.945 ;
        RECT 3026.675 360.665 3026.955 360.945 ;
        RECT 3027.385 360.665 3027.665 360.945 ;
        RECT 3028.095 360.665 3028.375 360.945 ;
        RECT 3028.805 360.665 3029.085 360.945 ;
        RECT 3029.515 360.665 3029.795 360.945 ;
        RECT 3030.225 360.665 3030.505 360.945 ;
        RECT 3030.935 360.665 3031.215 360.945 ;
        RECT 3031.645 360.665 3031.925 360.945 ;
        RECT 3032.355 360.665 3032.635 360.945 ;
        RECT 3033.065 360.665 3033.345 360.945 ;
        RECT 3033.775 360.665 3034.055 360.945 ;
        RECT 3034.485 360.665 3034.765 360.945 ;
        RECT 3035.195 360.665 3035.475 360.945 ;
        RECT 3039.495 369.895 3039.775 370.175 ;
        RECT 3040.205 369.895 3040.485 370.175 ;
        RECT 3040.915 369.895 3041.195 370.175 ;
        RECT 3041.625 369.895 3041.905 370.175 ;
        RECT 3042.335 369.895 3042.615 370.175 ;
        RECT 3046.595 369.895 3046.875 370.175 ;
        RECT 3047.305 369.895 3047.585 370.175 ;
        RECT 3048.015 369.895 3048.295 370.175 ;
        RECT 3048.725 369.895 3049.005 370.175 ;
        RECT 3039.495 369.185 3039.775 369.465 ;
        RECT 3040.205 369.185 3040.485 369.465 ;
        RECT 3040.915 369.185 3041.195 369.465 ;
        RECT 3041.625 369.185 3041.905 369.465 ;
        RECT 3042.335 369.185 3042.615 369.465 ;
        RECT 3046.595 369.185 3046.875 369.465 ;
        RECT 3047.305 369.185 3047.585 369.465 ;
        RECT 3048.015 369.185 3048.295 369.465 ;
        RECT 3048.725 369.185 3049.005 369.465 ;
        RECT 3039.495 368.475 3039.775 368.755 ;
        RECT 3040.205 368.475 3040.485 368.755 ;
        RECT 3040.915 368.475 3041.195 368.755 ;
        RECT 3041.625 368.475 3041.905 368.755 ;
        RECT 3042.335 368.475 3042.615 368.755 ;
        RECT 3046.595 368.475 3046.875 368.755 ;
        RECT 3047.305 368.475 3047.585 368.755 ;
        RECT 3048.015 368.475 3048.295 368.755 ;
        RECT 3048.725 368.475 3049.005 368.755 ;
        RECT 3039.495 367.765 3039.775 368.045 ;
        RECT 3040.205 367.765 3040.485 368.045 ;
        RECT 3040.915 367.765 3041.195 368.045 ;
        RECT 3041.625 367.765 3041.905 368.045 ;
        RECT 3042.335 367.765 3042.615 368.045 ;
        RECT 3046.595 367.765 3046.875 368.045 ;
        RECT 3047.305 367.765 3047.585 368.045 ;
        RECT 3048.015 367.765 3048.295 368.045 ;
        RECT 3048.725 367.765 3049.005 368.045 ;
        RECT 3039.495 367.055 3039.775 367.335 ;
        RECT 3040.205 367.055 3040.485 367.335 ;
        RECT 3040.915 367.055 3041.195 367.335 ;
        RECT 3041.625 367.055 3041.905 367.335 ;
        RECT 3042.335 367.055 3042.615 367.335 ;
        RECT 3046.595 367.055 3046.875 367.335 ;
        RECT 3047.305 367.055 3047.585 367.335 ;
        RECT 3048.015 367.055 3048.295 367.335 ;
        RECT 3048.725 367.055 3049.005 367.335 ;
        RECT 3039.495 366.345 3039.775 366.625 ;
        RECT 3040.205 366.345 3040.485 366.625 ;
        RECT 3040.915 366.345 3041.195 366.625 ;
        RECT 3041.625 366.345 3041.905 366.625 ;
        RECT 3042.335 366.345 3042.615 366.625 ;
        RECT 3046.595 366.345 3046.875 366.625 ;
        RECT 3047.305 366.345 3047.585 366.625 ;
        RECT 3048.015 366.345 3048.295 366.625 ;
        RECT 3048.725 366.345 3049.005 366.625 ;
        RECT 3039.495 365.635 3039.775 365.915 ;
        RECT 3040.205 365.635 3040.485 365.915 ;
        RECT 3040.915 365.635 3041.195 365.915 ;
        RECT 3041.625 365.635 3041.905 365.915 ;
        RECT 3042.335 365.635 3042.615 365.915 ;
        RECT 3046.595 365.635 3046.875 365.915 ;
        RECT 3047.305 365.635 3047.585 365.915 ;
        RECT 3048.015 365.635 3048.295 365.915 ;
        RECT 3048.725 365.635 3049.005 365.915 ;
        RECT 3039.495 364.925 3039.775 365.205 ;
        RECT 3040.205 364.925 3040.485 365.205 ;
        RECT 3040.915 364.925 3041.195 365.205 ;
        RECT 3041.625 364.925 3041.905 365.205 ;
        RECT 3042.335 364.925 3042.615 365.205 ;
        RECT 3046.595 364.925 3046.875 365.205 ;
        RECT 3047.305 364.925 3047.585 365.205 ;
        RECT 3048.015 364.925 3048.295 365.205 ;
        RECT 3048.725 364.925 3049.005 365.205 ;
        RECT 3039.495 364.215 3039.775 364.495 ;
        RECT 3040.205 364.215 3040.485 364.495 ;
        RECT 3040.915 364.215 3041.195 364.495 ;
        RECT 3041.625 364.215 3041.905 364.495 ;
        RECT 3042.335 364.215 3042.615 364.495 ;
        RECT 3046.595 364.215 3046.875 364.495 ;
        RECT 3047.305 364.215 3047.585 364.495 ;
        RECT 3048.015 364.215 3048.295 364.495 ;
        RECT 3048.725 364.215 3049.005 364.495 ;
        RECT 3039.495 363.505 3039.775 363.785 ;
        RECT 3040.205 363.505 3040.485 363.785 ;
        RECT 3040.915 363.505 3041.195 363.785 ;
        RECT 3041.625 363.505 3041.905 363.785 ;
        RECT 3042.335 363.505 3042.615 363.785 ;
        RECT 3046.595 363.505 3046.875 363.785 ;
        RECT 3047.305 363.505 3047.585 363.785 ;
        RECT 3048.015 363.505 3048.295 363.785 ;
        RECT 3048.725 363.505 3049.005 363.785 ;
        RECT 3039.495 362.795 3039.775 363.075 ;
        RECT 3040.205 362.795 3040.485 363.075 ;
        RECT 3040.915 362.795 3041.195 363.075 ;
        RECT 3041.625 362.795 3041.905 363.075 ;
        RECT 3042.335 362.795 3042.615 363.075 ;
        RECT 3046.595 362.795 3046.875 363.075 ;
        RECT 3047.305 362.795 3047.585 363.075 ;
        RECT 3048.015 362.795 3048.295 363.075 ;
        RECT 3048.725 362.795 3049.005 363.075 ;
        RECT 3039.495 362.085 3039.775 362.365 ;
        RECT 3040.205 362.085 3040.485 362.365 ;
        RECT 3040.915 362.085 3041.195 362.365 ;
        RECT 3041.625 362.085 3041.905 362.365 ;
        RECT 3042.335 362.085 3042.615 362.365 ;
        RECT 3046.595 362.085 3046.875 362.365 ;
        RECT 3047.305 362.085 3047.585 362.365 ;
        RECT 3048.015 362.085 3048.295 362.365 ;
        RECT 3048.725 362.085 3049.005 362.365 ;
        RECT 3039.495 361.375 3039.775 361.655 ;
        RECT 3040.205 361.375 3040.485 361.655 ;
        RECT 3040.915 361.375 3041.195 361.655 ;
        RECT 3041.625 361.375 3041.905 361.655 ;
        RECT 3042.335 361.375 3042.615 361.655 ;
        RECT 3046.595 361.375 3046.875 361.655 ;
        RECT 3047.305 361.375 3047.585 361.655 ;
        RECT 3048.015 361.375 3048.295 361.655 ;
        RECT 3048.725 361.375 3049.005 361.655 ;
        RECT 3039.495 360.665 3039.775 360.945 ;
        RECT 3040.205 360.665 3040.485 360.945 ;
        RECT 3040.915 360.665 3041.195 360.945 ;
        RECT 3041.625 360.665 3041.905 360.945 ;
        RECT 3042.335 360.665 3042.615 360.945 ;
        RECT 3046.595 360.665 3046.875 360.945 ;
        RECT 3047.305 360.665 3047.585 360.945 ;
        RECT 3048.015 360.665 3048.295 360.945 ;
        RECT 3048.725 360.665 3049.005 360.945 ;
        RECT 3051.345 369.895 3051.625 370.175 ;
        RECT 3052.055 369.895 3052.335 370.175 ;
        RECT 3052.765 369.895 3053.045 370.175 ;
        RECT 3053.475 369.895 3053.755 370.175 ;
        RECT 3054.185 369.895 3054.465 370.175 ;
        RECT 3054.895 369.895 3055.175 370.175 ;
        RECT 3055.605 369.895 3055.885 370.175 ;
        RECT 3056.315 369.895 3056.595 370.175 ;
        RECT 3057.025 369.895 3057.305 370.175 ;
        RECT 3057.735 369.895 3058.015 370.175 ;
        RECT 3058.445 369.895 3058.725 370.175 ;
        RECT 3059.155 369.895 3059.435 370.175 ;
        RECT 3059.865 369.895 3060.145 370.175 ;
        RECT 3060.575 369.895 3060.855 370.175 ;
        RECT 3051.345 369.185 3051.625 369.465 ;
        RECT 3052.055 369.185 3052.335 369.465 ;
        RECT 3052.765 369.185 3053.045 369.465 ;
        RECT 3053.475 369.185 3053.755 369.465 ;
        RECT 3054.185 369.185 3054.465 369.465 ;
        RECT 3054.895 369.185 3055.175 369.465 ;
        RECT 3055.605 369.185 3055.885 369.465 ;
        RECT 3056.315 369.185 3056.595 369.465 ;
        RECT 3057.025 369.185 3057.305 369.465 ;
        RECT 3057.735 369.185 3058.015 369.465 ;
        RECT 3058.445 369.185 3058.725 369.465 ;
        RECT 3059.155 369.185 3059.435 369.465 ;
        RECT 3059.865 369.185 3060.145 369.465 ;
        RECT 3060.575 369.185 3060.855 369.465 ;
        RECT 3051.345 368.475 3051.625 368.755 ;
        RECT 3052.055 368.475 3052.335 368.755 ;
        RECT 3052.765 368.475 3053.045 368.755 ;
        RECT 3053.475 368.475 3053.755 368.755 ;
        RECT 3054.185 368.475 3054.465 368.755 ;
        RECT 3054.895 368.475 3055.175 368.755 ;
        RECT 3055.605 368.475 3055.885 368.755 ;
        RECT 3056.315 368.475 3056.595 368.755 ;
        RECT 3057.025 368.475 3057.305 368.755 ;
        RECT 3057.735 368.475 3058.015 368.755 ;
        RECT 3058.445 368.475 3058.725 368.755 ;
        RECT 3059.155 368.475 3059.435 368.755 ;
        RECT 3059.865 368.475 3060.145 368.755 ;
        RECT 3060.575 368.475 3060.855 368.755 ;
        RECT 3051.345 367.765 3051.625 368.045 ;
        RECT 3052.055 367.765 3052.335 368.045 ;
        RECT 3052.765 367.765 3053.045 368.045 ;
        RECT 3053.475 367.765 3053.755 368.045 ;
        RECT 3054.185 367.765 3054.465 368.045 ;
        RECT 3054.895 367.765 3055.175 368.045 ;
        RECT 3055.605 367.765 3055.885 368.045 ;
        RECT 3056.315 367.765 3056.595 368.045 ;
        RECT 3057.025 367.765 3057.305 368.045 ;
        RECT 3057.735 367.765 3058.015 368.045 ;
        RECT 3058.445 367.765 3058.725 368.045 ;
        RECT 3059.155 367.765 3059.435 368.045 ;
        RECT 3059.865 367.765 3060.145 368.045 ;
        RECT 3060.575 367.765 3060.855 368.045 ;
        RECT 3051.345 367.055 3051.625 367.335 ;
        RECT 3052.055 367.055 3052.335 367.335 ;
        RECT 3052.765 367.055 3053.045 367.335 ;
        RECT 3053.475 367.055 3053.755 367.335 ;
        RECT 3054.185 367.055 3054.465 367.335 ;
        RECT 3054.895 367.055 3055.175 367.335 ;
        RECT 3055.605 367.055 3055.885 367.335 ;
        RECT 3056.315 367.055 3056.595 367.335 ;
        RECT 3057.025 367.055 3057.305 367.335 ;
        RECT 3057.735 367.055 3058.015 367.335 ;
        RECT 3058.445 367.055 3058.725 367.335 ;
        RECT 3059.155 367.055 3059.435 367.335 ;
        RECT 3059.865 367.055 3060.145 367.335 ;
        RECT 3060.575 367.055 3060.855 367.335 ;
        RECT 3051.345 366.345 3051.625 366.625 ;
        RECT 3052.055 366.345 3052.335 366.625 ;
        RECT 3052.765 366.345 3053.045 366.625 ;
        RECT 3053.475 366.345 3053.755 366.625 ;
        RECT 3054.185 366.345 3054.465 366.625 ;
        RECT 3054.895 366.345 3055.175 366.625 ;
        RECT 3055.605 366.345 3055.885 366.625 ;
        RECT 3056.315 366.345 3056.595 366.625 ;
        RECT 3057.025 366.345 3057.305 366.625 ;
        RECT 3057.735 366.345 3058.015 366.625 ;
        RECT 3058.445 366.345 3058.725 366.625 ;
        RECT 3059.155 366.345 3059.435 366.625 ;
        RECT 3059.865 366.345 3060.145 366.625 ;
        RECT 3060.575 366.345 3060.855 366.625 ;
        RECT 3051.345 365.635 3051.625 365.915 ;
        RECT 3052.055 365.635 3052.335 365.915 ;
        RECT 3052.765 365.635 3053.045 365.915 ;
        RECT 3053.475 365.635 3053.755 365.915 ;
        RECT 3054.185 365.635 3054.465 365.915 ;
        RECT 3054.895 365.635 3055.175 365.915 ;
        RECT 3055.605 365.635 3055.885 365.915 ;
        RECT 3056.315 365.635 3056.595 365.915 ;
        RECT 3057.025 365.635 3057.305 365.915 ;
        RECT 3057.735 365.635 3058.015 365.915 ;
        RECT 3058.445 365.635 3058.725 365.915 ;
        RECT 3059.155 365.635 3059.435 365.915 ;
        RECT 3059.865 365.635 3060.145 365.915 ;
        RECT 3060.575 365.635 3060.855 365.915 ;
        RECT 3051.345 364.925 3051.625 365.205 ;
        RECT 3052.055 364.925 3052.335 365.205 ;
        RECT 3052.765 364.925 3053.045 365.205 ;
        RECT 3053.475 364.925 3053.755 365.205 ;
        RECT 3054.185 364.925 3054.465 365.205 ;
        RECT 3054.895 364.925 3055.175 365.205 ;
        RECT 3055.605 364.925 3055.885 365.205 ;
        RECT 3056.315 364.925 3056.595 365.205 ;
        RECT 3057.025 364.925 3057.305 365.205 ;
        RECT 3057.735 364.925 3058.015 365.205 ;
        RECT 3058.445 364.925 3058.725 365.205 ;
        RECT 3059.155 364.925 3059.435 365.205 ;
        RECT 3059.865 364.925 3060.145 365.205 ;
        RECT 3060.575 364.925 3060.855 365.205 ;
        RECT 3051.345 364.215 3051.625 364.495 ;
        RECT 3052.055 364.215 3052.335 364.495 ;
        RECT 3052.765 364.215 3053.045 364.495 ;
        RECT 3053.475 364.215 3053.755 364.495 ;
        RECT 3054.185 364.215 3054.465 364.495 ;
        RECT 3054.895 364.215 3055.175 364.495 ;
        RECT 3055.605 364.215 3055.885 364.495 ;
        RECT 3056.315 364.215 3056.595 364.495 ;
        RECT 3057.025 364.215 3057.305 364.495 ;
        RECT 3057.735 364.215 3058.015 364.495 ;
        RECT 3058.445 364.215 3058.725 364.495 ;
        RECT 3059.155 364.215 3059.435 364.495 ;
        RECT 3059.865 364.215 3060.145 364.495 ;
        RECT 3060.575 364.215 3060.855 364.495 ;
        RECT 3051.345 363.505 3051.625 363.785 ;
        RECT 3052.055 363.505 3052.335 363.785 ;
        RECT 3052.765 363.505 3053.045 363.785 ;
        RECT 3053.475 363.505 3053.755 363.785 ;
        RECT 3054.185 363.505 3054.465 363.785 ;
        RECT 3054.895 363.505 3055.175 363.785 ;
        RECT 3055.605 363.505 3055.885 363.785 ;
        RECT 3056.315 363.505 3056.595 363.785 ;
        RECT 3057.025 363.505 3057.305 363.785 ;
        RECT 3057.735 363.505 3058.015 363.785 ;
        RECT 3058.445 363.505 3058.725 363.785 ;
        RECT 3059.155 363.505 3059.435 363.785 ;
        RECT 3059.865 363.505 3060.145 363.785 ;
        RECT 3060.575 363.505 3060.855 363.785 ;
        RECT 3051.345 362.795 3051.625 363.075 ;
        RECT 3052.055 362.795 3052.335 363.075 ;
        RECT 3052.765 362.795 3053.045 363.075 ;
        RECT 3053.475 362.795 3053.755 363.075 ;
        RECT 3054.185 362.795 3054.465 363.075 ;
        RECT 3054.895 362.795 3055.175 363.075 ;
        RECT 3055.605 362.795 3055.885 363.075 ;
        RECT 3056.315 362.795 3056.595 363.075 ;
        RECT 3057.025 362.795 3057.305 363.075 ;
        RECT 3057.735 362.795 3058.015 363.075 ;
        RECT 3058.445 362.795 3058.725 363.075 ;
        RECT 3059.155 362.795 3059.435 363.075 ;
        RECT 3059.865 362.795 3060.145 363.075 ;
        RECT 3060.575 362.795 3060.855 363.075 ;
        RECT 3051.345 362.085 3051.625 362.365 ;
        RECT 3052.055 362.085 3052.335 362.365 ;
        RECT 3052.765 362.085 3053.045 362.365 ;
        RECT 3053.475 362.085 3053.755 362.365 ;
        RECT 3054.185 362.085 3054.465 362.365 ;
        RECT 3054.895 362.085 3055.175 362.365 ;
        RECT 3055.605 362.085 3055.885 362.365 ;
        RECT 3056.315 362.085 3056.595 362.365 ;
        RECT 3057.025 362.085 3057.305 362.365 ;
        RECT 3057.735 362.085 3058.015 362.365 ;
        RECT 3058.445 362.085 3058.725 362.365 ;
        RECT 3059.155 362.085 3059.435 362.365 ;
        RECT 3059.865 362.085 3060.145 362.365 ;
        RECT 3060.575 362.085 3060.855 362.365 ;
        RECT 3051.345 361.375 3051.625 361.655 ;
        RECT 3052.055 361.375 3052.335 361.655 ;
        RECT 3052.765 361.375 3053.045 361.655 ;
        RECT 3053.475 361.375 3053.755 361.655 ;
        RECT 3054.185 361.375 3054.465 361.655 ;
        RECT 3054.895 361.375 3055.175 361.655 ;
        RECT 3055.605 361.375 3055.885 361.655 ;
        RECT 3056.315 361.375 3056.595 361.655 ;
        RECT 3057.025 361.375 3057.305 361.655 ;
        RECT 3057.735 361.375 3058.015 361.655 ;
        RECT 3058.445 361.375 3058.725 361.655 ;
        RECT 3059.155 361.375 3059.435 361.655 ;
        RECT 3059.865 361.375 3060.145 361.655 ;
        RECT 3060.575 361.375 3060.855 361.655 ;
        RECT 3051.345 360.665 3051.625 360.945 ;
        RECT 3052.055 360.665 3052.335 360.945 ;
        RECT 3052.765 360.665 3053.045 360.945 ;
        RECT 3053.475 360.665 3053.755 360.945 ;
        RECT 3054.185 360.665 3054.465 360.945 ;
        RECT 3054.895 360.665 3055.175 360.945 ;
        RECT 3055.605 360.665 3055.885 360.945 ;
        RECT 3056.315 360.665 3056.595 360.945 ;
        RECT 3057.025 360.665 3057.305 360.945 ;
        RECT 3057.735 360.665 3058.015 360.945 ;
        RECT 3058.445 360.665 3058.725 360.945 ;
        RECT 3059.155 360.665 3059.435 360.945 ;
        RECT 3059.865 360.665 3060.145 360.945 ;
        RECT 3060.575 360.665 3060.855 360.945 ;
        RECT 3064.495 369.895 3064.775 370.175 ;
        RECT 3065.205 369.895 3065.485 370.175 ;
        RECT 3065.915 369.895 3066.195 370.175 ;
        RECT 3066.625 369.895 3066.905 370.175 ;
        RECT 3067.335 369.895 3067.615 370.175 ;
        RECT 3068.045 369.895 3068.325 370.175 ;
        RECT 3068.755 369.895 3069.035 370.175 ;
        RECT 3069.465 369.895 3069.745 370.175 ;
        RECT 3070.175 369.895 3070.455 370.175 ;
        RECT 3070.885 369.895 3071.165 370.175 ;
        RECT 3071.595 369.895 3071.875 370.175 ;
        RECT 3072.305 369.895 3072.585 370.175 ;
        RECT 3073.015 369.895 3073.295 370.175 ;
        RECT 3064.495 369.185 3064.775 369.465 ;
        RECT 3065.205 369.185 3065.485 369.465 ;
        RECT 3065.915 369.185 3066.195 369.465 ;
        RECT 3066.625 369.185 3066.905 369.465 ;
        RECT 3067.335 369.185 3067.615 369.465 ;
        RECT 3068.045 369.185 3068.325 369.465 ;
        RECT 3068.755 369.185 3069.035 369.465 ;
        RECT 3069.465 369.185 3069.745 369.465 ;
        RECT 3070.175 369.185 3070.455 369.465 ;
        RECT 3070.885 369.185 3071.165 369.465 ;
        RECT 3071.595 369.185 3071.875 369.465 ;
        RECT 3072.305 369.185 3072.585 369.465 ;
        RECT 3073.015 369.185 3073.295 369.465 ;
        RECT 3064.495 368.475 3064.775 368.755 ;
        RECT 3065.205 368.475 3065.485 368.755 ;
        RECT 3065.915 368.475 3066.195 368.755 ;
        RECT 3066.625 368.475 3066.905 368.755 ;
        RECT 3067.335 368.475 3067.615 368.755 ;
        RECT 3068.045 368.475 3068.325 368.755 ;
        RECT 3068.755 368.475 3069.035 368.755 ;
        RECT 3069.465 368.475 3069.745 368.755 ;
        RECT 3070.175 368.475 3070.455 368.755 ;
        RECT 3070.885 368.475 3071.165 368.755 ;
        RECT 3071.595 368.475 3071.875 368.755 ;
        RECT 3072.305 368.475 3072.585 368.755 ;
        RECT 3073.015 368.475 3073.295 368.755 ;
        RECT 3064.495 367.765 3064.775 368.045 ;
        RECT 3065.205 367.765 3065.485 368.045 ;
        RECT 3065.915 367.765 3066.195 368.045 ;
        RECT 3066.625 367.765 3066.905 368.045 ;
        RECT 3067.335 367.765 3067.615 368.045 ;
        RECT 3068.045 367.765 3068.325 368.045 ;
        RECT 3068.755 367.765 3069.035 368.045 ;
        RECT 3069.465 367.765 3069.745 368.045 ;
        RECT 3070.175 367.765 3070.455 368.045 ;
        RECT 3070.885 367.765 3071.165 368.045 ;
        RECT 3071.595 367.765 3071.875 368.045 ;
        RECT 3072.305 367.765 3072.585 368.045 ;
        RECT 3073.015 367.765 3073.295 368.045 ;
        RECT 3064.495 367.055 3064.775 367.335 ;
        RECT 3065.205 367.055 3065.485 367.335 ;
        RECT 3065.915 367.055 3066.195 367.335 ;
        RECT 3066.625 367.055 3066.905 367.335 ;
        RECT 3067.335 367.055 3067.615 367.335 ;
        RECT 3068.045 367.055 3068.325 367.335 ;
        RECT 3068.755 367.055 3069.035 367.335 ;
        RECT 3069.465 367.055 3069.745 367.335 ;
        RECT 3070.175 367.055 3070.455 367.335 ;
        RECT 3070.885 367.055 3071.165 367.335 ;
        RECT 3071.595 367.055 3071.875 367.335 ;
        RECT 3072.305 367.055 3072.585 367.335 ;
        RECT 3073.015 367.055 3073.295 367.335 ;
        RECT 3064.495 366.345 3064.775 366.625 ;
        RECT 3065.205 366.345 3065.485 366.625 ;
        RECT 3065.915 366.345 3066.195 366.625 ;
        RECT 3066.625 366.345 3066.905 366.625 ;
        RECT 3067.335 366.345 3067.615 366.625 ;
        RECT 3068.045 366.345 3068.325 366.625 ;
        RECT 3068.755 366.345 3069.035 366.625 ;
        RECT 3069.465 366.345 3069.745 366.625 ;
        RECT 3070.175 366.345 3070.455 366.625 ;
        RECT 3070.885 366.345 3071.165 366.625 ;
        RECT 3071.595 366.345 3071.875 366.625 ;
        RECT 3072.305 366.345 3072.585 366.625 ;
        RECT 3073.015 366.345 3073.295 366.625 ;
        RECT 3064.495 365.635 3064.775 365.915 ;
        RECT 3065.205 365.635 3065.485 365.915 ;
        RECT 3065.915 365.635 3066.195 365.915 ;
        RECT 3066.625 365.635 3066.905 365.915 ;
        RECT 3067.335 365.635 3067.615 365.915 ;
        RECT 3068.045 365.635 3068.325 365.915 ;
        RECT 3068.755 365.635 3069.035 365.915 ;
        RECT 3069.465 365.635 3069.745 365.915 ;
        RECT 3070.175 365.635 3070.455 365.915 ;
        RECT 3070.885 365.635 3071.165 365.915 ;
        RECT 3071.595 365.635 3071.875 365.915 ;
        RECT 3072.305 365.635 3072.585 365.915 ;
        RECT 3073.015 365.635 3073.295 365.915 ;
        RECT 3064.495 364.925 3064.775 365.205 ;
        RECT 3065.205 364.925 3065.485 365.205 ;
        RECT 3065.915 364.925 3066.195 365.205 ;
        RECT 3066.625 364.925 3066.905 365.205 ;
        RECT 3067.335 364.925 3067.615 365.205 ;
        RECT 3068.045 364.925 3068.325 365.205 ;
        RECT 3068.755 364.925 3069.035 365.205 ;
        RECT 3069.465 364.925 3069.745 365.205 ;
        RECT 3070.175 364.925 3070.455 365.205 ;
        RECT 3070.885 364.925 3071.165 365.205 ;
        RECT 3071.595 364.925 3071.875 365.205 ;
        RECT 3072.305 364.925 3072.585 365.205 ;
        RECT 3073.015 364.925 3073.295 365.205 ;
        RECT 3064.495 364.215 3064.775 364.495 ;
        RECT 3065.205 364.215 3065.485 364.495 ;
        RECT 3065.915 364.215 3066.195 364.495 ;
        RECT 3066.625 364.215 3066.905 364.495 ;
        RECT 3067.335 364.215 3067.615 364.495 ;
        RECT 3068.045 364.215 3068.325 364.495 ;
        RECT 3068.755 364.215 3069.035 364.495 ;
        RECT 3069.465 364.215 3069.745 364.495 ;
        RECT 3070.175 364.215 3070.455 364.495 ;
        RECT 3070.885 364.215 3071.165 364.495 ;
        RECT 3071.595 364.215 3071.875 364.495 ;
        RECT 3072.305 364.215 3072.585 364.495 ;
        RECT 3073.015 364.215 3073.295 364.495 ;
        RECT 3064.495 363.505 3064.775 363.785 ;
        RECT 3065.205 363.505 3065.485 363.785 ;
        RECT 3065.915 363.505 3066.195 363.785 ;
        RECT 3066.625 363.505 3066.905 363.785 ;
        RECT 3067.335 363.505 3067.615 363.785 ;
        RECT 3068.045 363.505 3068.325 363.785 ;
        RECT 3068.755 363.505 3069.035 363.785 ;
        RECT 3069.465 363.505 3069.745 363.785 ;
        RECT 3070.175 363.505 3070.455 363.785 ;
        RECT 3070.885 363.505 3071.165 363.785 ;
        RECT 3071.595 363.505 3071.875 363.785 ;
        RECT 3072.305 363.505 3072.585 363.785 ;
        RECT 3073.015 363.505 3073.295 363.785 ;
        RECT 3064.495 362.795 3064.775 363.075 ;
        RECT 3065.205 362.795 3065.485 363.075 ;
        RECT 3065.915 362.795 3066.195 363.075 ;
        RECT 3066.625 362.795 3066.905 363.075 ;
        RECT 3067.335 362.795 3067.615 363.075 ;
        RECT 3068.045 362.795 3068.325 363.075 ;
        RECT 3068.755 362.795 3069.035 363.075 ;
        RECT 3069.465 362.795 3069.745 363.075 ;
        RECT 3070.175 362.795 3070.455 363.075 ;
        RECT 3070.885 362.795 3071.165 363.075 ;
        RECT 3071.595 362.795 3071.875 363.075 ;
        RECT 3072.305 362.795 3072.585 363.075 ;
        RECT 3073.015 362.795 3073.295 363.075 ;
        RECT 3064.495 362.085 3064.775 362.365 ;
        RECT 3065.205 362.085 3065.485 362.365 ;
        RECT 3065.915 362.085 3066.195 362.365 ;
        RECT 3066.625 362.085 3066.905 362.365 ;
        RECT 3067.335 362.085 3067.615 362.365 ;
        RECT 3068.045 362.085 3068.325 362.365 ;
        RECT 3068.755 362.085 3069.035 362.365 ;
        RECT 3069.465 362.085 3069.745 362.365 ;
        RECT 3070.175 362.085 3070.455 362.365 ;
        RECT 3070.885 362.085 3071.165 362.365 ;
        RECT 3071.595 362.085 3071.875 362.365 ;
        RECT 3072.305 362.085 3072.585 362.365 ;
        RECT 3073.015 362.085 3073.295 362.365 ;
        RECT 3064.495 361.375 3064.775 361.655 ;
        RECT 3065.205 361.375 3065.485 361.655 ;
        RECT 3065.915 361.375 3066.195 361.655 ;
        RECT 3066.625 361.375 3066.905 361.655 ;
        RECT 3067.335 361.375 3067.615 361.655 ;
        RECT 3068.045 361.375 3068.325 361.655 ;
        RECT 3068.755 361.375 3069.035 361.655 ;
        RECT 3069.465 361.375 3069.745 361.655 ;
        RECT 3070.175 361.375 3070.455 361.655 ;
        RECT 3070.885 361.375 3071.165 361.655 ;
        RECT 3071.595 361.375 3071.875 361.655 ;
        RECT 3072.305 361.375 3072.585 361.655 ;
        RECT 3073.015 361.375 3073.295 361.655 ;
        RECT 3064.495 360.665 3064.775 360.945 ;
        RECT 3065.205 360.665 3065.485 360.945 ;
        RECT 3065.915 360.665 3066.195 360.945 ;
        RECT 3066.625 360.665 3066.905 360.945 ;
        RECT 3067.335 360.665 3067.615 360.945 ;
        RECT 3068.045 360.665 3068.325 360.945 ;
        RECT 3068.755 360.665 3069.035 360.945 ;
        RECT 3069.465 360.665 3069.745 360.945 ;
        RECT 3070.175 360.665 3070.455 360.945 ;
        RECT 3070.885 360.665 3071.165 360.945 ;
        RECT 3071.595 360.665 3071.875 360.945 ;
        RECT 3072.305 360.665 3072.585 360.945 ;
        RECT 3073.015 360.665 3073.295 360.945 ;
      LAYER Metal5 ;
        RECT 1896.705 4708.095 1896.985 4708.375 ;
        RECT 1897.415 4708.095 1897.695 4708.375 ;
        RECT 1898.125 4708.095 1898.405 4708.375 ;
        RECT 1898.835 4708.095 1899.115 4708.375 ;
        RECT 1899.545 4708.095 1899.825 4708.375 ;
        RECT 1909.145 4708.095 1909.425 4708.375 ;
        RECT 1909.855 4708.095 1910.135 4708.375 ;
        RECT 1910.565 4708.095 1910.845 4708.375 ;
        RECT 1911.275 4708.095 1911.555 4708.375 ;
        RECT 1911.985 4708.095 1912.265 4708.375 ;
        RECT 1912.695 4708.095 1912.975 4708.375 ;
        RECT 1913.405 4708.095 1913.685 4708.375 ;
        RECT 1914.115 4708.095 1914.395 4708.375 ;
        RECT 1914.825 4708.095 1915.105 4708.375 ;
        RECT 1915.535 4708.095 1915.815 4708.375 ;
        RECT 1916.245 4708.095 1916.525 4708.375 ;
        RECT 1916.955 4708.095 1917.235 4708.375 ;
        RECT 1917.665 4708.095 1917.945 4708.375 ;
        RECT 1918.375 4708.095 1918.655 4708.375 ;
        RECT 1920.995 4708.095 1921.275 4708.375 ;
        RECT 1921.705 4708.095 1921.985 4708.375 ;
        RECT 1922.415 4708.095 1922.695 4708.375 ;
        RECT 1926.675 4708.095 1926.955 4708.375 ;
        RECT 1927.385 4708.095 1927.665 4708.375 ;
        RECT 1928.095 4708.095 1928.375 4708.375 ;
        RECT 1928.805 4708.095 1929.085 4708.375 ;
        RECT 1929.515 4708.095 1929.795 4708.375 ;
        RECT 1930.225 4708.095 1930.505 4708.375 ;
        RECT 1934.525 4708.095 1934.805 4708.375 ;
        RECT 1935.235 4708.095 1935.515 4708.375 ;
        RECT 1935.945 4708.095 1936.225 4708.375 ;
        RECT 1936.655 4708.095 1936.935 4708.375 ;
        RECT 1937.365 4708.095 1937.645 4708.375 ;
        RECT 1938.075 4708.095 1938.355 4708.375 ;
        RECT 1938.785 4708.095 1939.065 4708.375 ;
        RECT 1939.495 4708.095 1939.775 4708.375 ;
        RECT 1940.205 4708.095 1940.485 4708.375 ;
        RECT 1940.915 4708.095 1941.195 4708.375 ;
        RECT 1941.625 4708.095 1941.905 4708.375 ;
        RECT 1942.335 4708.095 1942.615 4708.375 ;
        RECT 1943.045 4708.095 1943.325 4708.375 ;
        RECT 1943.755 4708.095 1944.035 4708.375 ;
        RECT 1946.375 4708.095 1946.655 4708.375 ;
        RECT 1947.085 4708.095 1947.365 4708.375 ;
        RECT 1947.795 4708.095 1948.075 4708.375 ;
        RECT 1948.505 4708.095 1948.785 4708.375 ;
        RECT 1949.215 4708.095 1949.495 4708.375 ;
        RECT 1949.925 4708.095 1950.205 4708.375 ;
        RECT 1950.635 4708.095 1950.915 4708.375 ;
        RECT 1951.345 4708.095 1951.625 4708.375 ;
        RECT 1952.055 4708.095 1952.335 4708.375 ;
        RECT 1952.765 4708.095 1953.045 4708.375 ;
        RECT 1953.475 4708.095 1953.755 4708.375 ;
        RECT 1954.185 4708.095 1954.465 4708.375 ;
        RECT 1954.895 4708.095 1955.175 4708.375 ;
        RECT 1955.605 4708.095 1955.885 4708.375 ;
        RECT 1959.485 4708.095 1959.765 4708.375 ;
        RECT 1960.195 4708.095 1960.475 4708.375 ;
        RECT 1960.905 4708.095 1961.185 4708.375 ;
        RECT 1961.615 4708.095 1961.895 4708.375 ;
        RECT 1962.325 4708.095 1962.605 4708.375 ;
        RECT 1963.035 4708.095 1963.315 4708.375 ;
        RECT 1963.745 4708.095 1964.025 4708.375 ;
        RECT 1964.455 4708.095 1964.735 4708.375 ;
        RECT 1965.165 4708.095 1965.445 4708.375 ;
        RECT 1965.875 4708.095 1966.155 4708.375 ;
        RECT 1966.585 4708.095 1966.865 4708.375 ;
        RECT 1967.295 4708.095 1967.575 4708.375 ;
        RECT 1968.005 4708.095 1968.285 4708.375 ;
        RECT 2996.705 4708.095 2996.985 4708.375 ;
        RECT 2997.415 4708.095 2997.695 4708.375 ;
        RECT 2998.125 4708.095 2998.405 4708.375 ;
        RECT 2998.835 4708.095 2999.115 4708.375 ;
        RECT 2999.545 4708.095 2999.825 4708.375 ;
        RECT 3000.255 4708.095 3000.535 4708.375 ;
        RECT 3000.965 4708.095 3001.245 4708.375 ;
        RECT 3001.675 4708.095 3001.955 4708.375 ;
        RECT 3002.385 4708.095 3002.665 4708.375 ;
        RECT 3003.095 4708.095 3003.375 4708.375 ;
        RECT 3003.805 4708.095 3004.085 4708.375 ;
        RECT 3004.515 4708.095 3004.795 4708.375 ;
        RECT 3005.225 4708.095 3005.505 4708.375 ;
        RECT 3009.145 4708.095 3009.425 4708.375 ;
        RECT 3009.855 4708.095 3010.135 4708.375 ;
        RECT 3010.565 4708.095 3010.845 4708.375 ;
        RECT 3011.275 4708.095 3011.555 4708.375 ;
        RECT 3011.985 4708.095 3012.265 4708.375 ;
        RECT 3012.695 4708.095 3012.975 4708.375 ;
        RECT 3013.405 4708.095 3013.685 4708.375 ;
        RECT 3014.115 4708.095 3014.395 4708.375 ;
        RECT 3014.825 4708.095 3015.105 4708.375 ;
        RECT 3015.535 4708.095 3015.815 4708.375 ;
        RECT 3016.245 4708.095 3016.525 4708.375 ;
        RECT 3016.955 4708.095 3017.235 4708.375 ;
        RECT 3017.665 4708.095 3017.945 4708.375 ;
        RECT 3018.375 4708.095 3018.655 4708.375 ;
        RECT 3025.255 4708.095 3025.535 4708.375 ;
        RECT 3025.965 4708.095 3026.245 4708.375 ;
        RECT 3026.675 4708.095 3026.955 4708.375 ;
        RECT 3027.385 4708.095 3027.665 4708.375 ;
        RECT 3028.095 4708.095 3028.375 4708.375 ;
        RECT 3028.805 4708.095 3029.085 4708.375 ;
        RECT 3029.515 4708.095 3029.795 4708.375 ;
        RECT 3030.225 4708.095 3030.505 4708.375 ;
        RECT 3034.525 4708.095 3034.805 4708.375 ;
        RECT 3035.235 4708.095 3035.515 4708.375 ;
        RECT 3035.945 4708.095 3036.225 4708.375 ;
        RECT 3036.655 4708.095 3036.935 4708.375 ;
        RECT 3037.365 4708.095 3037.645 4708.375 ;
        RECT 3038.075 4708.095 3038.355 4708.375 ;
        RECT 3038.785 4708.095 3039.065 4708.375 ;
        RECT 3039.495 4708.095 3039.775 4708.375 ;
        RECT 3040.205 4708.095 3040.485 4708.375 ;
        RECT 3040.915 4708.095 3041.195 4708.375 ;
        RECT 3041.625 4708.095 3041.905 4708.375 ;
        RECT 3042.335 4708.095 3042.615 4708.375 ;
        RECT 3046.375 4708.095 3046.655 4708.375 ;
        RECT 3047.085 4708.095 3047.365 4708.375 ;
        RECT 3047.795 4708.095 3048.075 4708.375 ;
        RECT 3048.505 4708.095 3048.785 4708.375 ;
        RECT 3049.215 4708.095 3049.495 4708.375 ;
        RECT 3049.925 4708.095 3050.205 4708.375 ;
        RECT 3050.635 4708.095 3050.915 4708.375 ;
        RECT 3051.345 4708.095 3051.625 4708.375 ;
        RECT 3052.055 4708.095 3052.335 4708.375 ;
        RECT 3052.765 4708.095 3053.045 4708.375 ;
        RECT 3053.475 4708.095 3053.755 4708.375 ;
        RECT 3054.185 4708.095 3054.465 4708.375 ;
        RECT 3054.895 4708.095 3055.175 4708.375 ;
        RECT 3055.605 4708.095 3055.885 4708.375 ;
        RECT 3059.485 4708.095 3059.765 4708.375 ;
        RECT 3060.195 4708.095 3060.475 4708.375 ;
        RECT 3060.905 4708.095 3061.185 4708.375 ;
        RECT 3061.615 4708.095 3061.895 4708.375 ;
        RECT 3062.325 4708.095 3062.605 4708.375 ;
        RECT 3063.035 4708.095 3063.315 4708.375 ;
        RECT 3063.745 4708.095 3064.025 4708.375 ;
        RECT 3064.455 4708.095 3064.735 4708.375 ;
        RECT 3065.165 4708.095 3065.445 4708.375 ;
        RECT 3065.875 4708.095 3066.155 4708.375 ;
        RECT 3066.585 4708.095 3066.865 4708.375 ;
        RECT 3067.295 4708.095 3067.575 4708.375 ;
        RECT 3068.005 4708.095 3068.285 4708.375 ;
        RECT 1896.705 4707.385 1896.985 4707.665 ;
        RECT 1897.415 4707.385 1897.695 4707.665 ;
        RECT 1898.125 4707.385 1898.405 4707.665 ;
        RECT 1898.835 4707.385 1899.115 4707.665 ;
        RECT 1899.545 4707.385 1899.825 4707.665 ;
        RECT 1909.145 4707.385 1909.425 4707.665 ;
        RECT 1909.855 4707.385 1910.135 4707.665 ;
        RECT 1910.565 4707.385 1910.845 4707.665 ;
        RECT 1911.275 4707.385 1911.555 4707.665 ;
        RECT 1911.985 4707.385 1912.265 4707.665 ;
        RECT 1912.695 4707.385 1912.975 4707.665 ;
        RECT 1913.405 4707.385 1913.685 4707.665 ;
        RECT 1914.115 4707.385 1914.395 4707.665 ;
        RECT 1914.825 4707.385 1915.105 4707.665 ;
        RECT 1915.535 4707.385 1915.815 4707.665 ;
        RECT 1916.245 4707.385 1916.525 4707.665 ;
        RECT 1916.955 4707.385 1917.235 4707.665 ;
        RECT 1917.665 4707.385 1917.945 4707.665 ;
        RECT 1918.375 4707.385 1918.655 4707.665 ;
        RECT 1920.995 4707.385 1921.275 4707.665 ;
        RECT 1921.705 4707.385 1921.985 4707.665 ;
        RECT 1922.415 4707.385 1922.695 4707.665 ;
        RECT 1926.675 4707.385 1926.955 4707.665 ;
        RECT 1927.385 4707.385 1927.665 4707.665 ;
        RECT 1928.095 4707.385 1928.375 4707.665 ;
        RECT 1928.805 4707.385 1929.085 4707.665 ;
        RECT 1929.515 4707.385 1929.795 4707.665 ;
        RECT 1930.225 4707.385 1930.505 4707.665 ;
        RECT 1934.525 4707.385 1934.805 4707.665 ;
        RECT 1935.235 4707.385 1935.515 4707.665 ;
        RECT 1935.945 4707.385 1936.225 4707.665 ;
        RECT 1936.655 4707.385 1936.935 4707.665 ;
        RECT 1937.365 4707.385 1937.645 4707.665 ;
        RECT 1938.075 4707.385 1938.355 4707.665 ;
        RECT 1938.785 4707.385 1939.065 4707.665 ;
        RECT 1939.495 4707.385 1939.775 4707.665 ;
        RECT 1940.205 4707.385 1940.485 4707.665 ;
        RECT 1940.915 4707.385 1941.195 4707.665 ;
        RECT 1941.625 4707.385 1941.905 4707.665 ;
        RECT 1942.335 4707.385 1942.615 4707.665 ;
        RECT 1943.045 4707.385 1943.325 4707.665 ;
        RECT 1943.755 4707.385 1944.035 4707.665 ;
        RECT 1946.375 4707.385 1946.655 4707.665 ;
        RECT 1947.085 4707.385 1947.365 4707.665 ;
        RECT 1947.795 4707.385 1948.075 4707.665 ;
        RECT 1948.505 4707.385 1948.785 4707.665 ;
        RECT 1949.215 4707.385 1949.495 4707.665 ;
        RECT 1949.925 4707.385 1950.205 4707.665 ;
        RECT 1950.635 4707.385 1950.915 4707.665 ;
        RECT 1951.345 4707.385 1951.625 4707.665 ;
        RECT 1952.055 4707.385 1952.335 4707.665 ;
        RECT 1952.765 4707.385 1953.045 4707.665 ;
        RECT 1953.475 4707.385 1953.755 4707.665 ;
        RECT 1954.185 4707.385 1954.465 4707.665 ;
        RECT 1954.895 4707.385 1955.175 4707.665 ;
        RECT 1955.605 4707.385 1955.885 4707.665 ;
        RECT 1959.485 4707.385 1959.765 4707.665 ;
        RECT 1960.195 4707.385 1960.475 4707.665 ;
        RECT 1960.905 4707.385 1961.185 4707.665 ;
        RECT 1961.615 4707.385 1961.895 4707.665 ;
        RECT 1962.325 4707.385 1962.605 4707.665 ;
        RECT 1963.035 4707.385 1963.315 4707.665 ;
        RECT 1963.745 4707.385 1964.025 4707.665 ;
        RECT 1964.455 4707.385 1964.735 4707.665 ;
        RECT 1965.165 4707.385 1965.445 4707.665 ;
        RECT 1965.875 4707.385 1966.155 4707.665 ;
        RECT 1966.585 4707.385 1966.865 4707.665 ;
        RECT 1967.295 4707.385 1967.575 4707.665 ;
        RECT 1968.005 4707.385 1968.285 4707.665 ;
        RECT 2996.705 4707.385 2996.985 4707.665 ;
        RECT 2997.415 4707.385 2997.695 4707.665 ;
        RECT 2998.125 4707.385 2998.405 4707.665 ;
        RECT 2998.835 4707.385 2999.115 4707.665 ;
        RECT 2999.545 4707.385 2999.825 4707.665 ;
        RECT 3000.255 4707.385 3000.535 4707.665 ;
        RECT 3000.965 4707.385 3001.245 4707.665 ;
        RECT 3001.675 4707.385 3001.955 4707.665 ;
        RECT 3002.385 4707.385 3002.665 4707.665 ;
        RECT 3003.095 4707.385 3003.375 4707.665 ;
        RECT 3003.805 4707.385 3004.085 4707.665 ;
        RECT 3004.515 4707.385 3004.795 4707.665 ;
        RECT 3005.225 4707.385 3005.505 4707.665 ;
        RECT 3009.145 4707.385 3009.425 4707.665 ;
        RECT 3009.855 4707.385 3010.135 4707.665 ;
        RECT 3010.565 4707.385 3010.845 4707.665 ;
        RECT 3011.275 4707.385 3011.555 4707.665 ;
        RECT 3011.985 4707.385 3012.265 4707.665 ;
        RECT 3012.695 4707.385 3012.975 4707.665 ;
        RECT 3013.405 4707.385 3013.685 4707.665 ;
        RECT 3014.115 4707.385 3014.395 4707.665 ;
        RECT 3014.825 4707.385 3015.105 4707.665 ;
        RECT 3015.535 4707.385 3015.815 4707.665 ;
        RECT 3016.245 4707.385 3016.525 4707.665 ;
        RECT 3016.955 4707.385 3017.235 4707.665 ;
        RECT 3017.665 4707.385 3017.945 4707.665 ;
        RECT 3018.375 4707.385 3018.655 4707.665 ;
        RECT 3025.255 4707.385 3025.535 4707.665 ;
        RECT 3025.965 4707.385 3026.245 4707.665 ;
        RECT 3026.675 4707.385 3026.955 4707.665 ;
        RECT 3027.385 4707.385 3027.665 4707.665 ;
        RECT 3028.095 4707.385 3028.375 4707.665 ;
        RECT 3028.805 4707.385 3029.085 4707.665 ;
        RECT 3029.515 4707.385 3029.795 4707.665 ;
        RECT 3030.225 4707.385 3030.505 4707.665 ;
        RECT 3034.525 4707.385 3034.805 4707.665 ;
        RECT 3035.235 4707.385 3035.515 4707.665 ;
        RECT 3035.945 4707.385 3036.225 4707.665 ;
        RECT 3036.655 4707.385 3036.935 4707.665 ;
        RECT 3037.365 4707.385 3037.645 4707.665 ;
        RECT 3038.075 4707.385 3038.355 4707.665 ;
        RECT 3038.785 4707.385 3039.065 4707.665 ;
        RECT 3039.495 4707.385 3039.775 4707.665 ;
        RECT 3040.205 4707.385 3040.485 4707.665 ;
        RECT 3040.915 4707.385 3041.195 4707.665 ;
        RECT 3041.625 4707.385 3041.905 4707.665 ;
        RECT 3042.335 4707.385 3042.615 4707.665 ;
        RECT 3046.375 4707.385 3046.655 4707.665 ;
        RECT 3047.085 4707.385 3047.365 4707.665 ;
        RECT 3047.795 4707.385 3048.075 4707.665 ;
        RECT 3048.505 4707.385 3048.785 4707.665 ;
        RECT 3049.215 4707.385 3049.495 4707.665 ;
        RECT 3049.925 4707.385 3050.205 4707.665 ;
        RECT 3050.635 4707.385 3050.915 4707.665 ;
        RECT 3051.345 4707.385 3051.625 4707.665 ;
        RECT 3052.055 4707.385 3052.335 4707.665 ;
        RECT 3052.765 4707.385 3053.045 4707.665 ;
        RECT 3053.475 4707.385 3053.755 4707.665 ;
        RECT 3054.185 4707.385 3054.465 4707.665 ;
        RECT 3054.895 4707.385 3055.175 4707.665 ;
        RECT 3055.605 4707.385 3055.885 4707.665 ;
        RECT 3059.485 4707.385 3059.765 4707.665 ;
        RECT 3060.195 4707.385 3060.475 4707.665 ;
        RECT 3060.905 4707.385 3061.185 4707.665 ;
        RECT 3061.615 4707.385 3061.895 4707.665 ;
        RECT 3062.325 4707.385 3062.605 4707.665 ;
        RECT 3063.035 4707.385 3063.315 4707.665 ;
        RECT 3063.745 4707.385 3064.025 4707.665 ;
        RECT 3064.455 4707.385 3064.735 4707.665 ;
        RECT 3065.165 4707.385 3065.445 4707.665 ;
        RECT 3065.875 4707.385 3066.155 4707.665 ;
        RECT 3066.585 4707.385 3066.865 4707.665 ;
        RECT 3067.295 4707.385 3067.575 4707.665 ;
        RECT 3068.005 4707.385 3068.285 4707.665 ;
        RECT 1896.705 4706.675 1896.985 4706.955 ;
        RECT 1897.415 4706.675 1897.695 4706.955 ;
        RECT 1898.125 4706.675 1898.405 4706.955 ;
        RECT 1898.835 4706.675 1899.115 4706.955 ;
        RECT 1899.545 4706.675 1899.825 4706.955 ;
        RECT 1909.145 4706.675 1909.425 4706.955 ;
        RECT 1909.855 4706.675 1910.135 4706.955 ;
        RECT 1910.565 4706.675 1910.845 4706.955 ;
        RECT 1911.275 4706.675 1911.555 4706.955 ;
        RECT 1911.985 4706.675 1912.265 4706.955 ;
        RECT 1912.695 4706.675 1912.975 4706.955 ;
        RECT 1913.405 4706.675 1913.685 4706.955 ;
        RECT 1914.115 4706.675 1914.395 4706.955 ;
        RECT 1914.825 4706.675 1915.105 4706.955 ;
        RECT 1915.535 4706.675 1915.815 4706.955 ;
        RECT 1916.245 4706.675 1916.525 4706.955 ;
        RECT 1916.955 4706.675 1917.235 4706.955 ;
        RECT 1917.665 4706.675 1917.945 4706.955 ;
        RECT 1918.375 4706.675 1918.655 4706.955 ;
        RECT 1920.995 4706.675 1921.275 4706.955 ;
        RECT 1921.705 4706.675 1921.985 4706.955 ;
        RECT 1922.415 4706.675 1922.695 4706.955 ;
        RECT 1926.675 4706.675 1926.955 4706.955 ;
        RECT 1927.385 4706.675 1927.665 4706.955 ;
        RECT 1928.095 4706.675 1928.375 4706.955 ;
        RECT 1928.805 4706.675 1929.085 4706.955 ;
        RECT 1929.515 4706.675 1929.795 4706.955 ;
        RECT 1930.225 4706.675 1930.505 4706.955 ;
        RECT 1934.525 4706.675 1934.805 4706.955 ;
        RECT 1935.235 4706.675 1935.515 4706.955 ;
        RECT 1935.945 4706.675 1936.225 4706.955 ;
        RECT 1936.655 4706.675 1936.935 4706.955 ;
        RECT 1937.365 4706.675 1937.645 4706.955 ;
        RECT 1938.075 4706.675 1938.355 4706.955 ;
        RECT 1938.785 4706.675 1939.065 4706.955 ;
        RECT 1939.495 4706.675 1939.775 4706.955 ;
        RECT 1940.205 4706.675 1940.485 4706.955 ;
        RECT 1940.915 4706.675 1941.195 4706.955 ;
        RECT 1941.625 4706.675 1941.905 4706.955 ;
        RECT 1942.335 4706.675 1942.615 4706.955 ;
        RECT 1943.045 4706.675 1943.325 4706.955 ;
        RECT 1943.755 4706.675 1944.035 4706.955 ;
        RECT 1946.375 4706.675 1946.655 4706.955 ;
        RECT 1947.085 4706.675 1947.365 4706.955 ;
        RECT 1947.795 4706.675 1948.075 4706.955 ;
        RECT 1948.505 4706.675 1948.785 4706.955 ;
        RECT 1949.215 4706.675 1949.495 4706.955 ;
        RECT 1949.925 4706.675 1950.205 4706.955 ;
        RECT 1950.635 4706.675 1950.915 4706.955 ;
        RECT 1951.345 4706.675 1951.625 4706.955 ;
        RECT 1952.055 4706.675 1952.335 4706.955 ;
        RECT 1952.765 4706.675 1953.045 4706.955 ;
        RECT 1953.475 4706.675 1953.755 4706.955 ;
        RECT 1954.185 4706.675 1954.465 4706.955 ;
        RECT 1954.895 4706.675 1955.175 4706.955 ;
        RECT 1955.605 4706.675 1955.885 4706.955 ;
        RECT 1959.485 4706.675 1959.765 4706.955 ;
        RECT 1960.195 4706.675 1960.475 4706.955 ;
        RECT 1960.905 4706.675 1961.185 4706.955 ;
        RECT 1961.615 4706.675 1961.895 4706.955 ;
        RECT 1962.325 4706.675 1962.605 4706.955 ;
        RECT 1963.035 4706.675 1963.315 4706.955 ;
        RECT 1963.745 4706.675 1964.025 4706.955 ;
        RECT 1964.455 4706.675 1964.735 4706.955 ;
        RECT 1965.165 4706.675 1965.445 4706.955 ;
        RECT 1965.875 4706.675 1966.155 4706.955 ;
        RECT 1966.585 4706.675 1966.865 4706.955 ;
        RECT 1967.295 4706.675 1967.575 4706.955 ;
        RECT 1968.005 4706.675 1968.285 4706.955 ;
        RECT 2996.705 4706.675 2996.985 4706.955 ;
        RECT 2997.415 4706.675 2997.695 4706.955 ;
        RECT 2998.125 4706.675 2998.405 4706.955 ;
        RECT 2998.835 4706.675 2999.115 4706.955 ;
        RECT 2999.545 4706.675 2999.825 4706.955 ;
        RECT 3000.255 4706.675 3000.535 4706.955 ;
        RECT 3000.965 4706.675 3001.245 4706.955 ;
        RECT 3001.675 4706.675 3001.955 4706.955 ;
        RECT 3002.385 4706.675 3002.665 4706.955 ;
        RECT 3003.095 4706.675 3003.375 4706.955 ;
        RECT 3003.805 4706.675 3004.085 4706.955 ;
        RECT 3004.515 4706.675 3004.795 4706.955 ;
        RECT 3005.225 4706.675 3005.505 4706.955 ;
        RECT 3009.145 4706.675 3009.425 4706.955 ;
        RECT 3009.855 4706.675 3010.135 4706.955 ;
        RECT 3010.565 4706.675 3010.845 4706.955 ;
        RECT 3011.275 4706.675 3011.555 4706.955 ;
        RECT 3011.985 4706.675 3012.265 4706.955 ;
        RECT 3012.695 4706.675 3012.975 4706.955 ;
        RECT 3013.405 4706.675 3013.685 4706.955 ;
        RECT 3014.115 4706.675 3014.395 4706.955 ;
        RECT 3014.825 4706.675 3015.105 4706.955 ;
        RECT 3015.535 4706.675 3015.815 4706.955 ;
        RECT 3016.245 4706.675 3016.525 4706.955 ;
        RECT 3016.955 4706.675 3017.235 4706.955 ;
        RECT 3017.665 4706.675 3017.945 4706.955 ;
        RECT 3018.375 4706.675 3018.655 4706.955 ;
        RECT 3025.255 4706.675 3025.535 4706.955 ;
        RECT 3025.965 4706.675 3026.245 4706.955 ;
        RECT 3026.675 4706.675 3026.955 4706.955 ;
        RECT 3027.385 4706.675 3027.665 4706.955 ;
        RECT 3028.095 4706.675 3028.375 4706.955 ;
        RECT 3028.805 4706.675 3029.085 4706.955 ;
        RECT 3029.515 4706.675 3029.795 4706.955 ;
        RECT 3030.225 4706.675 3030.505 4706.955 ;
        RECT 3034.525 4706.675 3034.805 4706.955 ;
        RECT 3035.235 4706.675 3035.515 4706.955 ;
        RECT 3035.945 4706.675 3036.225 4706.955 ;
        RECT 3036.655 4706.675 3036.935 4706.955 ;
        RECT 3037.365 4706.675 3037.645 4706.955 ;
        RECT 3038.075 4706.675 3038.355 4706.955 ;
        RECT 3038.785 4706.675 3039.065 4706.955 ;
        RECT 3039.495 4706.675 3039.775 4706.955 ;
        RECT 3040.205 4706.675 3040.485 4706.955 ;
        RECT 3040.915 4706.675 3041.195 4706.955 ;
        RECT 3041.625 4706.675 3041.905 4706.955 ;
        RECT 3042.335 4706.675 3042.615 4706.955 ;
        RECT 3046.375 4706.675 3046.655 4706.955 ;
        RECT 3047.085 4706.675 3047.365 4706.955 ;
        RECT 3047.795 4706.675 3048.075 4706.955 ;
        RECT 3048.505 4706.675 3048.785 4706.955 ;
        RECT 3049.215 4706.675 3049.495 4706.955 ;
        RECT 3049.925 4706.675 3050.205 4706.955 ;
        RECT 3050.635 4706.675 3050.915 4706.955 ;
        RECT 3051.345 4706.675 3051.625 4706.955 ;
        RECT 3052.055 4706.675 3052.335 4706.955 ;
        RECT 3052.765 4706.675 3053.045 4706.955 ;
        RECT 3053.475 4706.675 3053.755 4706.955 ;
        RECT 3054.185 4706.675 3054.465 4706.955 ;
        RECT 3054.895 4706.675 3055.175 4706.955 ;
        RECT 3055.605 4706.675 3055.885 4706.955 ;
        RECT 3059.485 4706.675 3059.765 4706.955 ;
        RECT 3060.195 4706.675 3060.475 4706.955 ;
        RECT 3060.905 4706.675 3061.185 4706.955 ;
        RECT 3061.615 4706.675 3061.895 4706.955 ;
        RECT 3062.325 4706.675 3062.605 4706.955 ;
        RECT 3063.035 4706.675 3063.315 4706.955 ;
        RECT 3063.745 4706.675 3064.025 4706.955 ;
        RECT 3064.455 4706.675 3064.735 4706.955 ;
        RECT 3065.165 4706.675 3065.445 4706.955 ;
        RECT 3065.875 4706.675 3066.155 4706.955 ;
        RECT 3066.585 4706.675 3066.865 4706.955 ;
        RECT 3067.295 4706.675 3067.575 4706.955 ;
        RECT 3068.005 4706.675 3068.285 4706.955 ;
        RECT 1896.705 4705.965 1896.985 4706.245 ;
        RECT 1897.415 4705.965 1897.695 4706.245 ;
        RECT 1898.125 4705.965 1898.405 4706.245 ;
        RECT 1898.835 4705.965 1899.115 4706.245 ;
        RECT 1899.545 4705.965 1899.825 4706.245 ;
        RECT 1909.145 4705.965 1909.425 4706.245 ;
        RECT 1909.855 4705.965 1910.135 4706.245 ;
        RECT 1910.565 4705.965 1910.845 4706.245 ;
        RECT 1911.275 4705.965 1911.555 4706.245 ;
        RECT 1911.985 4705.965 1912.265 4706.245 ;
        RECT 1912.695 4705.965 1912.975 4706.245 ;
        RECT 1913.405 4705.965 1913.685 4706.245 ;
        RECT 1914.115 4705.965 1914.395 4706.245 ;
        RECT 1914.825 4705.965 1915.105 4706.245 ;
        RECT 1915.535 4705.965 1915.815 4706.245 ;
        RECT 1916.245 4705.965 1916.525 4706.245 ;
        RECT 1916.955 4705.965 1917.235 4706.245 ;
        RECT 1917.665 4705.965 1917.945 4706.245 ;
        RECT 1918.375 4705.965 1918.655 4706.245 ;
        RECT 1920.995 4705.965 1921.275 4706.245 ;
        RECT 1921.705 4705.965 1921.985 4706.245 ;
        RECT 1922.415 4705.965 1922.695 4706.245 ;
        RECT 1926.675 4705.965 1926.955 4706.245 ;
        RECT 1927.385 4705.965 1927.665 4706.245 ;
        RECT 1928.095 4705.965 1928.375 4706.245 ;
        RECT 1928.805 4705.965 1929.085 4706.245 ;
        RECT 1929.515 4705.965 1929.795 4706.245 ;
        RECT 1930.225 4705.965 1930.505 4706.245 ;
        RECT 1934.525 4705.965 1934.805 4706.245 ;
        RECT 1935.235 4705.965 1935.515 4706.245 ;
        RECT 1935.945 4705.965 1936.225 4706.245 ;
        RECT 1936.655 4705.965 1936.935 4706.245 ;
        RECT 1937.365 4705.965 1937.645 4706.245 ;
        RECT 1938.075 4705.965 1938.355 4706.245 ;
        RECT 1938.785 4705.965 1939.065 4706.245 ;
        RECT 1939.495 4705.965 1939.775 4706.245 ;
        RECT 1940.205 4705.965 1940.485 4706.245 ;
        RECT 1940.915 4705.965 1941.195 4706.245 ;
        RECT 1941.625 4705.965 1941.905 4706.245 ;
        RECT 1942.335 4705.965 1942.615 4706.245 ;
        RECT 1943.045 4705.965 1943.325 4706.245 ;
        RECT 1943.755 4705.965 1944.035 4706.245 ;
        RECT 1946.375 4705.965 1946.655 4706.245 ;
        RECT 1947.085 4705.965 1947.365 4706.245 ;
        RECT 1947.795 4705.965 1948.075 4706.245 ;
        RECT 1948.505 4705.965 1948.785 4706.245 ;
        RECT 1949.215 4705.965 1949.495 4706.245 ;
        RECT 1949.925 4705.965 1950.205 4706.245 ;
        RECT 1950.635 4705.965 1950.915 4706.245 ;
        RECT 1951.345 4705.965 1951.625 4706.245 ;
        RECT 1952.055 4705.965 1952.335 4706.245 ;
        RECT 1952.765 4705.965 1953.045 4706.245 ;
        RECT 1953.475 4705.965 1953.755 4706.245 ;
        RECT 1954.185 4705.965 1954.465 4706.245 ;
        RECT 1954.895 4705.965 1955.175 4706.245 ;
        RECT 1955.605 4705.965 1955.885 4706.245 ;
        RECT 1959.485 4705.965 1959.765 4706.245 ;
        RECT 1960.195 4705.965 1960.475 4706.245 ;
        RECT 1960.905 4705.965 1961.185 4706.245 ;
        RECT 1961.615 4705.965 1961.895 4706.245 ;
        RECT 1962.325 4705.965 1962.605 4706.245 ;
        RECT 1963.035 4705.965 1963.315 4706.245 ;
        RECT 1963.745 4705.965 1964.025 4706.245 ;
        RECT 1964.455 4705.965 1964.735 4706.245 ;
        RECT 1965.165 4705.965 1965.445 4706.245 ;
        RECT 1965.875 4705.965 1966.155 4706.245 ;
        RECT 1966.585 4705.965 1966.865 4706.245 ;
        RECT 1967.295 4705.965 1967.575 4706.245 ;
        RECT 1968.005 4705.965 1968.285 4706.245 ;
        RECT 2996.705 4705.965 2996.985 4706.245 ;
        RECT 2997.415 4705.965 2997.695 4706.245 ;
        RECT 2998.125 4705.965 2998.405 4706.245 ;
        RECT 2998.835 4705.965 2999.115 4706.245 ;
        RECT 2999.545 4705.965 2999.825 4706.245 ;
        RECT 3000.255 4705.965 3000.535 4706.245 ;
        RECT 3000.965 4705.965 3001.245 4706.245 ;
        RECT 3001.675 4705.965 3001.955 4706.245 ;
        RECT 3002.385 4705.965 3002.665 4706.245 ;
        RECT 3003.095 4705.965 3003.375 4706.245 ;
        RECT 3003.805 4705.965 3004.085 4706.245 ;
        RECT 3004.515 4705.965 3004.795 4706.245 ;
        RECT 3005.225 4705.965 3005.505 4706.245 ;
        RECT 3009.145 4705.965 3009.425 4706.245 ;
        RECT 3009.855 4705.965 3010.135 4706.245 ;
        RECT 3010.565 4705.965 3010.845 4706.245 ;
        RECT 3011.275 4705.965 3011.555 4706.245 ;
        RECT 3011.985 4705.965 3012.265 4706.245 ;
        RECT 3012.695 4705.965 3012.975 4706.245 ;
        RECT 3013.405 4705.965 3013.685 4706.245 ;
        RECT 3014.115 4705.965 3014.395 4706.245 ;
        RECT 3014.825 4705.965 3015.105 4706.245 ;
        RECT 3015.535 4705.965 3015.815 4706.245 ;
        RECT 3016.245 4705.965 3016.525 4706.245 ;
        RECT 3016.955 4705.965 3017.235 4706.245 ;
        RECT 3017.665 4705.965 3017.945 4706.245 ;
        RECT 3018.375 4705.965 3018.655 4706.245 ;
        RECT 3025.255 4705.965 3025.535 4706.245 ;
        RECT 3025.965 4705.965 3026.245 4706.245 ;
        RECT 3026.675 4705.965 3026.955 4706.245 ;
        RECT 3027.385 4705.965 3027.665 4706.245 ;
        RECT 3028.095 4705.965 3028.375 4706.245 ;
        RECT 3028.805 4705.965 3029.085 4706.245 ;
        RECT 3029.515 4705.965 3029.795 4706.245 ;
        RECT 3030.225 4705.965 3030.505 4706.245 ;
        RECT 3034.525 4705.965 3034.805 4706.245 ;
        RECT 3035.235 4705.965 3035.515 4706.245 ;
        RECT 3035.945 4705.965 3036.225 4706.245 ;
        RECT 3036.655 4705.965 3036.935 4706.245 ;
        RECT 3037.365 4705.965 3037.645 4706.245 ;
        RECT 3038.075 4705.965 3038.355 4706.245 ;
        RECT 3038.785 4705.965 3039.065 4706.245 ;
        RECT 3039.495 4705.965 3039.775 4706.245 ;
        RECT 3040.205 4705.965 3040.485 4706.245 ;
        RECT 3040.915 4705.965 3041.195 4706.245 ;
        RECT 3041.625 4705.965 3041.905 4706.245 ;
        RECT 3042.335 4705.965 3042.615 4706.245 ;
        RECT 3046.375 4705.965 3046.655 4706.245 ;
        RECT 3047.085 4705.965 3047.365 4706.245 ;
        RECT 3047.795 4705.965 3048.075 4706.245 ;
        RECT 3048.505 4705.965 3048.785 4706.245 ;
        RECT 3049.215 4705.965 3049.495 4706.245 ;
        RECT 3049.925 4705.965 3050.205 4706.245 ;
        RECT 3050.635 4705.965 3050.915 4706.245 ;
        RECT 3051.345 4705.965 3051.625 4706.245 ;
        RECT 3052.055 4705.965 3052.335 4706.245 ;
        RECT 3052.765 4705.965 3053.045 4706.245 ;
        RECT 3053.475 4705.965 3053.755 4706.245 ;
        RECT 3054.185 4705.965 3054.465 4706.245 ;
        RECT 3054.895 4705.965 3055.175 4706.245 ;
        RECT 3055.605 4705.965 3055.885 4706.245 ;
        RECT 3059.485 4705.965 3059.765 4706.245 ;
        RECT 3060.195 4705.965 3060.475 4706.245 ;
        RECT 3060.905 4705.965 3061.185 4706.245 ;
        RECT 3061.615 4705.965 3061.895 4706.245 ;
        RECT 3062.325 4705.965 3062.605 4706.245 ;
        RECT 3063.035 4705.965 3063.315 4706.245 ;
        RECT 3063.745 4705.965 3064.025 4706.245 ;
        RECT 3064.455 4705.965 3064.735 4706.245 ;
        RECT 3065.165 4705.965 3065.445 4706.245 ;
        RECT 3065.875 4705.965 3066.155 4706.245 ;
        RECT 3066.585 4705.965 3066.865 4706.245 ;
        RECT 3067.295 4705.965 3067.575 4706.245 ;
        RECT 3068.005 4705.965 3068.285 4706.245 ;
        RECT 1896.705 4705.255 1896.985 4705.535 ;
        RECT 1897.415 4705.255 1897.695 4705.535 ;
        RECT 1898.125 4705.255 1898.405 4705.535 ;
        RECT 1898.835 4705.255 1899.115 4705.535 ;
        RECT 1899.545 4705.255 1899.825 4705.535 ;
        RECT 1909.145 4705.255 1909.425 4705.535 ;
        RECT 1909.855 4705.255 1910.135 4705.535 ;
        RECT 1910.565 4705.255 1910.845 4705.535 ;
        RECT 1911.275 4705.255 1911.555 4705.535 ;
        RECT 1911.985 4705.255 1912.265 4705.535 ;
        RECT 1912.695 4705.255 1912.975 4705.535 ;
        RECT 1913.405 4705.255 1913.685 4705.535 ;
        RECT 1914.115 4705.255 1914.395 4705.535 ;
        RECT 1914.825 4705.255 1915.105 4705.535 ;
        RECT 1915.535 4705.255 1915.815 4705.535 ;
        RECT 1916.245 4705.255 1916.525 4705.535 ;
        RECT 1916.955 4705.255 1917.235 4705.535 ;
        RECT 1917.665 4705.255 1917.945 4705.535 ;
        RECT 1918.375 4705.255 1918.655 4705.535 ;
        RECT 1920.995 4705.255 1921.275 4705.535 ;
        RECT 1921.705 4705.255 1921.985 4705.535 ;
        RECT 1922.415 4705.255 1922.695 4705.535 ;
        RECT 1926.675 4705.255 1926.955 4705.535 ;
        RECT 1927.385 4705.255 1927.665 4705.535 ;
        RECT 1928.095 4705.255 1928.375 4705.535 ;
        RECT 1928.805 4705.255 1929.085 4705.535 ;
        RECT 1929.515 4705.255 1929.795 4705.535 ;
        RECT 1930.225 4705.255 1930.505 4705.535 ;
        RECT 1934.525 4705.255 1934.805 4705.535 ;
        RECT 1935.235 4705.255 1935.515 4705.535 ;
        RECT 1935.945 4705.255 1936.225 4705.535 ;
        RECT 1936.655 4705.255 1936.935 4705.535 ;
        RECT 1937.365 4705.255 1937.645 4705.535 ;
        RECT 1938.075 4705.255 1938.355 4705.535 ;
        RECT 1938.785 4705.255 1939.065 4705.535 ;
        RECT 1939.495 4705.255 1939.775 4705.535 ;
        RECT 1940.205 4705.255 1940.485 4705.535 ;
        RECT 1940.915 4705.255 1941.195 4705.535 ;
        RECT 1941.625 4705.255 1941.905 4705.535 ;
        RECT 1942.335 4705.255 1942.615 4705.535 ;
        RECT 1943.045 4705.255 1943.325 4705.535 ;
        RECT 1943.755 4705.255 1944.035 4705.535 ;
        RECT 1946.375 4705.255 1946.655 4705.535 ;
        RECT 1947.085 4705.255 1947.365 4705.535 ;
        RECT 1947.795 4705.255 1948.075 4705.535 ;
        RECT 1948.505 4705.255 1948.785 4705.535 ;
        RECT 1949.215 4705.255 1949.495 4705.535 ;
        RECT 1949.925 4705.255 1950.205 4705.535 ;
        RECT 1950.635 4705.255 1950.915 4705.535 ;
        RECT 1951.345 4705.255 1951.625 4705.535 ;
        RECT 1952.055 4705.255 1952.335 4705.535 ;
        RECT 1952.765 4705.255 1953.045 4705.535 ;
        RECT 1953.475 4705.255 1953.755 4705.535 ;
        RECT 1954.185 4705.255 1954.465 4705.535 ;
        RECT 1954.895 4705.255 1955.175 4705.535 ;
        RECT 1955.605 4705.255 1955.885 4705.535 ;
        RECT 1959.485 4705.255 1959.765 4705.535 ;
        RECT 1960.195 4705.255 1960.475 4705.535 ;
        RECT 1960.905 4705.255 1961.185 4705.535 ;
        RECT 1961.615 4705.255 1961.895 4705.535 ;
        RECT 1962.325 4705.255 1962.605 4705.535 ;
        RECT 1963.035 4705.255 1963.315 4705.535 ;
        RECT 1963.745 4705.255 1964.025 4705.535 ;
        RECT 1964.455 4705.255 1964.735 4705.535 ;
        RECT 1965.165 4705.255 1965.445 4705.535 ;
        RECT 1965.875 4705.255 1966.155 4705.535 ;
        RECT 1966.585 4705.255 1966.865 4705.535 ;
        RECT 1967.295 4705.255 1967.575 4705.535 ;
        RECT 1968.005 4705.255 1968.285 4705.535 ;
        RECT 2996.705 4705.255 2996.985 4705.535 ;
        RECT 2997.415 4705.255 2997.695 4705.535 ;
        RECT 2998.125 4705.255 2998.405 4705.535 ;
        RECT 2998.835 4705.255 2999.115 4705.535 ;
        RECT 2999.545 4705.255 2999.825 4705.535 ;
        RECT 3000.255 4705.255 3000.535 4705.535 ;
        RECT 3000.965 4705.255 3001.245 4705.535 ;
        RECT 3001.675 4705.255 3001.955 4705.535 ;
        RECT 3002.385 4705.255 3002.665 4705.535 ;
        RECT 3003.095 4705.255 3003.375 4705.535 ;
        RECT 3003.805 4705.255 3004.085 4705.535 ;
        RECT 3004.515 4705.255 3004.795 4705.535 ;
        RECT 3005.225 4705.255 3005.505 4705.535 ;
        RECT 3009.145 4705.255 3009.425 4705.535 ;
        RECT 3009.855 4705.255 3010.135 4705.535 ;
        RECT 3010.565 4705.255 3010.845 4705.535 ;
        RECT 3011.275 4705.255 3011.555 4705.535 ;
        RECT 3011.985 4705.255 3012.265 4705.535 ;
        RECT 3012.695 4705.255 3012.975 4705.535 ;
        RECT 3013.405 4705.255 3013.685 4705.535 ;
        RECT 3014.115 4705.255 3014.395 4705.535 ;
        RECT 3014.825 4705.255 3015.105 4705.535 ;
        RECT 3015.535 4705.255 3015.815 4705.535 ;
        RECT 3016.245 4705.255 3016.525 4705.535 ;
        RECT 3016.955 4705.255 3017.235 4705.535 ;
        RECT 3017.665 4705.255 3017.945 4705.535 ;
        RECT 3018.375 4705.255 3018.655 4705.535 ;
        RECT 3025.255 4705.255 3025.535 4705.535 ;
        RECT 3025.965 4705.255 3026.245 4705.535 ;
        RECT 3026.675 4705.255 3026.955 4705.535 ;
        RECT 3027.385 4705.255 3027.665 4705.535 ;
        RECT 3028.095 4705.255 3028.375 4705.535 ;
        RECT 3028.805 4705.255 3029.085 4705.535 ;
        RECT 3029.515 4705.255 3029.795 4705.535 ;
        RECT 3030.225 4705.255 3030.505 4705.535 ;
        RECT 3034.525 4705.255 3034.805 4705.535 ;
        RECT 3035.235 4705.255 3035.515 4705.535 ;
        RECT 3035.945 4705.255 3036.225 4705.535 ;
        RECT 3036.655 4705.255 3036.935 4705.535 ;
        RECT 3037.365 4705.255 3037.645 4705.535 ;
        RECT 3038.075 4705.255 3038.355 4705.535 ;
        RECT 3038.785 4705.255 3039.065 4705.535 ;
        RECT 3039.495 4705.255 3039.775 4705.535 ;
        RECT 3040.205 4705.255 3040.485 4705.535 ;
        RECT 3040.915 4705.255 3041.195 4705.535 ;
        RECT 3041.625 4705.255 3041.905 4705.535 ;
        RECT 3042.335 4705.255 3042.615 4705.535 ;
        RECT 3046.375 4705.255 3046.655 4705.535 ;
        RECT 3047.085 4705.255 3047.365 4705.535 ;
        RECT 3047.795 4705.255 3048.075 4705.535 ;
        RECT 3048.505 4705.255 3048.785 4705.535 ;
        RECT 3049.215 4705.255 3049.495 4705.535 ;
        RECT 3049.925 4705.255 3050.205 4705.535 ;
        RECT 3050.635 4705.255 3050.915 4705.535 ;
        RECT 3051.345 4705.255 3051.625 4705.535 ;
        RECT 3052.055 4705.255 3052.335 4705.535 ;
        RECT 3052.765 4705.255 3053.045 4705.535 ;
        RECT 3053.475 4705.255 3053.755 4705.535 ;
        RECT 3054.185 4705.255 3054.465 4705.535 ;
        RECT 3054.895 4705.255 3055.175 4705.535 ;
        RECT 3055.605 4705.255 3055.885 4705.535 ;
        RECT 3059.485 4705.255 3059.765 4705.535 ;
        RECT 3060.195 4705.255 3060.475 4705.535 ;
        RECT 3060.905 4705.255 3061.185 4705.535 ;
        RECT 3061.615 4705.255 3061.895 4705.535 ;
        RECT 3062.325 4705.255 3062.605 4705.535 ;
        RECT 3063.035 4705.255 3063.315 4705.535 ;
        RECT 3063.745 4705.255 3064.025 4705.535 ;
        RECT 3064.455 4705.255 3064.735 4705.535 ;
        RECT 3065.165 4705.255 3065.445 4705.535 ;
        RECT 3065.875 4705.255 3066.155 4705.535 ;
        RECT 3066.585 4705.255 3066.865 4705.535 ;
        RECT 3067.295 4705.255 3067.575 4705.535 ;
        RECT 3068.005 4705.255 3068.285 4705.535 ;
        RECT 1896.705 4704.545 1896.985 4704.825 ;
        RECT 1897.415 4704.545 1897.695 4704.825 ;
        RECT 1898.125 4704.545 1898.405 4704.825 ;
        RECT 1898.835 4704.545 1899.115 4704.825 ;
        RECT 1899.545 4704.545 1899.825 4704.825 ;
        RECT 1909.145 4704.545 1909.425 4704.825 ;
        RECT 1909.855 4704.545 1910.135 4704.825 ;
        RECT 1910.565 4704.545 1910.845 4704.825 ;
        RECT 1911.275 4704.545 1911.555 4704.825 ;
        RECT 1911.985 4704.545 1912.265 4704.825 ;
        RECT 1912.695 4704.545 1912.975 4704.825 ;
        RECT 1913.405 4704.545 1913.685 4704.825 ;
        RECT 1914.115 4704.545 1914.395 4704.825 ;
        RECT 1914.825 4704.545 1915.105 4704.825 ;
        RECT 1915.535 4704.545 1915.815 4704.825 ;
        RECT 1916.245 4704.545 1916.525 4704.825 ;
        RECT 1916.955 4704.545 1917.235 4704.825 ;
        RECT 1917.665 4704.545 1917.945 4704.825 ;
        RECT 1918.375 4704.545 1918.655 4704.825 ;
        RECT 1920.995 4704.545 1921.275 4704.825 ;
        RECT 1921.705 4704.545 1921.985 4704.825 ;
        RECT 1922.415 4704.545 1922.695 4704.825 ;
        RECT 1926.675 4704.545 1926.955 4704.825 ;
        RECT 1927.385 4704.545 1927.665 4704.825 ;
        RECT 1928.095 4704.545 1928.375 4704.825 ;
        RECT 1928.805 4704.545 1929.085 4704.825 ;
        RECT 1929.515 4704.545 1929.795 4704.825 ;
        RECT 1930.225 4704.545 1930.505 4704.825 ;
        RECT 1934.525 4704.545 1934.805 4704.825 ;
        RECT 1935.235 4704.545 1935.515 4704.825 ;
        RECT 1935.945 4704.545 1936.225 4704.825 ;
        RECT 1936.655 4704.545 1936.935 4704.825 ;
        RECT 1937.365 4704.545 1937.645 4704.825 ;
        RECT 1938.075 4704.545 1938.355 4704.825 ;
        RECT 1938.785 4704.545 1939.065 4704.825 ;
        RECT 1939.495 4704.545 1939.775 4704.825 ;
        RECT 1940.205 4704.545 1940.485 4704.825 ;
        RECT 1940.915 4704.545 1941.195 4704.825 ;
        RECT 1941.625 4704.545 1941.905 4704.825 ;
        RECT 1942.335 4704.545 1942.615 4704.825 ;
        RECT 1943.045 4704.545 1943.325 4704.825 ;
        RECT 1943.755 4704.545 1944.035 4704.825 ;
        RECT 1946.375 4704.545 1946.655 4704.825 ;
        RECT 1947.085 4704.545 1947.365 4704.825 ;
        RECT 1947.795 4704.545 1948.075 4704.825 ;
        RECT 1948.505 4704.545 1948.785 4704.825 ;
        RECT 1949.215 4704.545 1949.495 4704.825 ;
        RECT 1949.925 4704.545 1950.205 4704.825 ;
        RECT 1950.635 4704.545 1950.915 4704.825 ;
        RECT 1951.345 4704.545 1951.625 4704.825 ;
        RECT 1952.055 4704.545 1952.335 4704.825 ;
        RECT 1952.765 4704.545 1953.045 4704.825 ;
        RECT 1953.475 4704.545 1953.755 4704.825 ;
        RECT 1954.185 4704.545 1954.465 4704.825 ;
        RECT 1954.895 4704.545 1955.175 4704.825 ;
        RECT 1955.605 4704.545 1955.885 4704.825 ;
        RECT 1959.485 4704.545 1959.765 4704.825 ;
        RECT 1960.195 4704.545 1960.475 4704.825 ;
        RECT 1960.905 4704.545 1961.185 4704.825 ;
        RECT 1961.615 4704.545 1961.895 4704.825 ;
        RECT 1962.325 4704.545 1962.605 4704.825 ;
        RECT 1963.035 4704.545 1963.315 4704.825 ;
        RECT 1963.745 4704.545 1964.025 4704.825 ;
        RECT 1964.455 4704.545 1964.735 4704.825 ;
        RECT 1965.165 4704.545 1965.445 4704.825 ;
        RECT 1965.875 4704.545 1966.155 4704.825 ;
        RECT 1966.585 4704.545 1966.865 4704.825 ;
        RECT 1967.295 4704.545 1967.575 4704.825 ;
        RECT 1968.005 4704.545 1968.285 4704.825 ;
        RECT 2996.705 4704.545 2996.985 4704.825 ;
        RECT 2997.415 4704.545 2997.695 4704.825 ;
        RECT 2998.125 4704.545 2998.405 4704.825 ;
        RECT 2998.835 4704.545 2999.115 4704.825 ;
        RECT 2999.545 4704.545 2999.825 4704.825 ;
        RECT 3000.255 4704.545 3000.535 4704.825 ;
        RECT 3000.965 4704.545 3001.245 4704.825 ;
        RECT 3001.675 4704.545 3001.955 4704.825 ;
        RECT 3002.385 4704.545 3002.665 4704.825 ;
        RECT 3003.095 4704.545 3003.375 4704.825 ;
        RECT 3003.805 4704.545 3004.085 4704.825 ;
        RECT 3004.515 4704.545 3004.795 4704.825 ;
        RECT 3005.225 4704.545 3005.505 4704.825 ;
        RECT 3009.145 4704.545 3009.425 4704.825 ;
        RECT 3009.855 4704.545 3010.135 4704.825 ;
        RECT 3010.565 4704.545 3010.845 4704.825 ;
        RECT 3011.275 4704.545 3011.555 4704.825 ;
        RECT 3011.985 4704.545 3012.265 4704.825 ;
        RECT 3012.695 4704.545 3012.975 4704.825 ;
        RECT 3013.405 4704.545 3013.685 4704.825 ;
        RECT 3014.115 4704.545 3014.395 4704.825 ;
        RECT 3014.825 4704.545 3015.105 4704.825 ;
        RECT 3015.535 4704.545 3015.815 4704.825 ;
        RECT 3016.245 4704.545 3016.525 4704.825 ;
        RECT 3016.955 4704.545 3017.235 4704.825 ;
        RECT 3017.665 4704.545 3017.945 4704.825 ;
        RECT 3018.375 4704.545 3018.655 4704.825 ;
        RECT 3025.255 4704.545 3025.535 4704.825 ;
        RECT 3025.965 4704.545 3026.245 4704.825 ;
        RECT 3026.675 4704.545 3026.955 4704.825 ;
        RECT 3027.385 4704.545 3027.665 4704.825 ;
        RECT 3028.095 4704.545 3028.375 4704.825 ;
        RECT 3028.805 4704.545 3029.085 4704.825 ;
        RECT 3029.515 4704.545 3029.795 4704.825 ;
        RECT 3030.225 4704.545 3030.505 4704.825 ;
        RECT 3034.525 4704.545 3034.805 4704.825 ;
        RECT 3035.235 4704.545 3035.515 4704.825 ;
        RECT 3035.945 4704.545 3036.225 4704.825 ;
        RECT 3036.655 4704.545 3036.935 4704.825 ;
        RECT 3037.365 4704.545 3037.645 4704.825 ;
        RECT 3038.075 4704.545 3038.355 4704.825 ;
        RECT 3038.785 4704.545 3039.065 4704.825 ;
        RECT 3039.495 4704.545 3039.775 4704.825 ;
        RECT 3040.205 4704.545 3040.485 4704.825 ;
        RECT 3040.915 4704.545 3041.195 4704.825 ;
        RECT 3041.625 4704.545 3041.905 4704.825 ;
        RECT 3042.335 4704.545 3042.615 4704.825 ;
        RECT 3046.375 4704.545 3046.655 4704.825 ;
        RECT 3047.085 4704.545 3047.365 4704.825 ;
        RECT 3047.795 4704.545 3048.075 4704.825 ;
        RECT 3048.505 4704.545 3048.785 4704.825 ;
        RECT 3049.215 4704.545 3049.495 4704.825 ;
        RECT 3049.925 4704.545 3050.205 4704.825 ;
        RECT 3050.635 4704.545 3050.915 4704.825 ;
        RECT 3051.345 4704.545 3051.625 4704.825 ;
        RECT 3052.055 4704.545 3052.335 4704.825 ;
        RECT 3052.765 4704.545 3053.045 4704.825 ;
        RECT 3053.475 4704.545 3053.755 4704.825 ;
        RECT 3054.185 4704.545 3054.465 4704.825 ;
        RECT 3054.895 4704.545 3055.175 4704.825 ;
        RECT 3055.605 4704.545 3055.885 4704.825 ;
        RECT 3059.485 4704.545 3059.765 4704.825 ;
        RECT 3060.195 4704.545 3060.475 4704.825 ;
        RECT 3060.905 4704.545 3061.185 4704.825 ;
        RECT 3061.615 4704.545 3061.895 4704.825 ;
        RECT 3062.325 4704.545 3062.605 4704.825 ;
        RECT 3063.035 4704.545 3063.315 4704.825 ;
        RECT 3063.745 4704.545 3064.025 4704.825 ;
        RECT 3064.455 4704.545 3064.735 4704.825 ;
        RECT 3065.165 4704.545 3065.445 4704.825 ;
        RECT 3065.875 4704.545 3066.155 4704.825 ;
        RECT 3066.585 4704.545 3066.865 4704.825 ;
        RECT 3067.295 4704.545 3067.575 4704.825 ;
        RECT 3068.005 4704.545 3068.285 4704.825 ;
        RECT 1896.705 4703.835 1896.985 4704.115 ;
        RECT 1897.415 4703.835 1897.695 4704.115 ;
        RECT 1898.125 4703.835 1898.405 4704.115 ;
        RECT 1898.835 4703.835 1899.115 4704.115 ;
        RECT 1899.545 4703.835 1899.825 4704.115 ;
        RECT 1909.145 4703.835 1909.425 4704.115 ;
        RECT 1909.855 4703.835 1910.135 4704.115 ;
        RECT 1910.565 4703.835 1910.845 4704.115 ;
        RECT 1911.275 4703.835 1911.555 4704.115 ;
        RECT 1911.985 4703.835 1912.265 4704.115 ;
        RECT 1912.695 4703.835 1912.975 4704.115 ;
        RECT 1913.405 4703.835 1913.685 4704.115 ;
        RECT 1914.115 4703.835 1914.395 4704.115 ;
        RECT 1914.825 4703.835 1915.105 4704.115 ;
        RECT 1915.535 4703.835 1915.815 4704.115 ;
        RECT 1916.245 4703.835 1916.525 4704.115 ;
        RECT 1916.955 4703.835 1917.235 4704.115 ;
        RECT 1917.665 4703.835 1917.945 4704.115 ;
        RECT 1918.375 4703.835 1918.655 4704.115 ;
        RECT 1920.995 4703.835 1921.275 4704.115 ;
        RECT 1921.705 4703.835 1921.985 4704.115 ;
        RECT 1922.415 4703.835 1922.695 4704.115 ;
        RECT 1926.675 4703.835 1926.955 4704.115 ;
        RECT 1927.385 4703.835 1927.665 4704.115 ;
        RECT 1928.095 4703.835 1928.375 4704.115 ;
        RECT 1928.805 4703.835 1929.085 4704.115 ;
        RECT 1929.515 4703.835 1929.795 4704.115 ;
        RECT 1930.225 4703.835 1930.505 4704.115 ;
        RECT 1934.525 4703.835 1934.805 4704.115 ;
        RECT 1935.235 4703.835 1935.515 4704.115 ;
        RECT 1935.945 4703.835 1936.225 4704.115 ;
        RECT 1936.655 4703.835 1936.935 4704.115 ;
        RECT 1937.365 4703.835 1937.645 4704.115 ;
        RECT 1938.075 4703.835 1938.355 4704.115 ;
        RECT 1938.785 4703.835 1939.065 4704.115 ;
        RECT 1939.495 4703.835 1939.775 4704.115 ;
        RECT 1940.205 4703.835 1940.485 4704.115 ;
        RECT 1940.915 4703.835 1941.195 4704.115 ;
        RECT 1941.625 4703.835 1941.905 4704.115 ;
        RECT 1942.335 4703.835 1942.615 4704.115 ;
        RECT 1943.045 4703.835 1943.325 4704.115 ;
        RECT 1943.755 4703.835 1944.035 4704.115 ;
        RECT 1946.375 4703.835 1946.655 4704.115 ;
        RECT 1947.085 4703.835 1947.365 4704.115 ;
        RECT 1947.795 4703.835 1948.075 4704.115 ;
        RECT 1948.505 4703.835 1948.785 4704.115 ;
        RECT 1949.215 4703.835 1949.495 4704.115 ;
        RECT 1949.925 4703.835 1950.205 4704.115 ;
        RECT 1950.635 4703.835 1950.915 4704.115 ;
        RECT 1951.345 4703.835 1951.625 4704.115 ;
        RECT 1952.055 4703.835 1952.335 4704.115 ;
        RECT 1952.765 4703.835 1953.045 4704.115 ;
        RECT 1953.475 4703.835 1953.755 4704.115 ;
        RECT 1954.185 4703.835 1954.465 4704.115 ;
        RECT 1954.895 4703.835 1955.175 4704.115 ;
        RECT 1955.605 4703.835 1955.885 4704.115 ;
        RECT 1959.485 4703.835 1959.765 4704.115 ;
        RECT 1960.195 4703.835 1960.475 4704.115 ;
        RECT 1960.905 4703.835 1961.185 4704.115 ;
        RECT 1961.615 4703.835 1961.895 4704.115 ;
        RECT 1962.325 4703.835 1962.605 4704.115 ;
        RECT 1963.035 4703.835 1963.315 4704.115 ;
        RECT 1963.745 4703.835 1964.025 4704.115 ;
        RECT 1964.455 4703.835 1964.735 4704.115 ;
        RECT 1965.165 4703.835 1965.445 4704.115 ;
        RECT 1965.875 4703.835 1966.155 4704.115 ;
        RECT 1966.585 4703.835 1966.865 4704.115 ;
        RECT 1967.295 4703.835 1967.575 4704.115 ;
        RECT 1968.005 4703.835 1968.285 4704.115 ;
        RECT 2996.705 4703.835 2996.985 4704.115 ;
        RECT 2997.415 4703.835 2997.695 4704.115 ;
        RECT 2998.125 4703.835 2998.405 4704.115 ;
        RECT 2998.835 4703.835 2999.115 4704.115 ;
        RECT 2999.545 4703.835 2999.825 4704.115 ;
        RECT 3000.255 4703.835 3000.535 4704.115 ;
        RECT 3000.965 4703.835 3001.245 4704.115 ;
        RECT 3001.675 4703.835 3001.955 4704.115 ;
        RECT 3002.385 4703.835 3002.665 4704.115 ;
        RECT 3003.095 4703.835 3003.375 4704.115 ;
        RECT 3003.805 4703.835 3004.085 4704.115 ;
        RECT 3004.515 4703.835 3004.795 4704.115 ;
        RECT 3005.225 4703.835 3005.505 4704.115 ;
        RECT 3009.145 4703.835 3009.425 4704.115 ;
        RECT 3009.855 4703.835 3010.135 4704.115 ;
        RECT 3010.565 4703.835 3010.845 4704.115 ;
        RECT 3011.275 4703.835 3011.555 4704.115 ;
        RECT 3011.985 4703.835 3012.265 4704.115 ;
        RECT 3012.695 4703.835 3012.975 4704.115 ;
        RECT 3013.405 4703.835 3013.685 4704.115 ;
        RECT 3014.115 4703.835 3014.395 4704.115 ;
        RECT 3014.825 4703.835 3015.105 4704.115 ;
        RECT 3015.535 4703.835 3015.815 4704.115 ;
        RECT 3016.245 4703.835 3016.525 4704.115 ;
        RECT 3016.955 4703.835 3017.235 4704.115 ;
        RECT 3017.665 4703.835 3017.945 4704.115 ;
        RECT 3018.375 4703.835 3018.655 4704.115 ;
        RECT 3025.255 4703.835 3025.535 4704.115 ;
        RECT 3025.965 4703.835 3026.245 4704.115 ;
        RECT 3026.675 4703.835 3026.955 4704.115 ;
        RECT 3027.385 4703.835 3027.665 4704.115 ;
        RECT 3028.095 4703.835 3028.375 4704.115 ;
        RECT 3028.805 4703.835 3029.085 4704.115 ;
        RECT 3029.515 4703.835 3029.795 4704.115 ;
        RECT 3030.225 4703.835 3030.505 4704.115 ;
        RECT 3034.525 4703.835 3034.805 4704.115 ;
        RECT 3035.235 4703.835 3035.515 4704.115 ;
        RECT 3035.945 4703.835 3036.225 4704.115 ;
        RECT 3036.655 4703.835 3036.935 4704.115 ;
        RECT 3037.365 4703.835 3037.645 4704.115 ;
        RECT 3038.075 4703.835 3038.355 4704.115 ;
        RECT 3038.785 4703.835 3039.065 4704.115 ;
        RECT 3039.495 4703.835 3039.775 4704.115 ;
        RECT 3040.205 4703.835 3040.485 4704.115 ;
        RECT 3040.915 4703.835 3041.195 4704.115 ;
        RECT 3041.625 4703.835 3041.905 4704.115 ;
        RECT 3042.335 4703.835 3042.615 4704.115 ;
        RECT 3046.375 4703.835 3046.655 4704.115 ;
        RECT 3047.085 4703.835 3047.365 4704.115 ;
        RECT 3047.795 4703.835 3048.075 4704.115 ;
        RECT 3048.505 4703.835 3048.785 4704.115 ;
        RECT 3049.215 4703.835 3049.495 4704.115 ;
        RECT 3049.925 4703.835 3050.205 4704.115 ;
        RECT 3050.635 4703.835 3050.915 4704.115 ;
        RECT 3051.345 4703.835 3051.625 4704.115 ;
        RECT 3052.055 4703.835 3052.335 4704.115 ;
        RECT 3052.765 4703.835 3053.045 4704.115 ;
        RECT 3053.475 4703.835 3053.755 4704.115 ;
        RECT 3054.185 4703.835 3054.465 4704.115 ;
        RECT 3054.895 4703.835 3055.175 4704.115 ;
        RECT 3055.605 4703.835 3055.885 4704.115 ;
        RECT 3059.485 4703.835 3059.765 4704.115 ;
        RECT 3060.195 4703.835 3060.475 4704.115 ;
        RECT 3060.905 4703.835 3061.185 4704.115 ;
        RECT 3061.615 4703.835 3061.895 4704.115 ;
        RECT 3062.325 4703.835 3062.605 4704.115 ;
        RECT 3063.035 4703.835 3063.315 4704.115 ;
        RECT 3063.745 4703.835 3064.025 4704.115 ;
        RECT 3064.455 4703.835 3064.735 4704.115 ;
        RECT 3065.165 4703.835 3065.445 4704.115 ;
        RECT 3065.875 4703.835 3066.155 4704.115 ;
        RECT 3066.585 4703.835 3066.865 4704.115 ;
        RECT 3067.295 4703.835 3067.575 4704.115 ;
        RECT 3068.005 4703.835 3068.285 4704.115 ;
        RECT 1896.705 4703.125 1896.985 4703.405 ;
        RECT 1897.415 4703.125 1897.695 4703.405 ;
        RECT 1898.125 4703.125 1898.405 4703.405 ;
        RECT 1898.835 4703.125 1899.115 4703.405 ;
        RECT 1899.545 4703.125 1899.825 4703.405 ;
        RECT 1909.145 4703.125 1909.425 4703.405 ;
        RECT 1909.855 4703.125 1910.135 4703.405 ;
        RECT 1910.565 4703.125 1910.845 4703.405 ;
        RECT 1911.275 4703.125 1911.555 4703.405 ;
        RECT 1911.985 4703.125 1912.265 4703.405 ;
        RECT 1912.695 4703.125 1912.975 4703.405 ;
        RECT 1913.405 4703.125 1913.685 4703.405 ;
        RECT 1914.115 4703.125 1914.395 4703.405 ;
        RECT 1914.825 4703.125 1915.105 4703.405 ;
        RECT 1915.535 4703.125 1915.815 4703.405 ;
        RECT 1916.245 4703.125 1916.525 4703.405 ;
        RECT 1916.955 4703.125 1917.235 4703.405 ;
        RECT 1917.665 4703.125 1917.945 4703.405 ;
        RECT 1918.375 4703.125 1918.655 4703.405 ;
        RECT 1920.995 4703.125 1921.275 4703.405 ;
        RECT 1921.705 4703.125 1921.985 4703.405 ;
        RECT 1922.415 4703.125 1922.695 4703.405 ;
        RECT 1926.675 4703.125 1926.955 4703.405 ;
        RECT 1927.385 4703.125 1927.665 4703.405 ;
        RECT 1928.095 4703.125 1928.375 4703.405 ;
        RECT 1928.805 4703.125 1929.085 4703.405 ;
        RECT 1929.515 4703.125 1929.795 4703.405 ;
        RECT 1930.225 4703.125 1930.505 4703.405 ;
        RECT 1934.525 4703.125 1934.805 4703.405 ;
        RECT 1935.235 4703.125 1935.515 4703.405 ;
        RECT 1935.945 4703.125 1936.225 4703.405 ;
        RECT 1936.655 4703.125 1936.935 4703.405 ;
        RECT 1937.365 4703.125 1937.645 4703.405 ;
        RECT 1938.075 4703.125 1938.355 4703.405 ;
        RECT 1938.785 4703.125 1939.065 4703.405 ;
        RECT 1939.495 4703.125 1939.775 4703.405 ;
        RECT 1940.205 4703.125 1940.485 4703.405 ;
        RECT 1940.915 4703.125 1941.195 4703.405 ;
        RECT 1941.625 4703.125 1941.905 4703.405 ;
        RECT 1942.335 4703.125 1942.615 4703.405 ;
        RECT 1943.045 4703.125 1943.325 4703.405 ;
        RECT 1943.755 4703.125 1944.035 4703.405 ;
        RECT 1946.375 4703.125 1946.655 4703.405 ;
        RECT 1947.085 4703.125 1947.365 4703.405 ;
        RECT 1947.795 4703.125 1948.075 4703.405 ;
        RECT 1948.505 4703.125 1948.785 4703.405 ;
        RECT 1949.215 4703.125 1949.495 4703.405 ;
        RECT 1949.925 4703.125 1950.205 4703.405 ;
        RECT 1950.635 4703.125 1950.915 4703.405 ;
        RECT 1951.345 4703.125 1951.625 4703.405 ;
        RECT 1952.055 4703.125 1952.335 4703.405 ;
        RECT 1952.765 4703.125 1953.045 4703.405 ;
        RECT 1953.475 4703.125 1953.755 4703.405 ;
        RECT 1954.185 4703.125 1954.465 4703.405 ;
        RECT 1954.895 4703.125 1955.175 4703.405 ;
        RECT 1955.605 4703.125 1955.885 4703.405 ;
        RECT 1959.485 4703.125 1959.765 4703.405 ;
        RECT 1960.195 4703.125 1960.475 4703.405 ;
        RECT 1960.905 4703.125 1961.185 4703.405 ;
        RECT 1961.615 4703.125 1961.895 4703.405 ;
        RECT 1962.325 4703.125 1962.605 4703.405 ;
        RECT 1963.035 4703.125 1963.315 4703.405 ;
        RECT 1963.745 4703.125 1964.025 4703.405 ;
        RECT 1964.455 4703.125 1964.735 4703.405 ;
        RECT 1965.165 4703.125 1965.445 4703.405 ;
        RECT 1965.875 4703.125 1966.155 4703.405 ;
        RECT 1966.585 4703.125 1966.865 4703.405 ;
        RECT 1967.295 4703.125 1967.575 4703.405 ;
        RECT 1968.005 4703.125 1968.285 4703.405 ;
        RECT 2996.705 4703.125 2996.985 4703.405 ;
        RECT 2997.415 4703.125 2997.695 4703.405 ;
        RECT 2998.125 4703.125 2998.405 4703.405 ;
        RECT 2998.835 4703.125 2999.115 4703.405 ;
        RECT 2999.545 4703.125 2999.825 4703.405 ;
        RECT 3000.255 4703.125 3000.535 4703.405 ;
        RECT 3000.965 4703.125 3001.245 4703.405 ;
        RECT 3001.675 4703.125 3001.955 4703.405 ;
        RECT 3002.385 4703.125 3002.665 4703.405 ;
        RECT 3003.095 4703.125 3003.375 4703.405 ;
        RECT 3003.805 4703.125 3004.085 4703.405 ;
        RECT 3004.515 4703.125 3004.795 4703.405 ;
        RECT 3005.225 4703.125 3005.505 4703.405 ;
        RECT 3009.145 4703.125 3009.425 4703.405 ;
        RECT 3009.855 4703.125 3010.135 4703.405 ;
        RECT 3010.565 4703.125 3010.845 4703.405 ;
        RECT 3011.275 4703.125 3011.555 4703.405 ;
        RECT 3011.985 4703.125 3012.265 4703.405 ;
        RECT 3012.695 4703.125 3012.975 4703.405 ;
        RECT 3013.405 4703.125 3013.685 4703.405 ;
        RECT 3014.115 4703.125 3014.395 4703.405 ;
        RECT 3014.825 4703.125 3015.105 4703.405 ;
        RECT 3015.535 4703.125 3015.815 4703.405 ;
        RECT 3016.245 4703.125 3016.525 4703.405 ;
        RECT 3016.955 4703.125 3017.235 4703.405 ;
        RECT 3017.665 4703.125 3017.945 4703.405 ;
        RECT 3018.375 4703.125 3018.655 4703.405 ;
        RECT 3025.255 4703.125 3025.535 4703.405 ;
        RECT 3025.965 4703.125 3026.245 4703.405 ;
        RECT 3026.675 4703.125 3026.955 4703.405 ;
        RECT 3027.385 4703.125 3027.665 4703.405 ;
        RECT 3028.095 4703.125 3028.375 4703.405 ;
        RECT 3028.805 4703.125 3029.085 4703.405 ;
        RECT 3029.515 4703.125 3029.795 4703.405 ;
        RECT 3030.225 4703.125 3030.505 4703.405 ;
        RECT 3034.525 4703.125 3034.805 4703.405 ;
        RECT 3035.235 4703.125 3035.515 4703.405 ;
        RECT 3035.945 4703.125 3036.225 4703.405 ;
        RECT 3036.655 4703.125 3036.935 4703.405 ;
        RECT 3037.365 4703.125 3037.645 4703.405 ;
        RECT 3038.075 4703.125 3038.355 4703.405 ;
        RECT 3038.785 4703.125 3039.065 4703.405 ;
        RECT 3039.495 4703.125 3039.775 4703.405 ;
        RECT 3040.205 4703.125 3040.485 4703.405 ;
        RECT 3040.915 4703.125 3041.195 4703.405 ;
        RECT 3041.625 4703.125 3041.905 4703.405 ;
        RECT 3042.335 4703.125 3042.615 4703.405 ;
        RECT 3046.375 4703.125 3046.655 4703.405 ;
        RECT 3047.085 4703.125 3047.365 4703.405 ;
        RECT 3047.795 4703.125 3048.075 4703.405 ;
        RECT 3048.505 4703.125 3048.785 4703.405 ;
        RECT 3049.215 4703.125 3049.495 4703.405 ;
        RECT 3049.925 4703.125 3050.205 4703.405 ;
        RECT 3050.635 4703.125 3050.915 4703.405 ;
        RECT 3051.345 4703.125 3051.625 4703.405 ;
        RECT 3052.055 4703.125 3052.335 4703.405 ;
        RECT 3052.765 4703.125 3053.045 4703.405 ;
        RECT 3053.475 4703.125 3053.755 4703.405 ;
        RECT 3054.185 4703.125 3054.465 4703.405 ;
        RECT 3054.895 4703.125 3055.175 4703.405 ;
        RECT 3055.605 4703.125 3055.885 4703.405 ;
        RECT 3059.485 4703.125 3059.765 4703.405 ;
        RECT 3060.195 4703.125 3060.475 4703.405 ;
        RECT 3060.905 4703.125 3061.185 4703.405 ;
        RECT 3061.615 4703.125 3061.895 4703.405 ;
        RECT 3062.325 4703.125 3062.605 4703.405 ;
        RECT 3063.035 4703.125 3063.315 4703.405 ;
        RECT 3063.745 4703.125 3064.025 4703.405 ;
        RECT 3064.455 4703.125 3064.735 4703.405 ;
        RECT 3065.165 4703.125 3065.445 4703.405 ;
        RECT 3065.875 4703.125 3066.155 4703.405 ;
        RECT 3066.585 4703.125 3066.865 4703.405 ;
        RECT 3067.295 4703.125 3067.575 4703.405 ;
        RECT 3068.005 4703.125 3068.285 4703.405 ;
        RECT 1896.705 4702.415 1896.985 4702.695 ;
        RECT 1897.415 4702.415 1897.695 4702.695 ;
        RECT 1898.125 4702.415 1898.405 4702.695 ;
        RECT 1898.835 4702.415 1899.115 4702.695 ;
        RECT 1899.545 4702.415 1899.825 4702.695 ;
        RECT 1909.145 4702.415 1909.425 4702.695 ;
        RECT 1909.855 4702.415 1910.135 4702.695 ;
        RECT 1910.565 4702.415 1910.845 4702.695 ;
        RECT 1911.275 4702.415 1911.555 4702.695 ;
        RECT 1911.985 4702.415 1912.265 4702.695 ;
        RECT 1912.695 4702.415 1912.975 4702.695 ;
        RECT 1913.405 4702.415 1913.685 4702.695 ;
        RECT 1914.115 4702.415 1914.395 4702.695 ;
        RECT 1914.825 4702.415 1915.105 4702.695 ;
        RECT 1915.535 4702.415 1915.815 4702.695 ;
        RECT 1916.245 4702.415 1916.525 4702.695 ;
        RECT 1916.955 4702.415 1917.235 4702.695 ;
        RECT 1917.665 4702.415 1917.945 4702.695 ;
        RECT 1918.375 4702.415 1918.655 4702.695 ;
        RECT 1920.995 4702.415 1921.275 4702.695 ;
        RECT 1921.705 4702.415 1921.985 4702.695 ;
        RECT 1922.415 4702.415 1922.695 4702.695 ;
        RECT 1926.675 4702.415 1926.955 4702.695 ;
        RECT 1927.385 4702.415 1927.665 4702.695 ;
        RECT 1928.095 4702.415 1928.375 4702.695 ;
        RECT 1928.805 4702.415 1929.085 4702.695 ;
        RECT 1929.515 4702.415 1929.795 4702.695 ;
        RECT 1930.225 4702.415 1930.505 4702.695 ;
        RECT 1934.525 4702.415 1934.805 4702.695 ;
        RECT 1935.235 4702.415 1935.515 4702.695 ;
        RECT 1935.945 4702.415 1936.225 4702.695 ;
        RECT 1936.655 4702.415 1936.935 4702.695 ;
        RECT 1937.365 4702.415 1937.645 4702.695 ;
        RECT 1938.075 4702.415 1938.355 4702.695 ;
        RECT 1938.785 4702.415 1939.065 4702.695 ;
        RECT 1939.495 4702.415 1939.775 4702.695 ;
        RECT 1940.205 4702.415 1940.485 4702.695 ;
        RECT 1940.915 4702.415 1941.195 4702.695 ;
        RECT 1941.625 4702.415 1941.905 4702.695 ;
        RECT 1942.335 4702.415 1942.615 4702.695 ;
        RECT 1943.045 4702.415 1943.325 4702.695 ;
        RECT 1943.755 4702.415 1944.035 4702.695 ;
        RECT 1946.375 4702.415 1946.655 4702.695 ;
        RECT 1947.085 4702.415 1947.365 4702.695 ;
        RECT 1947.795 4702.415 1948.075 4702.695 ;
        RECT 1948.505 4702.415 1948.785 4702.695 ;
        RECT 1949.215 4702.415 1949.495 4702.695 ;
        RECT 1949.925 4702.415 1950.205 4702.695 ;
        RECT 1950.635 4702.415 1950.915 4702.695 ;
        RECT 1951.345 4702.415 1951.625 4702.695 ;
        RECT 1952.055 4702.415 1952.335 4702.695 ;
        RECT 1952.765 4702.415 1953.045 4702.695 ;
        RECT 1953.475 4702.415 1953.755 4702.695 ;
        RECT 1954.185 4702.415 1954.465 4702.695 ;
        RECT 1954.895 4702.415 1955.175 4702.695 ;
        RECT 1955.605 4702.415 1955.885 4702.695 ;
        RECT 1959.485 4702.415 1959.765 4702.695 ;
        RECT 1960.195 4702.415 1960.475 4702.695 ;
        RECT 1960.905 4702.415 1961.185 4702.695 ;
        RECT 1961.615 4702.415 1961.895 4702.695 ;
        RECT 1962.325 4702.415 1962.605 4702.695 ;
        RECT 1963.035 4702.415 1963.315 4702.695 ;
        RECT 1963.745 4702.415 1964.025 4702.695 ;
        RECT 1964.455 4702.415 1964.735 4702.695 ;
        RECT 1965.165 4702.415 1965.445 4702.695 ;
        RECT 1965.875 4702.415 1966.155 4702.695 ;
        RECT 1966.585 4702.415 1966.865 4702.695 ;
        RECT 1967.295 4702.415 1967.575 4702.695 ;
        RECT 1968.005 4702.415 1968.285 4702.695 ;
        RECT 2996.705 4702.415 2996.985 4702.695 ;
        RECT 2997.415 4702.415 2997.695 4702.695 ;
        RECT 2998.125 4702.415 2998.405 4702.695 ;
        RECT 2998.835 4702.415 2999.115 4702.695 ;
        RECT 2999.545 4702.415 2999.825 4702.695 ;
        RECT 3000.255 4702.415 3000.535 4702.695 ;
        RECT 3000.965 4702.415 3001.245 4702.695 ;
        RECT 3001.675 4702.415 3001.955 4702.695 ;
        RECT 3002.385 4702.415 3002.665 4702.695 ;
        RECT 3003.095 4702.415 3003.375 4702.695 ;
        RECT 3003.805 4702.415 3004.085 4702.695 ;
        RECT 3004.515 4702.415 3004.795 4702.695 ;
        RECT 3005.225 4702.415 3005.505 4702.695 ;
        RECT 3009.145 4702.415 3009.425 4702.695 ;
        RECT 3009.855 4702.415 3010.135 4702.695 ;
        RECT 3010.565 4702.415 3010.845 4702.695 ;
        RECT 3011.275 4702.415 3011.555 4702.695 ;
        RECT 3011.985 4702.415 3012.265 4702.695 ;
        RECT 3012.695 4702.415 3012.975 4702.695 ;
        RECT 3013.405 4702.415 3013.685 4702.695 ;
        RECT 3014.115 4702.415 3014.395 4702.695 ;
        RECT 3014.825 4702.415 3015.105 4702.695 ;
        RECT 3015.535 4702.415 3015.815 4702.695 ;
        RECT 3016.245 4702.415 3016.525 4702.695 ;
        RECT 3016.955 4702.415 3017.235 4702.695 ;
        RECT 3017.665 4702.415 3017.945 4702.695 ;
        RECT 3018.375 4702.415 3018.655 4702.695 ;
        RECT 3025.255 4702.415 3025.535 4702.695 ;
        RECT 3025.965 4702.415 3026.245 4702.695 ;
        RECT 3026.675 4702.415 3026.955 4702.695 ;
        RECT 3027.385 4702.415 3027.665 4702.695 ;
        RECT 3028.095 4702.415 3028.375 4702.695 ;
        RECT 3028.805 4702.415 3029.085 4702.695 ;
        RECT 3029.515 4702.415 3029.795 4702.695 ;
        RECT 3030.225 4702.415 3030.505 4702.695 ;
        RECT 3034.525 4702.415 3034.805 4702.695 ;
        RECT 3035.235 4702.415 3035.515 4702.695 ;
        RECT 3035.945 4702.415 3036.225 4702.695 ;
        RECT 3036.655 4702.415 3036.935 4702.695 ;
        RECT 3037.365 4702.415 3037.645 4702.695 ;
        RECT 3038.075 4702.415 3038.355 4702.695 ;
        RECT 3038.785 4702.415 3039.065 4702.695 ;
        RECT 3039.495 4702.415 3039.775 4702.695 ;
        RECT 3040.205 4702.415 3040.485 4702.695 ;
        RECT 3040.915 4702.415 3041.195 4702.695 ;
        RECT 3041.625 4702.415 3041.905 4702.695 ;
        RECT 3042.335 4702.415 3042.615 4702.695 ;
        RECT 3046.375 4702.415 3046.655 4702.695 ;
        RECT 3047.085 4702.415 3047.365 4702.695 ;
        RECT 3047.795 4702.415 3048.075 4702.695 ;
        RECT 3048.505 4702.415 3048.785 4702.695 ;
        RECT 3049.215 4702.415 3049.495 4702.695 ;
        RECT 3049.925 4702.415 3050.205 4702.695 ;
        RECT 3050.635 4702.415 3050.915 4702.695 ;
        RECT 3051.345 4702.415 3051.625 4702.695 ;
        RECT 3052.055 4702.415 3052.335 4702.695 ;
        RECT 3052.765 4702.415 3053.045 4702.695 ;
        RECT 3053.475 4702.415 3053.755 4702.695 ;
        RECT 3054.185 4702.415 3054.465 4702.695 ;
        RECT 3054.895 4702.415 3055.175 4702.695 ;
        RECT 3055.605 4702.415 3055.885 4702.695 ;
        RECT 3059.485 4702.415 3059.765 4702.695 ;
        RECT 3060.195 4702.415 3060.475 4702.695 ;
        RECT 3060.905 4702.415 3061.185 4702.695 ;
        RECT 3061.615 4702.415 3061.895 4702.695 ;
        RECT 3062.325 4702.415 3062.605 4702.695 ;
        RECT 3063.035 4702.415 3063.315 4702.695 ;
        RECT 3063.745 4702.415 3064.025 4702.695 ;
        RECT 3064.455 4702.415 3064.735 4702.695 ;
        RECT 3065.165 4702.415 3065.445 4702.695 ;
        RECT 3065.875 4702.415 3066.155 4702.695 ;
        RECT 3066.585 4702.415 3066.865 4702.695 ;
        RECT 3067.295 4702.415 3067.575 4702.695 ;
        RECT 3068.005 4702.415 3068.285 4702.695 ;
        RECT 1896.705 4701.705 1896.985 4701.985 ;
        RECT 1897.415 4701.705 1897.695 4701.985 ;
        RECT 1898.125 4701.705 1898.405 4701.985 ;
        RECT 1898.835 4701.705 1899.115 4701.985 ;
        RECT 1899.545 4701.705 1899.825 4701.985 ;
        RECT 1909.145 4701.705 1909.425 4701.985 ;
        RECT 1909.855 4701.705 1910.135 4701.985 ;
        RECT 1910.565 4701.705 1910.845 4701.985 ;
        RECT 1911.275 4701.705 1911.555 4701.985 ;
        RECT 1911.985 4701.705 1912.265 4701.985 ;
        RECT 1912.695 4701.705 1912.975 4701.985 ;
        RECT 1913.405 4701.705 1913.685 4701.985 ;
        RECT 1914.115 4701.705 1914.395 4701.985 ;
        RECT 1914.825 4701.705 1915.105 4701.985 ;
        RECT 1915.535 4701.705 1915.815 4701.985 ;
        RECT 1916.245 4701.705 1916.525 4701.985 ;
        RECT 1916.955 4701.705 1917.235 4701.985 ;
        RECT 1917.665 4701.705 1917.945 4701.985 ;
        RECT 1918.375 4701.705 1918.655 4701.985 ;
        RECT 1920.995 4701.705 1921.275 4701.985 ;
        RECT 1921.705 4701.705 1921.985 4701.985 ;
        RECT 1922.415 4701.705 1922.695 4701.985 ;
        RECT 1926.675 4701.705 1926.955 4701.985 ;
        RECT 1927.385 4701.705 1927.665 4701.985 ;
        RECT 1928.095 4701.705 1928.375 4701.985 ;
        RECT 1928.805 4701.705 1929.085 4701.985 ;
        RECT 1929.515 4701.705 1929.795 4701.985 ;
        RECT 1930.225 4701.705 1930.505 4701.985 ;
        RECT 1934.525 4701.705 1934.805 4701.985 ;
        RECT 1935.235 4701.705 1935.515 4701.985 ;
        RECT 1935.945 4701.705 1936.225 4701.985 ;
        RECT 1936.655 4701.705 1936.935 4701.985 ;
        RECT 1937.365 4701.705 1937.645 4701.985 ;
        RECT 1938.075 4701.705 1938.355 4701.985 ;
        RECT 1938.785 4701.705 1939.065 4701.985 ;
        RECT 1939.495 4701.705 1939.775 4701.985 ;
        RECT 1940.205 4701.705 1940.485 4701.985 ;
        RECT 1940.915 4701.705 1941.195 4701.985 ;
        RECT 1941.625 4701.705 1941.905 4701.985 ;
        RECT 1942.335 4701.705 1942.615 4701.985 ;
        RECT 1943.045 4701.705 1943.325 4701.985 ;
        RECT 1943.755 4701.705 1944.035 4701.985 ;
        RECT 1946.375 4701.705 1946.655 4701.985 ;
        RECT 1947.085 4701.705 1947.365 4701.985 ;
        RECT 1947.795 4701.705 1948.075 4701.985 ;
        RECT 1948.505 4701.705 1948.785 4701.985 ;
        RECT 1949.215 4701.705 1949.495 4701.985 ;
        RECT 1949.925 4701.705 1950.205 4701.985 ;
        RECT 1950.635 4701.705 1950.915 4701.985 ;
        RECT 1951.345 4701.705 1951.625 4701.985 ;
        RECT 1952.055 4701.705 1952.335 4701.985 ;
        RECT 1952.765 4701.705 1953.045 4701.985 ;
        RECT 1953.475 4701.705 1953.755 4701.985 ;
        RECT 1954.185 4701.705 1954.465 4701.985 ;
        RECT 1954.895 4701.705 1955.175 4701.985 ;
        RECT 1955.605 4701.705 1955.885 4701.985 ;
        RECT 1959.485 4701.705 1959.765 4701.985 ;
        RECT 1960.195 4701.705 1960.475 4701.985 ;
        RECT 1960.905 4701.705 1961.185 4701.985 ;
        RECT 1961.615 4701.705 1961.895 4701.985 ;
        RECT 1962.325 4701.705 1962.605 4701.985 ;
        RECT 1963.035 4701.705 1963.315 4701.985 ;
        RECT 1963.745 4701.705 1964.025 4701.985 ;
        RECT 1964.455 4701.705 1964.735 4701.985 ;
        RECT 1965.165 4701.705 1965.445 4701.985 ;
        RECT 1965.875 4701.705 1966.155 4701.985 ;
        RECT 1966.585 4701.705 1966.865 4701.985 ;
        RECT 1967.295 4701.705 1967.575 4701.985 ;
        RECT 1968.005 4701.705 1968.285 4701.985 ;
        RECT 2996.705 4701.705 2996.985 4701.985 ;
        RECT 2997.415 4701.705 2997.695 4701.985 ;
        RECT 2998.125 4701.705 2998.405 4701.985 ;
        RECT 2998.835 4701.705 2999.115 4701.985 ;
        RECT 2999.545 4701.705 2999.825 4701.985 ;
        RECT 3000.255 4701.705 3000.535 4701.985 ;
        RECT 3000.965 4701.705 3001.245 4701.985 ;
        RECT 3001.675 4701.705 3001.955 4701.985 ;
        RECT 3002.385 4701.705 3002.665 4701.985 ;
        RECT 3003.095 4701.705 3003.375 4701.985 ;
        RECT 3003.805 4701.705 3004.085 4701.985 ;
        RECT 3004.515 4701.705 3004.795 4701.985 ;
        RECT 3005.225 4701.705 3005.505 4701.985 ;
        RECT 3009.145 4701.705 3009.425 4701.985 ;
        RECT 3009.855 4701.705 3010.135 4701.985 ;
        RECT 3010.565 4701.705 3010.845 4701.985 ;
        RECT 3011.275 4701.705 3011.555 4701.985 ;
        RECT 3011.985 4701.705 3012.265 4701.985 ;
        RECT 3012.695 4701.705 3012.975 4701.985 ;
        RECT 3013.405 4701.705 3013.685 4701.985 ;
        RECT 3014.115 4701.705 3014.395 4701.985 ;
        RECT 3014.825 4701.705 3015.105 4701.985 ;
        RECT 3015.535 4701.705 3015.815 4701.985 ;
        RECT 3016.245 4701.705 3016.525 4701.985 ;
        RECT 3016.955 4701.705 3017.235 4701.985 ;
        RECT 3017.665 4701.705 3017.945 4701.985 ;
        RECT 3018.375 4701.705 3018.655 4701.985 ;
        RECT 3025.255 4701.705 3025.535 4701.985 ;
        RECT 3025.965 4701.705 3026.245 4701.985 ;
        RECT 3026.675 4701.705 3026.955 4701.985 ;
        RECT 3027.385 4701.705 3027.665 4701.985 ;
        RECT 3028.095 4701.705 3028.375 4701.985 ;
        RECT 3028.805 4701.705 3029.085 4701.985 ;
        RECT 3029.515 4701.705 3029.795 4701.985 ;
        RECT 3030.225 4701.705 3030.505 4701.985 ;
        RECT 3034.525 4701.705 3034.805 4701.985 ;
        RECT 3035.235 4701.705 3035.515 4701.985 ;
        RECT 3035.945 4701.705 3036.225 4701.985 ;
        RECT 3036.655 4701.705 3036.935 4701.985 ;
        RECT 3037.365 4701.705 3037.645 4701.985 ;
        RECT 3038.075 4701.705 3038.355 4701.985 ;
        RECT 3038.785 4701.705 3039.065 4701.985 ;
        RECT 3039.495 4701.705 3039.775 4701.985 ;
        RECT 3040.205 4701.705 3040.485 4701.985 ;
        RECT 3040.915 4701.705 3041.195 4701.985 ;
        RECT 3041.625 4701.705 3041.905 4701.985 ;
        RECT 3042.335 4701.705 3042.615 4701.985 ;
        RECT 3046.375 4701.705 3046.655 4701.985 ;
        RECT 3047.085 4701.705 3047.365 4701.985 ;
        RECT 3047.795 4701.705 3048.075 4701.985 ;
        RECT 3048.505 4701.705 3048.785 4701.985 ;
        RECT 3049.215 4701.705 3049.495 4701.985 ;
        RECT 3049.925 4701.705 3050.205 4701.985 ;
        RECT 3050.635 4701.705 3050.915 4701.985 ;
        RECT 3051.345 4701.705 3051.625 4701.985 ;
        RECT 3052.055 4701.705 3052.335 4701.985 ;
        RECT 3052.765 4701.705 3053.045 4701.985 ;
        RECT 3053.475 4701.705 3053.755 4701.985 ;
        RECT 3054.185 4701.705 3054.465 4701.985 ;
        RECT 3054.895 4701.705 3055.175 4701.985 ;
        RECT 3055.605 4701.705 3055.885 4701.985 ;
        RECT 3059.485 4701.705 3059.765 4701.985 ;
        RECT 3060.195 4701.705 3060.475 4701.985 ;
        RECT 3060.905 4701.705 3061.185 4701.985 ;
        RECT 3061.615 4701.705 3061.895 4701.985 ;
        RECT 3062.325 4701.705 3062.605 4701.985 ;
        RECT 3063.035 4701.705 3063.315 4701.985 ;
        RECT 3063.745 4701.705 3064.025 4701.985 ;
        RECT 3064.455 4701.705 3064.735 4701.985 ;
        RECT 3065.165 4701.705 3065.445 4701.985 ;
        RECT 3065.875 4701.705 3066.155 4701.985 ;
        RECT 3066.585 4701.705 3066.865 4701.985 ;
        RECT 3067.295 4701.705 3067.575 4701.985 ;
        RECT 3068.005 4701.705 3068.285 4701.985 ;
        RECT 1896.705 4700.995 1896.985 4701.275 ;
        RECT 1897.415 4700.995 1897.695 4701.275 ;
        RECT 1898.125 4700.995 1898.405 4701.275 ;
        RECT 1898.835 4700.995 1899.115 4701.275 ;
        RECT 1899.545 4700.995 1899.825 4701.275 ;
        RECT 1909.145 4700.995 1909.425 4701.275 ;
        RECT 1909.855 4700.995 1910.135 4701.275 ;
        RECT 1910.565 4700.995 1910.845 4701.275 ;
        RECT 1911.275 4700.995 1911.555 4701.275 ;
        RECT 1911.985 4700.995 1912.265 4701.275 ;
        RECT 1912.695 4700.995 1912.975 4701.275 ;
        RECT 1913.405 4700.995 1913.685 4701.275 ;
        RECT 1914.115 4700.995 1914.395 4701.275 ;
        RECT 1914.825 4700.995 1915.105 4701.275 ;
        RECT 1915.535 4700.995 1915.815 4701.275 ;
        RECT 1916.245 4700.995 1916.525 4701.275 ;
        RECT 1916.955 4700.995 1917.235 4701.275 ;
        RECT 1917.665 4700.995 1917.945 4701.275 ;
        RECT 1918.375 4700.995 1918.655 4701.275 ;
        RECT 1920.995 4700.995 1921.275 4701.275 ;
        RECT 1921.705 4700.995 1921.985 4701.275 ;
        RECT 1922.415 4700.995 1922.695 4701.275 ;
        RECT 1926.675 4700.995 1926.955 4701.275 ;
        RECT 1927.385 4700.995 1927.665 4701.275 ;
        RECT 1928.095 4700.995 1928.375 4701.275 ;
        RECT 1928.805 4700.995 1929.085 4701.275 ;
        RECT 1929.515 4700.995 1929.795 4701.275 ;
        RECT 1930.225 4700.995 1930.505 4701.275 ;
        RECT 1934.525 4700.995 1934.805 4701.275 ;
        RECT 1935.235 4700.995 1935.515 4701.275 ;
        RECT 1935.945 4700.995 1936.225 4701.275 ;
        RECT 1936.655 4700.995 1936.935 4701.275 ;
        RECT 1937.365 4700.995 1937.645 4701.275 ;
        RECT 1938.075 4700.995 1938.355 4701.275 ;
        RECT 1938.785 4700.995 1939.065 4701.275 ;
        RECT 1939.495 4700.995 1939.775 4701.275 ;
        RECT 1940.205 4700.995 1940.485 4701.275 ;
        RECT 1940.915 4700.995 1941.195 4701.275 ;
        RECT 1941.625 4700.995 1941.905 4701.275 ;
        RECT 1942.335 4700.995 1942.615 4701.275 ;
        RECT 1943.045 4700.995 1943.325 4701.275 ;
        RECT 1943.755 4700.995 1944.035 4701.275 ;
        RECT 1946.375 4700.995 1946.655 4701.275 ;
        RECT 1947.085 4700.995 1947.365 4701.275 ;
        RECT 1947.795 4700.995 1948.075 4701.275 ;
        RECT 1948.505 4700.995 1948.785 4701.275 ;
        RECT 1949.215 4700.995 1949.495 4701.275 ;
        RECT 1949.925 4700.995 1950.205 4701.275 ;
        RECT 1950.635 4700.995 1950.915 4701.275 ;
        RECT 1951.345 4700.995 1951.625 4701.275 ;
        RECT 1952.055 4700.995 1952.335 4701.275 ;
        RECT 1952.765 4700.995 1953.045 4701.275 ;
        RECT 1953.475 4700.995 1953.755 4701.275 ;
        RECT 1954.185 4700.995 1954.465 4701.275 ;
        RECT 1954.895 4700.995 1955.175 4701.275 ;
        RECT 1955.605 4700.995 1955.885 4701.275 ;
        RECT 1959.485 4700.995 1959.765 4701.275 ;
        RECT 1960.195 4700.995 1960.475 4701.275 ;
        RECT 1960.905 4700.995 1961.185 4701.275 ;
        RECT 1961.615 4700.995 1961.895 4701.275 ;
        RECT 1962.325 4700.995 1962.605 4701.275 ;
        RECT 1963.035 4700.995 1963.315 4701.275 ;
        RECT 1963.745 4700.995 1964.025 4701.275 ;
        RECT 1964.455 4700.995 1964.735 4701.275 ;
        RECT 1965.165 4700.995 1965.445 4701.275 ;
        RECT 1965.875 4700.995 1966.155 4701.275 ;
        RECT 1966.585 4700.995 1966.865 4701.275 ;
        RECT 1967.295 4700.995 1967.575 4701.275 ;
        RECT 1968.005 4700.995 1968.285 4701.275 ;
        RECT 2996.705 4700.995 2996.985 4701.275 ;
        RECT 2997.415 4700.995 2997.695 4701.275 ;
        RECT 2998.125 4700.995 2998.405 4701.275 ;
        RECT 2998.835 4700.995 2999.115 4701.275 ;
        RECT 2999.545 4700.995 2999.825 4701.275 ;
        RECT 3000.255 4700.995 3000.535 4701.275 ;
        RECT 3000.965 4700.995 3001.245 4701.275 ;
        RECT 3001.675 4700.995 3001.955 4701.275 ;
        RECT 3002.385 4700.995 3002.665 4701.275 ;
        RECT 3003.095 4700.995 3003.375 4701.275 ;
        RECT 3003.805 4700.995 3004.085 4701.275 ;
        RECT 3004.515 4700.995 3004.795 4701.275 ;
        RECT 3005.225 4700.995 3005.505 4701.275 ;
        RECT 3009.145 4700.995 3009.425 4701.275 ;
        RECT 3009.855 4700.995 3010.135 4701.275 ;
        RECT 3010.565 4700.995 3010.845 4701.275 ;
        RECT 3011.275 4700.995 3011.555 4701.275 ;
        RECT 3011.985 4700.995 3012.265 4701.275 ;
        RECT 3012.695 4700.995 3012.975 4701.275 ;
        RECT 3013.405 4700.995 3013.685 4701.275 ;
        RECT 3014.115 4700.995 3014.395 4701.275 ;
        RECT 3014.825 4700.995 3015.105 4701.275 ;
        RECT 3015.535 4700.995 3015.815 4701.275 ;
        RECT 3016.245 4700.995 3016.525 4701.275 ;
        RECT 3016.955 4700.995 3017.235 4701.275 ;
        RECT 3017.665 4700.995 3017.945 4701.275 ;
        RECT 3018.375 4700.995 3018.655 4701.275 ;
        RECT 3025.255 4700.995 3025.535 4701.275 ;
        RECT 3025.965 4700.995 3026.245 4701.275 ;
        RECT 3026.675 4700.995 3026.955 4701.275 ;
        RECT 3027.385 4700.995 3027.665 4701.275 ;
        RECT 3028.095 4700.995 3028.375 4701.275 ;
        RECT 3028.805 4700.995 3029.085 4701.275 ;
        RECT 3029.515 4700.995 3029.795 4701.275 ;
        RECT 3030.225 4700.995 3030.505 4701.275 ;
        RECT 3034.525 4700.995 3034.805 4701.275 ;
        RECT 3035.235 4700.995 3035.515 4701.275 ;
        RECT 3035.945 4700.995 3036.225 4701.275 ;
        RECT 3036.655 4700.995 3036.935 4701.275 ;
        RECT 3037.365 4700.995 3037.645 4701.275 ;
        RECT 3038.075 4700.995 3038.355 4701.275 ;
        RECT 3038.785 4700.995 3039.065 4701.275 ;
        RECT 3039.495 4700.995 3039.775 4701.275 ;
        RECT 3040.205 4700.995 3040.485 4701.275 ;
        RECT 3040.915 4700.995 3041.195 4701.275 ;
        RECT 3041.625 4700.995 3041.905 4701.275 ;
        RECT 3042.335 4700.995 3042.615 4701.275 ;
        RECT 3046.375 4700.995 3046.655 4701.275 ;
        RECT 3047.085 4700.995 3047.365 4701.275 ;
        RECT 3047.795 4700.995 3048.075 4701.275 ;
        RECT 3048.505 4700.995 3048.785 4701.275 ;
        RECT 3049.215 4700.995 3049.495 4701.275 ;
        RECT 3049.925 4700.995 3050.205 4701.275 ;
        RECT 3050.635 4700.995 3050.915 4701.275 ;
        RECT 3051.345 4700.995 3051.625 4701.275 ;
        RECT 3052.055 4700.995 3052.335 4701.275 ;
        RECT 3052.765 4700.995 3053.045 4701.275 ;
        RECT 3053.475 4700.995 3053.755 4701.275 ;
        RECT 3054.185 4700.995 3054.465 4701.275 ;
        RECT 3054.895 4700.995 3055.175 4701.275 ;
        RECT 3055.605 4700.995 3055.885 4701.275 ;
        RECT 3059.485 4700.995 3059.765 4701.275 ;
        RECT 3060.195 4700.995 3060.475 4701.275 ;
        RECT 3060.905 4700.995 3061.185 4701.275 ;
        RECT 3061.615 4700.995 3061.895 4701.275 ;
        RECT 3062.325 4700.995 3062.605 4701.275 ;
        RECT 3063.035 4700.995 3063.315 4701.275 ;
        RECT 3063.745 4700.995 3064.025 4701.275 ;
        RECT 3064.455 4700.995 3064.735 4701.275 ;
        RECT 3065.165 4700.995 3065.445 4701.275 ;
        RECT 3065.875 4700.995 3066.155 4701.275 ;
        RECT 3066.585 4700.995 3066.865 4701.275 ;
        RECT 3067.295 4700.995 3067.575 4701.275 ;
        RECT 3068.005 4700.995 3068.285 4701.275 ;
        RECT 1896.705 4700.285 1896.985 4700.565 ;
        RECT 1897.415 4700.285 1897.695 4700.565 ;
        RECT 1898.125 4700.285 1898.405 4700.565 ;
        RECT 1898.835 4700.285 1899.115 4700.565 ;
        RECT 1899.545 4700.285 1899.825 4700.565 ;
        RECT 1909.145 4700.285 1909.425 4700.565 ;
        RECT 1909.855 4700.285 1910.135 4700.565 ;
        RECT 1910.565 4700.285 1910.845 4700.565 ;
        RECT 1911.275 4700.285 1911.555 4700.565 ;
        RECT 1911.985 4700.285 1912.265 4700.565 ;
        RECT 1912.695 4700.285 1912.975 4700.565 ;
        RECT 1913.405 4700.285 1913.685 4700.565 ;
        RECT 1914.115 4700.285 1914.395 4700.565 ;
        RECT 1914.825 4700.285 1915.105 4700.565 ;
        RECT 1915.535 4700.285 1915.815 4700.565 ;
        RECT 1916.245 4700.285 1916.525 4700.565 ;
        RECT 1916.955 4700.285 1917.235 4700.565 ;
        RECT 1917.665 4700.285 1917.945 4700.565 ;
        RECT 1918.375 4700.285 1918.655 4700.565 ;
        RECT 1920.995 4700.285 1921.275 4700.565 ;
        RECT 1921.705 4700.285 1921.985 4700.565 ;
        RECT 1922.415 4700.285 1922.695 4700.565 ;
        RECT 1926.675 4700.285 1926.955 4700.565 ;
        RECT 1927.385 4700.285 1927.665 4700.565 ;
        RECT 1928.095 4700.285 1928.375 4700.565 ;
        RECT 1928.805 4700.285 1929.085 4700.565 ;
        RECT 1929.515 4700.285 1929.795 4700.565 ;
        RECT 1930.225 4700.285 1930.505 4700.565 ;
        RECT 1934.525 4700.285 1934.805 4700.565 ;
        RECT 1935.235 4700.285 1935.515 4700.565 ;
        RECT 1935.945 4700.285 1936.225 4700.565 ;
        RECT 1936.655 4700.285 1936.935 4700.565 ;
        RECT 1937.365 4700.285 1937.645 4700.565 ;
        RECT 1938.075 4700.285 1938.355 4700.565 ;
        RECT 1938.785 4700.285 1939.065 4700.565 ;
        RECT 1939.495 4700.285 1939.775 4700.565 ;
        RECT 1940.205 4700.285 1940.485 4700.565 ;
        RECT 1940.915 4700.285 1941.195 4700.565 ;
        RECT 1941.625 4700.285 1941.905 4700.565 ;
        RECT 1942.335 4700.285 1942.615 4700.565 ;
        RECT 1943.045 4700.285 1943.325 4700.565 ;
        RECT 1943.755 4700.285 1944.035 4700.565 ;
        RECT 1946.375 4700.285 1946.655 4700.565 ;
        RECT 1947.085 4700.285 1947.365 4700.565 ;
        RECT 1947.795 4700.285 1948.075 4700.565 ;
        RECT 1948.505 4700.285 1948.785 4700.565 ;
        RECT 1949.215 4700.285 1949.495 4700.565 ;
        RECT 1949.925 4700.285 1950.205 4700.565 ;
        RECT 1950.635 4700.285 1950.915 4700.565 ;
        RECT 1951.345 4700.285 1951.625 4700.565 ;
        RECT 1952.055 4700.285 1952.335 4700.565 ;
        RECT 1952.765 4700.285 1953.045 4700.565 ;
        RECT 1953.475 4700.285 1953.755 4700.565 ;
        RECT 1954.185 4700.285 1954.465 4700.565 ;
        RECT 1954.895 4700.285 1955.175 4700.565 ;
        RECT 1955.605 4700.285 1955.885 4700.565 ;
        RECT 1959.485 4700.285 1959.765 4700.565 ;
        RECT 1960.195 4700.285 1960.475 4700.565 ;
        RECT 1960.905 4700.285 1961.185 4700.565 ;
        RECT 1961.615 4700.285 1961.895 4700.565 ;
        RECT 1962.325 4700.285 1962.605 4700.565 ;
        RECT 1963.035 4700.285 1963.315 4700.565 ;
        RECT 1963.745 4700.285 1964.025 4700.565 ;
        RECT 1964.455 4700.285 1964.735 4700.565 ;
        RECT 1965.165 4700.285 1965.445 4700.565 ;
        RECT 1965.875 4700.285 1966.155 4700.565 ;
        RECT 1966.585 4700.285 1966.865 4700.565 ;
        RECT 1967.295 4700.285 1967.575 4700.565 ;
        RECT 1968.005 4700.285 1968.285 4700.565 ;
        RECT 2996.705 4700.285 2996.985 4700.565 ;
        RECT 2997.415 4700.285 2997.695 4700.565 ;
        RECT 2998.125 4700.285 2998.405 4700.565 ;
        RECT 2998.835 4700.285 2999.115 4700.565 ;
        RECT 2999.545 4700.285 2999.825 4700.565 ;
        RECT 3000.255 4700.285 3000.535 4700.565 ;
        RECT 3000.965 4700.285 3001.245 4700.565 ;
        RECT 3001.675 4700.285 3001.955 4700.565 ;
        RECT 3002.385 4700.285 3002.665 4700.565 ;
        RECT 3003.095 4700.285 3003.375 4700.565 ;
        RECT 3003.805 4700.285 3004.085 4700.565 ;
        RECT 3004.515 4700.285 3004.795 4700.565 ;
        RECT 3005.225 4700.285 3005.505 4700.565 ;
        RECT 3009.145 4700.285 3009.425 4700.565 ;
        RECT 3009.855 4700.285 3010.135 4700.565 ;
        RECT 3010.565 4700.285 3010.845 4700.565 ;
        RECT 3011.275 4700.285 3011.555 4700.565 ;
        RECT 3011.985 4700.285 3012.265 4700.565 ;
        RECT 3012.695 4700.285 3012.975 4700.565 ;
        RECT 3013.405 4700.285 3013.685 4700.565 ;
        RECT 3014.115 4700.285 3014.395 4700.565 ;
        RECT 3014.825 4700.285 3015.105 4700.565 ;
        RECT 3015.535 4700.285 3015.815 4700.565 ;
        RECT 3016.245 4700.285 3016.525 4700.565 ;
        RECT 3016.955 4700.285 3017.235 4700.565 ;
        RECT 3017.665 4700.285 3017.945 4700.565 ;
        RECT 3018.375 4700.285 3018.655 4700.565 ;
        RECT 3025.255 4700.285 3025.535 4700.565 ;
        RECT 3025.965 4700.285 3026.245 4700.565 ;
        RECT 3026.675 4700.285 3026.955 4700.565 ;
        RECT 3027.385 4700.285 3027.665 4700.565 ;
        RECT 3028.095 4700.285 3028.375 4700.565 ;
        RECT 3028.805 4700.285 3029.085 4700.565 ;
        RECT 3029.515 4700.285 3029.795 4700.565 ;
        RECT 3030.225 4700.285 3030.505 4700.565 ;
        RECT 3034.525 4700.285 3034.805 4700.565 ;
        RECT 3035.235 4700.285 3035.515 4700.565 ;
        RECT 3035.945 4700.285 3036.225 4700.565 ;
        RECT 3036.655 4700.285 3036.935 4700.565 ;
        RECT 3037.365 4700.285 3037.645 4700.565 ;
        RECT 3038.075 4700.285 3038.355 4700.565 ;
        RECT 3038.785 4700.285 3039.065 4700.565 ;
        RECT 3039.495 4700.285 3039.775 4700.565 ;
        RECT 3040.205 4700.285 3040.485 4700.565 ;
        RECT 3040.915 4700.285 3041.195 4700.565 ;
        RECT 3041.625 4700.285 3041.905 4700.565 ;
        RECT 3042.335 4700.285 3042.615 4700.565 ;
        RECT 3046.375 4700.285 3046.655 4700.565 ;
        RECT 3047.085 4700.285 3047.365 4700.565 ;
        RECT 3047.795 4700.285 3048.075 4700.565 ;
        RECT 3048.505 4700.285 3048.785 4700.565 ;
        RECT 3049.215 4700.285 3049.495 4700.565 ;
        RECT 3049.925 4700.285 3050.205 4700.565 ;
        RECT 3050.635 4700.285 3050.915 4700.565 ;
        RECT 3051.345 4700.285 3051.625 4700.565 ;
        RECT 3052.055 4700.285 3052.335 4700.565 ;
        RECT 3052.765 4700.285 3053.045 4700.565 ;
        RECT 3053.475 4700.285 3053.755 4700.565 ;
        RECT 3054.185 4700.285 3054.465 4700.565 ;
        RECT 3054.895 4700.285 3055.175 4700.565 ;
        RECT 3055.605 4700.285 3055.885 4700.565 ;
        RECT 3059.485 4700.285 3059.765 4700.565 ;
        RECT 3060.195 4700.285 3060.475 4700.565 ;
        RECT 3060.905 4700.285 3061.185 4700.565 ;
        RECT 3061.615 4700.285 3061.895 4700.565 ;
        RECT 3062.325 4700.285 3062.605 4700.565 ;
        RECT 3063.035 4700.285 3063.315 4700.565 ;
        RECT 3063.745 4700.285 3064.025 4700.565 ;
        RECT 3064.455 4700.285 3064.735 4700.565 ;
        RECT 3065.165 4700.285 3065.445 4700.565 ;
        RECT 3065.875 4700.285 3066.155 4700.565 ;
        RECT 3066.585 4700.285 3066.865 4700.565 ;
        RECT 3067.295 4700.285 3067.575 4700.565 ;
        RECT 3068.005 4700.285 3068.285 4700.565 ;
        RECT 1896.705 4699.575 1896.985 4699.855 ;
        RECT 1897.415 4699.575 1897.695 4699.855 ;
        RECT 1898.125 4699.575 1898.405 4699.855 ;
        RECT 1898.835 4699.575 1899.115 4699.855 ;
        RECT 1899.545 4699.575 1899.825 4699.855 ;
        RECT 1909.145 4699.575 1909.425 4699.855 ;
        RECT 1909.855 4699.575 1910.135 4699.855 ;
        RECT 1910.565 4699.575 1910.845 4699.855 ;
        RECT 1911.275 4699.575 1911.555 4699.855 ;
        RECT 1911.985 4699.575 1912.265 4699.855 ;
        RECT 1912.695 4699.575 1912.975 4699.855 ;
        RECT 1913.405 4699.575 1913.685 4699.855 ;
        RECT 1914.115 4699.575 1914.395 4699.855 ;
        RECT 1914.825 4699.575 1915.105 4699.855 ;
        RECT 1915.535 4699.575 1915.815 4699.855 ;
        RECT 1916.245 4699.575 1916.525 4699.855 ;
        RECT 1916.955 4699.575 1917.235 4699.855 ;
        RECT 1917.665 4699.575 1917.945 4699.855 ;
        RECT 1918.375 4699.575 1918.655 4699.855 ;
        RECT 1920.995 4699.575 1921.275 4699.855 ;
        RECT 1921.705 4699.575 1921.985 4699.855 ;
        RECT 1922.415 4699.575 1922.695 4699.855 ;
        RECT 1926.675 4699.575 1926.955 4699.855 ;
        RECT 1927.385 4699.575 1927.665 4699.855 ;
        RECT 1928.095 4699.575 1928.375 4699.855 ;
        RECT 1928.805 4699.575 1929.085 4699.855 ;
        RECT 1929.515 4699.575 1929.795 4699.855 ;
        RECT 1930.225 4699.575 1930.505 4699.855 ;
        RECT 1934.525 4699.575 1934.805 4699.855 ;
        RECT 1935.235 4699.575 1935.515 4699.855 ;
        RECT 1935.945 4699.575 1936.225 4699.855 ;
        RECT 1936.655 4699.575 1936.935 4699.855 ;
        RECT 1937.365 4699.575 1937.645 4699.855 ;
        RECT 1938.075 4699.575 1938.355 4699.855 ;
        RECT 1938.785 4699.575 1939.065 4699.855 ;
        RECT 1939.495 4699.575 1939.775 4699.855 ;
        RECT 1940.205 4699.575 1940.485 4699.855 ;
        RECT 1940.915 4699.575 1941.195 4699.855 ;
        RECT 1941.625 4699.575 1941.905 4699.855 ;
        RECT 1942.335 4699.575 1942.615 4699.855 ;
        RECT 1943.045 4699.575 1943.325 4699.855 ;
        RECT 1943.755 4699.575 1944.035 4699.855 ;
        RECT 1946.375 4699.575 1946.655 4699.855 ;
        RECT 1947.085 4699.575 1947.365 4699.855 ;
        RECT 1947.795 4699.575 1948.075 4699.855 ;
        RECT 1948.505 4699.575 1948.785 4699.855 ;
        RECT 1949.215 4699.575 1949.495 4699.855 ;
        RECT 1949.925 4699.575 1950.205 4699.855 ;
        RECT 1950.635 4699.575 1950.915 4699.855 ;
        RECT 1951.345 4699.575 1951.625 4699.855 ;
        RECT 1952.055 4699.575 1952.335 4699.855 ;
        RECT 1952.765 4699.575 1953.045 4699.855 ;
        RECT 1953.475 4699.575 1953.755 4699.855 ;
        RECT 1954.185 4699.575 1954.465 4699.855 ;
        RECT 1954.895 4699.575 1955.175 4699.855 ;
        RECT 1955.605 4699.575 1955.885 4699.855 ;
        RECT 1959.485 4699.575 1959.765 4699.855 ;
        RECT 1960.195 4699.575 1960.475 4699.855 ;
        RECT 1960.905 4699.575 1961.185 4699.855 ;
        RECT 1961.615 4699.575 1961.895 4699.855 ;
        RECT 1962.325 4699.575 1962.605 4699.855 ;
        RECT 1963.035 4699.575 1963.315 4699.855 ;
        RECT 1963.745 4699.575 1964.025 4699.855 ;
        RECT 1964.455 4699.575 1964.735 4699.855 ;
        RECT 1965.165 4699.575 1965.445 4699.855 ;
        RECT 1965.875 4699.575 1966.155 4699.855 ;
        RECT 1966.585 4699.575 1966.865 4699.855 ;
        RECT 1967.295 4699.575 1967.575 4699.855 ;
        RECT 1968.005 4699.575 1968.285 4699.855 ;
        RECT 2996.705 4699.575 2996.985 4699.855 ;
        RECT 2997.415 4699.575 2997.695 4699.855 ;
        RECT 2998.125 4699.575 2998.405 4699.855 ;
        RECT 2998.835 4699.575 2999.115 4699.855 ;
        RECT 2999.545 4699.575 2999.825 4699.855 ;
        RECT 3000.255 4699.575 3000.535 4699.855 ;
        RECT 3000.965 4699.575 3001.245 4699.855 ;
        RECT 3001.675 4699.575 3001.955 4699.855 ;
        RECT 3002.385 4699.575 3002.665 4699.855 ;
        RECT 3003.095 4699.575 3003.375 4699.855 ;
        RECT 3003.805 4699.575 3004.085 4699.855 ;
        RECT 3004.515 4699.575 3004.795 4699.855 ;
        RECT 3005.225 4699.575 3005.505 4699.855 ;
        RECT 3009.145 4699.575 3009.425 4699.855 ;
        RECT 3009.855 4699.575 3010.135 4699.855 ;
        RECT 3010.565 4699.575 3010.845 4699.855 ;
        RECT 3011.275 4699.575 3011.555 4699.855 ;
        RECT 3011.985 4699.575 3012.265 4699.855 ;
        RECT 3012.695 4699.575 3012.975 4699.855 ;
        RECT 3013.405 4699.575 3013.685 4699.855 ;
        RECT 3014.115 4699.575 3014.395 4699.855 ;
        RECT 3014.825 4699.575 3015.105 4699.855 ;
        RECT 3015.535 4699.575 3015.815 4699.855 ;
        RECT 3016.245 4699.575 3016.525 4699.855 ;
        RECT 3016.955 4699.575 3017.235 4699.855 ;
        RECT 3017.665 4699.575 3017.945 4699.855 ;
        RECT 3018.375 4699.575 3018.655 4699.855 ;
        RECT 3025.255 4699.575 3025.535 4699.855 ;
        RECT 3025.965 4699.575 3026.245 4699.855 ;
        RECT 3026.675 4699.575 3026.955 4699.855 ;
        RECT 3027.385 4699.575 3027.665 4699.855 ;
        RECT 3028.095 4699.575 3028.375 4699.855 ;
        RECT 3028.805 4699.575 3029.085 4699.855 ;
        RECT 3029.515 4699.575 3029.795 4699.855 ;
        RECT 3030.225 4699.575 3030.505 4699.855 ;
        RECT 3034.525 4699.575 3034.805 4699.855 ;
        RECT 3035.235 4699.575 3035.515 4699.855 ;
        RECT 3035.945 4699.575 3036.225 4699.855 ;
        RECT 3036.655 4699.575 3036.935 4699.855 ;
        RECT 3037.365 4699.575 3037.645 4699.855 ;
        RECT 3038.075 4699.575 3038.355 4699.855 ;
        RECT 3038.785 4699.575 3039.065 4699.855 ;
        RECT 3039.495 4699.575 3039.775 4699.855 ;
        RECT 3040.205 4699.575 3040.485 4699.855 ;
        RECT 3040.915 4699.575 3041.195 4699.855 ;
        RECT 3041.625 4699.575 3041.905 4699.855 ;
        RECT 3042.335 4699.575 3042.615 4699.855 ;
        RECT 3046.375 4699.575 3046.655 4699.855 ;
        RECT 3047.085 4699.575 3047.365 4699.855 ;
        RECT 3047.795 4699.575 3048.075 4699.855 ;
        RECT 3048.505 4699.575 3048.785 4699.855 ;
        RECT 3049.215 4699.575 3049.495 4699.855 ;
        RECT 3049.925 4699.575 3050.205 4699.855 ;
        RECT 3050.635 4699.575 3050.915 4699.855 ;
        RECT 3051.345 4699.575 3051.625 4699.855 ;
        RECT 3052.055 4699.575 3052.335 4699.855 ;
        RECT 3052.765 4699.575 3053.045 4699.855 ;
        RECT 3053.475 4699.575 3053.755 4699.855 ;
        RECT 3054.185 4699.575 3054.465 4699.855 ;
        RECT 3054.895 4699.575 3055.175 4699.855 ;
        RECT 3055.605 4699.575 3055.885 4699.855 ;
        RECT 3059.485 4699.575 3059.765 4699.855 ;
        RECT 3060.195 4699.575 3060.475 4699.855 ;
        RECT 3060.905 4699.575 3061.185 4699.855 ;
        RECT 3061.615 4699.575 3061.895 4699.855 ;
        RECT 3062.325 4699.575 3062.605 4699.855 ;
        RECT 3063.035 4699.575 3063.315 4699.855 ;
        RECT 3063.745 4699.575 3064.025 4699.855 ;
        RECT 3064.455 4699.575 3064.735 4699.855 ;
        RECT 3065.165 4699.575 3065.445 4699.855 ;
        RECT 3065.875 4699.575 3066.155 4699.855 ;
        RECT 3066.585 4699.575 3066.865 4699.855 ;
        RECT 3067.295 4699.575 3067.575 4699.855 ;
        RECT 3068.005 4699.575 3068.285 4699.855 ;
        RECT 1896.705 4698.865 1896.985 4699.145 ;
        RECT 1897.415 4698.865 1897.695 4699.145 ;
        RECT 1898.125 4698.865 1898.405 4699.145 ;
        RECT 1898.835 4698.865 1899.115 4699.145 ;
        RECT 1899.545 4698.865 1899.825 4699.145 ;
        RECT 1909.145 4698.865 1909.425 4699.145 ;
        RECT 1909.855 4698.865 1910.135 4699.145 ;
        RECT 1910.565 4698.865 1910.845 4699.145 ;
        RECT 1911.275 4698.865 1911.555 4699.145 ;
        RECT 1911.985 4698.865 1912.265 4699.145 ;
        RECT 1912.695 4698.865 1912.975 4699.145 ;
        RECT 1913.405 4698.865 1913.685 4699.145 ;
        RECT 1914.115 4698.865 1914.395 4699.145 ;
        RECT 1914.825 4698.865 1915.105 4699.145 ;
        RECT 1915.535 4698.865 1915.815 4699.145 ;
        RECT 1916.245 4698.865 1916.525 4699.145 ;
        RECT 1916.955 4698.865 1917.235 4699.145 ;
        RECT 1917.665 4698.865 1917.945 4699.145 ;
        RECT 1918.375 4698.865 1918.655 4699.145 ;
        RECT 1920.995 4698.865 1921.275 4699.145 ;
        RECT 1921.705 4698.865 1921.985 4699.145 ;
        RECT 1922.415 4698.865 1922.695 4699.145 ;
        RECT 1926.675 4698.865 1926.955 4699.145 ;
        RECT 1927.385 4698.865 1927.665 4699.145 ;
        RECT 1928.095 4698.865 1928.375 4699.145 ;
        RECT 1928.805 4698.865 1929.085 4699.145 ;
        RECT 1929.515 4698.865 1929.795 4699.145 ;
        RECT 1930.225 4698.865 1930.505 4699.145 ;
        RECT 1934.525 4698.865 1934.805 4699.145 ;
        RECT 1935.235 4698.865 1935.515 4699.145 ;
        RECT 1935.945 4698.865 1936.225 4699.145 ;
        RECT 1936.655 4698.865 1936.935 4699.145 ;
        RECT 1937.365 4698.865 1937.645 4699.145 ;
        RECT 1938.075 4698.865 1938.355 4699.145 ;
        RECT 1938.785 4698.865 1939.065 4699.145 ;
        RECT 1939.495 4698.865 1939.775 4699.145 ;
        RECT 1940.205 4698.865 1940.485 4699.145 ;
        RECT 1940.915 4698.865 1941.195 4699.145 ;
        RECT 1941.625 4698.865 1941.905 4699.145 ;
        RECT 1942.335 4698.865 1942.615 4699.145 ;
        RECT 1943.045 4698.865 1943.325 4699.145 ;
        RECT 1943.755 4698.865 1944.035 4699.145 ;
        RECT 1946.375 4698.865 1946.655 4699.145 ;
        RECT 1947.085 4698.865 1947.365 4699.145 ;
        RECT 1947.795 4698.865 1948.075 4699.145 ;
        RECT 1948.505 4698.865 1948.785 4699.145 ;
        RECT 1949.215 4698.865 1949.495 4699.145 ;
        RECT 1949.925 4698.865 1950.205 4699.145 ;
        RECT 1950.635 4698.865 1950.915 4699.145 ;
        RECT 1951.345 4698.865 1951.625 4699.145 ;
        RECT 1952.055 4698.865 1952.335 4699.145 ;
        RECT 1952.765 4698.865 1953.045 4699.145 ;
        RECT 1953.475 4698.865 1953.755 4699.145 ;
        RECT 1954.185 4698.865 1954.465 4699.145 ;
        RECT 1954.895 4698.865 1955.175 4699.145 ;
        RECT 1955.605 4698.865 1955.885 4699.145 ;
        RECT 1959.485 4698.865 1959.765 4699.145 ;
        RECT 1960.195 4698.865 1960.475 4699.145 ;
        RECT 1960.905 4698.865 1961.185 4699.145 ;
        RECT 1961.615 4698.865 1961.895 4699.145 ;
        RECT 1962.325 4698.865 1962.605 4699.145 ;
        RECT 1963.035 4698.865 1963.315 4699.145 ;
        RECT 1963.745 4698.865 1964.025 4699.145 ;
        RECT 1964.455 4698.865 1964.735 4699.145 ;
        RECT 1965.165 4698.865 1965.445 4699.145 ;
        RECT 1965.875 4698.865 1966.155 4699.145 ;
        RECT 1966.585 4698.865 1966.865 4699.145 ;
        RECT 1967.295 4698.865 1967.575 4699.145 ;
        RECT 1968.005 4698.865 1968.285 4699.145 ;
        RECT 2996.705 4698.865 2996.985 4699.145 ;
        RECT 2997.415 4698.865 2997.695 4699.145 ;
        RECT 2998.125 4698.865 2998.405 4699.145 ;
        RECT 2998.835 4698.865 2999.115 4699.145 ;
        RECT 2999.545 4698.865 2999.825 4699.145 ;
        RECT 3000.255 4698.865 3000.535 4699.145 ;
        RECT 3000.965 4698.865 3001.245 4699.145 ;
        RECT 3001.675 4698.865 3001.955 4699.145 ;
        RECT 3002.385 4698.865 3002.665 4699.145 ;
        RECT 3003.095 4698.865 3003.375 4699.145 ;
        RECT 3003.805 4698.865 3004.085 4699.145 ;
        RECT 3004.515 4698.865 3004.795 4699.145 ;
        RECT 3005.225 4698.865 3005.505 4699.145 ;
        RECT 3009.145 4698.865 3009.425 4699.145 ;
        RECT 3009.855 4698.865 3010.135 4699.145 ;
        RECT 3010.565 4698.865 3010.845 4699.145 ;
        RECT 3011.275 4698.865 3011.555 4699.145 ;
        RECT 3011.985 4698.865 3012.265 4699.145 ;
        RECT 3012.695 4698.865 3012.975 4699.145 ;
        RECT 3013.405 4698.865 3013.685 4699.145 ;
        RECT 3014.115 4698.865 3014.395 4699.145 ;
        RECT 3014.825 4698.865 3015.105 4699.145 ;
        RECT 3015.535 4698.865 3015.815 4699.145 ;
        RECT 3016.245 4698.865 3016.525 4699.145 ;
        RECT 3016.955 4698.865 3017.235 4699.145 ;
        RECT 3017.665 4698.865 3017.945 4699.145 ;
        RECT 3018.375 4698.865 3018.655 4699.145 ;
        RECT 3025.255 4698.865 3025.535 4699.145 ;
        RECT 3025.965 4698.865 3026.245 4699.145 ;
        RECT 3026.675 4698.865 3026.955 4699.145 ;
        RECT 3027.385 4698.865 3027.665 4699.145 ;
        RECT 3028.095 4698.865 3028.375 4699.145 ;
        RECT 3028.805 4698.865 3029.085 4699.145 ;
        RECT 3029.515 4698.865 3029.795 4699.145 ;
        RECT 3030.225 4698.865 3030.505 4699.145 ;
        RECT 3034.525 4698.865 3034.805 4699.145 ;
        RECT 3035.235 4698.865 3035.515 4699.145 ;
        RECT 3035.945 4698.865 3036.225 4699.145 ;
        RECT 3036.655 4698.865 3036.935 4699.145 ;
        RECT 3037.365 4698.865 3037.645 4699.145 ;
        RECT 3038.075 4698.865 3038.355 4699.145 ;
        RECT 3038.785 4698.865 3039.065 4699.145 ;
        RECT 3039.495 4698.865 3039.775 4699.145 ;
        RECT 3040.205 4698.865 3040.485 4699.145 ;
        RECT 3040.915 4698.865 3041.195 4699.145 ;
        RECT 3041.625 4698.865 3041.905 4699.145 ;
        RECT 3042.335 4698.865 3042.615 4699.145 ;
        RECT 3046.375 4698.865 3046.655 4699.145 ;
        RECT 3047.085 4698.865 3047.365 4699.145 ;
        RECT 3047.795 4698.865 3048.075 4699.145 ;
        RECT 3048.505 4698.865 3048.785 4699.145 ;
        RECT 3049.215 4698.865 3049.495 4699.145 ;
        RECT 3049.925 4698.865 3050.205 4699.145 ;
        RECT 3050.635 4698.865 3050.915 4699.145 ;
        RECT 3051.345 4698.865 3051.625 4699.145 ;
        RECT 3052.055 4698.865 3052.335 4699.145 ;
        RECT 3052.765 4698.865 3053.045 4699.145 ;
        RECT 3053.475 4698.865 3053.755 4699.145 ;
        RECT 3054.185 4698.865 3054.465 4699.145 ;
        RECT 3054.895 4698.865 3055.175 4699.145 ;
        RECT 3055.605 4698.865 3055.885 4699.145 ;
        RECT 3059.485 4698.865 3059.765 4699.145 ;
        RECT 3060.195 4698.865 3060.475 4699.145 ;
        RECT 3060.905 4698.865 3061.185 4699.145 ;
        RECT 3061.615 4698.865 3061.895 4699.145 ;
        RECT 3062.325 4698.865 3062.605 4699.145 ;
        RECT 3063.035 4698.865 3063.315 4699.145 ;
        RECT 3063.745 4698.865 3064.025 4699.145 ;
        RECT 3064.455 4698.865 3064.735 4699.145 ;
        RECT 3065.165 4698.865 3065.445 4699.145 ;
        RECT 3065.875 4698.865 3066.155 4699.145 ;
        RECT 3066.585 4698.865 3066.865 4699.145 ;
        RECT 3067.295 4698.865 3067.575 4699.145 ;
        RECT 3068.005 4698.865 3068.285 4699.145 ;
        RECT 3276.715 379.895 3276.995 380.175 ;
        RECT 3277.425 379.895 3277.705 380.175 ;
        RECT 3278.135 379.895 3278.415 380.175 ;
        RECT 3278.845 379.895 3279.125 380.175 ;
        RECT 3279.555 379.895 3279.835 380.175 ;
        RECT 3280.265 379.895 3280.545 380.175 ;
        RECT 3280.975 379.895 3281.255 380.175 ;
        RECT 3281.685 379.895 3281.965 380.175 ;
        RECT 3289.115 379.895 3289.395 380.175 ;
        RECT 3289.825 379.895 3290.105 380.175 ;
        RECT 3290.535 379.895 3290.815 380.175 ;
        RECT 3291.245 379.895 3291.525 380.175 ;
        RECT 3291.955 379.895 3292.235 380.175 ;
        RECT 3292.665 379.895 3292.945 380.175 ;
        RECT 3293.375 379.895 3293.655 380.175 ;
        RECT 3294.085 379.895 3294.365 380.175 ;
        RECT 3294.795 379.895 3295.075 380.175 ;
        RECT 3295.505 379.895 3295.785 380.175 ;
        RECT 3296.215 379.895 3296.495 380.175 ;
        RECT 3296.925 379.895 3297.205 380.175 ;
        RECT 3297.635 379.895 3297.915 380.175 ;
        RECT 3298.345 379.895 3298.625 380.175 ;
        RECT 3300.965 379.895 3301.245 380.175 ;
        RECT 3301.675 379.895 3301.955 380.175 ;
        RECT 3302.385 379.895 3302.665 380.175 ;
        RECT 3303.095 379.895 3303.375 380.175 ;
        RECT 3303.805 379.895 3304.085 380.175 ;
        RECT 3304.515 379.895 3304.795 380.175 ;
        RECT 3305.225 379.895 3305.505 380.175 ;
        RECT 3305.935 379.895 3306.215 380.175 ;
        RECT 3306.645 379.895 3306.925 380.175 ;
        RECT 3307.355 379.895 3307.635 380.175 ;
        RECT 3308.065 379.895 3308.345 380.175 ;
        RECT 3308.775 379.895 3309.055 380.175 ;
        RECT 3309.485 379.895 3309.765 380.175 ;
        RECT 3310.195 379.895 3310.475 380.175 ;
        RECT 3314.495 379.895 3314.775 380.175 ;
        RECT 3315.205 379.895 3315.485 380.175 ;
        RECT 3315.915 379.895 3316.195 380.175 ;
        RECT 3316.625 379.895 3316.905 380.175 ;
        RECT 3317.335 379.895 3317.615 380.175 ;
        RECT 3318.045 379.895 3318.325 380.175 ;
        RECT 3318.755 379.895 3319.035 380.175 ;
        RECT 3319.465 379.895 3319.745 380.175 ;
        RECT 3320.175 379.895 3320.455 380.175 ;
        RECT 3320.885 379.895 3321.165 380.175 ;
        RECT 3321.595 379.895 3321.875 380.175 ;
        RECT 3322.305 379.895 3322.585 380.175 ;
        RECT 3323.015 379.895 3323.295 380.175 ;
        RECT 3323.725 379.895 3324.005 380.175 ;
        RECT 3326.345 379.895 3326.625 380.175 ;
        RECT 3327.055 379.895 3327.335 380.175 ;
        RECT 3327.765 379.895 3328.045 380.175 ;
        RECT 3328.475 379.895 3328.755 380.175 ;
        RECT 3329.185 379.895 3329.465 380.175 ;
        RECT 3329.895 379.895 3330.175 380.175 ;
        RECT 3330.605 379.895 3330.885 380.175 ;
        RECT 3331.315 379.895 3331.595 380.175 ;
        RECT 3332.025 379.895 3332.305 380.175 ;
        RECT 3332.735 379.895 3333.015 380.175 ;
        RECT 3333.445 379.895 3333.725 380.175 ;
        RECT 3334.155 379.895 3334.435 380.175 ;
        RECT 3334.865 379.895 3335.145 380.175 ;
        RECT 3335.575 379.895 3335.855 380.175 ;
        RECT 3339.495 379.895 3339.775 380.175 ;
        RECT 3340.205 379.895 3340.485 380.175 ;
        RECT 3344.465 379.895 3344.745 380.175 ;
        RECT 3345.175 379.895 3345.455 380.175 ;
        RECT 3345.885 379.895 3346.165 380.175 ;
        RECT 3346.595 379.895 3346.875 380.175 ;
        RECT 3347.305 379.895 3347.585 380.175 ;
        RECT 3348.015 379.895 3348.295 380.175 ;
        RECT 3276.715 379.185 3276.995 379.465 ;
        RECT 3277.425 379.185 3277.705 379.465 ;
        RECT 3278.135 379.185 3278.415 379.465 ;
        RECT 3278.845 379.185 3279.125 379.465 ;
        RECT 3279.555 379.185 3279.835 379.465 ;
        RECT 3280.265 379.185 3280.545 379.465 ;
        RECT 3280.975 379.185 3281.255 379.465 ;
        RECT 3281.685 379.185 3281.965 379.465 ;
        RECT 3289.115 379.185 3289.395 379.465 ;
        RECT 3289.825 379.185 3290.105 379.465 ;
        RECT 3290.535 379.185 3290.815 379.465 ;
        RECT 3291.245 379.185 3291.525 379.465 ;
        RECT 3291.955 379.185 3292.235 379.465 ;
        RECT 3292.665 379.185 3292.945 379.465 ;
        RECT 3293.375 379.185 3293.655 379.465 ;
        RECT 3294.085 379.185 3294.365 379.465 ;
        RECT 3294.795 379.185 3295.075 379.465 ;
        RECT 3295.505 379.185 3295.785 379.465 ;
        RECT 3296.215 379.185 3296.495 379.465 ;
        RECT 3296.925 379.185 3297.205 379.465 ;
        RECT 3297.635 379.185 3297.915 379.465 ;
        RECT 3298.345 379.185 3298.625 379.465 ;
        RECT 3300.965 379.185 3301.245 379.465 ;
        RECT 3301.675 379.185 3301.955 379.465 ;
        RECT 3302.385 379.185 3302.665 379.465 ;
        RECT 3303.095 379.185 3303.375 379.465 ;
        RECT 3303.805 379.185 3304.085 379.465 ;
        RECT 3304.515 379.185 3304.795 379.465 ;
        RECT 3305.225 379.185 3305.505 379.465 ;
        RECT 3305.935 379.185 3306.215 379.465 ;
        RECT 3306.645 379.185 3306.925 379.465 ;
        RECT 3307.355 379.185 3307.635 379.465 ;
        RECT 3308.065 379.185 3308.345 379.465 ;
        RECT 3308.775 379.185 3309.055 379.465 ;
        RECT 3309.485 379.185 3309.765 379.465 ;
        RECT 3310.195 379.185 3310.475 379.465 ;
        RECT 3314.495 379.185 3314.775 379.465 ;
        RECT 3315.205 379.185 3315.485 379.465 ;
        RECT 3315.915 379.185 3316.195 379.465 ;
        RECT 3316.625 379.185 3316.905 379.465 ;
        RECT 3317.335 379.185 3317.615 379.465 ;
        RECT 3318.045 379.185 3318.325 379.465 ;
        RECT 3318.755 379.185 3319.035 379.465 ;
        RECT 3319.465 379.185 3319.745 379.465 ;
        RECT 3320.175 379.185 3320.455 379.465 ;
        RECT 3320.885 379.185 3321.165 379.465 ;
        RECT 3321.595 379.185 3321.875 379.465 ;
        RECT 3322.305 379.185 3322.585 379.465 ;
        RECT 3323.015 379.185 3323.295 379.465 ;
        RECT 3323.725 379.185 3324.005 379.465 ;
        RECT 3326.345 379.185 3326.625 379.465 ;
        RECT 3327.055 379.185 3327.335 379.465 ;
        RECT 3327.765 379.185 3328.045 379.465 ;
        RECT 3328.475 379.185 3328.755 379.465 ;
        RECT 3329.185 379.185 3329.465 379.465 ;
        RECT 3329.895 379.185 3330.175 379.465 ;
        RECT 3330.605 379.185 3330.885 379.465 ;
        RECT 3331.315 379.185 3331.595 379.465 ;
        RECT 3332.025 379.185 3332.305 379.465 ;
        RECT 3332.735 379.185 3333.015 379.465 ;
        RECT 3333.445 379.185 3333.725 379.465 ;
        RECT 3334.155 379.185 3334.435 379.465 ;
        RECT 3334.865 379.185 3335.145 379.465 ;
        RECT 3335.575 379.185 3335.855 379.465 ;
        RECT 3339.495 379.185 3339.775 379.465 ;
        RECT 3340.205 379.185 3340.485 379.465 ;
        RECT 3344.465 379.185 3344.745 379.465 ;
        RECT 3345.175 379.185 3345.455 379.465 ;
        RECT 3345.885 379.185 3346.165 379.465 ;
        RECT 3346.595 379.185 3346.875 379.465 ;
        RECT 3347.305 379.185 3347.585 379.465 ;
        RECT 3348.015 379.185 3348.295 379.465 ;
        RECT 3276.715 378.475 3276.995 378.755 ;
        RECT 3277.425 378.475 3277.705 378.755 ;
        RECT 3278.135 378.475 3278.415 378.755 ;
        RECT 3278.845 378.475 3279.125 378.755 ;
        RECT 3279.555 378.475 3279.835 378.755 ;
        RECT 3280.265 378.475 3280.545 378.755 ;
        RECT 3280.975 378.475 3281.255 378.755 ;
        RECT 3281.685 378.475 3281.965 378.755 ;
        RECT 3289.115 378.475 3289.395 378.755 ;
        RECT 3289.825 378.475 3290.105 378.755 ;
        RECT 3290.535 378.475 3290.815 378.755 ;
        RECT 3291.245 378.475 3291.525 378.755 ;
        RECT 3291.955 378.475 3292.235 378.755 ;
        RECT 3292.665 378.475 3292.945 378.755 ;
        RECT 3293.375 378.475 3293.655 378.755 ;
        RECT 3294.085 378.475 3294.365 378.755 ;
        RECT 3294.795 378.475 3295.075 378.755 ;
        RECT 3295.505 378.475 3295.785 378.755 ;
        RECT 3296.215 378.475 3296.495 378.755 ;
        RECT 3296.925 378.475 3297.205 378.755 ;
        RECT 3297.635 378.475 3297.915 378.755 ;
        RECT 3298.345 378.475 3298.625 378.755 ;
        RECT 3300.965 378.475 3301.245 378.755 ;
        RECT 3301.675 378.475 3301.955 378.755 ;
        RECT 3302.385 378.475 3302.665 378.755 ;
        RECT 3303.095 378.475 3303.375 378.755 ;
        RECT 3303.805 378.475 3304.085 378.755 ;
        RECT 3304.515 378.475 3304.795 378.755 ;
        RECT 3305.225 378.475 3305.505 378.755 ;
        RECT 3305.935 378.475 3306.215 378.755 ;
        RECT 3306.645 378.475 3306.925 378.755 ;
        RECT 3307.355 378.475 3307.635 378.755 ;
        RECT 3308.065 378.475 3308.345 378.755 ;
        RECT 3308.775 378.475 3309.055 378.755 ;
        RECT 3309.485 378.475 3309.765 378.755 ;
        RECT 3310.195 378.475 3310.475 378.755 ;
        RECT 3314.495 378.475 3314.775 378.755 ;
        RECT 3315.205 378.475 3315.485 378.755 ;
        RECT 3315.915 378.475 3316.195 378.755 ;
        RECT 3316.625 378.475 3316.905 378.755 ;
        RECT 3317.335 378.475 3317.615 378.755 ;
        RECT 3318.045 378.475 3318.325 378.755 ;
        RECT 3318.755 378.475 3319.035 378.755 ;
        RECT 3319.465 378.475 3319.745 378.755 ;
        RECT 3320.175 378.475 3320.455 378.755 ;
        RECT 3320.885 378.475 3321.165 378.755 ;
        RECT 3321.595 378.475 3321.875 378.755 ;
        RECT 3322.305 378.475 3322.585 378.755 ;
        RECT 3323.015 378.475 3323.295 378.755 ;
        RECT 3323.725 378.475 3324.005 378.755 ;
        RECT 3326.345 378.475 3326.625 378.755 ;
        RECT 3327.055 378.475 3327.335 378.755 ;
        RECT 3327.765 378.475 3328.045 378.755 ;
        RECT 3328.475 378.475 3328.755 378.755 ;
        RECT 3329.185 378.475 3329.465 378.755 ;
        RECT 3329.895 378.475 3330.175 378.755 ;
        RECT 3330.605 378.475 3330.885 378.755 ;
        RECT 3331.315 378.475 3331.595 378.755 ;
        RECT 3332.025 378.475 3332.305 378.755 ;
        RECT 3332.735 378.475 3333.015 378.755 ;
        RECT 3333.445 378.475 3333.725 378.755 ;
        RECT 3334.155 378.475 3334.435 378.755 ;
        RECT 3334.865 378.475 3335.145 378.755 ;
        RECT 3335.575 378.475 3335.855 378.755 ;
        RECT 3339.495 378.475 3339.775 378.755 ;
        RECT 3340.205 378.475 3340.485 378.755 ;
        RECT 3344.465 378.475 3344.745 378.755 ;
        RECT 3345.175 378.475 3345.455 378.755 ;
        RECT 3345.885 378.475 3346.165 378.755 ;
        RECT 3346.595 378.475 3346.875 378.755 ;
        RECT 3347.305 378.475 3347.585 378.755 ;
        RECT 3348.015 378.475 3348.295 378.755 ;
        RECT 3276.715 377.765 3276.995 378.045 ;
        RECT 3277.425 377.765 3277.705 378.045 ;
        RECT 3278.135 377.765 3278.415 378.045 ;
        RECT 3278.845 377.765 3279.125 378.045 ;
        RECT 3279.555 377.765 3279.835 378.045 ;
        RECT 3280.265 377.765 3280.545 378.045 ;
        RECT 3280.975 377.765 3281.255 378.045 ;
        RECT 3281.685 377.765 3281.965 378.045 ;
        RECT 3289.115 377.765 3289.395 378.045 ;
        RECT 3289.825 377.765 3290.105 378.045 ;
        RECT 3290.535 377.765 3290.815 378.045 ;
        RECT 3291.245 377.765 3291.525 378.045 ;
        RECT 3291.955 377.765 3292.235 378.045 ;
        RECT 3292.665 377.765 3292.945 378.045 ;
        RECT 3293.375 377.765 3293.655 378.045 ;
        RECT 3294.085 377.765 3294.365 378.045 ;
        RECT 3294.795 377.765 3295.075 378.045 ;
        RECT 3295.505 377.765 3295.785 378.045 ;
        RECT 3296.215 377.765 3296.495 378.045 ;
        RECT 3296.925 377.765 3297.205 378.045 ;
        RECT 3297.635 377.765 3297.915 378.045 ;
        RECT 3298.345 377.765 3298.625 378.045 ;
        RECT 3300.965 377.765 3301.245 378.045 ;
        RECT 3301.675 377.765 3301.955 378.045 ;
        RECT 3302.385 377.765 3302.665 378.045 ;
        RECT 3303.095 377.765 3303.375 378.045 ;
        RECT 3303.805 377.765 3304.085 378.045 ;
        RECT 3304.515 377.765 3304.795 378.045 ;
        RECT 3305.225 377.765 3305.505 378.045 ;
        RECT 3305.935 377.765 3306.215 378.045 ;
        RECT 3306.645 377.765 3306.925 378.045 ;
        RECT 3307.355 377.765 3307.635 378.045 ;
        RECT 3308.065 377.765 3308.345 378.045 ;
        RECT 3308.775 377.765 3309.055 378.045 ;
        RECT 3309.485 377.765 3309.765 378.045 ;
        RECT 3310.195 377.765 3310.475 378.045 ;
        RECT 3314.495 377.765 3314.775 378.045 ;
        RECT 3315.205 377.765 3315.485 378.045 ;
        RECT 3315.915 377.765 3316.195 378.045 ;
        RECT 3316.625 377.765 3316.905 378.045 ;
        RECT 3317.335 377.765 3317.615 378.045 ;
        RECT 3318.045 377.765 3318.325 378.045 ;
        RECT 3318.755 377.765 3319.035 378.045 ;
        RECT 3319.465 377.765 3319.745 378.045 ;
        RECT 3320.175 377.765 3320.455 378.045 ;
        RECT 3320.885 377.765 3321.165 378.045 ;
        RECT 3321.595 377.765 3321.875 378.045 ;
        RECT 3322.305 377.765 3322.585 378.045 ;
        RECT 3323.015 377.765 3323.295 378.045 ;
        RECT 3323.725 377.765 3324.005 378.045 ;
        RECT 3326.345 377.765 3326.625 378.045 ;
        RECT 3327.055 377.765 3327.335 378.045 ;
        RECT 3327.765 377.765 3328.045 378.045 ;
        RECT 3328.475 377.765 3328.755 378.045 ;
        RECT 3329.185 377.765 3329.465 378.045 ;
        RECT 3329.895 377.765 3330.175 378.045 ;
        RECT 3330.605 377.765 3330.885 378.045 ;
        RECT 3331.315 377.765 3331.595 378.045 ;
        RECT 3332.025 377.765 3332.305 378.045 ;
        RECT 3332.735 377.765 3333.015 378.045 ;
        RECT 3333.445 377.765 3333.725 378.045 ;
        RECT 3334.155 377.765 3334.435 378.045 ;
        RECT 3334.865 377.765 3335.145 378.045 ;
        RECT 3335.575 377.765 3335.855 378.045 ;
        RECT 3339.495 377.765 3339.775 378.045 ;
        RECT 3340.205 377.765 3340.485 378.045 ;
        RECT 3344.465 377.765 3344.745 378.045 ;
        RECT 3345.175 377.765 3345.455 378.045 ;
        RECT 3345.885 377.765 3346.165 378.045 ;
        RECT 3346.595 377.765 3346.875 378.045 ;
        RECT 3347.305 377.765 3347.585 378.045 ;
        RECT 3348.015 377.765 3348.295 378.045 ;
        RECT 3276.715 377.055 3276.995 377.335 ;
        RECT 3277.425 377.055 3277.705 377.335 ;
        RECT 3278.135 377.055 3278.415 377.335 ;
        RECT 3278.845 377.055 3279.125 377.335 ;
        RECT 3279.555 377.055 3279.835 377.335 ;
        RECT 3280.265 377.055 3280.545 377.335 ;
        RECT 3280.975 377.055 3281.255 377.335 ;
        RECT 3281.685 377.055 3281.965 377.335 ;
        RECT 3289.115 377.055 3289.395 377.335 ;
        RECT 3289.825 377.055 3290.105 377.335 ;
        RECT 3290.535 377.055 3290.815 377.335 ;
        RECT 3291.245 377.055 3291.525 377.335 ;
        RECT 3291.955 377.055 3292.235 377.335 ;
        RECT 3292.665 377.055 3292.945 377.335 ;
        RECT 3293.375 377.055 3293.655 377.335 ;
        RECT 3294.085 377.055 3294.365 377.335 ;
        RECT 3294.795 377.055 3295.075 377.335 ;
        RECT 3295.505 377.055 3295.785 377.335 ;
        RECT 3296.215 377.055 3296.495 377.335 ;
        RECT 3296.925 377.055 3297.205 377.335 ;
        RECT 3297.635 377.055 3297.915 377.335 ;
        RECT 3298.345 377.055 3298.625 377.335 ;
        RECT 3300.965 377.055 3301.245 377.335 ;
        RECT 3301.675 377.055 3301.955 377.335 ;
        RECT 3302.385 377.055 3302.665 377.335 ;
        RECT 3303.095 377.055 3303.375 377.335 ;
        RECT 3303.805 377.055 3304.085 377.335 ;
        RECT 3304.515 377.055 3304.795 377.335 ;
        RECT 3305.225 377.055 3305.505 377.335 ;
        RECT 3305.935 377.055 3306.215 377.335 ;
        RECT 3306.645 377.055 3306.925 377.335 ;
        RECT 3307.355 377.055 3307.635 377.335 ;
        RECT 3308.065 377.055 3308.345 377.335 ;
        RECT 3308.775 377.055 3309.055 377.335 ;
        RECT 3309.485 377.055 3309.765 377.335 ;
        RECT 3310.195 377.055 3310.475 377.335 ;
        RECT 3314.495 377.055 3314.775 377.335 ;
        RECT 3315.205 377.055 3315.485 377.335 ;
        RECT 3315.915 377.055 3316.195 377.335 ;
        RECT 3316.625 377.055 3316.905 377.335 ;
        RECT 3317.335 377.055 3317.615 377.335 ;
        RECT 3318.045 377.055 3318.325 377.335 ;
        RECT 3318.755 377.055 3319.035 377.335 ;
        RECT 3319.465 377.055 3319.745 377.335 ;
        RECT 3320.175 377.055 3320.455 377.335 ;
        RECT 3320.885 377.055 3321.165 377.335 ;
        RECT 3321.595 377.055 3321.875 377.335 ;
        RECT 3322.305 377.055 3322.585 377.335 ;
        RECT 3323.015 377.055 3323.295 377.335 ;
        RECT 3323.725 377.055 3324.005 377.335 ;
        RECT 3326.345 377.055 3326.625 377.335 ;
        RECT 3327.055 377.055 3327.335 377.335 ;
        RECT 3327.765 377.055 3328.045 377.335 ;
        RECT 3328.475 377.055 3328.755 377.335 ;
        RECT 3329.185 377.055 3329.465 377.335 ;
        RECT 3329.895 377.055 3330.175 377.335 ;
        RECT 3330.605 377.055 3330.885 377.335 ;
        RECT 3331.315 377.055 3331.595 377.335 ;
        RECT 3332.025 377.055 3332.305 377.335 ;
        RECT 3332.735 377.055 3333.015 377.335 ;
        RECT 3333.445 377.055 3333.725 377.335 ;
        RECT 3334.155 377.055 3334.435 377.335 ;
        RECT 3334.865 377.055 3335.145 377.335 ;
        RECT 3335.575 377.055 3335.855 377.335 ;
        RECT 3339.495 377.055 3339.775 377.335 ;
        RECT 3340.205 377.055 3340.485 377.335 ;
        RECT 3344.465 377.055 3344.745 377.335 ;
        RECT 3345.175 377.055 3345.455 377.335 ;
        RECT 3345.885 377.055 3346.165 377.335 ;
        RECT 3346.595 377.055 3346.875 377.335 ;
        RECT 3347.305 377.055 3347.585 377.335 ;
        RECT 3348.015 377.055 3348.295 377.335 ;
        RECT 3276.715 376.345 3276.995 376.625 ;
        RECT 3277.425 376.345 3277.705 376.625 ;
        RECT 3278.135 376.345 3278.415 376.625 ;
        RECT 3278.845 376.345 3279.125 376.625 ;
        RECT 3279.555 376.345 3279.835 376.625 ;
        RECT 3280.265 376.345 3280.545 376.625 ;
        RECT 3280.975 376.345 3281.255 376.625 ;
        RECT 3281.685 376.345 3281.965 376.625 ;
        RECT 3289.115 376.345 3289.395 376.625 ;
        RECT 3289.825 376.345 3290.105 376.625 ;
        RECT 3290.535 376.345 3290.815 376.625 ;
        RECT 3291.245 376.345 3291.525 376.625 ;
        RECT 3291.955 376.345 3292.235 376.625 ;
        RECT 3292.665 376.345 3292.945 376.625 ;
        RECT 3293.375 376.345 3293.655 376.625 ;
        RECT 3294.085 376.345 3294.365 376.625 ;
        RECT 3294.795 376.345 3295.075 376.625 ;
        RECT 3295.505 376.345 3295.785 376.625 ;
        RECT 3296.215 376.345 3296.495 376.625 ;
        RECT 3296.925 376.345 3297.205 376.625 ;
        RECT 3297.635 376.345 3297.915 376.625 ;
        RECT 3298.345 376.345 3298.625 376.625 ;
        RECT 3300.965 376.345 3301.245 376.625 ;
        RECT 3301.675 376.345 3301.955 376.625 ;
        RECT 3302.385 376.345 3302.665 376.625 ;
        RECT 3303.095 376.345 3303.375 376.625 ;
        RECT 3303.805 376.345 3304.085 376.625 ;
        RECT 3304.515 376.345 3304.795 376.625 ;
        RECT 3305.225 376.345 3305.505 376.625 ;
        RECT 3305.935 376.345 3306.215 376.625 ;
        RECT 3306.645 376.345 3306.925 376.625 ;
        RECT 3307.355 376.345 3307.635 376.625 ;
        RECT 3308.065 376.345 3308.345 376.625 ;
        RECT 3308.775 376.345 3309.055 376.625 ;
        RECT 3309.485 376.345 3309.765 376.625 ;
        RECT 3310.195 376.345 3310.475 376.625 ;
        RECT 3314.495 376.345 3314.775 376.625 ;
        RECT 3315.205 376.345 3315.485 376.625 ;
        RECT 3315.915 376.345 3316.195 376.625 ;
        RECT 3316.625 376.345 3316.905 376.625 ;
        RECT 3317.335 376.345 3317.615 376.625 ;
        RECT 3318.045 376.345 3318.325 376.625 ;
        RECT 3318.755 376.345 3319.035 376.625 ;
        RECT 3319.465 376.345 3319.745 376.625 ;
        RECT 3320.175 376.345 3320.455 376.625 ;
        RECT 3320.885 376.345 3321.165 376.625 ;
        RECT 3321.595 376.345 3321.875 376.625 ;
        RECT 3322.305 376.345 3322.585 376.625 ;
        RECT 3323.015 376.345 3323.295 376.625 ;
        RECT 3323.725 376.345 3324.005 376.625 ;
        RECT 3326.345 376.345 3326.625 376.625 ;
        RECT 3327.055 376.345 3327.335 376.625 ;
        RECT 3327.765 376.345 3328.045 376.625 ;
        RECT 3328.475 376.345 3328.755 376.625 ;
        RECT 3329.185 376.345 3329.465 376.625 ;
        RECT 3329.895 376.345 3330.175 376.625 ;
        RECT 3330.605 376.345 3330.885 376.625 ;
        RECT 3331.315 376.345 3331.595 376.625 ;
        RECT 3332.025 376.345 3332.305 376.625 ;
        RECT 3332.735 376.345 3333.015 376.625 ;
        RECT 3333.445 376.345 3333.725 376.625 ;
        RECT 3334.155 376.345 3334.435 376.625 ;
        RECT 3334.865 376.345 3335.145 376.625 ;
        RECT 3335.575 376.345 3335.855 376.625 ;
        RECT 3339.495 376.345 3339.775 376.625 ;
        RECT 3340.205 376.345 3340.485 376.625 ;
        RECT 3344.465 376.345 3344.745 376.625 ;
        RECT 3345.175 376.345 3345.455 376.625 ;
        RECT 3345.885 376.345 3346.165 376.625 ;
        RECT 3346.595 376.345 3346.875 376.625 ;
        RECT 3347.305 376.345 3347.585 376.625 ;
        RECT 3348.015 376.345 3348.295 376.625 ;
        RECT 3276.715 375.635 3276.995 375.915 ;
        RECT 3277.425 375.635 3277.705 375.915 ;
        RECT 3278.135 375.635 3278.415 375.915 ;
        RECT 3278.845 375.635 3279.125 375.915 ;
        RECT 3279.555 375.635 3279.835 375.915 ;
        RECT 3280.265 375.635 3280.545 375.915 ;
        RECT 3280.975 375.635 3281.255 375.915 ;
        RECT 3281.685 375.635 3281.965 375.915 ;
        RECT 3289.115 375.635 3289.395 375.915 ;
        RECT 3289.825 375.635 3290.105 375.915 ;
        RECT 3290.535 375.635 3290.815 375.915 ;
        RECT 3291.245 375.635 3291.525 375.915 ;
        RECT 3291.955 375.635 3292.235 375.915 ;
        RECT 3292.665 375.635 3292.945 375.915 ;
        RECT 3293.375 375.635 3293.655 375.915 ;
        RECT 3294.085 375.635 3294.365 375.915 ;
        RECT 3294.795 375.635 3295.075 375.915 ;
        RECT 3295.505 375.635 3295.785 375.915 ;
        RECT 3296.215 375.635 3296.495 375.915 ;
        RECT 3296.925 375.635 3297.205 375.915 ;
        RECT 3297.635 375.635 3297.915 375.915 ;
        RECT 3298.345 375.635 3298.625 375.915 ;
        RECT 3300.965 375.635 3301.245 375.915 ;
        RECT 3301.675 375.635 3301.955 375.915 ;
        RECT 3302.385 375.635 3302.665 375.915 ;
        RECT 3303.095 375.635 3303.375 375.915 ;
        RECT 3303.805 375.635 3304.085 375.915 ;
        RECT 3304.515 375.635 3304.795 375.915 ;
        RECT 3305.225 375.635 3305.505 375.915 ;
        RECT 3305.935 375.635 3306.215 375.915 ;
        RECT 3306.645 375.635 3306.925 375.915 ;
        RECT 3307.355 375.635 3307.635 375.915 ;
        RECT 3308.065 375.635 3308.345 375.915 ;
        RECT 3308.775 375.635 3309.055 375.915 ;
        RECT 3309.485 375.635 3309.765 375.915 ;
        RECT 3310.195 375.635 3310.475 375.915 ;
        RECT 3314.495 375.635 3314.775 375.915 ;
        RECT 3315.205 375.635 3315.485 375.915 ;
        RECT 3315.915 375.635 3316.195 375.915 ;
        RECT 3316.625 375.635 3316.905 375.915 ;
        RECT 3317.335 375.635 3317.615 375.915 ;
        RECT 3318.045 375.635 3318.325 375.915 ;
        RECT 3318.755 375.635 3319.035 375.915 ;
        RECT 3319.465 375.635 3319.745 375.915 ;
        RECT 3320.175 375.635 3320.455 375.915 ;
        RECT 3320.885 375.635 3321.165 375.915 ;
        RECT 3321.595 375.635 3321.875 375.915 ;
        RECT 3322.305 375.635 3322.585 375.915 ;
        RECT 3323.015 375.635 3323.295 375.915 ;
        RECT 3323.725 375.635 3324.005 375.915 ;
        RECT 3326.345 375.635 3326.625 375.915 ;
        RECT 3327.055 375.635 3327.335 375.915 ;
        RECT 3327.765 375.635 3328.045 375.915 ;
        RECT 3328.475 375.635 3328.755 375.915 ;
        RECT 3329.185 375.635 3329.465 375.915 ;
        RECT 3329.895 375.635 3330.175 375.915 ;
        RECT 3330.605 375.635 3330.885 375.915 ;
        RECT 3331.315 375.635 3331.595 375.915 ;
        RECT 3332.025 375.635 3332.305 375.915 ;
        RECT 3332.735 375.635 3333.015 375.915 ;
        RECT 3333.445 375.635 3333.725 375.915 ;
        RECT 3334.155 375.635 3334.435 375.915 ;
        RECT 3334.865 375.635 3335.145 375.915 ;
        RECT 3335.575 375.635 3335.855 375.915 ;
        RECT 3339.495 375.635 3339.775 375.915 ;
        RECT 3340.205 375.635 3340.485 375.915 ;
        RECT 3344.465 375.635 3344.745 375.915 ;
        RECT 3345.175 375.635 3345.455 375.915 ;
        RECT 3345.885 375.635 3346.165 375.915 ;
        RECT 3346.595 375.635 3346.875 375.915 ;
        RECT 3347.305 375.635 3347.585 375.915 ;
        RECT 3348.015 375.635 3348.295 375.915 ;
        RECT 3276.715 374.925 3276.995 375.205 ;
        RECT 3277.425 374.925 3277.705 375.205 ;
        RECT 3278.135 374.925 3278.415 375.205 ;
        RECT 3278.845 374.925 3279.125 375.205 ;
        RECT 3279.555 374.925 3279.835 375.205 ;
        RECT 3280.265 374.925 3280.545 375.205 ;
        RECT 3280.975 374.925 3281.255 375.205 ;
        RECT 3281.685 374.925 3281.965 375.205 ;
        RECT 3289.115 374.925 3289.395 375.205 ;
        RECT 3289.825 374.925 3290.105 375.205 ;
        RECT 3290.535 374.925 3290.815 375.205 ;
        RECT 3291.245 374.925 3291.525 375.205 ;
        RECT 3291.955 374.925 3292.235 375.205 ;
        RECT 3292.665 374.925 3292.945 375.205 ;
        RECT 3293.375 374.925 3293.655 375.205 ;
        RECT 3294.085 374.925 3294.365 375.205 ;
        RECT 3294.795 374.925 3295.075 375.205 ;
        RECT 3295.505 374.925 3295.785 375.205 ;
        RECT 3296.215 374.925 3296.495 375.205 ;
        RECT 3296.925 374.925 3297.205 375.205 ;
        RECT 3297.635 374.925 3297.915 375.205 ;
        RECT 3298.345 374.925 3298.625 375.205 ;
        RECT 3300.965 374.925 3301.245 375.205 ;
        RECT 3301.675 374.925 3301.955 375.205 ;
        RECT 3302.385 374.925 3302.665 375.205 ;
        RECT 3303.095 374.925 3303.375 375.205 ;
        RECT 3303.805 374.925 3304.085 375.205 ;
        RECT 3304.515 374.925 3304.795 375.205 ;
        RECT 3305.225 374.925 3305.505 375.205 ;
        RECT 3305.935 374.925 3306.215 375.205 ;
        RECT 3306.645 374.925 3306.925 375.205 ;
        RECT 3307.355 374.925 3307.635 375.205 ;
        RECT 3308.065 374.925 3308.345 375.205 ;
        RECT 3308.775 374.925 3309.055 375.205 ;
        RECT 3309.485 374.925 3309.765 375.205 ;
        RECT 3310.195 374.925 3310.475 375.205 ;
        RECT 3314.495 374.925 3314.775 375.205 ;
        RECT 3315.205 374.925 3315.485 375.205 ;
        RECT 3315.915 374.925 3316.195 375.205 ;
        RECT 3316.625 374.925 3316.905 375.205 ;
        RECT 3317.335 374.925 3317.615 375.205 ;
        RECT 3318.045 374.925 3318.325 375.205 ;
        RECT 3318.755 374.925 3319.035 375.205 ;
        RECT 3319.465 374.925 3319.745 375.205 ;
        RECT 3320.175 374.925 3320.455 375.205 ;
        RECT 3320.885 374.925 3321.165 375.205 ;
        RECT 3321.595 374.925 3321.875 375.205 ;
        RECT 3322.305 374.925 3322.585 375.205 ;
        RECT 3323.015 374.925 3323.295 375.205 ;
        RECT 3323.725 374.925 3324.005 375.205 ;
        RECT 3326.345 374.925 3326.625 375.205 ;
        RECT 3327.055 374.925 3327.335 375.205 ;
        RECT 3327.765 374.925 3328.045 375.205 ;
        RECT 3328.475 374.925 3328.755 375.205 ;
        RECT 3329.185 374.925 3329.465 375.205 ;
        RECT 3329.895 374.925 3330.175 375.205 ;
        RECT 3330.605 374.925 3330.885 375.205 ;
        RECT 3331.315 374.925 3331.595 375.205 ;
        RECT 3332.025 374.925 3332.305 375.205 ;
        RECT 3332.735 374.925 3333.015 375.205 ;
        RECT 3333.445 374.925 3333.725 375.205 ;
        RECT 3334.155 374.925 3334.435 375.205 ;
        RECT 3334.865 374.925 3335.145 375.205 ;
        RECT 3335.575 374.925 3335.855 375.205 ;
        RECT 3339.495 374.925 3339.775 375.205 ;
        RECT 3340.205 374.925 3340.485 375.205 ;
        RECT 3344.465 374.925 3344.745 375.205 ;
        RECT 3345.175 374.925 3345.455 375.205 ;
        RECT 3345.885 374.925 3346.165 375.205 ;
        RECT 3346.595 374.925 3346.875 375.205 ;
        RECT 3347.305 374.925 3347.585 375.205 ;
        RECT 3348.015 374.925 3348.295 375.205 ;
        RECT 3276.715 374.215 3276.995 374.495 ;
        RECT 3277.425 374.215 3277.705 374.495 ;
        RECT 3278.135 374.215 3278.415 374.495 ;
        RECT 3278.845 374.215 3279.125 374.495 ;
        RECT 3279.555 374.215 3279.835 374.495 ;
        RECT 3280.265 374.215 3280.545 374.495 ;
        RECT 3280.975 374.215 3281.255 374.495 ;
        RECT 3281.685 374.215 3281.965 374.495 ;
        RECT 3289.115 374.215 3289.395 374.495 ;
        RECT 3289.825 374.215 3290.105 374.495 ;
        RECT 3290.535 374.215 3290.815 374.495 ;
        RECT 3291.245 374.215 3291.525 374.495 ;
        RECT 3291.955 374.215 3292.235 374.495 ;
        RECT 3292.665 374.215 3292.945 374.495 ;
        RECT 3293.375 374.215 3293.655 374.495 ;
        RECT 3294.085 374.215 3294.365 374.495 ;
        RECT 3294.795 374.215 3295.075 374.495 ;
        RECT 3295.505 374.215 3295.785 374.495 ;
        RECT 3296.215 374.215 3296.495 374.495 ;
        RECT 3296.925 374.215 3297.205 374.495 ;
        RECT 3297.635 374.215 3297.915 374.495 ;
        RECT 3298.345 374.215 3298.625 374.495 ;
        RECT 3300.965 374.215 3301.245 374.495 ;
        RECT 3301.675 374.215 3301.955 374.495 ;
        RECT 3302.385 374.215 3302.665 374.495 ;
        RECT 3303.095 374.215 3303.375 374.495 ;
        RECT 3303.805 374.215 3304.085 374.495 ;
        RECT 3304.515 374.215 3304.795 374.495 ;
        RECT 3305.225 374.215 3305.505 374.495 ;
        RECT 3305.935 374.215 3306.215 374.495 ;
        RECT 3306.645 374.215 3306.925 374.495 ;
        RECT 3307.355 374.215 3307.635 374.495 ;
        RECT 3308.065 374.215 3308.345 374.495 ;
        RECT 3308.775 374.215 3309.055 374.495 ;
        RECT 3309.485 374.215 3309.765 374.495 ;
        RECT 3310.195 374.215 3310.475 374.495 ;
        RECT 3314.495 374.215 3314.775 374.495 ;
        RECT 3315.205 374.215 3315.485 374.495 ;
        RECT 3315.915 374.215 3316.195 374.495 ;
        RECT 3316.625 374.215 3316.905 374.495 ;
        RECT 3317.335 374.215 3317.615 374.495 ;
        RECT 3318.045 374.215 3318.325 374.495 ;
        RECT 3318.755 374.215 3319.035 374.495 ;
        RECT 3319.465 374.215 3319.745 374.495 ;
        RECT 3320.175 374.215 3320.455 374.495 ;
        RECT 3320.885 374.215 3321.165 374.495 ;
        RECT 3321.595 374.215 3321.875 374.495 ;
        RECT 3322.305 374.215 3322.585 374.495 ;
        RECT 3323.015 374.215 3323.295 374.495 ;
        RECT 3323.725 374.215 3324.005 374.495 ;
        RECT 3326.345 374.215 3326.625 374.495 ;
        RECT 3327.055 374.215 3327.335 374.495 ;
        RECT 3327.765 374.215 3328.045 374.495 ;
        RECT 3328.475 374.215 3328.755 374.495 ;
        RECT 3329.185 374.215 3329.465 374.495 ;
        RECT 3329.895 374.215 3330.175 374.495 ;
        RECT 3330.605 374.215 3330.885 374.495 ;
        RECT 3331.315 374.215 3331.595 374.495 ;
        RECT 3332.025 374.215 3332.305 374.495 ;
        RECT 3332.735 374.215 3333.015 374.495 ;
        RECT 3333.445 374.215 3333.725 374.495 ;
        RECT 3334.155 374.215 3334.435 374.495 ;
        RECT 3334.865 374.215 3335.145 374.495 ;
        RECT 3335.575 374.215 3335.855 374.495 ;
        RECT 3339.495 374.215 3339.775 374.495 ;
        RECT 3340.205 374.215 3340.485 374.495 ;
        RECT 3344.465 374.215 3344.745 374.495 ;
        RECT 3345.175 374.215 3345.455 374.495 ;
        RECT 3345.885 374.215 3346.165 374.495 ;
        RECT 3346.595 374.215 3346.875 374.495 ;
        RECT 3347.305 374.215 3347.585 374.495 ;
        RECT 3348.015 374.215 3348.295 374.495 ;
        RECT 3276.715 373.505 3276.995 373.785 ;
        RECT 3277.425 373.505 3277.705 373.785 ;
        RECT 3278.135 373.505 3278.415 373.785 ;
        RECT 3278.845 373.505 3279.125 373.785 ;
        RECT 3279.555 373.505 3279.835 373.785 ;
        RECT 3280.265 373.505 3280.545 373.785 ;
        RECT 3280.975 373.505 3281.255 373.785 ;
        RECT 3281.685 373.505 3281.965 373.785 ;
        RECT 3289.115 373.505 3289.395 373.785 ;
        RECT 3289.825 373.505 3290.105 373.785 ;
        RECT 3290.535 373.505 3290.815 373.785 ;
        RECT 3291.245 373.505 3291.525 373.785 ;
        RECT 3291.955 373.505 3292.235 373.785 ;
        RECT 3292.665 373.505 3292.945 373.785 ;
        RECT 3293.375 373.505 3293.655 373.785 ;
        RECT 3294.085 373.505 3294.365 373.785 ;
        RECT 3294.795 373.505 3295.075 373.785 ;
        RECT 3295.505 373.505 3295.785 373.785 ;
        RECT 3296.215 373.505 3296.495 373.785 ;
        RECT 3296.925 373.505 3297.205 373.785 ;
        RECT 3297.635 373.505 3297.915 373.785 ;
        RECT 3298.345 373.505 3298.625 373.785 ;
        RECT 3300.965 373.505 3301.245 373.785 ;
        RECT 3301.675 373.505 3301.955 373.785 ;
        RECT 3302.385 373.505 3302.665 373.785 ;
        RECT 3303.095 373.505 3303.375 373.785 ;
        RECT 3303.805 373.505 3304.085 373.785 ;
        RECT 3304.515 373.505 3304.795 373.785 ;
        RECT 3305.225 373.505 3305.505 373.785 ;
        RECT 3305.935 373.505 3306.215 373.785 ;
        RECT 3306.645 373.505 3306.925 373.785 ;
        RECT 3307.355 373.505 3307.635 373.785 ;
        RECT 3308.065 373.505 3308.345 373.785 ;
        RECT 3308.775 373.505 3309.055 373.785 ;
        RECT 3309.485 373.505 3309.765 373.785 ;
        RECT 3310.195 373.505 3310.475 373.785 ;
        RECT 3314.495 373.505 3314.775 373.785 ;
        RECT 3315.205 373.505 3315.485 373.785 ;
        RECT 3315.915 373.505 3316.195 373.785 ;
        RECT 3316.625 373.505 3316.905 373.785 ;
        RECT 3317.335 373.505 3317.615 373.785 ;
        RECT 3318.045 373.505 3318.325 373.785 ;
        RECT 3318.755 373.505 3319.035 373.785 ;
        RECT 3319.465 373.505 3319.745 373.785 ;
        RECT 3320.175 373.505 3320.455 373.785 ;
        RECT 3320.885 373.505 3321.165 373.785 ;
        RECT 3321.595 373.505 3321.875 373.785 ;
        RECT 3322.305 373.505 3322.585 373.785 ;
        RECT 3323.015 373.505 3323.295 373.785 ;
        RECT 3323.725 373.505 3324.005 373.785 ;
        RECT 3326.345 373.505 3326.625 373.785 ;
        RECT 3327.055 373.505 3327.335 373.785 ;
        RECT 3327.765 373.505 3328.045 373.785 ;
        RECT 3328.475 373.505 3328.755 373.785 ;
        RECT 3329.185 373.505 3329.465 373.785 ;
        RECT 3329.895 373.505 3330.175 373.785 ;
        RECT 3330.605 373.505 3330.885 373.785 ;
        RECT 3331.315 373.505 3331.595 373.785 ;
        RECT 3332.025 373.505 3332.305 373.785 ;
        RECT 3332.735 373.505 3333.015 373.785 ;
        RECT 3333.445 373.505 3333.725 373.785 ;
        RECT 3334.155 373.505 3334.435 373.785 ;
        RECT 3334.865 373.505 3335.145 373.785 ;
        RECT 3335.575 373.505 3335.855 373.785 ;
        RECT 3339.495 373.505 3339.775 373.785 ;
        RECT 3340.205 373.505 3340.485 373.785 ;
        RECT 3344.465 373.505 3344.745 373.785 ;
        RECT 3345.175 373.505 3345.455 373.785 ;
        RECT 3345.885 373.505 3346.165 373.785 ;
        RECT 3346.595 373.505 3346.875 373.785 ;
        RECT 3347.305 373.505 3347.585 373.785 ;
        RECT 3348.015 373.505 3348.295 373.785 ;
        RECT 3276.715 372.795 3276.995 373.075 ;
        RECT 3277.425 372.795 3277.705 373.075 ;
        RECT 3278.135 372.795 3278.415 373.075 ;
        RECT 3278.845 372.795 3279.125 373.075 ;
        RECT 3279.555 372.795 3279.835 373.075 ;
        RECT 3280.265 372.795 3280.545 373.075 ;
        RECT 3280.975 372.795 3281.255 373.075 ;
        RECT 3281.685 372.795 3281.965 373.075 ;
        RECT 3289.115 372.795 3289.395 373.075 ;
        RECT 3289.825 372.795 3290.105 373.075 ;
        RECT 3290.535 372.795 3290.815 373.075 ;
        RECT 3291.245 372.795 3291.525 373.075 ;
        RECT 3291.955 372.795 3292.235 373.075 ;
        RECT 3292.665 372.795 3292.945 373.075 ;
        RECT 3293.375 372.795 3293.655 373.075 ;
        RECT 3294.085 372.795 3294.365 373.075 ;
        RECT 3294.795 372.795 3295.075 373.075 ;
        RECT 3295.505 372.795 3295.785 373.075 ;
        RECT 3296.215 372.795 3296.495 373.075 ;
        RECT 3296.925 372.795 3297.205 373.075 ;
        RECT 3297.635 372.795 3297.915 373.075 ;
        RECT 3298.345 372.795 3298.625 373.075 ;
        RECT 3300.965 372.795 3301.245 373.075 ;
        RECT 3301.675 372.795 3301.955 373.075 ;
        RECT 3302.385 372.795 3302.665 373.075 ;
        RECT 3303.095 372.795 3303.375 373.075 ;
        RECT 3303.805 372.795 3304.085 373.075 ;
        RECT 3304.515 372.795 3304.795 373.075 ;
        RECT 3305.225 372.795 3305.505 373.075 ;
        RECT 3305.935 372.795 3306.215 373.075 ;
        RECT 3306.645 372.795 3306.925 373.075 ;
        RECT 3307.355 372.795 3307.635 373.075 ;
        RECT 3308.065 372.795 3308.345 373.075 ;
        RECT 3308.775 372.795 3309.055 373.075 ;
        RECT 3309.485 372.795 3309.765 373.075 ;
        RECT 3310.195 372.795 3310.475 373.075 ;
        RECT 3314.495 372.795 3314.775 373.075 ;
        RECT 3315.205 372.795 3315.485 373.075 ;
        RECT 3315.915 372.795 3316.195 373.075 ;
        RECT 3316.625 372.795 3316.905 373.075 ;
        RECT 3317.335 372.795 3317.615 373.075 ;
        RECT 3318.045 372.795 3318.325 373.075 ;
        RECT 3318.755 372.795 3319.035 373.075 ;
        RECT 3319.465 372.795 3319.745 373.075 ;
        RECT 3320.175 372.795 3320.455 373.075 ;
        RECT 3320.885 372.795 3321.165 373.075 ;
        RECT 3321.595 372.795 3321.875 373.075 ;
        RECT 3322.305 372.795 3322.585 373.075 ;
        RECT 3323.015 372.795 3323.295 373.075 ;
        RECT 3323.725 372.795 3324.005 373.075 ;
        RECT 3326.345 372.795 3326.625 373.075 ;
        RECT 3327.055 372.795 3327.335 373.075 ;
        RECT 3327.765 372.795 3328.045 373.075 ;
        RECT 3328.475 372.795 3328.755 373.075 ;
        RECT 3329.185 372.795 3329.465 373.075 ;
        RECT 3329.895 372.795 3330.175 373.075 ;
        RECT 3330.605 372.795 3330.885 373.075 ;
        RECT 3331.315 372.795 3331.595 373.075 ;
        RECT 3332.025 372.795 3332.305 373.075 ;
        RECT 3332.735 372.795 3333.015 373.075 ;
        RECT 3333.445 372.795 3333.725 373.075 ;
        RECT 3334.155 372.795 3334.435 373.075 ;
        RECT 3334.865 372.795 3335.145 373.075 ;
        RECT 3335.575 372.795 3335.855 373.075 ;
        RECT 3339.495 372.795 3339.775 373.075 ;
        RECT 3340.205 372.795 3340.485 373.075 ;
        RECT 3344.465 372.795 3344.745 373.075 ;
        RECT 3345.175 372.795 3345.455 373.075 ;
        RECT 3345.885 372.795 3346.165 373.075 ;
        RECT 3346.595 372.795 3346.875 373.075 ;
        RECT 3347.305 372.795 3347.585 373.075 ;
        RECT 3348.015 372.795 3348.295 373.075 ;
        RECT 526.715 369.895 526.995 370.175 ;
        RECT 527.425 369.895 527.705 370.175 ;
        RECT 528.135 369.895 528.415 370.175 ;
        RECT 528.845 369.895 529.125 370.175 ;
        RECT 529.555 369.895 529.835 370.175 ;
        RECT 530.265 369.895 530.545 370.175 ;
        RECT 530.975 369.895 531.255 370.175 ;
        RECT 531.685 369.895 531.965 370.175 ;
        RECT 532.395 369.895 532.675 370.175 ;
        RECT 533.105 369.895 533.385 370.175 ;
        RECT 533.815 369.895 534.095 370.175 ;
        RECT 534.525 369.895 534.805 370.175 ;
        RECT 535.235 369.895 535.515 370.175 ;
        RECT 544.975 369.895 545.255 370.175 ;
        RECT 545.685 369.895 545.965 370.175 ;
        RECT 546.395 369.895 546.675 370.175 ;
        RECT 547.105 369.895 547.385 370.175 ;
        RECT 547.815 369.895 548.095 370.175 ;
        RECT 548.525 369.895 548.805 370.175 ;
        RECT 550.965 369.895 551.245 370.175 ;
        RECT 551.675 369.895 551.955 370.175 ;
        RECT 552.385 369.895 552.665 370.175 ;
        RECT 553.095 369.895 553.375 370.175 ;
        RECT 553.805 369.895 554.085 370.175 ;
        RECT 554.515 369.895 554.795 370.175 ;
        RECT 555.225 369.895 555.505 370.175 ;
        RECT 555.935 369.895 556.215 370.175 ;
        RECT 556.645 369.895 556.925 370.175 ;
        RECT 557.355 369.895 557.635 370.175 ;
        RECT 558.065 369.895 558.345 370.175 ;
        RECT 558.775 369.895 559.055 370.175 ;
        RECT 559.485 369.895 559.765 370.175 ;
        RECT 560.195 369.895 560.475 370.175 ;
        RECT 566.625 369.895 566.905 370.175 ;
        RECT 567.335 369.895 567.615 370.175 ;
        RECT 568.045 369.895 568.325 370.175 ;
        RECT 568.755 369.895 569.035 370.175 ;
        RECT 569.465 369.895 569.745 370.175 ;
        RECT 570.175 369.895 570.455 370.175 ;
        RECT 570.885 369.895 571.165 370.175 ;
        RECT 571.595 369.895 571.875 370.175 ;
        RECT 572.305 369.895 572.585 370.175 ;
        RECT 573.015 369.895 573.295 370.175 ;
        RECT 573.725 369.895 574.005 370.175 ;
        RECT 576.345 369.895 576.625 370.175 ;
        RECT 577.055 369.895 577.335 370.175 ;
        RECT 577.765 369.895 578.045 370.175 ;
        RECT 578.475 369.895 578.755 370.175 ;
        RECT 579.185 369.895 579.465 370.175 ;
        RECT 579.895 369.895 580.175 370.175 ;
        RECT 580.605 369.895 580.885 370.175 ;
        RECT 581.315 369.895 581.595 370.175 ;
        RECT 582.025 369.895 582.305 370.175 ;
        RECT 582.735 369.895 583.015 370.175 ;
        RECT 583.445 369.895 583.725 370.175 ;
        RECT 584.155 369.895 584.435 370.175 ;
        RECT 584.865 369.895 585.145 370.175 ;
        RECT 585.575 369.895 585.855 370.175 ;
        RECT 589.495 369.895 589.775 370.175 ;
        RECT 590.205 369.895 590.485 370.175 ;
        RECT 590.915 369.895 591.195 370.175 ;
        RECT 591.625 369.895 591.905 370.175 ;
        RECT 592.335 369.895 592.615 370.175 ;
        RECT 593.045 369.895 593.325 370.175 ;
        RECT 593.755 369.895 594.035 370.175 ;
        RECT 594.465 369.895 594.745 370.175 ;
        RECT 595.175 369.895 595.455 370.175 ;
        RECT 595.885 369.895 596.165 370.175 ;
        RECT 596.595 369.895 596.875 370.175 ;
        RECT 597.305 369.895 597.585 370.175 ;
        RECT 598.015 369.895 598.295 370.175 ;
        RECT 1351.715 369.895 1351.995 370.175 ;
        RECT 1352.425 369.895 1352.705 370.175 ;
        RECT 1353.135 369.895 1353.415 370.175 ;
        RECT 1353.845 369.895 1354.125 370.175 ;
        RECT 1354.555 369.895 1354.835 370.175 ;
        RECT 1355.265 369.895 1355.545 370.175 ;
        RECT 1355.975 369.895 1356.255 370.175 ;
        RECT 1356.685 369.895 1356.965 370.175 ;
        RECT 1357.395 369.895 1357.675 370.175 ;
        RECT 1358.105 369.895 1358.385 370.175 ;
        RECT 1358.815 369.895 1359.095 370.175 ;
        RECT 1359.525 369.895 1359.805 370.175 ;
        RECT 1360.235 369.895 1360.515 370.175 ;
        RECT 1366.245 369.895 1366.525 370.175 ;
        RECT 1366.955 369.895 1367.235 370.175 ;
        RECT 1367.665 369.895 1367.945 370.175 ;
        RECT 1368.375 369.895 1368.655 370.175 ;
        RECT 1369.085 369.895 1369.365 370.175 ;
        RECT 1369.795 369.895 1370.075 370.175 ;
        RECT 1370.505 369.895 1370.785 370.175 ;
        RECT 1371.215 369.895 1371.495 370.175 ;
        RECT 1371.925 369.895 1372.205 370.175 ;
        RECT 1372.635 369.895 1372.915 370.175 ;
        RECT 1373.345 369.895 1373.625 370.175 ;
        RECT 1375.965 369.895 1376.245 370.175 ;
        RECT 1376.675 369.895 1376.955 370.175 ;
        RECT 1377.385 369.895 1377.665 370.175 ;
        RECT 1378.095 369.895 1378.375 370.175 ;
        RECT 1378.805 369.895 1379.085 370.175 ;
        RECT 1379.515 369.895 1379.795 370.175 ;
        RECT 1380.225 369.895 1380.505 370.175 ;
        RECT 1380.935 369.895 1381.215 370.175 ;
        RECT 1381.645 369.895 1381.925 370.175 ;
        RECT 1382.355 369.895 1382.635 370.175 ;
        RECT 1383.065 369.895 1383.345 370.175 ;
        RECT 1383.775 369.895 1384.055 370.175 ;
        RECT 1384.485 369.895 1384.765 370.175 ;
        RECT 1385.195 369.895 1385.475 370.175 ;
        RECT 1389.495 369.895 1389.775 370.175 ;
        RECT 1390.205 369.895 1390.485 370.175 ;
        RECT 1390.915 369.895 1391.195 370.175 ;
        RECT 1391.625 369.895 1391.905 370.175 ;
        RECT 1392.335 369.895 1392.615 370.175 ;
        RECT 1393.045 369.895 1393.325 370.175 ;
        RECT 1393.755 369.895 1394.035 370.175 ;
        RECT 1394.465 369.895 1394.745 370.175 ;
        RECT 1395.175 369.895 1395.455 370.175 ;
        RECT 1395.885 369.895 1396.165 370.175 ;
        RECT 1396.595 369.895 1396.875 370.175 ;
        RECT 1397.305 369.895 1397.585 370.175 ;
        RECT 1398.015 369.895 1398.295 370.175 ;
        RECT 1398.725 369.895 1399.005 370.175 ;
        RECT 1401.345 369.895 1401.625 370.175 ;
        RECT 1402.055 369.895 1402.335 370.175 ;
        RECT 1402.765 369.895 1403.045 370.175 ;
        RECT 1403.475 369.895 1403.755 370.175 ;
        RECT 1404.185 369.895 1404.465 370.175 ;
        RECT 1404.895 369.895 1405.175 370.175 ;
        RECT 1405.605 369.895 1405.885 370.175 ;
        RECT 1406.315 369.895 1406.595 370.175 ;
        RECT 1407.025 369.895 1407.305 370.175 ;
        RECT 1407.735 369.895 1408.015 370.175 ;
        RECT 1408.445 369.895 1408.725 370.175 ;
        RECT 1409.155 369.895 1409.435 370.175 ;
        RECT 1409.865 369.895 1410.145 370.175 ;
        RECT 1410.575 369.895 1410.855 370.175 ;
        RECT 1414.495 369.895 1414.775 370.175 ;
        RECT 1415.205 369.895 1415.485 370.175 ;
        RECT 1415.915 369.895 1416.195 370.175 ;
        RECT 1416.625 369.895 1416.905 370.175 ;
        RECT 1417.335 369.895 1417.615 370.175 ;
        RECT 1418.045 369.895 1418.325 370.175 ;
        RECT 1418.755 369.895 1419.035 370.175 ;
        RECT 1419.465 369.895 1419.745 370.175 ;
        RECT 3001.715 369.895 3001.995 370.175 ;
        RECT 3002.425 369.895 3002.705 370.175 ;
        RECT 3003.135 369.895 3003.415 370.175 ;
        RECT 3003.845 369.895 3004.125 370.175 ;
        RECT 3004.555 369.895 3004.835 370.175 ;
        RECT 3005.265 369.895 3005.545 370.175 ;
        RECT 3005.975 369.895 3006.255 370.175 ;
        RECT 3006.685 369.895 3006.965 370.175 ;
        RECT 3007.395 369.895 3007.675 370.175 ;
        RECT 3008.105 369.895 3008.385 370.175 ;
        RECT 3008.815 369.895 3009.095 370.175 ;
        RECT 3009.525 369.895 3009.805 370.175 ;
        RECT 3010.235 369.895 3010.515 370.175 ;
        RECT 3014.115 369.895 3014.395 370.175 ;
        RECT 3014.825 369.895 3015.105 370.175 ;
        RECT 3015.535 369.895 3015.815 370.175 ;
        RECT 3016.245 369.895 3016.525 370.175 ;
        RECT 3016.955 369.895 3017.235 370.175 ;
        RECT 3017.665 369.895 3017.945 370.175 ;
        RECT 3018.375 369.895 3018.655 370.175 ;
        RECT 3019.085 369.895 3019.365 370.175 ;
        RECT 3019.795 369.895 3020.075 370.175 ;
        RECT 3025.965 369.895 3026.245 370.175 ;
        RECT 3026.675 369.895 3026.955 370.175 ;
        RECT 3027.385 369.895 3027.665 370.175 ;
        RECT 3028.095 369.895 3028.375 370.175 ;
        RECT 3028.805 369.895 3029.085 370.175 ;
        RECT 3029.515 369.895 3029.795 370.175 ;
        RECT 3030.225 369.895 3030.505 370.175 ;
        RECT 3030.935 369.895 3031.215 370.175 ;
        RECT 3031.645 369.895 3031.925 370.175 ;
        RECT 3032.355 369.895 3032.635 370.175 ;
        RECT 3033.065 369.895 3033.345 370.175 ;
        RECT 3033.775 369.895 3034.055 370.175 ;
        RECT 3034.485 369.895 3034.765 370.175 ;
        RECT 3035.195 369.895 3035.475 370.175 ;
        RECT 3039.495 369.895 3039.775 370.175 ;
        RECT 3040.205 369.895 3040.485 370.175 ;
        RECT 3040.915 369.895 3041.195 370.175 ;
        RECT 3041.625 369.895 3041.905 370.175 ;
        RECT 3042.335 369.895 3042.615 370.175 ;
        RECT 3046.595 369.895 3046.875 370.175 ;
        RECT 3047.305 369.895 3047.585 370.175 ;
        RECT 3048.015 369.895 3048.295 370.175 ;
        RECT 3048.725 369.895 3049.005 370.175 ;
        RECT 3051.345 369.895 3051.625 370.175 ;
        RECT 3052.055 369.895 3052.335 370.175 ;
        RECT 3052.765 369.895 3053.045 370.175 ;
        RECT 3053.475 369.895 3053.755 370.175 ;
        RECT 3054.185 369.895 3054.465 370.175 ;
        RECT 3054.895 369.895 3055.175 370.175 ;
        RECT 3055.605 369.895 3055.885 370.175 ;
        RECT 3056.315 369.895 3056.595 370.175 ;
        RECT 3057.025 369.895 3057.305 370.175 ;
        RECT 3057.735 369.895 3058.015 370.175 ;
        RECT 3058.445 369.895 3058.725 370.175 ;
        RECT 3059.155 369.895 3059.435 370.175 ;
        RECT 3059.865 369.895 3060.145 370.175 ;
        RECT 3060.575 369.895 3060.855 370.175 ;
        RECT 3064.495 369.895 3064.775 370.175 ;
        RECT 3065.205 369.895 3065.485 370.175 ;
        RECT 3065.915 369.895 3066.195 370.175 ;
        RECT 3066.625 369.895 3066.905 370.175 ;
        RECT 3067.335 369.895 3067.615 370.175 ;
        RECT 3068.045 369.895 3068.325 370.175 ;
        RECT 3068.755 369.895 3069.035 370.175 ;
        RECT 3069.465 369.895 3069.745 370.175 ;
        RECT 3070.175 369.895 3070.455 370.175 ;
        RECT 3070.885 369.895 3071.165 370.175 ;
        RECT 3071.595 369.895 3071.875 370.175 ;
        RECT 3072.305 369.895 3072.585 370.175 ;
        RECT 3073.015 369.895 3073.295 370.175 ;
        RECT 526.715 369.185 526.995 369.465 ;
        RECT 527.425 369.185 527.705 369.465 ;
        RECT 528.135 369.185 528.415 369.465 ;
        RECT 528.845 369.185 529.125 369.465 ;
        RECT 529.555 369.185 529.835 369.465 ;
        RECT 530.265 369.185 530.545 369.465 ;
        RECT 530.975 369.185 531.255 369.465 ;
        RECT 531.685 369.185 531.965 369.465 ;
        RECT 532.395 369.185 532.675 369.465 ;
        RECT 533.105 369.185 533.385 369.465 ;
        RECT 533.815 369.185 534.095 369.465 ;
        RECT 534.525 369.185 534.805 369.465 ;
        RECT 535.235 369.185 535.515 369.465 ;
        RECT 544.975 369.185 545.255 369.465 ;
        RECT 545.685 369.185 545.965 369.465 ;
        RECT 546.395 369.185 546.675 369.465 ;
        RECT 547.105 369.185 547.385 369.465 ;
        RECT 547.815 369.185 548.095 369.465 ;
        RECT 548.525 369.185 548.805 369.465 ;
        RECT 550.965 369.185 551.245 369.465 ;
        RECT 551.675 369.185 551.955 369.465 ;
        RECT 552.385 369.185 552.665 369.465 ;
        RECT 553.095 369.185 553.375 369.465 ;
        RECT 553.805 369.185 554.085 369.465 ;
        RECT 554.515 369.185 554.795 369.465 ;
        RECT 555.225 369.185 555.505 369.465 ;
        RECT 555.935 369.185 556.215 369.465 ;
        RECT 556.645 369.185 556.925 369.465 ;
        RECT 557.355 369.185 557.635 369.465 ;
        RECT 558.065 369.185 558.345 369.465 ;
        RECT 558.775 369.185 559.055 369.465 ;
        RECT 559.485 369.185 559.765 369.465 ;
        RECT 560.195 369.185 560.475 369.465 ;
        RECT 566.625 369.185 566.905 369.465 ;
        RECT 567.335 369.185 567.615 369.465 ;
        RECT 568.045 369.185 568.325 369.465 ;
        RECT 568.755 369.185 569.035 369.465 ;
        RECT 569.465 369.185 569.745 369.465 ;
        RECT 570.175 369.185 570.455 369.465 ;
        RECT 570.885 369.185 571.165 369.465 ;
        RECT 571.595 369.185 571.875 369.465 ;
        RECT 572.305 369.185 572.585 369.465 ;
        RECT 573.015 369.185 573.295 369.465 ;
        RECT 573.725 369.185 574.005 369.465 ;
        RECT 576.345 369.185 576.625 369.465 ;
        RECT 577.055 369.185 577.335 369.465 ;
        RECT 577.765 369.185 578.045 369.465 ;
        RECT 578.475 369.185 578.755 369.465 ;
        RECT 579.185 369.185 579.465 369.465 ;
        RECT 579.895 369.185 580.175 369.465 ;
        RECT 580.605 369.185 580.885 369.465 ;
        RECT 581.315 369.185 581.595 369.465 ;
        RECT 582.025 369.185 582.305 369.465 ;
        RECT 582.735 369.185 583.015 369.465 ;
        RECT 583.445 369.185 583.725 369.465 ;
        RECT 584.155 369.185 584.435 369.465 ;
        RECT 584.865 369.185 585.145 369.465 ;
        RECT 585.575 369.185 585.855 369.465 ;
        RECT 589.495 369.185 589.775 369.465 ;
        RECT 590.205 369.185 590.485 369.465 ;
        RECT 590.915 369.185 591.195 369.465 ;
        RECT 591.625 369.185 591.905 369.465 ;
        RECT 592.335 369.185 592.615 369.465 ;
        RECT 593.045 369.185 593.325 369.465 ;
        RECT 593.755 369.185 594.035 369.465 ;
        RECT 594.465 369.185 594.745 369.465 ;
        RECT 595.175 369.185 595.455 369.465 ;
        RECT 595.885 369.185 596.165 369.465 ;
        RECT 596.595 369.185 596.875 369.465 ;
        RECT 597.305 369.185 597.585 369.465 ;
        RECT 598.015 369.185 598.295 369.465 ;
        RECT 1351.715 369.185 1351.995 369.465 ;
        RECT 1352.425 369.185 1352.705 369.465 ;
        RECT 1353.135 369.185 1353.415 369.465 ;
        RECT 1353.845 369.185 1354.125 369.465 ;
        RECT 1354.555 369.185 1354.835 369.465 ;
        RECT 1355.265 369.185 1355.545 369.465 ;
        RECT 1355.975 369.185 1356.255 369.465 ;
        RECT 1356.685 369.185 1356.965 369.465 ;
        RECT 1357.395 369.185 1357.675 369.465 ;
        RECT 1358.105 369.185 1358.385 369.465 ;
        RECT 1358.815 369.185 1359.095 369.465 ;
        RECT 1359.525 369.185 1359.805 369.465 ;
        RECT 1360.235 369.185 1360.515 369.465 ;
        RECT 1366.245 369.185 1366.525 369.465 ;
        RECT 1366.955 369.185 1367.235 369.465 ;
        RECT 1367.665 369.185 1367.945 369.465 ;
        RECT 1368.375 369.185 1368.655 369.465 ;
        RECT 1369.085 369.185 1369.365 369.465 ;
        RECT 1369.795 369.185 1370.075 369.465 ;
        RECT 1370.505 369.185 1370.785 369.465 ;
        RECT 1371.215 369.185 1371.495 369.465 ;
        RECT 1371.925 369.185 1372.205 369.465 ;
        RECT 1372.635 369.185 1372.915 369.465 ;
        RECT 1373.345 369.185 1373.625 369.465 ;
        RECT 1375.965 369.185 1376.245 369.465 ;
        RECT 1376.675 369.185 1376.955 369.465 ;
        RECT 1377.385 369.185 1377.665 369.465 ;
        RECT 1378.095 369.185 1378.375 369.465 ;
        RECT 1378.805 369.185 1379.085 369.465 ;
        RECT 1379.515 369.185 1379.795 369.465 ;
        RECT 1380.225 369.185 1380.505 369.465 ;
        RECT 1380.935 369.185 1381.215 369.465 ;
        RECT 1381.645 369.185 1381.925 369.465 ;
        RECT 1382.355 369.185 1382.635 369.465 ;
        RECT 1383.065 369.185 1383.345 369.465 ;
        RECT 1383.775 369.185 1384.055 369.465 ;
        RECT 1384.485 369.185 1384.765 369.465 ;
        RECT 1385.195 369.185 1385.475 369.465 ;
        RECT 1389.495 369.185 1389.775 369.465 ;
        RECT 1390.205 369.185 1390.485 369.465 ;
        RECT 1390.915 369.185 1391.195 369.465 ;
        RECT 1391.625 369.185 1391.905 369.465 ;
        RECT 1392.335 369.185 1392.615 369.465 ;
        RECT 1393.045 369.185 1393.325 369.465 ;
        RECT 1393.755 369.185 1394.035 369.465 ;
        RECT 1394.465 369.185 1394.745 369.465 ;
        RECT 1395.175 369.185 1395.455 369.465 ;
        RECT 1395.885 369.185 1396.165 369.465 ;
        RECT 1396.595 369.185 1396.875 369.465 ;
        RECT 1397.305 369.185 1397.585 369.465 ;
        RECT 1398.015 369.185 1398.295 369.465 ;
        RECT 1398.725 369.185 1399.005 369.465 ;
        RECT 1401.345 369.185 1401.625 369.465 ;
        RECT 1402.055 369.185 1402.335 369.465 ;
        RECT 1402.765 369.185 1403.045 369.465 ;
        RECT 1403.475 369.185 1403.755 369.465 ;
        RECT 1404.185 369.185 1404.465 369.465 ;
        RECT 1404.895 369.185 1405.175 369.465 ;
        RECT 1405.605 369.185 1405.885 369.465 ;
        RECT 1406.315 369.185 1406.595 369.465 ;
        RECT 1407.025 369.185 1407.305 369.465 ;
        RECT 1407.735 369.185 1408.015 369.465 ;
        RECT 1408.445 369.185 1408.725 369.465 ;
        RECT 1409.155 369.185 1409.435 369.465 ;
        RECT 1409.865 369.185 1410.145 369.465 ;
        RECT 1410.575 369.185 1410.855 369.465 ;
        RECT 1414.495 369.185 1414.775 369.465 ;
        RECT 1415.205 369.185 1415.485 369.465 ;
        RECT 1415.915 369.185 1416.195 369.465 ;
        RECT 1416.625 369.185 1416.905 369.465 ;
        RECT 1417.335 369.185 1417.615 369.465 ;
        RECT 1418.045 369.185 1418.325 369.465 ;
        RECT 1418.755 369.185 1419.035 369.465 ;
        RECT 1419.465 369.185 1419.745 369.465 ;
        RECT 3001.715 369.185 3001.995 369.465 ;
        RECT 3002.425 369.185 3002.705 369.465 ;
        RECT 3003.135 369.185 3003.415 369.465 ;
        RECT 3003.845 369.185 3004.125 369.465 ;
        RECT 3004.555 369.185 3004.835 369.465 ;
        RECT 3005.265 369.185 3005.545 369.465 ;
        RECT 3005.975 369.185 3006.255 369.465 ;
        RECT 3006.685 369.185 3006.965 369.465 ;
        RECT 3007.395 369.185 3007.675 369.465 ;
        RECT 3008.105 369.185 3008.385 369.465 ;
        RECT 3008.815 369.185 3009.095 369.465 ;
        RECT 3009.525 369.185 3009.805 369.465 ;
        RECT 3010.235 369.185 3010.515 369.465 ;
        RECT 3014.115 369.185 3014.395 369.465 ;
        RECT 3014.825 369.185 3015.105 369.465 ;
        RECT 3015.535 369.185 3015.815 369.465 ;
        RECT 3016.245 369.185 3016.525 369.465 ;
        RECT 3016.955 369.185 3017.235 369.465 ;
        RECT 3017.665 369.185 3017.945 369.465 ;
        RECT 3018.375 369.185 3018.655 369.465 ;
        RECT 3019.085 369.185 3019.365 369.465 ;
        RECT 3019.795 369.185 3020.075 369.465 ;
        RECT 3025.965 369.185 3026.245 369.465 ;
        RECT 3026.675 369.185 3026.955 369.465 ;
        RECT 3027.385 369.185 3027.665 369.465 ;
        RECT 3028.095 369.185 3028.375 369.465 ;
        RECT 3028.805 369.185 3029.085 369.465 ;
        RECT 3029.515 369.185 3029.795 369.465 ;
        RECT 3030.225 369.185 3030.505 369.465 ;
        RECT 3030.935 369.185 3031.215 369.465 ;
        RECT 3031.645 369.185 3031.925 369.465 ;
        RECT 3032.355 369.185 3032.635 369.465 ;
        RECT 3033.065 369.185 3033.345 369.465 ;
        RECT 3033.775 369.185 3034.055 369.465 ;
        RECT 3034.485 369.185 3034.765 369.465 ;
        RECT 3035.195 369.185 3035.475 369.465 ;
        RECT 3039.495 369.185 3039.775 369.465 ;
        RECT 3040.205 369.185 3040.485 369.465 ;
        RECT 3040.915 369.185 3041.195 369.465 ;
        RECT 3041.625 369.185 3041.905 369.465 ;
        RECT 3042.335 369.185 3042.615 369.465 ;
        RECT 3046.595 369.185 3046.875 369.465 ;
        RECT 3047.305 369.185 3047.585 369.465 ;
        RECT 3048.015 369.185 3048.295 369.465 ;
        RECT 3048.725 369.185 3049.005 369.465 ;
        RECT 3051.345 369.185 3051.625 369.465 ;
        RECT 3052.055 369.185 3052.335 369.465 ;
        RECT 3052.765 369.185 3053.045 369.465 ;
        RECT 3053.475 369.185 3053.755 369.465 ;
        RECT 3054.185 369.185 3054.465 369.465 ;
        RECT 3054.895 369.185 3055.175 369.465 ;
        RECT 3055.605 369.185 3055.885 369.465 ;
        RECT 3056.315 369.185 3056.595 369.465 ;
        RECT 3057.025 369.185 3057.305 369.465 ;
        RECT 3057.735 369.185 3058.015 369.465 ;
        RECT 3058.445 369.185 3058.725 369.465 ;
        RECT 3059.155 369.185 3059.435 369.465 ;
        RECT 3059.865 369.185 3060.145 369.465 ;
        RECT 3060.575 369.185 3060.855 369.465 ;
        RECT 3064.495 369.185 3064.775 369.465 ;
        RECT 3065.205 369.185 3065.485 369.465 ;
        RECT 3065.915 369.185 3066.195 369.465 ;
        RECT 3066.625 369.185 3066.905 369.465 ;
        RECT 3067.335 369.185 3067.615 369.465 ;
        RECT 3068.045 369.185 3068.325 369.465 ;
        RECT 3068.755 369.185 3069.035 369.465 ;
        RECT 3069.465 369.185 3069.745 369.465 ;
        RECT 3070.175 369.185 3070.455 369.465 ;
        RECT 3070.885 369.185 3071.165 369.465 ;
        RECT 3071.595 369.185 3071.875 369.465 ;
        RECT 3072.305 369.185 3072.585 369.465 ;
        RECT 3073.015 369.185 3073.295 369.465 ;
        RECT 526.715 368.475 526.995 368.755 ;
        RECT 527.425 368.475 527.705 368.755 ;
        RECT 528.135 368.475 528.415 368.755 ;
        RECT 528.845 368.475 529.125 368.755 ;
        RECT 529.555 368.475 529.835 368.755 ;
        RECT 530.265 368.475 530.545 368.755 ;
        RECT 530.975 368.475 531.255 368.755 ;
        RECT 531.685 368.475 531.965 368.755 ;
        RECT 532.395 368.475 532.675 368.755 ;
        RECT 533.105 368.475 533.385 368.755 ;
        RECT 533.815 368.475 534.095 368.755 ;
        RECT 534.525 368.475 534.805 368.755 ;
        RECT 535.235 368.475 535.515 368.755 ;
        RECT 544.975 368.475 545.255 368.755 ;
        RECT 545.685 368.475 545.965 368.755 ;
        RECT 546.395 368.475 546.675 368.755 ;
        RECT 547.105 368.475 547.385 368.755 ;
        RECT 547.815 368.475 548.095 368.755 ;
        RECT 548.525 368.475 548.805 368.755 ;
        RECT 550.965 368.475 551.245 368.755 ;
        RECT 551.675 368.475 551.955 368.755 ;
        RECT 552.385 368.475 552.665 368.755 ;
        RECT 553.095 368.475 553.375 368.755 ;
        RECT 553.805 368.475 554.085 368.755 ;
        RECT 554.515 368.475 554.795 368.755 ;
        RECT 555.225 368.475 555.505 368.755 ;
        RECT 555.935 368.475 556.215 368.755 ;
        RECT 556.645 368.475 556.925 368.755 ;
        RECT 557.355 368.475 557.635 368.755 ;
        RECT 558.065 368.475 558.345 368.755 ;
        RECT 558.775 368.475 559.055 368.755 ;
        RECT 559.485 368.475 559.765 368.755 ;
        RECT 560.195 368.475 560.475 368.755 ;
        RECT 566.625 368.475 566.905 368.755 ;
        RECT 567.335 368.475 567.615 368.755 ;
        RECT 568.045 368.475 568.325 368.755 ;
        RECT 568.755 368.475 569.035 368.755 ;
        RECT 569.465 368.475 569.745 368.755 ;
        RECT 570.175 368.475 570.455 368.755 ;
        RECT 570.885 368.475 571.165 368.755 ;
        RECT 571.595 368.475 571.875 368.755 ;
        RECT 572.305 368.475 572.585 368.755 ;
        RECT 573.015 368.475 573.295 368.755 ;
        RECT 573.725 368.475 574.005 368.755 ;
        RECT 576.345 368.475 576.625 368.755 ;
        RECT 577.055 368.475 577.335 368.755 ;
        RECT 577.765 368.475 578.045 368.755 ;
        RECT 578.475 368.475 578.755 368.755 ;
        RECT 579.185 368.475 579.465 368.755 ;
        RECT 579.895 368.475 580.175 368.755 ;
        RECT 580.605 368.475 580.885 368.755 ;
        RECT 581.315 368.475 581.595 368.755 ;
        RECT 582.025 368.475 582.305 368.755 ;
        RECT 582.735 368.475 583.015 368.755 ;
        RECT 583.445 368.475 583.725 368.755 ;
        RECT 584.155 368.475 584.435 368.755 ;
        RECT 584.865 368.475 585.145 368.755 ;
        RECT 585.575 368.475 585.855 368.755 ;
        RECT 589.495 368.475 589.775 368.755 ;
        RECT 590.205 368.475 590.485 368.755 ;
        RECT 590.915 368.475 591.195 368.755 ;
        RECT 591.625 368.475 591.905 368.755 ;
        RECT 592.335 368.475 592.615 368.755 ;
        RECT 593.045 368.475 593.325 368.755 ;
        RECT 593.755 368.475 594.035 368.755 ;
        RECT 594.465 368.475 594.745 368.755 ;
        RECT 595.175 368.475 595.455 368.755 ;
        RECT 595.885 368.475 596.165 368.755 ;
        RECT 596.595 368.475 596.875 368.755 ;
        RECT 597.305 368.475 597.585 368.755 ;
        RECT 598.015 368.475 598.295 368.755 ;
        RECT 1351.715 368.475 1351.995 368.755 ;
        RECT 1352.425 368.475 1352.705 368.755 ;
        RECT 1353.135 368.475 1353.415 368.755 ;
        RECT 1353.845 368.475 1354.125 368.755 ;
        RECT 1354.555 368.475 1354.835 368.755 ;
        RECT 1355.265 368.475 1355.545 368.755 ;
        RECT 1355.975 368.475 1356.255 368.755 ;
        RECT 1356.685 368.475 1356.965 368.755 ;
        RECT 1357.395 368.475 1357.675 368.755 ;
        RECT 1358.105 368.475 1358.385 368.755 ;
        RECT 1358.815 368.475 1359.095 368.755 ;
        RECT 1359.525 368.475 1359.805 368.755 ;
        RECT 1360.235 368.475 1360.515 368.755 ;
        RECT 1366.245 368.475 1366.525 368.755 ;
        RECT 1366.955 368.475 1367.235 368.755 ;
        RECT 1367.665 368.475 1367.945 368.755 ;
        RECT 1368.375 368.475 1368.655 368.755 ;
        RECT 1369.085 368.475 1369.365 368.755 ;
        RECT 1369.795 368.475 1370.075 368.755 ;
        RECT 1370.505 368.475 1370.785 368.755 ;
        RECT 1371.215 368.475 1371.495 368.755 ;
        RECT 1371.925 368.475 1372.205 368.755 ;
        RECT 1372.635 368.475 1372.915 368.755 ;
        RECT 1373.345 368.475 1373.625 368.755 ;
        RECT 1375.965 368.475 1376.245 368.755 ;
        RECT 1376.675 368.475 1376.955 368.755 ;
        RECT 1377.385 368.475 1377.665 368.755 ;
        RECT 1378.095 368.475 1378.375 368.755 ;
        RECT 1378.805 368.475 1379.085 368.755 ;
        RECT 1379.515 368.475 1379.795 368.755 ;
        RECT 1380.225 368.475 1380.505 368.755 ;
        RECT 1380.935 368.475 1381.215 368.755 ;
        RECT 1381.645 368.475 1381.925 368.755 ;
        RECT 1382.355 368.475 1382.635 368.755 ;
        RECT 1383.065 368.475 1383.345 368.755 ;
        RECT 1383.775 368.475 1384.055 368.755 ;
        RECT 1384.485 368.475 1384.765 368.755 ;
        RECT 1385.195 368.475 1385.475 368.755 ;
        RECT 1389.495 368.475 1389.775 368.755 ;
        RECT 1390.205 368.475 1390.485 368.755 ;
        RECT 1390.915 368.475 1391.195 368.755 ;
        RECT 1391.625 368.475 1391.905 368.755 ;
        RECT 1392.335 368.475 1392.615 368.755 ;
        RECT 1393.045 368.475 1393.325 368.755 ;
        RECT 1393.755 368.475 1394.035 368.755 ;
        RECT 1394.465 368.475 1394.745 368.755 ;
        RECT 1395.175 368.475 1395.455 368.755 ;
        RECT 1395.885 368.475 1396.165 368.755 ;
        RECT 1396.595 368.475 1396.875 368.755 ;
        RECT 1397.305 368.475 1397.585 368.755 ;
        RECT 1398.015 368.475 1398.295 368.755 ;
        RECT 1398.725 368.475 1399.005 368.755 ;
        RECT 1401.345 368.475 1401.625 368.755 ;
        RECT 1402.055 368.475 1402.335 368.755 ;
        RECT 1402.765 368.475 1403.045 368.755 ;
        RECT 1403.475 368.475 1403.755 368.755 ;
        RECT 1404.185 368.475 1404.465 368.755 ;
        RECT 1404.895 368.475 1405.175 368.755 ;
        RECT 1405.605 368.475 1405.885 368.755 ;
        RECT 1406.315 368.475 1406.595 368.755 ;
        RECT 1407.025 368.475 1407.305 368.755 ;
        RECT 1407.735 368.475 1408.015 368.755 ;
        RECT 1408.445 368.475 1408.725 368.755 ;
        RECT 1409.155 368.475 1409.435 368.755 ;
        RECT 1409.865 368.475 1410.145 368.755 ;
        RECT 1410.575 368.475 1410.855 368.755 ;
        RECT 1414.495 368.475 1414.775 368.755 ;
        RECT 1415.205 368.475 1415.485 368.755 ;
        RECT 1415.915 368.475 1416.195 368.755 ;
        RECT 1416.625 368.475 1416.905 368.755 ;
        RECT 1417.335 368.475 1417.615 368.755 ;
        RECT 1418.045 368.475 1418.325 368.755 ;
        RECT 1418.755 368.475 1419.035 368.755 ;
        RECT 1419.465 368.475 1419.745 368.755 ;
        RECT 3001.715 368.475 3001.995 368.755 ;
        RECT 3002.425 368.475 3002.705 368.755 ;
        RECT 3003.135 368.475 3003.415 368.755 ;
        RECT 3003.845 368.475 3004.125 368.755 ;
        RECT 3004.555 368.475 3004.835 368.755 ;
        RECT 3005.265 368.475 3005.545 368.755 ;
        RECT 3005.975 368.475 3006.255 368.755 ;
        RECT 3006.685 368.475 3006.965 368.755 ;
        RECT 3007.395 368.475 3007.675 368.755 ;
        RECT 3008.105 368.475 3008.385 368.755 ;
        RECT 3008.815 368.475 3009.095 368.755 ;
        RECT 3009.525 368.475 3009.805 368.755 ;
        RECT 3010.235 368.475 3010.515 368.755 ;
        RECT 3014.115 368.475 3014.395 368.755 ;
        RECT 3014.825 368.475 3015.105 368.755 ;
        RECT 3015.535 368.475 3015.815 368.755 ;
        RECT 3016.245 368.475 3016.525 368.755 ;
        RECT 3016.955 368.475 3017.235 368.755 ;
        RECT 3017.665 368.475 3017.945 368.755 ;
        RECT 3018.375 368.475 3018.655 368.755 ;
        RECT 3019.085 368.475 3019.365 368.755 ;
        RECT 3019.795 368.475 3020.075 368.755 ;
        RECT 3025.965 368.475 3026.245 368.755 ;
        RECT 3026.675 368.475 3026.955 368.755 ;
        RECT 3027.385 368.475 3027.665 368.755 ;
        RECT 3028.095 368.475 3028.375 368.755 ;
        RECT 3028.805 368.475 3029.085 368.755 ;
        RECT 3029.515 368.475 3029.795 368.755 ;
        RECT 3030.225 368.475 3030.505 368.755 ;
        RECT 3030.935 368.475 3031.215 368.755 ;
        RECT 3031.645 368.475 3031.925 368.755 ;
        RECT 3032.355 368.475 3032.635 368.755 ;
        RECT 3033.065 368.475 3033.345 368.755 ;
        RECT 3033.775 368.475 3034.055 368.755 ;
        RECT 3034.485 368.475 3034.765 368.755 ;
        RECT 3035.195 368.475 3035.475 368.755 ;
        RECT 3039.495 368.475 3039.775 368.755 ;
        RECT 3040.205 368.475 3040.485 368.755 ;
        RECT 3040.915 368.475 3041.195 368.755 ;
        RECT 3041.625 368.475 3041.905 368.755 ;
        RECT 3042.335 368.475 3042.615 368.755 ;
        RECT 3046.595 368.475 3046.875 368.755 ;
        RECT 3047.305 368.475 3047.585 368.755 ;
        RECT 3048.015 368.475 3048.295 368.755 ;
        RECT 3048.725 368.475 3049.005 368.755 ;
        RECT 3051.345 368.475 3051.625 368.755 ;
        RECT 3052.055 368.475 3052.335 368.755 ;
        RECT 3052.765 368.475 3053.045 368.755 ;
        RECT 3053.475 368.475 3053.755 368.755 ;
        RECT 3054.185 368.475 3054.465 368.755 ;
        RECT 3054.895 368.475 3055.175 368.755 ;
        RECT 3055.605 368.475 3055.885 368.755 ;
        RECT 3056.315 368.475 3056.595 368.755 ;
        RECT 3057.025 368.475 3057.305 368.755 ;
        RECT 3057.735 368.475 3058.015 368.755 ;
        RECT 3058.445 368.475 3058.725 368.755 ;
        RECT 3059.155 368.475 3059.435 368.755 ;
        RECT 3059.865 368.475 3060.145 368.755 ;
        RECT 3060.575 368.475 3060.855 368.755 ;
        RECT 3064.495 368.475 3064.775 368.755 ;
        RECT 3065.205 368.475 3065.485 368.755 ;
        RECT 3065.915 368.475 3066.195 368.755 ;
        RECT 3066.625 368.475 3066.905 368.755 ;
        RECT 3067.335 368.475 3067.615 368.755 ;
        RECT 3068.045 368.475 3068.325 368.755 ;
        RECT 3068.755 368.475 3069.035 368.755 ;
        RECT 3069.465 368.475 3069.745 368.755 ;
        RECT 3070.175 368.475 3070.455 368.755 ;
        RECT 3070.885 368.475 3071.165 368.755 ;
        RECT 3071.595 368.475 3071.875 368.755 ;
        RECT 3072.305 368.475 3072.585 368.755 ;
        RECT 3073.015 368.475 3073.295 368.755 ;
        RECT 526.715 367.765 526.995 368.045 ;
        RECT 527.425 367.765 527.705 368.045 ;
        RECT 528.135 367.765 528.415 368.045 ;
        RECT 528.845 367.765 529.125 368.045 ;
        RECT 529.555 367.765 529.835 368.045 ;
        RECT 530.265 367.765 530.545 368.045 ;
        RECT 530.975 367.765 531.255 368.045 ;
        RECT 531.685 367.765 531.965 368.045 ;
        RECT 532.395 367.765 532.675 368.045 ;
        RECT 533.105 367.765 533.385 368.045 ;
        RECT 533.815 367.765 534.095 368.045 ;
        RECT 534.525 367.765 534.805 368.045 ;
        RECT 535.235 367.765 535.515 368.045 ;
        RECT 544.975 367.765 545.255 368.045 ;
        RECT 545.685 367.765 545.965 368.045 ;
        RECT 546.395 367.765 546.675 368.045 ;
        RECT 547.105 367.765 547.385 368.045 ;
        RECT 547.815 367.765 548.095 368.045 ;
        RECT 548.525 367.765 548.805 368.045 ;
        RECT 550.965 367.765 551.245 368.045 ;
        RECT 551.675 367.765 551.955 368.045 ;
        RECT 552.385 367.765 552.665 368.045 ;
        RECT 553.095 367.765 553.375 368.045 ;
        RECT 553.805 367.765 554.085 368.045 ;
        RECT 554.515 367.765 554.795 368.045 ;
        RECT 555.225 367.765 555.505 368.045 ;
        RECT 555.935 367.765 556.215 368.045 ;
        RECT 556.645 367.765 556.925 368.045 ;
        RECT 557.355 367.765 557.635 368.045 ;
        RECT 558.065 367.765 558.345 368.045 ;
        RECT 558.775 367.765 559.055 368.045 ;
        RECT 559.485 367.765 559.765 368.045 ;
        RECT 560.195 367.765 560.475 368.045 ;
        RECT 566.625 367.765 566.905 368.045 ;
        RECT 567.335 367.765 567.615 368.045 ;
        RECT 568.045 367.765 568.325 368.045 ;
        RECT 568.755 367.765 569.035 368.045 ;
        RECT 569.465 367.765 569.745 368.045 ;
        RECT 570.175 367.765 570.455 368.045 ;
        RECT 570.885 367.765 571.165 368.045 ;
        RECT 571.595 367.765 571.875 368.045 ;
        RECT 572.305 367.765 572.585 368.045 ;
        RECT 573.015 367.765 573.295 368.045 ;
        RECT 573.725 367.765 574.005 368.045 ;
        RECT 576.345 367.765 576.625 368.045 ;
        RECT 577.055 367.765 577.335 368.045 ;
        RECT 577.765 367.765 578.045 368.045 ;
        RECT 578.475 367.765 578.755 368.045 ;
        RECT 579.185 367.765 579.465 368.045 ;
        RECT 579.895 367.765 580.175 368.045 ;
        RECT 580.605 367.765 580.885 368.045 ;
        RECT 581.315 367.765 581.595 368.045 ;
        RECT 582.025 367.765 582.305 368.045 ;
        RECT 582.735 367.765 583.015 368.045 ;
        RECT 583.445 367.765 583.725 368.045 ;
        RECT 584.155 367.765 584.435 368.045 ;
        RECT 584.865 367.765 585.145 368.045 ;
        RECT 585.575 367.765 585.855 368.045 ;
        RECT 589.495 367.765 589.775 368.045 ;
        RECT 590.205 367.765 590.485 368.045 ;
        RECT 590.915 367.765 591.195 368.045 ;
        RECT 591.625 367.765 591.905 368.045 ;
        RECT 592.335 367.765 592.615 368.045 ;
        RECT 593.045 367.765 593.325 368.045 ;
        RECT 593.755 367.765 594.035 368.045 ;
        RECT 594.465 367.765 594.745 368.045 ;
        RECT 595.175 367.765 595.455 368.045 ;
        RECT 595.885 367.765 596.165 368.045 ;
        RECT 596.595 367.765 596.875 368.045 ;
        RECT 597.305 367.765 597.585 368.045 ;
        RECT 598.015 367.765 598.295 368.045 ;
        RECT 1351.715 367.765 1351.995 368.045 ;
        RECT 1352.425 367.765 1352.705 368.045 ;
        RECT 1353.135 367.765 1353.415 368.045 ;
        RECT 1353.845 367.765 1354.125 368.045 ;
        RECT 1354.555 367.765 1354.835 368.045 ;
        RECT 1355.265 367.765 1355.545 368.045 ;
        RECT 1355.975 367.765 1356.255 368.045 ;
        RECT 1356.685 367.765 1356.965 368.045 ;
        RECT 1357.395 367.765 1357.675 368.045 ;
        RECT 1358.105 367.765 1358.385 368.045 ;
        RECT 1358.815 367.765 1359.095 368.045 ;
        RECT 1359.525 367.765 1359.805 368.045 ;
        RECT 1360.235 367.765 1360.515 368.045 ;
        RECT 1366.245 367.765 1366.525 368.045 ;
        RECT 1366.955 367.765 1367.235 368.045 ;
        RECT 1367.665 367.765 1367.945 368.045 ;
        RECT 1368.375 367.765 1368.655 368.045 ;
        RECT 1369.085 367.765 1369.365 368.045 ;
        RECT 1369.795 367.765 1370.075 368.045 ;
        RECT 1370.505 367.765 1370.785 368.045 ;
        RECT 1371.215 367.765 1371.495 368.045 ;
        RECT 1371.925 367.765 1372.205 368.045 ;
        RECT 1372.635 367.765 1372.915 368.045 ;
        RECT 1373.345 367.765 1373.625 368.045 ;
        RECT 1375.965 367.765 1376.245 368.045 ;
        RECT 1376.675 367.765 1376.955 368.045 ;
        RECT 1377.385 367.765 1377.665 368.045 ;
        RECT 1378.095 367.765 1378.375 368.045 ;
        RECT 1378.805 367.765 1379.085 368.045 ;
        RECT 1379.515 367.765 1379.795 368.045 ;
        RECT 1380.225 367.765 1380.505 368.045 ;
        RECT 1380.935 367.765 1381.215 368.045 ;
        RECT 1381.645 367.765 1381.925 368.045 ;
        RECT 1382.355 367.765 1382.635 368.045 ;
        RECT 1383.065 367.765 1383.345 368.045 ;
        RECT 1383.775 367.765 1384.055 368.045 ;
        RECT 1384.485 367.765 1384.765 368.045 ;
        RECT 1385.195 367.765 1385.475 368.045 ;
        RECT 1389.495 367.765 1389.775 368.045 ;
        RECT 1390.205 367.765 1390.485 368.045 ;
        RECT 1390.915 367.765 1391.195 368.045 ;
        RECT 1391.625 367.765 1391.905 368.045 ;
        RECT 1392.335 367.765 1392.615 368.045 ;
        RECT 1393.045 367.765 1393.325 368.045 ;
        RECT 1393.755 367.765 1394.035 368.045 ;
        RECT 1394.465 367.765 1394.745 368.045 ;
        RECT 1395.175 367.765 1395.455 368.045 ;
        RECT 1395.885 367.765 1396.165 368.045 ;
        RECT 1396.595 367.765 1396.875 368.045 ;
        RECT 1397.305 367.765 1397.585 368.045 ;
        RECT 1398.015 367.765 1398.295 368.045 ;
        RECT 1398.725 367.765 1399.005 368.045 ;
        RECT 1401.345 367.765 1401.625 368.045 ;
        RECT 1402.055 367.765 1402.335 368.045 ;
        RECT 1402.765 367.765 1403.045 368.045 ;
        RECT 1403.475 367.765 1403.755 368.045 ;
        RECT 1404.185 367.765 1404.465 368.045 ;
        RECT 1404.895 367.765 1405.175 368.045 ;
        RECT 1405.605 367.765 1405.885 368.045 ;
        RECT 1406.315 367.765 1406.595 368.045 ;
        RECT 1407.025 367.765 1407.305 368.045 ;
        RECT 1407.735 367.765 1408.015 368.045 ;
        RECT 1408.445 367.765 1408.725 368.045 ;
        RECT 1409.155 367.765 1409.435 368.045 ;
        RECT 1409.865 367.765 1410.145 368.045 ;
        RECT 1410.575 367.765 1410.855 368.045 ;
        RECT 1414.495 367.765 1414.775 368.045 ;
        RECT 1415.205 367.765 1415.485 368.045 ;
        RECT 1415.915 367.765 1416.195 368.045 ;
        RECT 1416.625 367.765 1416.905 368.045 ;
        RECT 1417.335 367.765 1417.615 368.045 ;
        RECT 1418.045 367.765 1418.325 368.045 ;
        RECT 1418.755 367.765 1419.035 368.045 ;
        RECT 1419.465 367.765 1419.745 368.045 ;
        RECT 3001.715 367.765 3001.995 368.045 ;
        RECT 3002.425 367.765 3002.705 368.045 ;
        RECT 3003.135 367.765 3003.415 368.045 ;
        RECT 3003.845 367.765 3004.125 368.045 ;
        RECT 3004.555 367.765 3004.835 368.045 ;
        RECT 3005.265 367.765 3005.545 368.045 ;
        RECT 3005.975 367.765 3006.255 368.045 ;
        RECT 3006.685 367.765 3006.965 368.045 ;
        RECT 3007.395 367.765 3007.675 368.045 ;
        RECT 3008.105 367.765 3008.385 368.045 ;
        RECT 3008.815 367.765 3009.095 368.045 ;
        RECT 3009.525 367.765 3009.805 368.045 ;
        RECT 3010.235 367.765 3010.515 368.045 ;
        RECT 3014.115 367.765 3014.395 368.045 ;
        RECT 3014.825 367.765 3015.105 368.045 ;
        RECT 3015.535 367.765 3015.815 368.045 ;
        RECT 3016.245 367.765 3016.525 368.045 ;
        RECT 3016.955 367.765 3017.235 368.045 ;
        RECT 3017.665 367.765 3017.945 368.045 ;
        RECT 3018.375 367.765 3018.655 368.045 ;
        RECT 3019.085 367.765 3019.365 368.045 ;
        RECT 3019.795 367.765 3020.075 368.045 ;
        RECT 3025.965 367.765 3026.245 368.045 ;
        RECT 3026.675 367.765 3026.955 368.045 ;
        RECT 3027.385 367.765 3027.665 368.045 ;
        RECT 3028.095 367.765 3028.375 368.045 ;
        RECT 3028.805 367.765 3029.085 368.045 ;
        RECT 3029.515 367.765 3029.795 368.045 ;
        RECT 3030.225 367.765 3030.505 368.045 ;
        RECT 3030.935 367.765 3031.215 368.045 ;
        RECT 3031.645 367.765 3031.925 368.045 ;
        RECT 3032.355 367.765 3032.635 368.045 ;
        RECT 3033.065 367.765 3033.345 368.045 ;
        RECT 3033.775 367.765 3034.055 368.045 ;
        RECT 3034.485 367.765 3034.765 368.045 ;
        RECT 3035.195 367.765 3035.475 368.045 ;
        RECT 3039.495 367.765 3039.775 368.045 ;
        RECT 3040.205 367.765 3040.485 368.045 ;
        RECT 3040.915 367.765 3041.195 368.045 ;
        RECT 3041.625 367.765 3041.905 368.045 ;
        RECT 3042.335 367.765 3042.615 368.045 ;
        RECT 3046.595 367.765 3046.875 368.045 ;
        RECT 3047.305 367.765 3047.585 368.045 ;
        RECT 3048.015 367.765 3048.295 368.045 ;
        RECT 3048.725 367.765 3049.005 368.045 ;
        RECT 3051.345 367.765 3051.625 368.045 ;
        RECT 3052.055 367.765 3052.335 368.045 ;
        RECT 3052.765 367.765 3053.045 368.045 ;
        RECT 3053.475 367.765 3053.755 368.045 ;
        RECT 3054.185 367.765 3054.465 368.045 ;
        RECT 3054.895 367.765 3055.175 368.045 ;
        RECT 3055.605 367.765 3055.885 368.045 ;
        RECT 3056.315 367.765 3056.595 368.045 ;
        RECT 3057.025 367.765 3057.305 368.045 ;
        RECT 3057.735 367.765 3058.015 368.045 ;
        RECT 3058.445 367.765 3058.725 368.045 ;
        RECT 3059.155 367.765 3059.435 368.045 ;
        RECT 3059.865 367.765 3060.145 368.045 ;
        RECT 3060.575 367.765 3060.855 368.045 ;
        RECT 3064.495 367.765 3064.775 368.045 ;
        RECT 3065.205 367.765 3065.485 368.045 ;
        RECT 3065.915 367.765 3066.195 368.045 ;
        RECT 3066.625 367.765 3066.905 368.045 ;
        RECT 3067.335 367.765 3067.615 368.045 ;
        RECT 3068.045 367.765 3068.325 368.045 ;
        RECT 3068.755 367.765 3069.035 368.045 ;
        RECT 3069.465 367.765 3069.745 368.045 ;
        RECT 3070.175 367.765 3070.455 368.045 ;
        RECT 3070.885 367.765 3071.165 368.045 ;
        RECT 3071.595 367.765 3071.875 368.045 ;
        RECT 3072.305 367.765 3072.585 368.045 ;
        RECT 3073.015 367.765 3073.295 368.045 ;
        RECT 526.715 367.055 526.995 367.335 ;
        RECT 527.425 367.055 527.705 367.335 ;
        RECT 528.135 367.055 528.415 367.335 ;
        RECT 528.845 367.055 529.125 367.335 ;
        RECT 529.555 367.055 529.835 367.335 ;
        RECT 530.265 367.055 530.545 367.335 ;
        RECT 530.975 367.055 531.255 367.335 ;
        RECT 531.685 367.055 531.965 367.335 ;
        RECT 532.395 367.055 532.675 367.335 ;
        RECT 533.105 367.055 533.385 367.335 ;
        RECT 533.815 367.055 534.095 367.335 ;
        RECT 534.525 367.055 534.805 367.335 ;
        RECT 535.235 367.055 535.515 367.335 ;
        RECT 544.975 367.055 545.255 367.335 ;
        RECT 545.685 367.055 545.965 367.335 ;
        RECT 546.395 367.055 546.675 367.335 ;
        RECT 547.105 367.055 547.385 367.335 ;
        RECT 547.815 367.055 548.095 367.335 ;
        RECT 548.525 367.055 548.805 367.335 ;
        RECT 550.965 367.055 551.245 367.335 ;
        RECT 551.675 367.055 551.955 367.335 ;
        RECT 552.385 367.055 552.665 367.335 ;
        RECT 553.095 367.055 553.375 367.335 ;
        RECT 553.805 367.055 554.085 367.335 ;
        RECT 554.515 367.055 554.795 367.335 ;
        RECT 555.225 367.055 555.505 367.335 ;
        RECT 555.935 367.055 556.215 367.335 ;
        RECT 556.645 367.055 556.925 367.335 ;
        RECT 557.355 367.055 557.635 367.335 ;
        RECT 558.065 367.055 558.345 367.335 ;
        RECT 558.775 367.055 559.055 367.335 ;
        RECT 559.485 367.055 559.765 367.335 ;
        RECT 560.195 367.055 560.475 367.335 ;
        RECT 566.625 367.055 566.905 367.335 ;
        RECT 567.335 367.055 567.615 367.335 ;
        RECT 568.045 367.055 568.325 367.335 ;
        RECT 568.755 367.055 569.035 367.335 ;
        RECT 569.465 367.055 569.745 367.335 ;
        RECT 570.175 367.055 570.455 367.335 ;
        RECT 570.885 367.055 571.165 367.335 ;
        RECT 571.595 367.055 571.875 367.335 ;
        RECT 572.305 367.055 572.585 367.335 ;
        RECT 573.015 367.055 573.295 367.335 ;
        RECT 573.725 367.055 574.005 367.335 ;
        RECT 576.345 367.055 576.625 367.335 ;
        RECT 577.055 367.055 577.335 367.335 ;
        RECT 577.765 367.055 578.045 367.335 ;
        RECT 578.475 367.055 578.755 367.335 ;
        RECT 579.185 367.055 579.465 367.335 ;
        RECT 579.895 367.055 580.175 367.335 ;
        RECT 580.605 367.055 580.885 367.335 ;
        RECT 581.315 367.055 581.595 367.335 ;
        RECT 582.025 367.055 582.305 367.335 ;
        RECT 582.735 367.055 583.015 367.335 ;
        RECT 583.445 367.055 583.725 367.335 ;
        RECT 584.155 367.055 584.435 367.335 ;
        RECT 584.865 367.055 585.145 367.335 ;
        RECT 585.575 367.055 585.855 367.335 ;
        RECT 589.495 367.055 589.775 367.335 ;
        RECT 590.205 367.055 590.485 367.335 ;
        RECT 590.915 367.055 591.195 367.335 ;
        RECT 591.625 367.055 591.905 367.335 ;
        RECT 592.335 367.055 592.615 367.335 ;
        RECT 593.045 367.055 593.325 367.335 ;
        RECT 593.755 367.055 594.035 367.335 ;
        RECT 594.465 367.055 594.745 367.335 ;
        RECT 595.175 367.055 595.455 367.335 ;
        RECT 595.885 367.055 596.165 367.335 ;
        RECT 596.595 367.055 596.875 367.335 ;
        RECT 597.305 367.055 597.585 367.335 ;
        RECT 598.015 367.055 598.295 367.335 ;
        RECT 1351.715 367.055 1351.995 367.335 ;
        RECT 1352.425 367.055 1352.705 367.335 ;
        RECT 1353.135 367.055 1353.415 367.335 ;
        RECT 1353.845 367.055 1354.125 367.335 ;
        RECT 1354.555 367.055 1354.835 367.335 ;
        RECT 1355.265 367.055 1355.545 367.335 ;
        RECT 1355.975 367.055 1356.255 367.335 ;
        RECT 1356.685 367.055 1356.965 367.335 ;
        RECT 1357.395 367.055 1357.675 367.335 ;
        RECT 1358.105 367.055 1358.385 367.335 ;
        RECT 1358.815 367.055 1359.095 367.335 ;
        RECT 1359.525 367.055 1359.805 367.335 ;
        RECT 1360.235 367.055 1360.515 367.335 ;
        RECT 1366.245 367.055 1366.525 367.335 ;
        RECT 1366.955 367.055 1367.235 367.335 ;
        RECT 1367.665 367.055 1367.945 367.335 ;
        RECT 1368.375 367.055 1368.655 367.335 ;
        RECT 1369.085 367.055 1369.365 367.335 ;
        RECT 1369.795 367.055 1370.075 367.335 ;
        RECT 1370.505 367.055 1370.785 367.335 ;
        RECT 1371.215 367.055 1371.495 367.335 ;
        RECT 1371.925 367.055 1372.205 367.335 ;
        RECT 1372.635 367.055 1372.915 367.335 ;
        RECT 1373.345 367.055 1373.625 367.335 ;
        RECT 1375.965 367.055 1376.245 367.335 ;
        RECT 1376.675 367.055 1376.955 367.335 ;
        RECT 1377.385 367.055 1377.665 367.335 ;
        RECT 1378.095 367.055 1378.375 367.335 ;
        RECT 1378.805 367.055 1379.085 367.335 ;
        RECT 1379.515 367.055 1379.795 367.335 ;
        RECT 1380.225 367.055 1380.505 367.335 ;
        RECT 1380.935 367.055 1381.215 367.335 ;
        RECT 1381.645 367.055 1381.925 367.335 ;
        RECT 1382.355 367.055 1382.635 367.335 ;
        RECT 1383.065 367.055 1383.345 367.335 ;
        RECT 1383.775 367.055 1384.055 367.335 ;
        RECT 1384.485 367.055 1384.765 367.335 ;
        RECT 1385.195 367.055 1385.475 367.335 ;
        RECT 1389.495 367.055 1389.775 367.335 ;
        RECT 1390.205 367.055 1390.485 367.335 ;
        RECT 1390.915 367.055 1391.195 367.335 ;
        RECT 1391.625 367.055 1391.905 367.335 ;
        RECT 1392.335 367.055 1392.615 367.335 ;
        RECT 1393.045 367.055 1393.325 367.335 ;
        RECT 1393.755 367.055 1394.035 367.335 ;
        RECT 1394.465 367.055 1394.745 367.335 ;
        RECT 1395.175 367.055 1395.455 367.335 ;
        RECT 1395.885 367.055 1396.165 367.335 ;
        RECT 1396.595 367.055 1396.875 367.335 ;
        RECT 1397.305 367.055 1397.585 367.335 ;
        RECT 1398.015 367.055 1398.295 367.335 ;
        RECT 1398.725 367.055 1399.005 367.335 ;
        RECT 1401.345 367.055 1401.625 367.335 ;
        RECT 1402.055 367.055 1402.335 367.335 ;
        RECT 1402.765 367.055 1403.045 367.335 ;
        RECT 1403.475 367.055 1403.755 367.335 ;
        RECT 1404.185 367.055 1404.465 367.335 ;
        RECT 1404.895 367.055 1405.175 367.335 ;
        RECT 1405.605 367.055 1405.885 367.335 ;
        RECT 1406.315 367.055 1406.595 367.335 ;
        RECT 1407.025 367.055 1407.305 367.335 ;
        RECT 1407.735 367.055 1408.015 367.335 ;
        RECT 1408.445 367.055 1408.725 367.335 ;
        RECT 1409.155 367.055 1409.435 367.335 ;
        RECT 1409.865 367.055 1410.145 367.335 ;
        RECT 1410.575 367.055 1410.855 367.335 ;
        RECT 1414.495 367.055 1414.775 367.335 ;
        RECT 1415.205 367.055 1415.485 367.335 ;
        RECT 1415.915 367.055 1416.195 367.335 ;
        RECT 1416.625 367.055 1416.905 367.335 ;
        RECT 1417.335 367.055 1417.615 367.335 ;
        RECT 1418.045 367.055 1418.325 367.335 ;
        RECT 1418.755 367.055 1419.035 367.335 ;
        RECT 1419.465 367.055 1419.745 367.335 ;
        RECT 3001.715 367.055 3001.995 367.335 ;
        RECT 3002.425 367.055 3002.705 367.335 ;
        RECT 3003.135 367.055 3003.415 367.335 ;
        RECT 3003.845 367.055 3004.125 367.335 ;
        RECT 3004.555 367.055 3004.835 367.335 ;
        RECT 3005.265 367.055 3005.545 367.335 ;
        RECT 3005.975 367.055 3006.255 367.335 ;
        RECT 3006.685 367.055 3006.965 367.335 ;
        RECT 3007.395 367.055 3007.675 367.335 ;
        RECT 3008.105 367.055 3008.385 367.335 ;
        RECT 3008.815 367.055 3009.095 367.335 ;
        RECT 3009.525 367.055 3009.805 367.335 ;
        RECT 3010.235 367.055 3010.515 367.335 ;
        RECT 3014.115 367.055 3014.395 367.335 ;
        RECT 3014.825 367.055 3015.105 367.335 ;
        RECT 3015.535 367.055 3015.815 367.335 ;
        RECT 3016.245 367.055 3016.525 367.335 ;
        RECT 3016.955 367.055 3017.235 367.335 ;
        RECT 3017.665 367.055 3017.945 367.335 ;
        RECT 3018.375 367.055 3018.655 367.335 ;
        RECT 3019.085 367.055 3019.365 367.335 ;
        RECT 3019.795 367.055 3020.075 367.335 ;
        RECT 3025.965 367.055 3026.245 367.335 ;
        RECT 3026.675 367.055 3026.955 367.335 ;
        RECT 3027.385 367.055 3027.665 367.335 ;
        RECT 3028.095 367.055 3028.375 367.335 ;
        RECT 3028.805 367.055 3029.085 367.335 ;
        RECT 3029.515 367.055 3029.795 367.335 ;
        RECT 3030.225 367.055 3030.505 367.335 ;
        RECT 3030.935 367.055 3031.215 367.335 ;
        RECT 3031.645 367.055 3031.925 367.335 ;
        RECT 3032.355 367.055 3032.635 367.335 ;
        RECT 3033.065 367.055 3033.345 367.335 ;
        RECT 3033.775 367.055 3034.055 367.335 ;
        RECT 3034.485 367.055 3034.765 367.335 ;
        RECT 3035.195 367.055 3035.475 367.335 ;
        RECT 3039.495 367.055 3039.775 367.335 ;
        RECT 3040.205 367.055 3040.485 367.335 ;
        RECT 3040.915 367.055 3041.195 367.335 ;
        RECT 3041.625 367.055 3041.905 367.335 ;
        RECT 3042.335 367.055 3042.615 367.335 ;
        RECT 3046.595 367.055 3046.875 367.335 ;
        RECT 3047.305 367.055 3047.585 367.335 ;
        RECT 3048.015 367.055 3048.295 367.335 ;
        RECT 3048.725 367.055 3049.005 367.335 ;
        RECT 3051.345 367.055 3051.625 367.335 ;
        RECT 3052.055 367.055 3052.335 367.335 ;
        RECT 3052.765 367.055 3053.045 367.335 ;
        RECT 3053.475 367.055 3053.755 367.335 ;
        RECT 3054.185 367.055 3054.465 367.335 ;
        RECT 3054.895 367.055 3055.175 367.335 ;
        RECT 3055.605 367.055 3055.885 367.335 ;
        RECT 3056.315 367.055 3056.595 367.335 ;
        RECT 3057.025 367.055 3057.305 367.335 ;
        RECT 3057.735 367.055 3058.015 367.335 ;
        RECT 3058.445 367.055 3058.725 367.335 ;
        RECT 3059.155 367.055 3059.435 367.335 ;
        RECT 3059.865 367.055 3060.145 367.335 ;
        RECT 3060.575 367.055 3060.855 367.335 ;
        RECT 3064.495 367.055 3064.775 367.335 ;
        RECT 3065.205 367.055 3065.485 367.335 ;
        RECT 3065.915 367.055 3066.195 367.335 ;
        RECT 3066.625 367.055 3066.905 367.335 ;
        RECT 3067.335 367.055 3067.615 367.335 ;
        RECT 3068.045 367.055 3068.325 367.335 ;
        RECT 3068.755 367.055 3069.035 367.335 ;
        RECT 3069.465 367.055 3069.745 367.335 ;
        RECT 3070.175 367.055 3070.455 367.335 ;
        RECT 3070.885 367.055 3071.165 367.335 ;
        RECT 3071.595 367.055 3071.875 367.335 ;
        RECT 3072.305 367.055 3072.585 367.335 ;
        RECT 3073.015 367.055 3073.295 367.335 ;
        RECT 526.715 366.345 526.995 366.625 ;
        RECT 527.425 366.345 527.705 366.625 ;
        RECT 528.135 366.345 528.415 366.625 ;
        RECT 528.845 366.345 529.125 366.625 ;
        RECT 529.555 366.345 529.835 366.625 ;
        RECT 530.265 366.345 530.545 366.625 ;
        RECT 530.975 366.345 531.255 366.625 ;
        RECT 531.685 366.345 531.965 366.625 ;
        RECT 532.395 366.345 532.675 366.625 ;
        RECT 533.105 366.345 533.385 366.625 ;
        RECT 533.815 366.345 534.095 366.625 ;
        RECT 534.525 366.345 534.805 366.625 ;
        RECT 535.235 366.345 535.515 366.625 ;
        RECT 544.975 366.345 545.255 366.625 ;
        RECT 545.685 366.345 545.965 366.625 ;
        RECT 546.395 366.345 546.675 366.625 ;
        RECT 547.105 366.345 547.385 366.625 ;
        RECT 547.815 366.345 548.095 366.625 ;
        RECT 548.525 366.345 548.805 366.625 ;
        RECT 550.965 366.345 551.245 366.625 ;
        RECT 551.675 366.345 551.955 366.625 ;
        RECT 552.385 366.345 552.665 366.625 ;
        RECT 553.095 366.345 553.375 366.625 ;
        RECT 553.805 366.345 554.085 366.625 ;
        RECT 554.515 366.345 554.795 366.625 ;
        RECT 555.225 366.345 555.505 366.625 ;
        RECT 555.935 366.345 556.215 366.625 ;
        RECT 556.645 366.345 556.925 366.625 ;
        RECT 557.355 366.345 557.635 366.625 ;
        RECT 558.065 366.345 558.345 366.625 ;
        RECT 558.775 366.345 559.055 366.625 ;
        RECT 559.485 366.345 559.765 366.625 ;
        RECT 560.195 366.345 560.475 366.625 ;
        RECT 566.625 366.345 566.905 366.625 ;
        RECT 567.335 366.345 567.615 366.625 ;
        RECT 568.045 366.345 568.325 366.625 ;
        RECT 568.755 366.345 569.035 366.625 ;
        RECT 569.465 366.345 569.745 366.625 ;
        RECT 570.175 366.345 570.455 366.625 ;
        RECT 570.885 366.345 571.165 366.625 ;
        RECT 571.595 366.345 571.875 366.625 ;
        RECT 572.305 366.345 572.585 366.625 ;
        RECT 573.015 366.345 573.295 366.625 ;
        RECT 573.725 366.345 574.005 366.625 ;
        RECT 576.345 366.345 576.625 366.625 ;
        RECT 577.055 366.345 577.335 366.625 ;
        RECT 577.765 366.345 578.045 366.625 ;
        RECT 578.475 366.345 578.755 366.625 ;
        RECT 579.185 366.345 579.465 366.625 ;
        RECT 579.895 366.345 580.175 366.625 ;
        RECT 580.605 366.345 580.885 366.625 ;
        RECT 581.315 366.345 581.595 366.625 ;
        RECT 582.025 366.345 582.305 366.625 ;
        RECT 582.735 366.345 583.015 366.625 ;
        RECT 583.445 366.345 583.725 366.625 ;
        RECT 584.155 366.345 584.435 366.625 ;
        RECT 584.865 366.345 585.145 366.625 ;
        RECT 585.575 366.345 585.855 366.625 ;
        RECT 589.495 366.345 589.775 366.625 ;
        RECT 590.205 366.345 590.485 366.625 ;
        RECT 590.915 366.345 591.195 366.625 ;
        RECT 591.625 366.345 591.905 366.625 ;
        RECT 592.335 366.345 592.615 366.625 ;
        RECT 593.045 366.345 593.325 366.625 ;
        RECT 593.755 366.345 594.035 366.625 ;
        RECT 594.465 366.345 594.745 366.625 ;
        RECT 595.175 366.345 595.455 366.625 ;
        RECT 595.885 366.345 596.165 366.625 ;
        RECT 596.595 366.345 596.875 366.625 ;
        RECT 597.305 366.345 597.585 366.625 ;
        RECT 598.015 366.345 598.295 366.625 ;
        RECT 1351.715 366.345 1351.995 366.625 ;
        RECT 1352.425 366.345 1352.705 366.625 ;
        RECT 1353.135 366.345 1353.415 366.625 ;
        RECT 1353.845 366.345 1354.125 366.625 ;
        RECT 1354.555 366.345 1354.835 366.625 ;
        RECT 1355.265 366.345 1355.545 366.625 ;
        RECT 1355.975 366.345 1356.255 366.625 ;
        RECT 1356.685 366.345 1356.965 366.625 ;
        RECT 1357.395 366.345 1357.675 366.625 ;
        RECT 1358.105 366.345 1358.385 366.625 ;
        RECT 1358.815 366.345 1359.095 366.625 ;
        RECT 1359.525 366.345 1359.805 366.625 ;
        RECT 1360.235 366.345 1360.515 366.625 ;
        RECT 1366.245 366.345 1366.525 366.625 ;
        RECT 1366.955 366.345 1367.235 366.625 ;
        RECT 1367.665 366.345 1367.945 366.625 ;
        RECT 1368.375 366.345 1368.655 366.625 ;
        RECT 1369.085 366.345 1369.365 366.625 ;
        RECT 1369.795 366.345 1370.075 366.625 ;
        RECT 1370.505 366.345 1370.785 366.625 ;
        RECT 1371.215 366.345 1371.495 366.625 ;
        RECT 1371.925 366.345 1372.205 366.625 ;
        RECT 1372.635 366.345 1372.915 366.625 ;
        RECT 1373.345 366.345 1373.625 366.625 ;
        RECT 1375.965 366.345 1376.245 366.625 ;
        RECT 1376.675 366.345 1376.955 366.625 ;
        RECT 1377.385 366.345 1377.665 366.625 ;
        RECT 1378.095 366.345 1378.375 366.625 ;
        RECT 1378.805 366.345 1379.085 366.625 ;
        RECT 1379.515 366.345 1379.795 366.625 ;
        RECT 1380.225 366.345 1380.505 366.625 ;
        RECT 1380.935 366.345 1381.215 366.625 ;
        RECT 1381.645 366.345 1381.925 366.625 ;
        RECT 1382.355 366.345 1382.635 366.625 ;
        RECT 1383.065 366.345 1383.345 366.625 ;
        RECT 1383.775 366.345 1384.055 366.625 ;
        RECT 1384.485 366.345 1384.765 366.625 ;
        RECT 1385.195 366.345 1385.475 366.625 ;
        RECT 1389.495 366.345 1389.775 366.625 ;
        RECT 1390.205 366.345 1390.485 366.625 ;
        RECT 1390.915 366.345 1391.195 366.625 ;
        RECT 1391.625 366.345 1391.905 366.625 ;
        RECT 1392.335 366.345 1392.615 366.625 ;
        RECT 1393.045 366.345 1393.325 366.625 ;
        RECT 1393.755 366.345 1394.035 366.625 ;
        RECT 1394.465 366.345 1394.745 366.625 ;
        RECT 1395.175 366.345 1395.455 366.625 ;
        RECT 1395.885 366.345 1396.165 366.625 ;
        RECT 1396.595 366.345 1396.875 366.625 ;
        RECT 1397.305 366.345 1397.585 366.625 ;
        RECT 1398.015 366.345 1398.295 366.625 ;
        RECT 1398.725 366.345 1399.005 366.625 ;
        RECT 1401.345 366.345 1401.625 366.625 ;
        RECT 1402.055 366.345 1402.335 366.625 ;
        RECT 1402.765 366.345 1403.045 366.625 ;
        RECT 1403.475 366.345 1403.755 366.625 ;
        RECT 1404.185 366.345 1404.465 366.625 ;
        RECT 1404.895 366.345 1405.175 366.625 ;
        RECT 1405.605 366.345 1405.885 366.625 ;
        RECT 1406.315 366.345 1406.595 366.625 ;
        RECT 1407.025 366.345 1407.305 366.625 ;
        RECT 1407.735 366.345 1408.015 366.625 ;
        RECT 1408.445 366.345 1408.725 366.625 ;
        RECT 1409.155 366.345 1409.435 366.625 ;
        RECT 1409.865 366.345 1410.145 366.625 ;
        RECT 1410.575 366.345 1410.855 366.625 ;
        RECT 1414.495 366.345 1414.775 366.625 ;
        RECT 1415.205 366.345 1415.485 366.625 ;
        RECT 1415.915 366.345 1416.195 366.625 ;
        RECT 1416.625 366.345 1416.905 366.625 ;
        RECT 1417.335 366.345 1417.615 366.625 ;
        RECT 1418.045 366.345 1418.325 366.625 ;
        RECT 1418.755 366.345 1419.035 366.625 ;
        RECT 1419.465 366.345 1419.745 366.625 ;
        RECT 3001.715 366.345 3001.995 366.625 ;
        RECT 3002.425 366.345 3002.705 366.625 ;
        RECT 3003.135 366.345 3003.415 366.625 ;
        RECT 3003.845 366.345 3004.125 366.625 ;
        RECT 3004.555 366.345 3004.835 366.625 ;
        RECT 3005.265 366.345 3005.545 366.625 ;
        RECT 3005.975 366.345 3006.255 366.625 ;
        RECT 3006.685 366.345 3006.965 366.625 ;
        RECT 3007.395 366.345 3007.675 366.625 ;
        RECT 3008.105 366.345 3008.385 366.625 ;
        RECT 3008.815 366.345 3009.095 366.625 ;
        RECT 3009.525 366.345 3009.805 366.625 ;
        RECT 3010.235 366.345 3010.515 366.625 ;
        RECT 3014.115 366.345 3014.395 366.625 ;
        RECT 3014.825 366.345 3015.105 366.625 ;
        RECT 3015.535 366.345 3015.815 366.625 ;
        RECT 3016.245 366.345 3016.525 366.625 ;
        RECT 3016.955 366.345 3017.235 366.625 ;
        RECT 3017.665 366.345 3017.945 366.625 ;
        RECT 3018.375 366.345 3018.655 366.625 ;
        RECT 3019.085 366.345 3019.365 366.625 ;
        RECT 3019.795 366.345 3020.075 366.625 ;
        RECT 3025.965 366.345 3026.245 366.625 ;
        RECT 3026.675 366.345 3026.955 366.625 ;
        RECT 3027.385 366.345 3027.665 366.625 ;
        RECT 3028.095 366.345 3028.375 366.625 ;
        RECT 3028.805 366.345 3029.085 366.625 ;
        RECT 3029.515 366.345 3029.795 366.625 ;
        RECT 3030.225 366.345 3030.505 366.625 ;
        RECT 3030.935 366.345 3031.215 366.625 ;
        RECT 3031.645 366.345 3031.925 366.625 ;
        RECT 3032.355 366.345 3032.635 366.625 ;
        RECT 3033.065 366.345 3033.345 366.625 ;
        RECT 3033.775 366.345 3034.055 366.625 ;
        RECT 3034.485 366.345 3034.765 366.625 ;
        RECT 3035.195 366.345 3035.475 366.625 ;
        RECT 3039.495 366.345 3039.775 366.625 ;
        RECT 3040.205 366.345 3040.485 366.625 ;
        RECT 3040.915 366.345 3041.195 366.625 ;
        RECT 3041.625 366.345 3041.905 366.625 ;
        RECT 3042.335 366.345 3042.615 366.625 ;
        RECT 3046.595 366.345 3046.875 366.625 ;
        RECT 3047.305 366.345 3047.585 366.625 ;
        RECT 3048.015 366.345 3048.295 366.625 ;
        RECT 3048.725 366.345 3049.005 366.625 ;
        RECT 3051.345 366.345 3051.625 366.625 ;
        RECT 3052.055 366.345 3052.335 366.625 ;
        RECT 3052.765 366.345 3053.045 366.625 ;
        RECT 3053.475 366.345 3053.755 366.625 ;
        RECT 3054.185 366.345 3054.465 366.625 ;
        RECT 3054.895 366.345 3055.175 366.625 ;
        RECT 3055.605 366.345 3055.885 366.625 ;
        RECT 3056.315 366.345 3056.595 366.625 ;
        RECT 3057.025 366.345 3057.305 366.625 ;
        RECT 3057.735 366.345 3058.015 366.625 ;
        RECT 3058.445 366.345 3058.725 366.625 ;
        RECT 3059.155 366.345 3059.435 366.625 ;
        RECT 3059.865 366.345 3060.145 366.625 ;
        RECT 3060.575 366.345 3060.855 366.625 ;
        RECT 3064.495 366.345 3064.775 366.625 ;
        RECT 3065.205 366.345 3065.485 366.625 ;
        RECT 3065.915 366.345 3066.195 366.625 ;
        RECT 3066.625 366.345 3066.905 366.625 ;
        RECT 3067.335 366.345 3067.615 366.625 ;
        RECT 3068.045 366.345 3068.325 366.625 ;
        RECT 3068.755 366.345 3069.035 366.625 ;
        RECT 3069.465 366.345 3069.745 366.625 ;
        RECT 3070.175 366.345 3070.455 366.625 ;
        RECT 3070.885 366.345 3071.165 366.625 ;
        RECT 3071.595 366.345 3071.875 366.625 ;
        RECT 3072.305 366.345 3072.585 366.625 ;
        RECT 3073.015 366.345 3073.295 366.625 ;
        RECT 526.715 365.635 526.995 365.915 ;
        RECT 527.425 365.635 527.705 365.915 ;
        RECT 528.135 365.635 528.415 365.915 ;
        RECT 528.845 365.635 529.125 365.915 ;
        RECT 529.555 365.635 529.835 365.915 ;
        RECT 530.265 365.635 530.545 365.915 ;
        RECT 530.975 365.635 531.255 365.915 ;
        RECT 531.685 365.635 531.965 365.915 ;
        RECT 532.395 365.635 532.675 365.915 ;
        RECT 533.105 365.635 533.385 365.915 ;
        RECT 533.815 365.635 534.095 365.915 ;
        RECT 534.525 365.635 534.805 365.915 ;
        RECT 535.235 365.635 535.515 365.915 ;
        RECT 544.975 365.635 545.255 365.915 ;
        RECT 545.685 365.635 545.965 365.915 ;
        RECT 546.395 365.635 546.675 365.915 ;
        RECT 547.105 365.635 547.385 365.915 ;
        RECT 547.815 365.635 548.095 365.915 ;
        RECT 548.525 365.635 548.805 365.915 ;
        RECT 550.965 365.635 551.245 365.915 ;
        RECT 551.675 365.635 551.955 365.915 ;
        RECT 552.385 365.635 552.665 365.915 ;
        RECT 553.095 365.635 553.375 365.915 ;
        RECT 553.805 365.635 554.085 365.915 ;
        RECT 554.515 365.635 554.795 365.915 ;
        RECT 555.225 365.635 555.505 365.915 ;
        RECT 555.935 365.635 556.215 365.915 ;
        RECT 556.645 365.635 556.925 365.915 ;
        RECT 557.355 365.635 557.635 365.915 ;
        RECT 558.065 365.635 558.345 365.915 ;
        RECT 558.775 365.635 559.055 365.915 ;
        RECT 559.485 365.635 559.765 365.915 ;
        RECT 560.195 365.635 560.475 365.915 ;
        RECT 566.625 365.635 566.905 365.915 ;
        RECT 567.335 365.635 567.615 365.915 ;
        RECT 568.045 365.635 568.325 365.915 ;
        RECT 568.755 365.635 569.035 365.915 ;
        RECT 569.465 365.635 569.745 365.915 ;
        RECT 570.175 365.635 570.455 365.915 ;
        RECT 570.885 365.635 571.165 365.915 ;
        RECT 571.595 365.635 571.875 365.915 ;
        RECT 572.305 365.635 572.585 365.915 ;
        RECT 573.015 365.635 573.295 365.915 ;
        RECT 573.725 365.635 574.005 365.915 ;
        RECT 576.345 365.635 576.625 365.915 ;
        RECT 577.055 365.635 577.335 365.915 ;
        RECT 577.765 365.635 578.045 365.915 ;
        RECT 578.475 365.635 578.755 365.915 ;
        RECT 579.185 365.635 579.465 365.915 ;
        RECT 579.895 365.635 580.175 365.915 ;
        RECT 580.605 365.635 580.885 365.915 ;
        RECT 581.315 365.635 581.595 365.915 ;
        RECT 582.025 365.635 582.305 365.915 ;
        RECT 582.735 365.635 583.015 365.915 ;
        RECT 583.445 365.635 583.725 365.915 ;
        RECT 584.155 365.635 584.435 365.915 ;
        RECT 584.865 365.635 585.145 365.915 ;
        RECT 585.575 365.635 585.855 365.915 ;
        RECT 589.495 365.635 589.775 365.915 ;
        RECT 590.205 365.635 590.485 365.915 ;
        RECT 590.915 365.635 591.195 365.915 ;
        RECT 591.625 365.635 591.905 365.915 ;
        RECT 592.335 365.635 592.615 365.915 ;
        RECT 593.045 365.635 593.325 365.915 ;
        RECT 593.755 365.635 594.035 365.915 ;
        RECT 594.465 365.635 594.745 365.915 ;
        RECT 595.175 365.635 595.455 365.915 ;
        RECT 595.885 365.635 596.165 365.915 ;
        RECT 596.595 365.635 596.875 365.915 ;
        RECT 597.305 365.635 597.585 365.915 ;
        RECT 598.015 365.635 598.295 365.915 ;
        RECT 1351.715 365.635 1351.995 365.915 ;
        RECT 1352.425 365.635 1352.705 365.915 ;
        RECT 1353.135 365.635 1353.415 365.915 ;
        RECT 1353.845 365.635 1354.125 365.915 ;
        RECT 1354.555 365.635 1354.835 365.915 ;
        RECT 1355.265 365.635 1355.545 365.915 ;
        RECT 1355.975 365.635 1356.255 365.915 ;
        RECT 1356.685 365.635 1356.965 365.915 ;
        RECT 1357.395 365.635 1357.675 365.915 ;
        RECT 1358.105 365.635 1358.385 365.915 ;
        RECT 1358.815 365.635 1359.095 365.915 ;
        RECT 1359.525 365.635 1359.805 365.915 ;
        RECT 1360.235 365.635 1360.515 365.915 ;
        RECT 1366.245 365.635 1366.525 365.915 ;
        RECT 1366.955 365.635 1367.235 365.915 ;
        RECT 1367.665 365.635 1367.945 365.915 ;
        RECT 1368.375 365.635 1368.655 365.915 ;
        RECT 1369.085 365.635 1369.365 365.915 ;
        RECT 1369.795 365.635 1370.075 365.915 ;
        RECT 1370.505 365.635 1370.785 365.915 ;
        RECT 1371.215 365.635 1371.495 365.915 ;
        RECT 1371.925 365.635 1372.205 365.915 ;
        RECT 1372.635 365.635 1372.915 365.915 ;
        RECT 1373.345 365.635 1373.625 365.915 ;
        RECT 1375.965 365.635 1376.245 365.915 ;
        RECT 1376.675 365.635 1376.955 365.915 ;
        RECT 1377.385 365.635 1377.665 365.915 ;
        RECT 1378.095 365.635 1378.375 365.915 ;
        RECT 1378.805 365.635 1379.085 365.915 ;
        RECT 1379.515 365.635 1379.795 365.915 ;
        RECT 1380.225 365.635 1380.505 365.915 ;
        RECT 1380.935 365.635 1381.215 365.915 ;
        RECT 1381.645 365.635 1381.925 365.915 ;
        RECT 1382.355 365.635 1382.635 365.915 ;
        RECT 1383.065 365.635 1383.345 365.915 ;
        RECT 1383.775 365.635 1384.055 365.915 ;
        RECT 1384.485 365.635 1384.765 365.915 ;
        RECT 1385.195 365.635 1385.475 365.915 ;
        RECT 1389.495 365.635 1389.775 365.915 ;
        RECT 1390.205 365.635 1390.485 365.915 ;
        RECT 1390.915 365.635 1391.195 365.915 ;
        RECT 1391.625 365.635 1391.905 365.915 ;
        RECT 1392.335 365.635 1392.615 365.915 ;
        RECT 1393.045 365.635 1393.325 365.915 ;
        RECT 1393.755 365.635 1394.035 365.915 ;
        RECT 1394.465 365.635 1394.745 365.915 ;
        RECT 1395.175 365.635 1395.455 365.915 ;
        RECT 1395.885 365.635 1396.165 365.915 ;
        RECT 1396.595 365.635 1396.875 365.915 ;
        RECT 1397.305 365.635 1397.585 365.915 ;
        RECT 1398.015 365.635 1398.295 365.915 ;
        RECT 1398.725 365.635 1399.005 365.915 ;
        RECT 1401.345 365.635 1401.625 365.915 ;
        RECT 1402.055 365.635 1402.335 365.915 ;
        RECT 1402.765 365.635 1403.045 365.915 ;
        RECT 1403.475 365.635 1403.755 365.915 ;
        RECT 1404.185 365.635 1404.465 365.915 ;
        RECT 1404.895 365.635 1405.175 365.915 ;
        RECT 1405.605 365.635 1405.885 365.915 ;
        RECT 1406.315 365.635 1406.595 365.915 ;
        RECT 1407.025 365.635 1407.305 365.915 ;
        RECT 1407.735 365.635 1408.015 365.915 ;
        RECT 1408.445 365.635 1408.725 365.915 ;
        RECT 1409.155 365.635 1409.435 365.915 ;
        RECT 1409.865 365.635 1410.145 365.915 ;
        RECT 1410.575 365.635 1410.855 365.915 ;
        RECT 1414.495 365.635 1414.775 365.915 ;
        RECT 1415.205 365.635 1415.485 365.915 ;
        RECT 1415.915 365.635 1416.195 365.915 ;
        RECT 1416.625 365.635 1416.905 365.915 ;
        RECT 1417.335 365.635 1417.615 365.915 ;
        RECT 1418.045 365.635 1418.325 365.915 ;
        RECT 1418.755 365.635 1419.035 365.915 ;
        RECT 1419.465 365.635 1419.745 365.915 ;
        RECT 3001.715 365.635 3001.995 365.915 ;
        RECT 3002.425 365.635 3002.705 365.915 ;
        RECT 3003.135 365.635 3003.415 365.915 ;
        RECT 3003.845 365.635 3004.125 365.915 ;
        RECT 3004.555 365.635 3004.835 365.915 ;
        RECT 3005.265 365.635 3005.545 365.915 ;
        RECT 3005.975 365.635 3006.255 365.915 ;
        RECT 3006.685 365.635 3006.965 365.915 ;
        RECT 3007.395 365.635 3007.675 365.915 ;
        RECT 3008.105 365.635 3008.385 365.915 ;
        RECT 3008.815 365.635 3009.095 365.915 ;
        RECT 3009.525 365.635 3009.805 365.915 ;
        RECT 3010.235 365.635 3010.515 365.915 ;
        RECT 3014.115 365.635 3014.395 365.915 ;
        RECT 3014.825 365.635 3015.105 365.915 ;
        RECT 3015.535 365.635 3015.815 365.915 ;
        RECT 3016.245 365.635 3016.525 365.915 ;
        RECT 3016.955 365.635 3017.235 365.915 ;
        RECT 3017.665 365.635 3017.945 365.915 ;
        RECT 3018.375 365.635 3018.655 365.915 ;
        RECT 3019.085 365.635 3019.365 365.915 ;
        RECT 3019.795 365.635 3020.075 365.915 ;
        RECT 3025.965 365.635 3026.245 365.915 ;
        RECT 3026.675 365.635 3026.955 365.915 ;
        RECT 3027.385 365.635 3027.665 365.915 ;
        RECT 3028.095 365.635 3028.375 365.915 ;
        RECT 3028.805 365.635 3029.085 365.915 ;
        RECT 3029.515 365.635 3029.795 365.915 ;
        RECT 3030.225 365.635 3030.505 365.915 ;
        RECT 3030.935 365.635 3031.215 365.915 ;
        RECT 3031.645 365.635 3031.925 365.915 ;
        RECT 3032.355 365.635 3032.635 365.915 ;
        RECT 3033.065 365.635 3033.345 365.915 ;
        RECT 3033.775 365.635 3034.055 365.915 ;
        RECT 3034.485 365.635 3034.765 365.915 ;
        RECT 3035.195 365.635 3035.475 365.915 ;
        RECT 3039.495 365.635 3039.775 365.915 ;
        RECT 3040.205 365.635 3040.485 365.915 ;
        RECT 3040.915 365.635 3041.195 365.915 ;
        RECT 3041.625 365.635 3041.905 365.915 ;
        RECT 3042.335 365.635 3042.615 365.915 ;
        RECT 3046.595 365.635 3046.875 365.915 ;
        RECT 3047.305 365.635 3047.585 365.915 ;
        RECT 3048.015 365.635 3048.295 365.915 ;
        RECT 3048.725 365.635 3049.005 365.915 ;
        RECT 3051.345 365.635 3051.625 365.915 ;
        RECT 3052.055 365.635 3052.335 365.915 ;
        RECT 3052.765 365.635 3053.045 365.915 ;
        RECT 3053.475 365.635 3053.755 365.915 ;
        RECT 3054.185 365.635 3054.465 365.915 ;
        RECT 3054.895 365.635 3055.175 365.915 ;
        RECT 3055.605 365.635 3055.885 365.915 ;
        RECT 3056.315 365.635 3056.595 365.915 ;
        RECT 3057.025 365.635 3057.305 365.915 ;
        RECT 3057.735 365.635 3058.015 365.915 ;
        RECT 3058.445 365.635 3058.725 365.915 ;
        RECT 3059.155 365.635 3059.435 365.915 ;
        RECT 3059.865 365.635 3060.145 365.915 ;
        RECT 3060.575 365.635 3060.855 365.915 ;
        RECT 3064.495 365.635 3064.775 365.915 ;
        RECT 3065.205 365.635 3065.485 365.915 ;
        RECT 3065.915 365.635 3066.195 365.915 ;
        RECT 3066.625 365.635 3066.905 365.915 ;
        RECT 3067.335 365.635 3067.615 365.915 ;
        RECT 3068.045 365.635 3068.325 365.915 ;
        RECT 3068.755 365.635 3069.035 365.915 ;
        RECT 3069.465 365.635 3069.745 365.915 ;
        RECT 3070.175 365.635 3070.455 365.915 ;
        RECT 3070.885 365.635 3071.165 365.915 ;
        RECT 3071.595 365.635 3071.875 365.915 ;
        RECT 3072.305 365.635 3072.585 365.915 ;
        RECT 3073.015 365.635 3073.295 365.915 ;
        RECT 526.715 364.925 526.995 365.205 ;
        RECT 527.425 364.925 527.705 365.205 ;
        RECT 528.135 364.925 528.415 365.205 ;
        RECT 528.845 364.925 529.125 365.205 ;
        RECT 529.555 364.925 529.835 365.205 ;
        RECT 530.265 364.925 530.545 365.205 ;
        RECT 530.975 364.925 531.255 365.205 ;
        RECT 531.685 364.925 531.965 365.205 ;
        RECT 532.395 364.925 532.675 365.205 ;
        RECT 533.105 364.925 533.385 365.205 ;
        RECT 533.815 364.925 534.095 365.205 ;
        RECT 534.525 364.925 534.805 365.205 ;
        RECT 535.235 364.925 535.515 365.205 ;
        RECT 544.975 364.925 545.255 365.205 ;
        RECT 545.685 364.925 545.965 365.205 ;
        RECT 546.395 364.925 546.675 365.205 ;
        RECT 547.105 364.925 547.385 365.205 ;
        RECT 547.815 364.925 548.095 365.205 ;
        RECT 548.525 364.925 548.805 365.205 ;
        RECT 550.965 364.925 551.245 365.205 ;
        RECT 551.675 364.925 551.955 365.205 ;
        RECT 552.385 364.925 552.665 365.205 ;
        RECT 553.095 364.925 553.375 365.205 ;
        RECT 553.805 364.925 554.085 365.205 ;
        RECT 554.515 364.925 554.795 365.205 ;
        RECT 555.225 364.925 555.505 365.205 ;
        RECT 555.935 364.925 556.215 365.205 ;
        RECT 556.645 364.925 556.925 365.205 ;
        RECT 557.355 364.925 557.635 365.205 ;
        RECT 558.065 364.925 558.345 365.205 ;
        RECT 558.775 364.925 559.055 365.205 ;
        RECT 559.485 364.925 559.765 365.205 ;
        RECT 560.195 364.925 560.475 365.205 ;
        RECT 566.625 364.925 566.905 365.205 ;
        RECT 567.335 364.925 567.615 365.205 ;
        RECT 568.045 364.925 568.325 365.205 ;
        RECT 568.755 364.925 569.035 365.205 ;
        RECT 569.465 364.925 569.745 365.205 ;
        RECT 570.175 364.925 570.455 365.205 ;
        RECT 570.885 364.925 571.165 365.205 ;
        RECT 571.595 364.925 571.875 365.205 ;
        RECT 572.305 364.925 572.585 365.205 ;
        RECT 573.015 364.925 573.295 365.205 ;
        RECT 573.725 364.925 574.005 365.205 ;
        RECT 576.345 364.925 576.625 365.205 ;
        RECT 577.055 364.925 577.335 365.205 ;
        RECT 577.765 364.925 578.045 365.205 ;
        RECT 578.475 364.925 578.755 365.205 ;
        RECT 579.185 364.925 579.465 365.205 ;
        RECT 579.895 364.925 580.175 365.205 ;
        RECT 580.605 364.925 580.885 365.205 ;
        RECT 581.315 364.925 581.595 365.205 ;
        RECT 582.025 364.925 582.305 365.205 ;
        RECT 582.735 364.925 583.015 365.205 ;
        RECT 583.445 364.925 583.725 365.205 ;
        RECT 584.155 364.925 584.435 365.205 ;
        RECT 584.865 364.925 585.145 365.205 ;
        RECT 585.575 364.925 585.855 365.205 ;
        RECT 589.495 364.925 589.775 365.205 ;
        RECT 590.205 364.925 590.485 365.205 ;
        RECT 590.915 364.925 591.195 365.205 ;
        RECT 591.625 364.925 591.905 365.205 ;
        RECT 592.335 364.925 592.615 365.205 ;
        RECT 593.045 364.925 593.325 365.205 ;
        RECT 593.755 364.925 594.035 365.205 ;
        RECT 594.465 364.925 594.745 365.205 ;
        RECT 595.175 364.925 595.455 365.205 ;
        RECT 595.885 364.925 596.165 365.205 ;
        RECT 596.595 364.925 596.875 365.205 ;
        RECT 597.305 364.925 597.585 365.205 ;
        RECT 598.015 364.925 598.295 365.205 ;
        RECT 1351.715 364.925 1351.995 365.205 ;
        RECT 1352.425 364.925 1352.705 365.205 ;
        RECT 1353.135 364.925 1353.415 365.205 ;
        RECT 1353.845 364.925 1354.125 365.205 ;
        RECT 1354.555 364.925 1354.835 365.205 ;
        RECT 1355.265 364.925 1355.545 365.205 ;
        RECT 1355.975 364.925 1356.255 365.205 ;
        RECT 1356.685 364.925 1356.965 365.205 ;
        RECT 1357.395 364.925 1357.675 365.205 ;
        RECT 1358.105 364.925 1358.385 365.205 ;
        RECT 1358.815 364.925 1359.095 365.205 ;
        RECT 1359.525 364.925 1359.805 365.205 ;
        RECT 1360.235 364.925 1360.515 365.205 ;
        RECT 1366.245 364.925 1366.525 365.205 ;
        RECT 1366.955 364.925 1367.235 365.205 ;
        RECT 1367.665 364.925 1367.945 365.205 ;
        RECT 1368.375 364.925 1368.655 365.205 ;
        RECT 1369.085 364.925 1369.365 365.205 ;
        RECT 1369.795 364.925 1370.075 365.205 ;
        RECT 1370.505 364.925 1370.785 365.205 ;
        RECT 1371.215 364.925 1371.495 365.205 ;
        RECT 1371.925 364.925 1372.205 365.205 ;
        RECT 1372.635 364.925 1372.915 365.205 ;
        RECT 1373.345 364.925 1373.625 365.205 ;
        RECT 1375.965 364.925 1376.245 365.205 ;
        RECT 1376.675 364.925 1376.955 365.205 ;
        RECT 1377.385 364.925 1377.665 365.205 ;
        RECT 1378.095 364.925 1378.375 365.205 ;
        RECT 1378.805 364.925 1379.085 365.205 ;
        RECT 1379.515 364.925 1379.795 365.205 ;
        RECT 1380.225 364.925 1380.505 365.205 ;
        RECT 1380.935 364.925 1381.215 365.205 ;
        RECT 1381.645 364.925 1381.925 365.205 ;
        RECT 1382.355 364.925 1382.635 365.205 ;
        RECT 1383.065 364.925 1383.345 365.205 ;
        RECT 1383.775 364.925 1384.055 365.205 ;
        RECT 1384.485 364.925 1384.765 365.205 ;
        RECT 1385.195 364.925 1385.475 365.205 ;
        RECT 1389.495 364.925 1389.775 365.205 ;
        RECT 1390.205 364.925 1390.485 365.205 ;
        RECT 1390.915 364.925 1391.195 365.205 ;
        RECT 1391.625 364.925 1391.905 365.205 ;
        RECT 1392.335 364.925 1392.615 365.205 ;
        RECT 1393.045 364.925 1393.325 365.205 ;
        RECT 1393.755 364.925 1394.035 365.205 ;
        RECT 1394.465 364.925 1394.745 365.205 ;
        RECT 1395.175 364.925 1395.455 365.205 ;
        RECT 1395.885 364.925 1396.165 365.205 ;
        RECT 1396.595 364.925 1396.875 365.205 ;
        RECT 1397.305 364.925 1397.585 365.205 ;
        RECT 1398.015 364.925 1398.295 365.205 ;
        RECT 1398.725 364.925 1399.005 365.205 ;
        RECT 1401.345 364.925 1401.625 365.205 ;
        RECT 1402.055 364.925 1402.335 365.205 ;
        RECT 1402.765 364.925 1403.045 365.205 ;
        RECT 1403.475 364.925 1403.755 365.205 ;
        RECT 1404.185 364.925 1404.465 365.205 ;
        RECT 1404.895 364.925 1405.175 365.205 ;
        RECT 1405.605 364.925 1405.885 365.205 ;
        RECT 1406.315 364.925 1406.595 365.205 ;
        RECT 1407.025 364.925 1407.305 365.205 ;
        RECT 1407.735 364.925 1408.015 365.205 ;
        RECT 1408.445 364.925 1408.725 365.205 ;
        RECT 1409.155 364.925 1409.435 365.205 ;
        RECT 1409.865 364.925 1410.145 365.205 ;
        RECT 1410.575 364.925 1410.855 365.205 ;
        RECT 1414.495 364.925 1414.775 365.205 ;
        RECT 1415.205 364.925 1415.485 365.205 ;
        RECT 1415.915 364.925 1416.195 365.205 ;
        RECT 1416.625 364.925 1416.905 365.205 ;
        RECT 1417.335 364.925 1417.615 365.205 ;
        RECT 1418.045 364.925 1418.325 365.205 ;
        RECT 1418.755 364.925 1419.035 365.205 ;
        RECT 1419.465 364.925 1419.745 365.205 ;
        RECT 3001.715 364.925 3001.995 365.205 ;
        RECT 3002.425 364.925 3002.705 365.205 ;
        RECT 3003.135 364.925 3003.415 365.205 ;
        RECT 3003.845 364.925 3004.125 365.205 ;
        RECT 3004.555 364.925 3004.835 365.205 ;
        RECT 3005.265 364.925 3005.545 365.205 ;
        RECT 3005.975 364.925 3006.255 365.205 ;
        RECT 3006.685 364.925 3006.965 365.205 ;
        RECT 3007.395 364.925 3007.675 365.205 ;
        RECT 3008.105 364.925 3008.385 365.205 ;
        RECT 3008.815 364.925 3009.095 365.205 ;
        RECT 3009.525 364.925 3009.805 365.205 ;
        RECT 3010.235 364.925 3010.515 365.205 ;
        RECT 3014.115 364.925 3014.395 365.205 ;
        RECT 3014.825 364.925 3015.105 365.205 ;
        RECT 3015.535 364.925 3015.815 365.205 ;
        RECT 3016.245 364.925 3016.525 365.205 ;
        RECT 3016.955 364.925 3017.235 365.205 ;
        RECT 3017.665 364.925 3017.945 365.205 ;
        RECT 3018.375 364.925 3018.655 365.205 ;
        RECT 3019.085 364.925 3019.365 365.205 ;
        RECT 3019.795 364.925 3020.075 365.205 ;
        RECT 3025.965 364.925 3026.245 365.205 ;
        RECT 3026.675 364.925 3026.955 365.205 ;
        RECT 3027.385 364.925 3027.665 365.205 ;
        RECT 3028.095 364.925 3028.375 365.205 ;
        RECT 3028.805 364.925 3029.085 365.205 ;
        RECT 3029.515 364.925 3029.795 365.205 ;
        RECT 3030.225 364.925 3030.505 365.205 ;
        RECT 3030.935 364.925 3031.215 365.205 ;
        RECT 3031.645 364.925 3031.925 365.205 ;
        RECT 3032.355 364.925 3032.635 365.205 ;
        RECT 3033.065 364.925 3033.345 365.205 ;
        RECT 3033.775 364.925 3034.055 365.205 ;
        RECT 3034.485 364.925 3034.765 365.205 ;
        RECT 3035.195 364.925 3035.475 365.205 ;
        RECT 3039.495 364.925 3039.775 365.205 ;
        RECT 3040.205 364.925 3040.485 365.205 ;
        RECT 3040.915 364.925 3041.195 365.205 ;
        RECT 3041.625 364.925 3041.905 365.205 ;
        RECT 3042.335 364.925 3042.615 365.205 ;
        RECT 3046.595 364.925 3046.875 365.205 ;
        RECT 3047.305 364.925 3047.585 365.205 ;
        RECT 3048.015 364.925 3048.295 365.205 ;
        RECT 3048.725 364.925 3049.005 365.205 ;
        RECT 3051.345 364.925 3051.625 365.205 ;
        RECT 3052.055 364.925 3052.335 365.205 ;
        RECT 3052.765 364.925 3053.045 365.205 ;
        RECT 3053.475 364.925 3053.755 365.205 ;
        RECT 3054.185 364.925 3054.465 365.205 ;
        RECT 3054.895 364.925 3055.175 365.205 ;
        RECT 3055.605 364.925 3055.885 365.205 ;
        RECT 3056.315 364.925 3056.595 365.205 ;
        RECT 3057.025 364.925 3057.305 365.205 ;
        RECT 3057.735 364.925 3058.015 365.205 ;
        RECT 3058.445 364.925 3058.725 365.205 ;
        RECT 3059.155 364.925 3059.435 365.205 ;
        RECT 3059.865 364.925 3060.145 365.205 ;
        RECT 3060.575 364.925 3060.855 365.205 ;
        RECT 3064.495 364.925 3064.775 365.205 ;
        RECT 3065.205 364.925 3065.485 365.205 ;
        RECT 3065.915 364.925 3066.195 365.205 ;
        RECT 3066.625 364.925 3066.905 365.205 ;
        RECT 3067.335 364.925 3067.615 365.205 ;
        RECT 3068.045 364.925 3068.325 365.205 ;
        RECT 3068.755 364.925 3069.035 365.205 ;
        RECT 3069.465 364.925 3069.745 365.205 ;
        RECT 3070.175 364.925 3070.455 365.205 ;
        RECT 3070.885 364.925 3071.165 365.205 ;
        RECT 3071.595 364.925 3071.875 365.205 ;
        RECT 3072.305 364.925 3072.585 365.205 ;
        RECT 3073.015 364.925 3073.295 365.205 ;
        RECT 526.715 364.215 526.995 364.495 ;
        RECT 527.425 364.215 527.705 364.495 ;
        RECT 528.135 364.215 528.415 364.495 ;
        RECT 528.845 364.215 529.125 364.495 ;
        RECT 529.555 364.215 529.835 364.495 ;
        RECT 530.265 364.215 530.545 364.495 ;
        RECT 530.975 364.215 531.255 364.495 ;
        RECT 531.685 364.215 531.965 364.495 ;
        RECT 532.395 364.215 532.675 364.495 ;
        RECT 533.105 364.215 533.385 364.495 ;
        RECT 533.815 364.215 534.095 364.495 ;
        RECT 534.525 364.215 534.805 364.495 ;
        RECT 535.235 364.215 535.515 364.495 ;
        RECT 544.975 364.215 545.255 364.495 ;
        RECT 545.685 364.215 545.965 364.495 ;
        RECT 546.395 364.215 546.675 364.495 ;
        RECT 547.105 364.215 547.385 364.495 ;
        RECT 547.815 364.215 548.095 364.495 ;
        RECT 548.525 364.215 548.805 364.495 ;
        RECT 550.965 364.215 551.245 364.495 ;
        RECT 551.675 364.215 551.955 364.495 ;
        RECT 552.385 364.215 552.665 364.495 ;
        RECT 553.095 364.215 553.375 364.495 ;
        RECT 553.805 364.215 554.085 364.495 ;
        RECT 554.515 364.215 554.795 364.495 ;
        RECT 555.225 364.215 555.505 364.495 ;
        RECT 555.935 364.215 556.215 364.495 ;
        RECT 556.645 364.215 556.925 364.495 ;
        RECT 557.355 364.215 557.635 364.495 ;
        RECT 558.065 364.215 558.345 364.495 ;
        RECT 558.775 364.215 559.055 364.495 ;
        RECT 559.485 364.215 559.765 364.495 ;
        RECT 560.195 364.215 560.475 364.495 ;
        RECT 566.625 364.215 566.905 364.495 ;
        RECT 567.335 364.215 567.615 364.495 ;
        RECT 568.045 364.215 568.325 364.495 ;
        RECT 568.755 364.215 569.035 364.495 ;
        RECT 569.465 364.215 569.745 364.495 ;
        RECT 570.175 364.215 570.455 364.495 ;
        RECT 570.885 364.215 571.165 364.495 ;
        RECT 571.595 364.215 571.875 364.495 ;
        RECT 572.305 364.215 572.585 364.495 ;
        RECT 573.015 364.215 573.295 364.495 ;
        RECT 573.725 364.215 574.005 364.495 ;
        RECT 576.345 364.215 576.625 364.495 ;
        RECT 577.055 364.215 577.335 364.495 ;
        RECT 577.765 364.215 578.045 364.495 ;
        RECT 578.475 364.215 578.755 364.495 ;
        RECT 579.185 364.215 579.465 364.495 ;
        RECT 579.895 364.215 580.175 364.495 ;
        RECT 580.605 364.215 580.885 364.495 ;
        RECT 581.315 364.215 581.595 364.495 ;
        RECT 582.025 364.215 582.305 364.495 ;
        RECT 582.735 364.215 583.015 364.495 ;
        RECT 583.445 364.215 583.725 364.495 ;
        RECT 584.155 364.215 584.435 364.495 ;
        RECT 584.865 364.215 585.145 364.495 ;
        RECT 585.575 364.215 585.855 364.495 ;
        RECT 589.495 364.215 589.775 364.495 ;
        RECT 590.205 364.215 590.485 364.495 ;
        RECT 590.915 364.215 591.195 364.495 ;
        RECT 591.625 364.215 591.905 364.495 ;
        RECT 592.335 364.215 592.615 364.495 ;
        RECT 593.045 364.215 593.325 364.495 ;
        RECT 593.755 364.215 594.035 364.495 ;
        RECT 594.465 364.215 594.745 364.495 ;
        RECT 595.175 364.215 595.455 364.495 ;
        RECT 595.885 364.215 596.165 364.495 ;
        RECT 596.595 364.215 596.875 364.495 ;
        RECT 597.305 364.215 597.585 364.495 ;
        RECT 598.015 364.215 598.295 364.495 ;
        RECT 1351.715 364.215 1351.995 364.495 ;
        RECT 1352.425 364.215 1352.705 364.495 ;
        RECT 1353.135 364.215 1353.415 364.495 ;
        RECT 1353.845 364.215 1354.125 364.495 ;
        RECT 1354.555 364.215 1354.835 364.495 ;
        RECT 1355.265 364.215 1355.545 364.495 ;
        RECT 1355.975 364.215 1356.255 364.495 ;
        RECT 1356.685 364.215 1356.965 364.495 ;
        RECT 1357.395 364.215 1357.675 364.495 ;
        RECT 1358.105 364.215 1358.385 364.495 ;
        RECT 1358.815 364.215 1359.095 364.495 ;
        RECT 1359.525 364.215 1359.805 364.495 ;
        RECT 1360.235 364.215 1360.515 364.495 ;
        RECT 1366.245 364.215 1366.525 364.495 ;
        RECT 1366.955 364.215 1367.235 364.495 ;
        RECT 1367.665 364.215 1367.945 364.495 ;
        RECT 1368.375 364.215 1368.655 364.495 ;
        RECT 1369.085 364.215 1369.365 364.495 ;
        RECT 1369.795 364.215 1370.075 364.495 ;
        RECT 1370.505 364.215 1370.785 364.495 ;
        RECT 1371.215 364.215 1371.495 364.495 ;
        RECT 1371.925 364.215 1372.205 364.495 ;
        RECT 1372.635 364.215 1372.915 364.495 ;
        RECT 1373.345 364.215 1373.625 364.495 ;
        RECT 1375.965 364.215 1376.245 364.495 ;
        RECT 1376.675 364.215 1376.955 364.495 ;
        RECT 1377.385 364.215 1377.665 364.495 ;
        RECT 1378.095 364.215 1378.375 364.495 ;
        RECT 1378.805 364.215 1379.085 364.495 ;
        RECT 1379.515 364.215 1379.795 364.495 ;
        RECT 1380.225 364.215 1380.505 364.495 ;
        RECT 1380.935 364.215 1381.215 364.495 ;
        RECT 1381.645 364.215 1381.925 364.495 ;
        RECT 1382.355 364.215 1382.635 364.495 ;
        RECT 1383.065 364.215 1383.345 364.495 ;
        RECT 1383.775 364.215 1384.055 364.495 ;
        RECT 1384.485 364.215 1384.765 364.495 ;
        RECT 1385.195 364.215 1385.475 364.495 ;
        RECT 1389.495 364.215 1389.775 364.495 ;
        RECT 1390.205 364.215 1390.485 364.495 ;
        RECT 1390.915 364.215 1391.195 364.495 ;
        RECT 1391.625 364.215 1391.905 364.495 ;
        RECT 1392.335 364.215 1392.615 364.495 ;
        RECT 1393.045 364.215 1393.325 364.495 ;
        RECT 1393.755 364.215 1394.035 364.495 ;
        RECT 1394.465 364.215 1394.745 364.495 ;
        RECT 1395.175 364.215 1395.455 364.495 ;
        RECT 1395.885 364.215 1396.165 364.495 ;
        RECT 1396.595 364.215 1396.875 364.495 ;
        RECT 1397.305 364.215 1397.585 364.495 ;
        RECT 1398.015 364.215 1398.295 364.495 ;
        RECT 1398.725 364.215 1399.005 364.495 ;
        RECT 1401.345 364.215 1401.625 364.495 ;
        RECT 1402.055 364.215 1402.335 364.495 ;
        RECT 1402.765 364.215 1403.045 364.495 ;
        RECT 1403.475 364.215 1403.755 364.495 ;
        RECT 1404.185 364.215 1404.465 364.495 ;
        RECT 1404.895 364.215 1405.175 364.495 ;
        RECT 1405.605 364.215 1405.885 364.495 ;
        RECT 1406.315 364.215 1406.595 364.495 ;
        RECT 1407.025 364.215 1407.305 364.495 ;
        RECT 1407.735 364.215 1408.015 364.495 ;
        RECT 1408.445 364.215 1408.725 364.495 ;
        RECT 1409.155 364.215 1409.435 364.495 ;
        RECT 1409.865 364.215 1410.145 364.495 ;
        RECT 1410.575 364.215 1410.855 364.495 ;
        RECT 1414.495 364.215 1414.775 364.495 ;
        RECT 1415.205 364.215 1415.485 364.495 ;
        RECT 1415.915 364.215 1416.195 364.495 ;
        RECT 1416.625 364.215 1416.905 364.495 ;
        RECT 1417.335 364.215 1417.615 364.495 ;
        RECT 1418.045 364.215 1418.325 364.495 ;
        RECT 1418.755 364.215 1419.035 364.495 ;
        RECT 1419.465 364.215 1419.745 364.495 ;
        RECT 3001.715 364.215 3001.995 364.495 ;
        RECT 3002.425 364.215 3002.705 364.495 ;
        RECT 3003.135 364.215 3003.415 364.495 ;
        RECT 3003.845 364.215 3004.125 364.495 ;
        RECT 3004.555 364.215 3004.835 364.495 ;
        RECT 3005.265 364.215 3005.545 364.495 ;
        RECT 3005.975 364.215 3006.255 364.495 ;
        RECT 3006.685 364.215 3006.965 364.495 ;
        RECT 3007.395 364.215 3007.675 364.495 ;
        RECT 3008.105 364.215 3008.385 364.495 ;
        RECT 3008.815 364.215 3009.095 364.495 ;
        RECT 3009.525 364.215 3009.805 364.495 ;
        RECT 3010.235 364.215 3010.515 364.495 ;
        RECT 3014.115 364.215 3014.395 364.495 ;
        RECT 3014.825 364.215 3015.105 364.495 ;
        RECT 3015.535 364.215 3015.815 364.495 ;
        RECT 3016.245 364.215 3016.525 364.495 ;
        RECT 3016.955 364.215 3017.235 364.495 ;
        RECT 3017.665 364.215 3017.945 364.495 ;
        RECT 3018.375 364.215 3018.655 364.495 ;
        RECT 3019.085 364.215 3019.365 364.495 ;
        RECT 3019.795 364.215 3020.075 364.495 ;
        RECT 3025.965 364.215 3026.245 364.495 ;
        RECT 3026.675 364.215 3026.955 364.495 ;
        RECT 3027.385 364.215 3027.665 364.495 ;
        RECT 3028.095 364.215 3028.375 364.495 ;
        RECT 3028.805 364.215 3029.085 364.495 ;
        RECT 3029.515 364.215 3029.795 364.495 ;
        RECT 3030.225 364.215 3030.505 364.495 ;
        RECT 3030.935 364.215 3031.215 364.495 ;
        RECT 3031.645 364.215 3031.925 364.495 ;
        RECT 3032.355 364.215 3032.635 364.495 ;
        RECT 3033.065 364.215 3033.345 364.495 ;
        RECT 3033.775 364.215 3034.055 364.495 ;
        RECT 3034.485 364.215 3034.765 364.495 ;
        RECT 3035.195 364.215 3035.475 364.495 ;
        RECT 3039.495 364.215 3039.775 364.495 ;
        RECT 3040.205 364.215 3040.485 364.495 ;
        RECT 3040.915 364.215 3041.195 364.495 ;
        RECT 3041.625 364.215 3041.905 364.495 ;
        RECT 3042.335 364.215 3042.615 364.495 ;
        RECT 3046.595 364.215 3046.875 364.495 ;
        RECT 3047.305 364.215 3047.585 364.495 ;
        RECT 3048.015 364.215 3048.295 364.495 ;
        RECT 3048.725 364.215 3049.005 364.495 ;
        RECT 3051.345 364.215 3051.625 364.495 ;
        RECT 3052.055 364.215 3052.335 364.495 ;
        RECT 3052.765 364.215 3053.045 364.495 ;
        RECT 3053.475 364.215 3053.755 364.495 ;
        RECT 3054.185 364.215 3054.465 364.495 ;
        RECT 3054.895 364.215 3055.175 364.495 ;
        RECT 3055.605 364.215 3055.885 364.495 ;
        RECT 3056.315 364.215 3056.595 364.495 ;
        RECT 3057.025 364.215 3057.305 364.495 ;
        RECT 3057.735 364.215 3058.015 364.495 ;
        RECT 3058.445 364.215 3058.725 364.495 ;
        RECT 3059.155 364.215 3059.435 364.495 ;
        RECT 3059.865 364.215 3060.145 364.495 ;
        RECT 3060.575 364.215 3060.855 364.495 ;
        RECT 3064.495 364.215 3064.775 364.495 ;
        RECT 3065.205 364.215 3065.485 364.495 ;
        RECT 3065.915 364.215 3066.195 364.495 ;
        RECT 3066.625 364.215 3066.905 364.495 ;
        RECT 3067.335 364.215 3067.615 364.495 ;
        RECT 3068.045 364.215 3068.325 364.495 ;
        RECT 3068.755 364.215 3069.035 364.495 ;
        RECT 3069.465 364.215 3069.745 364.495 ;
        RECT 3070.175 364.215 3070.455 364.495 ;
        RECT 3070.885 364.215 3071.165 364.495 ;
        RECT 3071.595 364.215 3071.875 364.495 ;
        RECT 3072.305 364.215 3072.585 364.495 ;
        RECT 3073.015 364.215 3073.295 364.495 ;
        RECT 526.715 363.505 526.995 363.785 ;
        RECT 527.425 363.505 527.705 363.785 ;
        RECT 528.135 363.505 528.415 363.785 ;
        RECT 528.845 363.505 529.125 363.785 ;
        RECT 529.555 363.505 529.835 363.785 ;
        RECT 530.265 363.505 530.545 363.785 ;
        RECT 530.975 363.505 531.255 363.785 ;
        RECT 531.685 363.505 531.965 363.785 ;
        RECT 532.395 363.505 532.675 363.785 ;
        RECT 533.105 363.505 533.385 363.785 ;
        RECT 533.815 363.505 534.095 363.785 ;
        RECT 534.525 363.505 534.805 363.785 ;
        RECT 535.235 363.505 535.515 363.785 ;
        RECT 544.975 363.505 545.255 363.785 ;
        RECT 545.685 363.505 545.965 363.785 ;
        RECT 546.395 363.505 546.675 363.785 ;
        RECT 547.105 363.505 547.385 363.785 ;
        RECT 547.815 363.505 548.095 363.785 ;
        RECT 548.525 363.505 548.805 363.785 ;
        RECT 550.965 363.505 551.245 363.785 ;
        RECT 551.675 363.505 551.955 363.785 ;
        RECT 552.385 363.505 552.665 363.785 ;
        RECT 553.095 363.505 553.375 363.785 ;
        RECT 553.805 363.505 554.085 363.785 ;
        RECT 554.515 363.505 554.795 363.785 ;
        RECT 555.225 363.505 555.505 363.785 ;
        RECT 555.935 363.505 556.215 363.785 ;
        RECT 556.645 363.505 556.925 363.785 ;
        RECT 557.355 363.505 557.635 363.785 ;
        RECT 558.065 363.505 558.345 363.785 ;
        RECT 558.775 363.505 559.055 363.785 ;
        RECT 559.485 363.505 559.765 363.785 ;
        RECT 560.195 363.505 560.475 363.785 ;
        RECT 566.625 363.505 566.905 363.785 ;
        RECT 567.335 363.505 567.615 363.785 ;
        RECT 568.045 363.505 568.325 363.785 ;
        RECT 568.755 363.505 569.035 363.785 ;
        RECT 569.465 363.505 569.745 363.785 ;
        RECT 570.175 363.505 570.455 363.785 ;
        RECT 570.885 363.505 571.165 363.785 ;
        RECT 571.595 363.505 571.875 363.785 ;
        RECT 572.305 363.505 572.585 363.785 ;
        RECT 573.015 363.505 573.295 363.785 ;
        RECT 573.725 363.505 574.005 363.785 ;
        RECT 576.345 363.505 576.625 363.785 ;
        RECT 577.055 363.505 577.335 363.785 ;
        RECT 577.765 363.505 578.045 363.785 ;
        RECT 578.475 363.505 578.755 363.785 ;
        RECT 579.185 363.505 579.465 363.785 ;
        RECT 579.895 363.505 580.175 363.785 ;
        RECT 580.605 363.505 580.885 363.785 ;
        RECT 581.315 363.505 581.595 363.785 ;
        RECT 582.025 363.505 582.305 363.785 ;
        RECT 582.735 363.505 583.015 363.785 ;
        RECT 583.445 363.505 583.725 363.785 ;
        RECT 584.155 363.505 584.435 363.785 ;
        RECT 584.865 363.505 585.145 363.785 ;
        RECT 585.575 363.505 585.855 363.785 ;
        RECT 589.495 363.505 589.775 363.785 ;
        RECT 590.205 363.505 590.485 363.785 ;
        RECT 590.915 363.505 591.195 363.785 ;
        RECT 591.625 363.505 591.905 363.785 ;
        RECT 592.335 363.505 592.615 363.785 ;
        RECT 593.045 363.505 593.325 363.785 ;
        RECT 593.755 363.505 594.035 363.785 ;
        RECT 594.465 363.505 594.745 363.785 ;
        RECT 595.175 363.505 595.455 363.785 ;
        RECT 595.885 363.505 596.165 363.785 ;
        RECT 596.595 363.505 596.875 363.785 ;
        RECT 597.305 363.505 597.585 363.785 ;
        RECT 598.015 363.505 598.295 363.785 ;
        RECT 1351.715 363.505 1351.995 363.785 ;
        RECT 1352.425 363.505 1352.705 363.785 ;
        RECT 1353.135 363.505 1353.415 363.785 ;
        RECT 1353.845 363.505 1354.125 363.785 ;
        RECT 1354.555 363.505 1354.835 363.785 ;
        RECT 1355.265 363.505 1355.545 363.785 ;
        RECT 1355.975 363.505 1356.255 363.785 ;
        RECT 1356.685 363.505 1356.965 363.785 ;
        RECT 1357.395 363.505 1357.675 363.785 ;
        RECT 1358.105 363.505 1358.385 363.785 ;
        RECT 1358.815 363.505 1359.095 363.785 ;
        RECT 1359.525 363.505 1359.805 363.785 ;
        RECT 1360.235 363.505 1360.515 363.785 ;
        RECT 1366.245 363.505 1366.525 363.785 ;
        RECT 1366.955 363.505 1367.235 363.785 ;
        RECT 1367.665 363.505 1367.945 363.785 ;
        RECT 1368.375 363.505 1368.655 363.785 ;
        RECT 1369.085 363.505 1369.365 363.785 ;
        RECT 1369.795 363.505 1370.075 363.785 ;
        RECT 1370.505 363.505 1370.785 363.785 ;
        RECT 1371.215 363.505 1371.495 363.785 ;
        RECT 1371.925 363.505 1372.205 363.785 ;
        RECT 1372.635 363.505 1372.915 363.785 ;
        RECT 1373.345 363.505 1373.625 363.785 ;
        RECT 1375.965 363.505 1376.245 363.785 ;
        RECT 1376.675 363.505 1376.955 363.785 ;
        RECT 1377.385 363.505 1377.665 363.785 ;
        RECT 1378.095 363.505 1378.375 363.785 ;
        RECT 1378.805 363.505 1379.085 363.785 ;
        RECT 1379.515 363.505 1379.795 363.785 ;
        RECT 1380.225 363.505 1380.505 363.785 ;
        RECT 1380.935 363.505 1381.215 363.785 ;
        RECT 1381.645 363.505 1381.925 363.785 ;
        RECT 1382.355 363.505 1382.635 363.785 ;
        RECT 1383.065 363.505 1383.345 363.785 ;
        RECT 1383.775 363.505 1384.055 363.785 ;
        RECT 1384.485 363.505 1384.765 363.785 ;
        RECT 1385.195 363.505 1385.475 363.785 ;
        RECT 1389.495 363.505 1389.775 363.785 ;
        RECT 1390.205 363.505 1390.485 363.785 ;
        RECT 1390.915 363.505 1391.195 363.785 ;
        RECT 1391.625 363.505 1391.905 363.785 ;
        RECT 1392.335 363.505 1392.615 363.785 ;
        RECT 1393.045 363.505 1393.325 363.785 ;
        RECT 1393.755 363.505 1394.035 363.785 ;
        RECT 1394.465 363.505 1394.745 363.785 ;
        RECT 1395.175 363.505 1395.455 363.785 ;
        RECT 1395.885 363.505 1396.165 363.785 ;
        RECT 1396.595 363.505 1396.875 363.785 ;
        RECT 1397.305 363.505 1397.585 363.785 ;
        RECT 1398.015 363.505 1398.295 363.785 ;
        RECT 1398.725 363.505 1399.005 363.785 ;
        RECT 1401.345 363.505 1401.625 363.785 ;
        RECT 1402.055 363.505 1402.335 363.785 ;
        RECT 1402.765 363.505 1403.045 363.785 ;
        RECT 1403.475 363.505 1403.755 363.785 ;
        RECT 1404.185 363.505 1404.465 363.785 ;
        RECT 1404.895 363.505 1405.175 363.785 ;
        RECT 1405.605 363.505 1405.885 363.785 ;
        RECT 1406.315 363.505 1406.595 363.785 ;
        RECT 1407.025 363.505 1407.305 363.785 ;
        RECT 1407.735 363.505 1408.015 363.785 ;
        RECT 1408.445 363.505 1408.725 363.785 ;
        RECT 1409.155 363.505 1409.435 363.785 ;
        RECT 1409.865 363.505 1410.145 363.785 ;
        RECT 1410.575 363.505 1410.855 363.785 ;
        RECT 1414.495 363.505 1414.775 363.785 ;
        RECT 1415.205 363.505 1415.485 363.785 ;
        RECT 1415.915 363.505 1416.195 363.785 ;
        RECT 1416.625 363.505 1416.905 363.785 ;
        RECT 1417.335 363.505 1417.615 363.785 ;
        RECT 1418.045 363.505 1418.325 363.785 ;
        RECT 1418.755 363.505 1419.035 363.785 ;
        RECT 1419.465 363.505 1419.745 363.785 ;
        RECT 3001.715 363.505 3001.995 363.785 ;
        RECT 3002.425 363.505 3002.705 363.785 ;
        RECT 3003.135 363.505 3003.415 363.785 ;
        RECT 3003.845 363.505 3004.125 363.785 ;
        RECT 3004.555 363.505 3004.835 363.785 ;
        RECT 3005.265 363.505 3005.545 363.785 ;
        RECT 3005.975 363.505 3006.255 363.785 ;
        RECT 3006.685 363.505 3006.965 363.785 ;
        RECT 3007.395 363.505 3007.675 363.785 ;
        RECT 3008.105 363.505 3008.385 363.785 ;
        RECT 3008.815 363.505 3009.095 363.785 ;
        RECT 3009.525 363.505 3009.805 363.785 ;
        RECT 3010.235 363.505 3010.515 363.785 ;
        RECT 3014.115 363.505 3014.395 363.785 ;
        RECT 3014.825 363.505 3015.105 363.785 ;
        RECT 3015.535 363.505 3015.815 363.785 ;
        RECT 3016.245 363.505 3016.525 363.785 ;
        RECT 3016.955 363.505 3017.235 363.785 ;
        RECT 3017.665 363.505 3017.945 363.785 ;
        RECT 3018.375 363.505 3018.655 363.785 ;
        RECT 3019.085 363.505 3019.365 363.785 ;
        RECT 3019.795 363.505 3020.075 363.785 ;
        RECT 3025.965 363.505 3026.245 363.785 ;
        RECT 3026.675 363.505 3026.955 363.785 ;
        RECT 3027.385 363.505 3027.665 363.785 ;
        RECT 3028.095 363.505 3028.375 363.785 ;
        RECT 3028.805 363.505 3029.085 363.785 ;
        RECT 3029.515 363.505 3029.795 363.785 ;
        RECT 3030.225 363.505 3030.505 363.785 ;
        RECT 3030.935 363.505 3031.215 363.785 ;
        RECT 3031.645 363.505 3031.925 363.785 ;
        RECT 3032.355 363.505 3032.635 363.785 ;
        RECT 3033.065 363.505 3033.345 363.785 ;
        RECT 3033.775 363.505 3034.055 363.785 ;
        RECT 3034.485 363.505 3034.765 363.785 ;
        RECT 3035.195 363.505 3035.475 363.785 ;
        RECT 3039.495 363.505 3039.775 363.785 ;
        RECT 3040.205 363.505 3040.485 363.785 ;
        RECT 3040.915 363.505 3041.195 363.785 ;
        RECT 3041.625 363.505 3041.905 363.785 ;
        RECT 3042.335 363.505 3042.615 363.785 ;
        RECT 3046.595 363.505 3046.875 363.785 ;
        RECT 3047.305 363.505 3047.585 363.785 ;
        RECT 3048.015 363.505 3048.295 363.785 ;
        RECT 3048.725 363.505 3049.005 363.785 ;
        RECT 3051.345 363.505 3051.625 363.785 ;
        RECT 3052.055 363.505 3052.335 363.785 ;
        RECT 3052.765 363.505 3053.045 363.785 ;
        RECT 3053.475 363.505 3053.755 363.785 ;
        RECT 3054.185 363.505 3054.465 363.785 ;
        RECT 3054.895 363.505 3055.175 363.785 ;
        RECT 3055.605 363.505 3055.885 363.785 ;
        RECT 3056.315 363.505 3056.595 363.785 ;
        RECT 3057.025 363.505 3057.305 363.785 ;
        RECT 3057.735 363.505 3058.015 363.785 ;
        RECT 3058.445 363.505 3058.725 363.785 ;
        RECT 3059.155 363.505 3059.435 363.785 ;
        RECT 3059.865 363.505 3060.145 363.785 ;
        RECT 3060.575 363.505 3060.855 363.785 ;
        RECT 3064.495 363.505 3064.775 363.785 ;
        RECT 3065.205 363.505 3065.485 363.785 ;
        RECT 3065.915 363.505 3066.195 363.785 ;
        RECT 3066.625 363.505 3066.905 363.785 ;
        RECT 3067.335 363.505 3067.615 363.785 ;
        RECT 3068.045 363.505 3068.325 363.785 ;
        RECT 3068.755 363.505 3069.035 363.785 ;
        RECT 3069.465 363.505 3069.745 363.785 ;
        RECT 3070.175 363.505 3070.455 363.785 ;
        RECT 3070.885 363.505 3071.165 363.785 ;
        RECT 3071.595 363.505 3071.875 363.785 ;
        RECT 3072.305 363.505 3072.585 363.785 ;
        RECT 3073.015 363.505 3073.295 363.785 ;
        RECT 526.715 362.795 526.995 363.075 ;
        RECT 527.425 362.795 527.705 363.075 ;
        RECT 528.135 362.795 528.415 363.075 ;
        RECT 528.845 362.795 529.125 363.075 ;
        RECT 529.555 362.795 529.835 363.075 ;
        RECT 530.265 362.795 530.545 363.075 ;
        RECT 530.975 362.795 531.255 363.075 ;
        RECT 531.685 362.795 531.965 363.075 ;
        RECT 532.395 362.795 532.675 363.075 ;
        RECT 533.105 362.795 533.385 363.075 ;
        RECT 533.815 362.795 534.095 363.075 ;
        RECT 534.525 362.795 534.805 363.075 ;
        RECT 535.235 362.795 535.515 363.075 ;
        RECT 544.975 362.795 545.255 363.075 ;
        RECT 545.685 362.795 545.965 363.075 ;
        RECT 546.395 362.795 546.675 363.075 ;
        RECT 547.105 362.795 547.385 363.075 ;
        RECT 547.815 362.795 548.095 363.075 ;
        RECT 548.525 362.795 548.805 363.075 ;
        RECT 550.965 362.795 551.245 363.075 ;
        RECT 551.675 362.795 551.955 363.075 ;
        RECT 552.385 362.795 552.665 363.075 ;
        RECT 553.095 362.795 553.375 363.075 ;
        RECT 553.805 362.795 554.085 363.075 ;
        RECT 554.515 362.795 554.795 363.075 ;
        RECT 555.225 362.795 555.505 363.075 ;
        RECT 555.935 362.795 556.215 363.075 ;
        RECT 556.645 362.795 556.925 363.075 ;
        RECT 557.355 362.795 557.635 363.075 ;
        RECT 558.065 362.795 558.345 363.075 ;
        RECT 558.775 362.795 559.055 363.075 ;
        RECT 559.485 362.795 559.765 363.075 ;
        RECT 560.195 362.795 560.475 363.075 ;
        RECT 566.625 362.795 566.905 363.075 ;
        RECT 567.335 362.795 567.615 363.075 ;
        RECT 568.045 362.795 568.325 363.075 ;
        RECT 568.755 362.795 569.035 363.075 ;
        RECT 569.465 362.795 569.745 363.075 ;
        RECT 570.175 362.795 570.455 363.075 ;
        RECT 570.885 362.795 571.165 363.075 ;
        RECT 571.595 362.795 571.875 363.075 ;
        RECT 572.305 362.795 572.585 363.075 ;
        RECT 573.015 362.795 573.295 363.075 ;
        RECT 573.725 362.795 574.005 363.075 ;
        RECT 576.345 362.795 576.625 363.075 ;
        RECT 577.055 362.795 577.335 363.075 ;
        RECT 577.765 362.795 578.045 363.075 ;
        RECT 578.475 362.795 578.755 363.075 ;
        RECT 579.185 362.795 579.465 363.075 ;
        RECT 579.895 362.795 580.175 363.075 ;
        RECT 580.605 362.795 580.885 363.075 ;
        RECT 581.315 362.795 581.595 363.075 ;
        RECT 582.025 362.795 582.305 363.075 ;
        RECT 582.735 362.795 583.015 363.075 ;
        RECT 583.445 362.795 583.725 363.075 ;
        RECT 584.155 362.795 584.435 363.075 ;
        RECT 584.865 362.795 585.145 363.075 ;
        RECT 585.575 362.795 585.855 363.075 ;
        RECT 589.495 362.795 589.775 363.075 ;
        RECT 590.205 362.795 590.485 363.075 ;
        RECT 590.915 362.795 591.195 363.075 ;
        RECT 591.625 362.795 591.905 363.075 ;
        RECT 592.335 362.795 592.615 363.075 ;
        RECT 593.045 362.795 593.325 363.075 ;
        RECT 593.755 362.795 594.035 363.075 ;
        RECT 594.465 362.795 594.745 363.075 ;
        RECT 595.175 362.795 595.455 363.075 ;
        RECT 595.885 362.795 596.165 363.075 ;
        RECT 596.595 362.795 596.875 363.075 ;
        RECT 597.305 362.795 597.585 363.075 ;
        RECT 598.015 362.795 598.295 363.075 ;
        RECT 1351.715 362.795 1351.995 363.075 ;
        RECT 1352.425 362.795 1352.705 363.075 ;
        RECT 1353.135 362.795 1353.415 363.075 ;
        RECT 1353.845 362.795 1354.125 363.075 ;
        RECT 1354.555 362.795 1354.835 363.075 ;
        RECT 1355.265 362.795 1355.545 363.075 ;
        RECT 1355.975 362.795 1356.255 363.075 ;
        RECT 1356.685 362.795 1356.965 363.075 ;
        RECT 1357.395 362.795 1357.675 363.075 ;
        RECT 1358.105 362.795 1358.385 363.075 ;
        RECT 1358.815 362.795 1359.095 363.075 ;
        RECT 1359.525 362.795 1359.805 363.075 ;
        RECT 1360.235 362.795 1360.515 363.075 ;
        RECT 1366.245 362.795 1366.525 363.075 ;
        RECT 1366.955 362.795 1367.235 363.075 ;
        RECT 1367.665 362.795 1367.945 363.075 ;
        RECT 1368.375 362.795 1368.655 363.075 ;
        RECT 1369.085 362.795 1369.365 363.075 ;
        RECT 1369.795 362.795 1370.075 363.075 ;
        RECT 1370.505 362.795 1370.785 363.075 ;
        RECT 1371.215 362.795 1371.495 363.075 ;
        RECT 1371.925 362.795 1372.205 363.075 ;
        RECT 1372.635 362.795 1372.915 363.075 ;
        RECT 1373.345 362.795 1373.625 363.075 ;
        RECT 1375.965 362.795 1376.245 363.075 ;
        RECT 1376.675 362.795 1376.955 363.075 ;
        RECT 1377.385 362.795 1377.665 363.075 ;
        RECT 1378.095 362.795 1378.375 363.075 ;
        RECT 1378.805 362.795 1379.085 363.075 ;
        RECT 1379.515 362.795 1379.795 363.075 ;
        RECT 1380.225 362.795 1380.505 363.075 ;
        RECT 1380.935 362.795 1381.215 363.075 ;
        RECT 1381.645 362.795 1381.925 363.075 ;
        RECT 1382.355 362.795 1382.635 363.075 ;
        RECT 1383.065 362.795 1383.345 363.075 ;
        RECT 1383.775 362.795 1384.055 363.075 ;
        RECT 1384.485 362.795 1384.765 363.075 ;
        RECT 1385.195 362.795 1385.475 363.075 ;
        RECT 1389.495 362.795 1389.775 363.075 ;
        RECT 1390.205 362.795 1390.485 363.075 ;
        RECT 1390.915 362.795 1391.195 363.075 ;
        RECT 1391.625 362.795 1391.905 363.075 ;
        RECT 1392.335 362.795 1392.615 363.075 ;
        RECT 1393.045 362.795 1393.325 363.075 ;
        RECT 1393.755 362.795 1394.035 363.075 ;
        RECT 1394.465 362.795 1394.745 363.075 ;
        RECT 1395.175 362.795 1395.455 363.075 ;
        RECT 1395.885 362.795 1396.165 363.075 ;
        RECT 1396.595 362.795 1396.875 363.075 ;
        RECT 1397.305 362.795 1397.585 363.075 ;
        RECT 1398.015 362.795 1398.295 363.075 ;
        RECT 1398.725 362.795 1399.005 363.075 ;
        RECT 1401.345 362.795 1401.625 363.075 ;
        RECT 1402.055 362.795 1402.335 363.075 ;
        RECT 1402.765 362.795 1403.045 363.075 ;
        RECT 1403.475 362.795 1403.755 363.075 ;
        RECT 1404.185 362.795 1404.465 363.075 ;
        RECT 1404.895 362.795 1405.175 363.075 ;
        RECT 1405.605 362.795 1405.885 363.075 ;
        RECT 1406.315 362.795 1406.595 363.075 ;
        RECT 1407.025 362.795 1407.305 363.075 ;
        RECT 1407.735 362.795 1408.015 363.075 ;
        RECT 1408.445 362.795 1408.725 363.075 ;
        RECT 1409.155 362.795 1409.435 363.075 ;
        RECT 1409.865 362.795 1410.145 363.075 ;
        RECT 1410.575 362.795 1410.855 363.075 ;
        RECT 1414.495 362.795 1414.775 363.075 ;
        RECT 1415.205 362.795 1415.485 363.075 ;
        RECT 1415.915 362.795 1416.195 363.075 ;
        RECT 1416.625 362.795 1416.905 363.075 ;
        RECT 1417.335 362.795 1417.615 363.075 ;
        RECT 1418.045 362.795 1418.325 363.075 ;
        RECT 1418.755 362.795 1419.035 363.075 ;
        RECT 1419.465 362.795 1419.745 363.075 ;
        RECT 3001.715 362.795 3001.995 363.075 ;
        RECT 3002.425 362.795 3002.705 363.075 ;
        RECT 3003.135 362.795 3003.415 363.075 ;
        RECT 3003.845 362.795 3004.125 363.075 ;
        RECT 3004.555 362.795 3004.835 363.075 ;
        RECT 3005.265 362.795 3005.545 363.075 ;
        RECT 3005.975 362.795 3006.255 363.075 ;
        RECT 3006.685 362.795 3006.965 363.075 ;
        RECT 3007.395 362.795 3007.675 363.075 ;
        RECT 3008.105 362.795 3008.385 363.075 ;
        RECT 3008.815 362.795 3009.095 363.075 ;
        RECT 3009.525 362.795 3009.805 363.075 ;
        RECT 3010.235 362.795 3010.515 363.075 ;
        RECT 3014.115 362.795 3014.395 363.075 ;
        RECT 3014.825 362.795 3015.105 363.075 ;
        RECT 3015.535 362.795 3015.815 363.075 ;
        RECT 3016.245 362.795 3016.525 363.075 ;
        RECT 3016.955 362.795 3017.235 363.075 ;
        RECT 3017.665 362.795 3017.945 363.075 ;
        RECT 3018.375 362.795 3018.655 363.075 ;
        RECT 3019.085 362.795 3019.365 363.075 ;
        RECT 3019.795 362.795 3020.075 363.075 ;
        RECT 3025.965 362.795 3026.245 363.075 ;
        RECT 3026.675 362.795 3026.955 363.075 ;
        RECT 3027.385 362.795 3027.665 363.075 ;
        RECT 3028.095 362.795 3028.375 363.075 ;
        RECT 3028.805 362.795 3029.085 363.075 ;
        RECT 3029.515 362.795 3029.795 363.075 ;
        RECT 3030.225 362.795 3030.505 363.075 ;
        RECT 3030.935 362.795 3031.215 363.075 ;
        RECT 3031.645 362.795 3031.925 363.075 ;
        RECT 3032.355 362.795 3032.635 363.075 ;
        RECT 3033.065 362.795 3033.345 363.075 ;
        RECT 3033.775 362.795 3034.055 363.075 ;
        RECT 3034.485 362.795 3034.765 363.075 ;
        RECT 3035.195 362.795 3035.475 363.075 ;
        RECT 3039.495 362.795 3039.775 363.075 ;
        RECT 3040.205 362.795 3040.485 363.075 ;
        RECT 3040.915 362.795 3041.195 363.075 ;
        RECT 3041.625 362.795 3041.905 363.075 ;
        RECT 3042.335 362.795 3042.615 363.075 ;
        RECT 3046.595 362.795 3046.875 363.075 ;
        RECT 3047.305 362.795 3047.585 363.075 ;
        RECT 3048.015 362.795 3048.295 363.075 ;
        RECT 3048.725 362.795 3049.005 363.075 ;
        RECT 3051.345 362.795 3051.625 363.075 ;
        RECT 3052.055 362.795 3052.335 363.075 ;
        RECT 3052.765 362.795 3053.045 363.075 ;
        RECT 3053.475 362.795 3053.755 363.075 ;
        RECT 3054.185 362.795 3054.465 363.075 ;
        RECT 3054.895 362.795 3055.175 363.075 ;
        RECT 3055.605 362.795 3055.885 363.075 ;
        RECT 3056.315 362.795 3056.595 363.075 ;
        RECT 3057.025 362.795 3057.305 363.075 ;
        RECT 3057.735 362.795 3058.015 363.075 ;
        RECT 3058.445 362.795 3058.725 363.075 ;
        RECT 3059.155 362.795 3059.435 363.075 ;
        RECT 3059.865 362.795 3060.145 363.075 ;
        RECT 3060.575 362.795 3060.855 363.075 ;
        RECT 3064.495 362.795 3064.775 363.075 ;
        RECT 3065.205 362.795 3065.485 363.075 ;
        RECT 3065.915 362.795 3066.195 363.075 ;
        RECT 3066.625 362.795 3066.905 363.075 ;
        RECT 3067.335 362.795 3067.615 363.075 ;
        RECT 3068.045 362.795 3068.325 363.075 ;
        RECT 3068.755 362.795 3069.035 363.075 ;
        RECT 3069.465 362.795 3069.745 363.075 ;
        RECT 3070.175 362.795 3070.455 363.075 ;
        RECT 3070.885 362.795 3071.165 363.075 ;
        RECT 3071.595 362.795 3071.875 363.075 ;
        RECT 3072.305 362.795 3072.585 363.075 ;
        RECT 3073.015 362.795 3073.295 363.075 ;
        RECT 526.715 362.085 526.995 362.365 ;
        RECT 527.425 362.085 527.705 362.365 ;
        RECT 528.135 362.085 528.415 362.365 ;
        RECT 528.845 362.085 529.125 362.365 ;
        RECT 529.555 362.085 529.835 362.365 ;
        RECT 530.265 362.085 530.545 362.365 ;
        RECT 530.975 362.085 531.255 362.365 ;
        RECT 531.685 362.085 531.965 362.365 ;
        RECT 532.395 362.085 532.675 362.365 ;
        RECT 533.105 362.085 533.385 362.365 ;
        RECT 533.815 362.085 534.095 362.365 ;
        RECT 534.525 362.085 534.805 362.365 ;
        RECT 535.235 362.085 535.515 362.365 ;
        RECT 544.975 362.085 545.255 362.365 ;
        RECT 545.685 362.085 545.965 362.365 ;
        RECT 546.395 362.085 546.675 362.365 ;
        RECT 547.105 362.085 547.385 362.365 ;
        RECT 547.815 362.085 548.095 362.365 ;
        RECT 548.525 362.085 548.805 362.365 ;
        RECT 550.965 362.085 551.245 362.365 ;
        RECT 551.675 362.085 551.955 362.365 ;
        RECT 552.385 362.085 552.665 362.365 ;
        RECT 553.095 362.085 553.375 362.365 ;
        RECT 553.805 362.085 554.085 362.365 ;
        RECT 554.515 362.085 554.795 362.365 ;
        RECT 555.225 362.085 555.505 362.365 ;
        RECT 555.935 362.085 556.215 362.365 ;
        RECT 556.645 362.085 556.925 362.365 ;
        RECT 557.355 362.085 557.635 362.365 ;
        RECT 558.065 362.085 558.345 362.365 ;
        RECT 558.775 362.085 559.055 362.365 ;
        RECT 559.485 362.085 559.765 362.365 ;
        RECT 560.195 362.085 560.475 362.365 ;
        RECT 566.625 362.085 566.905 362.365 ;
        RECT 567.335 362.085 567.615 362.365 ;
        RECT 568.045 362.085 568.325 362.365 ;
        RECT 568.755 362.085 569.035 362.365 ;
        RECT 569.465 362.085 569.745 362.365 ;
        RECT 570.175 362.085 570.455 362.365 ;
        RECT 570.885 362.085 571.165 362.365 ;
        RECT 571.595 362.085 571.875 362.365 ;
        RECT 572.305 362.085 572.585 362.365 ;
        RECT 573.015 362.085 573.295 362.365 ;
        RECT 573.725 362.085 574.005 362.365 ;
        RECT 576.345 362.085 576.625 362.365 ;
        RECT 577.055 362.085 577.335 362.365 ;
        RECT 577.765 362.085 578.045 362.365 ;
        RECT 578.475 362.085 578.755 362.365 ;
        RECT 579.185 362.085 579.465 362.365 ;
        RECT 579.895 362.085 580.175 362.365 ;
        RECT 580.605 362.085 580.885 362.365 ;
        RECT 581.315 362.085 581.595 362.365 ;
        RECT 582.025 362.085 582.305 362.365 ;
        RECT 582.735 362.085 583.015 362.365 ;
        RECT 583.445 362.085 583.725 362.365 ;
        RECT 584.155 362.085 584.435 362.365 ;
        RECT 584.865 362.085 585.145 362.365 ;
        RECT 585.575 362.085 585.855 362.365 ;
        RECT 589.495 362.085 589.775 362.365 ;
        RECT 590.205 362.085 590.485 362.365 ;
        RECT 590.915 362.085 591.195 362.365 ;
        RECT 591.625 362.085 591.905 362.365 ;
        RECT 592.335 362.085 592.615 362.365 ;
        RECT 593.045 362.085 593.325 362.365 ;
        RECT 593.755 362.085 594.035 362.365 ;
        RECT 594.465 362.085 594.745 362.365 ;
        RECT 595.175 362.085 595.455 362.365 ;
        RECT 595.885 362.085 596.165 362.365 ;
        RECT 596.595 362.085 596.875 362.365 ;
        RECT 597.305 362.085 597.585 362.365 ;
        RECT 598.015 362.085 598.295 362.365 ;
        RECT 1351.715 362.085 1351.995 362.365 ;
        RECT 1352.425 362.085 1352.705 362.365 ;
        RECT 1353.135 362.085 1353.415 362.365 ;
        RECT 1353.845 362.085 1354.125 362.365 ;
        RECT 1354.555 362.085 1354.835 362.365 ;
        RECT 1355.265 362.085 1355.545 362.365 ;
        RECT 1355.975 362.085 1356.255 362.365 ;
        RECT 1356.685 362.085 1356.965 362.365 ;
        RECT 1357.395 362.085 1357.675 362.365 ;
        RECT 1358.105 362.085 1358.385 362.365 ;
        RECT 1358.815 362.085 1359.095 362.365 ;
        RECT 1359.525 362.085 1359.805 362.365 ;
        RECT 1360.235 362.085 1360.515 362.365 ;
        RECT 1366.245 362.085 1366.525 362.365 ;
        RECT 1366.955 362.085 1367.235 362.365 ;
        RECT 1367.665 362.085 1367.945 362.365 ;
        RECT 1368.375 362.085 1368.655 362.365 ;
        RECT 1369.085 362.085 1369.365 362.365 ;
        RECT 1369.795 362.085 1370.075 362.365 ;
        RECT 1370.505 362.085 1370.785 362.365 ;
        RECT 1371.215 362.085 1371.495 362.365 ;
        RECT 1371.925 362.085 1372.205 362.365 ;
        RECT 1372.635 362.085 1372.915 362.365 ;
        RECT 1373.345 362.085 1373.625 362.365 ;
        RECT 1375.965 362.085 1376.245 362.365 ;
        RECT 1376.675 362.085 1376.955 362.365 ;
        RECT 1377.385 362.085 1377.665 362.365 ;
        RECT 1378.095 362.085 1378.375 362.365 ;
        RECT 1378.805 362.085 1379.085 362.365 ;
        RECT 1379.515 362.085 1379.795 362.365 ;
        RECT 1380.225 362.085 1380.505 362.365 ;
        RECT 1380.935 362.085 1381.215 362.365 ;
        RECT 1381.645 362.085 1381.925 362.365 ;
        RECT 1382.355 362.085 1382.635 362.365 ;
        RECT 1383.065 362.085 1383.345 362.365 ;
        RECT 1383.775 362.085 1384.055 362.365 ;
        RECT 1384.485 362.085 1384.765 362.365 ;
        RECT 1385.195 362.085 1385.475 362.365 ;
        RECT 1389.495 362.085 1389.775 362.365 ;
        RECT 1390.205 362.085 1390.485 362.365 ;
        RECT 1390.915 362.085 1391.195 362.365 ;
        RECT 1391.625 362.085 1391.905 362.365 ;
        RECT 1392.335 362.085 1392.615 362.365 ;
        RECT 1393.045 362.085 1393.325 362.365 ;
        RECT 1393.755 362.085 1394.035 362.365 ;
        RECT 1394.465 362.085 1394.745 362.365 ;
        RECT 1395.175 362.085 1395.455 362.365 ;
        RECT 1395.885 362.085 1396.165 362.365 ;
        RECT 1396.595 362.085 1396.875 362.365 ;
        RECT 1397.305 362.085 1397.585 362.365 ;
        RECT 1398.015 362.085 1398.295 362.365 ;
        RECT 1398.725 362.085 1399.005 362.365 ;
        RECT 1401.345 362.085 1401.625 362.365 ;
        RECT 1402.055 362.085 1402.335 362.365 ;
        RECT 1402.765 362.085 1403.045 362.365 ;
        RECT 1403.475 362.085 1403.755 362.365 ;
        RECT 1404.185 362.085 1404.465 362.365 ;
        RECT 1404.895 362.085 1405.175 362.365 ;
        RECT 1405.605 362.085 1405.885 362.365 ;
        RECT 1406.315 362.085 1406.595 362.365 ;
        RECT 1407.025 362.085 1407.305 362.365 ;
        RECT 1407.735 362.085 1408.015 362.365 ;
        RECT 1408.445 362.085 1408.725 362.365 ;
        RECT 1409.155 362.085 1409.435 362.365 ;
        RECT 1409.865 362.085 1410.145 362.365 ;
        RECT 1410.575 362.085 1410.855 362.365 ;
        RECT 1414.495 362.085 1414.775 362.365 ;
        RECT 1415.205 362.085 1415.485 362.365 ;
        RECT 1415.915 362.085 1416.195 362.365 ;
        RECT 1416.625 362.085 1416.905 362.365 ;
        RECT 1417.335 362.085 1417.615 362.365 ;
        RECT 1418.045 362.085 1418.325 362.365 ;
        RECT 1418.755 362.085 1419.035 362.365 ;
        RECT 1419.465 362.085 1419.745 362.365 ;
        RECT 3001.715 362.085 3001.995 362.365 ;
        RECT 3002.425 362.085 3002.705 362.365 ;
        RECT 3003.135 362.085 3003.415 362.365 ;
        RECT 3003.845 362.085 3004.125 362.365 ;
        RECT 3004.555 362.085 3004.835 362.365 ;
        RECT 3005.265 362.085 3005.545 362.365 ;
        RECT 3005.975 362.085 3006.255 362.365 ;
        RECT 3006.685 362.085 3006.965 362.365 ;
        RECT 3007.395 362.085 3007.675 362.365 ;
        RECT 3008.105 362.085 3008.385 362.365 ;
        RECT 3008.815 362.085 3009.095 362.365 ;
        RECT 3009.525 362.085 3009.805 362.365 ;
        RECT 3010.235 362.085 3010.515 362.365 ;
        RECT 3014.115 362.085 3014.395 362.365 ;
        RECT 3014.825 362.085 3015.105 362.365 ;
        RECT 3015.535 362.085 3015.815 362.365 ;
        RECT 3016.245 362.085 3016.525 362.365 ;
        RECT 3016.955 362.085 3017.235 362.365 ;
        RECT 3017.665 362.085 3017.945 362.365 ;
        RECT 3018.375 362.085 3018.655 362.365 ;
        RECT 3019.085 362.085 3019.365 362.365 ;
        RECT 3019.795 362.085 3020.075 362.365 ;
        RECT 3025.965 362.085 3026.245 362.365 ;
        RECT 3026.675 362.085 3026.955 362.365 ;
        RECT 3027.385 362.085 3027.665 362.365 ;
        RECT 3028.095 362.085 3028.375 362.365 ;
        RECT 3028.805 362.085 3029.085 362.365 ;
        RECT 3029.515 362.085 3029.795 362.365 ;
        RECT 3030.225 362.085 3030.505 362.365 ;
        RECT 3030.935 362.085 3031.215 362.365 ;
        RECT 3031.645 362.085 3031.925 362.365 ;
        RECT 3032.355 362.085 3032.635 362.365 ;
        RECT 3033.065 362.085 3033.345 362.365 ;
        RECT 3033.775 362.085 3034.055 362.365 ;
        RECT 3034.485 362.085 3034.765 362.365 ;
        RECT 3035.195 362.085 3035.475 362.365 ;
        RECT 3039.495 362.085 3039.775 362.365 ;
        RECT 3040.205 362.085 3040.485 362.365 ;
        RECT 3040.915 362.085 3041.195 362.365 ;
        RECT 3041.625 362.085 3041.905 362.365 ;
        RECT 3042.335 362.085 3042.615 362.365 ;
        RECT 3046.595 362.085 3046.875 362.365 ;
        RECT 3047.305 362.085 3047.585 362.365 ;
        RECT 3048.015 362.085 3048.295 362.365 ;
        RECT 3048.725 362.085 3049.005 362.365 ;
        RECT 3051.345 362.085 3051.625 362.365 ;
        RECT 3052.055 362.085 3052.335 362.365 ;
        RECT 3052.765 362.085 3053.045 362.365 ;
        RECT 3053.475 362.085 3053.755 362.365 ;
        RECT 3054.185 362.085 3054.465 362.365 ;
        RECT 3054.895 362.085 3055.175 362.365 ;
        RECT 3055.605 362.085 3055.885 362.365 ;
        RECT 3056.315 362.085 3056.595 362.365 ;
        RECT 3057.025 362.085 3057.305 362.365 ;
        RECT 3057.735 362.085 3058.015 362.365 ;
        RECT 3058.445 362.085 3058.725 362.365 ;
        RECT 3059.155 362.085 3059.435 362.365 ;
        RECT 3059.865 362.085 3060.145 362.365 ;
        RECT 3060.575 362.085 3060.855 362.365 ;
        RECT 3064.495 362.085 3064.775 362.365 ;
        RECT 3065.205 362.085 3065.485 362.365 ;
        RECT 3065.915 362.085 3066.195 362.365 ;
        RECT 3066.625 362.085 3066.905 362.365 ;
        RECT 3067.335 362.085 3067.615 362.365 ;
        RECT 3068.045 362.085 3068.325 362.365 ;
        RECT 3068.755 362.085 3069.035 362.365 ;
        RECT 3069.465 362.085 3069.745 362.365 ;
        RECT 3070.175 362.085 3070.455 362.365 ;
        RECT 3070.885 362.085 3071.165 362.365 ;
        RECT 3071.595 362.085 3071.875 362.365 ;
        RECT 3072.305 362.085 3072.585 362.365 ;
        RECT 3073.015 362.085 3073.295 362.365 ;
        RECT 526.715 361.375 526.995 361.655 ;
        RECT 527.425 361.375 527.705 361.655 ;
        RECT 528.135 361.375 528.415 361.655 ;
        RECT 528.845 361.375 529.125 361.655 ;
        RECT 529.555 361.375 529.835 361.655 ;
        RECT 530.265 361.375 530.545 361.655 ;
        RECT 530.975 361.375 531.255 361.655 ;
        RECT 531.685 361.375 531.965 361.655 ;
        RECT 532.395 361.375 532.675 361.655 ;
        RECT 533.105 361.375 533.385 361.655 ;
        RECT 533.815 361.375 534.095 361.655 ;
        RECT 534.525 361.375 534.805 361.655 ;
        RECT 535.235 361.375 535.515 361.655 ;
        RECT 544.975 361.375 545.255 361.655 ;
        RECT 545.685 361.375 545.965 361.655 ;
        RECT 546.395 361.375 546.675 361.655 ;
        RECT 547.105 361.375 547.385 361.655 ;
        RECT 547.815 361.375 548.095 361.655 ;
        RECT 548.525 361.375 548.805 361.655 ;
        RECT 550.965 361.375 551.245 361.655 ;
        RECT 551.675 361.375 551.955 361.655 ;
        RECT 552.385 361.375 552.665 361.655 ;
        RECT 553.095 361.375 553.375 361.655 ;
        RECT 553.805 361.375 554.085 361.655 ;
        RECT 554.515 361.375 554.795 361.655 ;
        RECT 555.225 361.375 555.505 361.655 ;
        RECT 555.935 361.375 556.215 361.655 ;
        RECT 556.645 361.375 556.925 361.655 ;
        RECT 557.355 361.375 557.635 361.655 ;
        RECT 558.065 361.375 558.345 361.655 ;
        RECT 558.775 361.375 559.055 361.655 ;
        RECT 559.485 361.375 559.765 361.655 ;
        RECT 560.195 361.375 560.475 361.655 ;
        RECT 566.625 361.375 566.905 361.655 ;
        RECT 567.335 361.375 567.615 361.655 ;
        RECT 568.045 361.375 568.325 361.655 ;
        RECT 568.755 361.375 569.035 361.655 ;
        RECT 569.465 361.375 569.745 361.655 ;
        RECT 570.175 361.375 570.455 361.655 ;
        RECT 570.885 361.375 571.165 361.655 ;
        RECT 571.595 361.375 571.875 361.655 ;
        RECT 572.305 361.375 572.585 361.655 ;
        RECT 573.015 361.375 573.295 361.655 ;
        RECT 573.725 361.375 574.005 361.655 ;
        RECT 576.345 361.375 576.625 361.655 ;
        RECT 577.055 361.375 577.335 361.655 ;
        RECT 577.765 361.375 578.045 361.655 ;
        RECT 578.475 361.375 578.755 361.655 ;
        RECT 579.185 361.375 579.465 361.655 ;
        RECT 579.895 361.375 580.175 361.655 ;
        RECT 580.605 361.375 580.885 361.655 ;
        RECT 581.315 361.375 581.595 361.655 ;
        RECT 582.025 361.375 582.305 361.655 ;
        RECT 582.735 361.375 583.015 361.655 ;
        RECT 583.445 361.375 583.725 361.655 ;
        RECT 584.155 361.375 584.435 361.655 ;
        RECT 584.865 361.375 585.145 361.655 ;
        RECT 585.575 361.375 585.855 361.655 ;
        RECT 589.495 361.375 589.775 361.655 ;
        RECT 590.205 361.375 590.485 361.655 ;
        RECT 590.915 361.375 591.195 361.655 ;
        RECT 591.625 361.375 591.905 361.655 ;
        RECT 592.335 361.375 592.615 361.655 ;
        RECT 593.045 361.375 593.325 361.655 ;
        RECT 593.755 361.375 594.035 361.655 ;
        RECT 594.465 361.375 594.745 361.655 ;
        RECT 595.175 361.375 595.455 361.655 ;
        RECT 595.885 361.375 596.165 361.655 ;
        RECT 596.595 361.375 596.875 361.655 ;
        RECT 597.305 361.375 597.585 361.655 ;
        RECT 598.015 361.375 598.295 361.655 ;
        RECT 1351.715 361.375 1351.995 361.655 ;
        RECT 1352.425 361.375 1352.705 361.655 ;
        RECT 1353.135 361.375 1353.415 361.655 ;
        RECT 1353.845 361.375 1354.125 361.655 ;
        RECT 1354.555 361.375 1354.835 361.655 ;
        RECT 1355.265 361.375 1355.545 361.655 ;
        RECT 1355.975 361.375 1356.255 361.655 ;
        RECT 1356.685 361.375 1356.965 361.655 ;
        RECT 1357.395 361.375 1357.675 361.655 ;
        RECT 1358.105 361.375 1358.385 361.655 ;
        RECT 1358.815 361.375 1359.095 361.655 ;
        RECT 1359.525 361.375 1359.805 361.655 ;
        RECT 1360.235 361.375 1360.515 361.655 ;
        RECT 1366.245 361.375 1366.525 361.655 ;
        RECT 1366.955 361.375 1367.235 361.655 ;
        RECT 1367.665 361.375 1367.945 361.655 ;
        RECT 1368.375 361.375 1368.655 361.655 ;
        RECT 1369.085 361.375 1369.365 361.655 ;
        RECT 1369.795 361.375 1370.075 361.655 ;
        RECT 1370.505 361.375 1370.785 361.655 ;
        RECT 1371.215 361.375 1371.495 361.655 ;
        RECT 1371.925 361.375 1372.205 361.655 ;
        RECT 1372.635 361.375 1372.915 361.655 ;
        RECT 1373.345 361.375 1373.625 361.655 ;
        RECT 1375.965 361.375 1376.245 361.655 ;
        RECT 1376.675 361.375 1376.955 361.655 ;
        RECT 1377.385 361.375 1377.665 361.655 ;
        RECT 1378.095 361.375 1378.375 361.655 ;
        RECT 1378.805 361.375 1379.085 361.655 ;
        RECT 1379.515 361.375 1379.795 361.655 ;
        RECT 1380.225 361.375 1380.505 361.655 ;
        RECT 1380.935 361.375 1381.215 361.655 ;
        RECT 1381.645 361.375 1381.925 361.655 ;
        RECT 1382.355 361.375 1382.635 361.655 ;
        RECT 1383.065 361.375 1383.345 361.655 ;
        RECT 1383.775 361.375 1384.055 361.655 ;
        RECT 1384.485 361.375 1384.765 361.655 ;
        RECT 1385.195 361.375 1385.475 361.655 ;
        RECT 1389.495 361.375 1389.775 361.655 ;
        RECT 1390.205 361.375 1390.485 361.655 ;
        RECT 1390.915 361.375 1391.195 361.655 ;
        RECT 1391.625 361.375 1391.905 361.655 ;
        RECT 1392.335 361.375 1392.615 361.655 ;
        RECT 1393.045 361.375 1393.325 361.655 ;
        RECT 1393.755 361.375 1394.035 361.655 ;
        RECT 1394.465 361.375 1394.745 361.655 ;
        RECT 1395.175 361.375 1395.455 361.655 ;
        RECT 1395.885 361.375 1396.165 361.655 ;
        RECT 1396.595 361.375 1396.875 361.655 ;
        RECT 1397.305 361.375 1397.585 361.655 ;
        RECT 1398.015 361.375 1398.295 361.655 ;
        RECT 1398.725 361.375 1399.005 361.655 ;
        RECT 1401.345 361.375 1401.625 361.655 ;
        RECT 1402.055 361.375 1402.335 361.655 ;
        RECT 1402.765 361.375 1403.045 361.655 ;
        RECT 1403.475 361.375 1403.755 361.655 ;
        RECT 1404.185 361.375 1404.465 361.655 ;
        RECT 1404.895 361.375 1405.175 361.655 ;
        RECT 1405.605 361.375 1405.885 361.655 ;
        RECT 1406.315 361.375 1406.595 361.655 ;
        RECT 1407.025 361.375 1407.305 361.655 ;
        RECT 1407.735 361.375 1408.015 361.655 ;
        RECT 1408.445 361.375 1408.725 361.655 ;
        RECT 1409.155 361.375 1409.435 361.655 ;
        RECT 1409.865 361.375 1410.145 361.655 ;
        RECT 1410.575 361.375 1410.855 361.655 ;
        RECT 1414.495 361.375 1414.775 361.655 ;
        RECT 1415.205 361.375 1415.485 361.655 ;
        RECT 1415.915 361.375 1416.195 361.655 ;
        RECT 1416.625 361.375 1416.905 361.655 ;
        RECT 1417.335 361.375 1417.615 361.655 ;
        RECT 1418.045 361.375 1418.325 361.655 ;
        RECT 1418.755 361.375 1419.035 361.655 ;
        RECT 1419.465 361.375 1419.745 361.655 ;
        RECT 3001.715 361.375 3001.995 361.655 ;
        RECT 3002.425 361.375 3002.705 361.655 ;
        RECT 3003.135 361.375 3003.415 361.655 ;
        RECT 3003.845 361.375 3004.125 361.655 ;
        RECT 3004.555 361.375 3004.835 361.655 ;
        RECT 3005.265 361.375 3005.545 361.655 ;
        RECT 3005.975 361.375 3006.255 361.655 ;
        RECT 3006.685 361.375 3006.965 361.655 ;
        RECT 3007.395 361.375 3007.675 361.655 ;
        RECT 3008.105 361.375 3008.385 361.655 ;
        RECT 3008.815 361.375 3009.095 361.655 ;
        RECT 3009.525 361.375 3009.805 361.655 ;
        RECT 3010.235 361.375 3010.515 361.655 ;
        RECT 3014.115 361.375 3014.395 361.655 ;
        RECT 3014.825 361.375 3015.105 361.655 ;
        RECT 3015.535 361.375 3015.815 361.655 ;
        RECT 3016.245 361.375 3016.525 361.655 ;
        RECT 3016.955 361.375 3017.235 361.655 ;
        RECT 3017.665 361.375 3017.945 361.655 ;
        RECT 3018.375 361.375 3018.655 361.655 ;
        RECT 3019.085 361.375 3019.365 361.655 ;
        RECT 3019.795 361.375 3020.075 361.655 ;
        RECT 3025.965 361.375 3026.245 361.655 ;
        RECT 3026.675 361.375 3026.955 361.655 ;
        RECT 3027.385 361.375 3027.665 361.655 ;
        RECT 3028.095 361.375 3028.375 361.655 ;
        RECT 3028.805 361.375 3029.085 361.655 ;
        RECT 3029.515 361.375 3029.795 361.655 ;
        RECT 3030.225 361.375 3030.505 361.655 ;
        RECT 3030.935 361.375 3031.215 361.655 ;
        RECT 3031.645 361.375 3031.925 361.655 ;
        RECT 3032.355 361.375 3032.635 361.655 ;
        RECT 3033.065 361.375 3033.345 361.655 ;
        RECT 3033.775 361.375 3034.055 361.655 ;
        RECT 3034.485 361.375 3034.765 361.655 ;
        RECT 3035.195 361.375 3035.475 361.655 ;
        RECT 3039.495 361.375 3039.775 361.655 ;
        RECT 3040.205 361.375 3040.485 361.655 ;
        RECT 3040.915 361.375 3041.195 361.655 ;
        RECT 3041.625 361.375 3041.905 361.655 ;
        RECT 3042.335 361.375 3042.615 361.655 ;
        RECT 3046.595 361.375 3046.875 361.655 ;
        RECT 3047.305 361.375 3047.585 361.655 ;
        RECT 3048.015 361.375 3048.295 361.655 ;
        RECT 3048.725 361.375 3049.005 361.655 ;
        RECT 3051.345 361.375 3051.625 361.655 ;
        RECT 3052.055 361.375 3052.335 361.655 ;
        RECT 3052.765 361.375 3053.045 361.655 ;
        RECT 3053.475 361.375 3053.755 361.655 ;
        RECT 3054.185 361.375 3054.465 361.655 ;
        RECT 3054.895 361.375 3055.175 361.655 ;
        RECT 3055.605 361.375 3055.885 361.655 ;
        RECT 3056.315 361.375 3056.595 361.655 ;
        RECT 3057.025 361.375 3057.305 361.655 ;
        RECT 3057.735 361.375 3058.015 361.655 ;
        RECT 3058.445 361.375 3058.725 361.655 ;
        RECT 3059.155 361.375 3059.435 361.655 ;
        RECT 3059.865 361.375 3060.145 361.655 ;
        RECT 3060.575 361.375 3060.855 361.655 ;
        RECT 3064.495 361.375 3064.775 361.655 ;
        RECT 3065.205 361.375 3065.485 361.655 ;
        RECT 3065.915 361.375 3066.195 361.655 ;
        RECT 3066.625 361.375 3066.905 361.655 ;
        RECT 3067.335 361.375 3067.615 361.655 ;
        RECT 3068.045 361.375 3068.325 361.655 ;
        RECT 3068.755 361.375 3069.035 361.655 ;
        RECT 3069.465 361.375 3069.745 361.655 ;
        RECT 3070.175 361.375 3070.455 361.655 ;
        RECT 3070.885 361.375 3071.165 361.655 ;
        RECT 3071.595 361.375 3071.875 361.655 ;
        RECT 3072.305 361.375 3072.585 361.655 ;
        RECT 3073.015 361.375 3073.295 361.655 ;
        RECT 526.715 360.665 526.995 360.945 ;
        RECT 527.425 360.665 527.705 360.945 ;
        RECT 528.135 360.665 528.415 360.945 ;
        RECT 528.845 360.665 529.125 360.945 ;
        RECT 529.555 360.665 529.835 360.945 ;
        RECT 530.265 360.665 530.545 360.945 ;
        RECT 530.975 360.665 531.255 360.945 ;
        RECT 531.685 360.665 531.965 360.945 ;
        RECT 532.395 360.665 532.675 360.945 ;
        RECT 533.105 360.665 533.385 360.945 ;
        RECT 533.815 360.665 534.095 360.945 ;
        RECT 534.525 360.665 534.805 360.945 ;
        RECT 535.235 360.665 535.515 360.945 ;
        RECT 544.975 360.665 545.255 360.945 ;
        RECT 545.685 360.665 545.965 360.945 ;
        RECT 546.395 360.665 546.675 360.945 ;
        RECT 547.105 360.665 547.385 360.945 ;
        RECT 547.815 360.665 548.095 360.945 ;
        RECT 548.525 360.665 548.805 360.945 ;
        RECT 550.965 360.665 551.245 360.945 ;
        RECT 551.675 360.665 551.955 360.945 ;
        RECT 552.385 360.665 552.665 360.945 ;
        RECT 553.095 360.665 553.375 360.945 ;
        RECT 553.805 360.665 554.085 360.945 ;
        RECT 554.515 360.665 554.795 360.945 ;
        RECT 555.225 360.665 555.505 360.945 ;
        RECT 555.935 360.665 556.215 360.945 ;
        RECT 556.645 360.665 556.925 360.945 ;
        RECT 557.355 360.665 557.635 360.945 ;
        RECT 558.065 360.665 558.345 360.945 ;
        RECT 558.775 360.665 559.055 360.945 ;
        RECT 559.485 360.665 559.765 360.945 ;
        RECT 560.195 360.665 560.475 360.945 ;
        RECT 566.625 360.665 566.905 360.945 ;
        RECT 567.335 360.665 567.615 360.945 ;
        RECT 568.045 360.665 568.325 360.945 ;
        RECT 568.755 360.665 569.035 360.945 ;
        RECT 569.465 360.665 569.745 360.945 ;
        RECT 570.175 360.665 570.455 360.945 ;
        RECT 570.885 360.665 571.165 360.945 ;
        RECT 571.595 360.665 571.875 360.945 ;
        RECT 572.305 360.665 572.585 360.945 ;
        RECT 573.015 360.665 573.295 360.945 ;
        RECT 573.725 360.665 574.005 360.945 ;
        RECT 576.345 360.665 576.625 360.945 ;
        RECT 577.055 360.665 577.335 360.945 ;
        RECT 577.765 360.665 578.045 360.945 ;
        RECT 578.475 360.665 578.755 360.945 ;
        RECT 579.185 360.665 579.465 360.945 ;
        RECT 579.895 360.665 580.175 360.945 ;
        RECT 580.605 360.665 580.885 360.945 ;
        RECT 581.315 360.665 581.595 360.945 ;
        RECT 582.025 360.665 582.305 360.945 ;
        RECT 582.735 360.665 583.015 360.945 ;
        RECT 583.445 360.665 583.725 360.945 ;
        RECT 584.155 360.665 584.435 360.945 ;
        RECT 584.865 360.665 585.145 360.945 ;
        RECT 585.575 360.665 585.855 360.945 ;
        RECT 589.495 360.665 589.775 360.945 ;
        RECT 590.205 360.665 590.485 360.945 ;
        RECT 590.915 360.665 591.195 360.945 ;
        RECT 591.625 360.665 591.905 360.945 ;
        RECT 592.335 360.665 592.615 360.945 ;
        RECT 593.045 360.665 593.325 360.945 ;
        RECT 593.755 360.665 594.035 360.945 ;
        RECT 594.465 360.665 594.745 360.945 ;
        RECT 595.175 360.665 595.455 360.945 ;
        RECT 595.885 360.665 596.165 360.945 ;
        RECT 596.595 360.665 596.875 360.945 ;
        RECT 597.305 360.665 597.585 360.945 ;
        RECT 598.015 360.665 598.295 360.945 ;
        RECT 1351.715 360.665 1351.995 360.945 ;
        RECT 1352.425 360.665 1352.705 360.945 ;
        RECT 1353.135 360.665 1353.415 360.945 ;
        RECT 1353.845 360.665 1354.125 360.945 ;
        RECT 1354.555 360.665 1354.835 360.945 ;
        RECT 1355.265 360.665 1355.545 360.945 ;
        RECT 1355.975 360.665 1356.255 360.945 ;
        RECT 1356.685 360.665 1356.965 360.945 ;
        RECT 1357.395 360.665 1357.675 360.945 ;
        RECT 1358.105 360.665 1358.385 360.945 ;
        RECT 1358.815 360.665 1359.095 360.945 ;
        RECT 1359.525 360.665 1359.805 360.945 ;
        RECT 1360.235 360.665 1360.515 360.945 ;
        RECT 1366.245 360.665 1366.525 360.945 ;
        RECT 1366.955 360.665 1367.235 360.945 ;
        RECT 1367.665 360.665 1367.945 360.945 ;
        RECT 1368.375 360.665 1368.655 360.945 ;
        RECT 1369.085 360.665 1369.365 360.945 ;
        RECT 1369.795 360.665 1370.075 360.945 ;
        RECT 1370.505 360.665 1370.785 360.945 ;
        RECT 1371.215 360.665 1371.495 360.945 ;
        RECT 1371.925 360.665 1372.205 360.945 ;
        RECT 1372.635 360.665 1372.915 360.945 ;
        RECT 1373.345 360.665 1373.625 360.945 ;
        RECT 1375.965 360.665 1376.245 360.945 ;
        RECT 1376.675 360.665 1376.955 360.945 ;
        RECT 1377.385 360.665 1377.665 360.945 ;
        RECT 1378.095 360.665 1378.375 360.945 ;
        RECT 1378.805 360.665 1379.085 360.945 ;
        RECT 1379.515 360.665 1379.795 360.945 ;
        RECT 1380.225 360.665 1380.505 360.945 ;
        RECT 1380.935 360.665 1381.215 360.945 ;
        RECT 1381.645 360.665 1381.925 360.945 ;
        RECT 1382.355 360.665 1382.635 360.945 ;
        RECT 1383.065 360.665 1383.345 360.945 ;
        RECT 1383.775 360.665 1384.055 360.945 ;
        RECT 1384.485 360.665 1384.765 360.945 ;
        RECT 1385.195 360.665 1385.475 360.945 ;
        RECT 1389.495 360.665 1389.775 360.945 ;
        RECT 1390.205 360.665 1390.485 360.945 ;
        RECT 1390.915 360.665 1391.195 360.945 ;
        RECT 1391.625 360.665 1391.905 360.945 ;
        RECT 1392.335 360.665 1392.615 360.945 ;
        RECT 1393.045 360.665 1393.325 360.945 ;
        RECT 1393.755 360.665 1394.035 360.945 ;
        RECT 1394.465 360.665 1394.745 360.945 ;
        RECT 1395.175 360.665 1395.455 360.945 ;
        RECT 1395.885 360.665 1396.165 360.945 ;
        RECT 1396.595 360.665 1396.875 360.945 ;
        RECT 1397.305 360.665 1397.585 360.945 ;
        RECT 1398.015 360.665 1398.295 360.945 ;
        RECT 1398.725 360.665 1399.005 360.945 ;
        RECT 1401.345 360.665 1401.625 360.945 ;
        RECT 1402.055 360.665 1402.335 360.945 ;
        RECT 1402.765 360.665 1403.045 360.945 ;
        RECT 1403.475 360.665 1403.755 360.945 ;
        RECT 1404.185 360.665 1404.465 360.945 ;
        RECT 1404.895 360.665 1405.175 360.945 ;
        RECT 1405.605 360.665 1405.885 360.945 ;
        RECT 1406.315 360.665 1406.595 360.945 ;
        RECT 1407.025 360.665 1407.305 360.945 ;
        RECT 1407.735 360.665 1408.015 360.945 ;
        RECT 1408.445 360.665 1408.725 360.945 ;
        RECT 1409.155 360.665 1409.435 360.945 ;
        RECT 1409.865 360.665 1410.145 360.945 ;
        RECT 1410.575 360.665 1410.855 360.945 ;
        RECT 1414.495 360.665 1414.775 360.945 ;
        RECT 1415.205 360.665 1415.485 360.945 ;
        RECT 1415.915 360.665 1416.195 360.945 ;
        RECT 1416.625 360.665 1416.905 360.945 ;
        RECT 1417.335 360.665 1417.615 360.945 ;
        RECT 1418.045 360.665 1418.325 360.945 ;
        RECT 1418.755 360.665 1419.035 360.945 ;
        RECT 1419.465 360.665 1419.745 360.945 ;
        RECT 3001.715 360.665 3001.995 360.945 ;
        RECT 3002.425 360.665 3002.705 360.945 ;
        RECT 3003.135 360.665 3003.415 360.945 ;
        RECT 3003.845 360.665 3004.125 360.945 ;
        RECT 3004.555 360.665 3004.835 360.945 ;
        RECT 3005.265 360.665 3005.545 360.945 ;
        RECT 3005.975 360.665 3006.255 360.945 ;
        RECT 3006.685 360.665 3006.965 360.945 ;
        RECT 3007.395 360.665 3007.675 360.945 ;
        RECT 3008.105 360.665 3008.385 360.945 ;
        RECT 3008.815 360.665 3009.095 360.945 ;
        RECT 3009.525 360.665 3009.805 360.945 ;
        RECT 3010.235 360.665 3010.515 360.945 ;
        RECT 3014.115 360.665 3014.395 360.945 ;
        RECT 3014.825 360.665 3015.105 360.945 ;
        RECT 3015.535 360.665 3015.815 360.945 ;
        RECT 3016.245 360.665 3016.525 360.945 ;
        RECT 3016.955 360.665 3017.235 360.945 ;
        RECT 3017.665 360.665 3017.945 360.945 ;
        RECT 3018.375 360.665 3018.655 360.945 ;
        RECT 3019.085 360.665 3019.365 360.945 ;
        RECT 3019.795 360.665 3020.075 360.945 ;
        RECT 3025.965 360.665 3026.245 360.945 ;
        RECT 3026.675 360.665 3026.955 360.945 ;
        RECT 3027.385 360.665 3027.665 360.945 ;
        RECT 3028.095 360.665 3028.375 360.945 ;
        RECT 3028.805 360.665 3029.085 360.945 ;
        RECT 3029.515 360.665 3029.795 360.945 ;
        RECT 3030.225 360.665 3030.505 360.945 ;
        RECT 3030.935 360.665 3031.215 360.945 ;
        RECT 3031.645 360.665 3031.925 360.945 ;
        RECT 3032.355 360.665 3032.635 360.945 ;
        RECT 3033.065 360.665 3033.345 360.945 ;
        RECT 3033.775 360.665 3034.055 360.945 ;
        RECT 3034.485 360.665 3034.765 360.945 ;
        RECT 3035.195 360.665 3035.475 360.945 ;
        RECT 3039.495 360.665 3039.775 360.945 ;
        RECT 3040.205 360.665 3040.485 360.945 ;
        RECT 3040.915 360.665 3041.195 360.945 ;
        RECT 3041.625 360.665 3041.905 360.945 ;
        RECT 3042.335 360.665 3042.615 360.945 ;
        RECT 3046.595 360.665 3046.875 360.945 ;
        RECT 3047.305 360.665 3047.585 360.945 ;
        RECT 3048.015 360.665 3048.295 360.945 ;
        RECT 3048.725 360.665 3049.005 360.945 ;
        RECT 3051.345 360.665 3051.625 360.945 ;
        RECT 3052.055 360.665 3052.335 360.945 ;
        RECT 3052.765 360.665 3053.045 360.945 ;
        RECT 3053.475 360.665 3053.755 360.945 ;
        RECT 3054.185 360.665 3054.465 360.945 ;
        RECT 3054.895 360.665 3055.175 360.945 ;
        RECT 3055.605 360.665 3055.885 360.945 ;
        RECT 3056.315 360.665 3056.595 360.945 ;
        RECT 3057.025 360.665 3057.305 360.945 ;
        RECT 3057.735 360.665 3058.015 360.945 ;
        RECT 3058.445 360.665 3058.725 360.945 ;
        RECT 3059.155 360.665 3059.435 360.945 ;
        RECT 3059.865 360.665 3060.145 360.945 ;
        RECT 3060.575 360.665 3060.855 360.945 ;
        RECT 3064.495 360.665 3064.775 360.945 ;
        RECT 3065.205 360.665 3065.485 360.945 ;
        RECT 3065.915 360.665 3066.195 360.945 ;
        RECT 3066.625 360.665 3066.905 360.945 ;
        RECT 3067.335 360.665 3067.615 360.945 ;
        RECT 3068.045 360.665 3068.325 360.945 ;
        RECT 3068.755 360.665 3069.035 360.945 ;
        RECT 3069.465 360.665 3069.745 360.945 ;
        RECT 3070.175 360.665 3070.455 360.945 ;
        RECT 3070.885 360.665 3071.165 360.945 ;
        RECT 3071.595 360.665 3071.875 360.945 ;
        RECT 3072.305 360.665 3072.585 360.945 ;
        RECT 3073.015 360.665 3073.295 360.945 ;
  END
END caravel_power_routing
END LIBRARY

