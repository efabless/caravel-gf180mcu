magic
tech gf180mcuD
magscale 1 10
timestamp 1655307388
<< pwell >>
rect -334 -432 334 432
<< mvnmos >>
rect -70 -224 70 176
<< mvndiff >>
rect -158 163 -70 176
rect -158 -211 -145 163
rect -99 -211 -70 163
rect -158 -224 -70 -211
rect 70 163 158 176
rect 70 -211 99 163
rect 145 -211 158 163
rect 70 -224 158 -211
<< mvndiffc >>
rect -145 -211 -99 163
rect 99 -211 145 163
<< mvpsubdiff >>
rect -302 328 302 400
rect -302 284 -230 328
rect -302 -284 -289 284
rect -243 -284 -230 284
rect 230 284 302 328
rect -302 -328 -230 -284
rect 230 -284 243 284
rect 289 -284 302 284
rect 230 -328 302 -284
rect -302 -341 302 -328
rect -302 -387 -186 -341
rect 186 -387 302 -341
rect -302 -400 302 -387
<< mvpsubdiffcont >>
rect -289 -284 -243 284
rect 243 -284 289 284
rect -186 -387 186 -341
<< polysilicon >>
rect -70 255 70 268
rect -70 209 -57 255
rect 57 209 70 255
rect -70 176 70 209
rect -70 -268 70 -224
<< polycontact >>
rect -57 209 57 255
<< metal1 >>
rect -289 341 289 387
rect -289 284 -243 341
rect 243 284 289 341
rect -68 209 -57 255
rect 57 209 68 255
rect -145 163 -99 174
rect -145 -222 -99 -211
rect 99 163 145 174
rect 99 -222 145 -211
rect -289 -341 -243 -284
rect 243 -341 289 -284
rect -289 -387 -186 -341
rect 186 -387 289 -341
<< properties >>
string FIXED_BBOX -266 -364 266 364
string gencell nmos_6p0
string library gf180mcu
string parameters w 2.0 l 0.7 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.6 wmin 0.3 full_metal 1 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
