magic
tech gf180mcuC
magscale 1 10
timestamp 1655302813
<< checkpaint >>
rect -2000 1008903 73000 1022000
rect 103968 1008903 123032 1022000
rect 158968 1008903 178032 1022000
rect 213968 1008903 233032 1022000
rect 268968 1008903 288032 1022000
rect 323968 1008903 343032 1022000
rect 378968 1008903 398032 1022000
rect 433968 1008903 453032 1022000
rect 488968 1008903 508032 1022000
rect 543968 1008903 563032 1022000
rect 598968 1008903 618032 1022000
rect 653968 1008903 673032 1022000
rect 705000 1008903 780000 1022000
rect -2000 948032 780000 1008903
rect -2000 947000 73000 948032
rect 103968 948000 123032 948032
rect 158968 948000 178032 948032
rect 213968 948000 233032 948032
rect 268968 948000 288032 948032
rect 323968 948000 343032 948032
rect 378968 948000 398032 948032
rect 433968 948000 453032 948032
rect 488968 948000 508032 948032
rect 543968 948000 563032 948032
rect 598968 948000 618032 948032
rect 653968 948000 673032 948032
rect 705000 947000 780000 948032
rect 11097 928032 71968 947000
rect 706032 929032 766903 947000
rect -2000 908968 72000 928032
rect 706000 909968 780000 929032
rect 11097 887032 71968 908968
rect -2000 867968 72000 887032
rect 706032 886032 766903 909968
rect 11097 846032 71968 867968
rect 706000 866968 780000 886032
rect -2000 826968 72000 846032
rect 706032 843032 766903 866968
rect 11097 805032 71968 826968
rect 706000 823968 780000 843032
rect -2000 785968 72000 805032
rect 706032 800032 766903 823968
rect 11097 764032 71968 785968
rect 706000 780968 780000 800032
rect -2000 744968 72000 764032
rect 706032 757032 766903 780968
rect 11097 723032 71968 744968
rect 706000 737968 780000 757032
rect -2000 703968 72000 723032
rect 706032 714032 766903 737968
rect 11097 682032 71968 703968
rect 706000 694968 780000 714032
rect -2000 662968 72000 682032
rect 706032 671032 766903 694968
rect 11097 641032 71968 662968
rect 706000 651968 780000 671032
rect -2000 621968 72000 641032
rect 706032 628032 766903 651968
rect 11097 600032 71968 621968
rect 706000 608968 780000 628032
rect -2000 580968 72000 600032
rect 706032 585032 766903 608968
rect 11097 559032 71968 580968
rect 706000 565968 780000 585032
rect -2000 539968 72000 559032
rect 706032 542032 766903 565968
rect 11097 518032 71968 539968
rect 706000 522968 780000 542032
rect -2000 498968 72000 518032
rect 706032 499032 766903 522968
rect 11097 477032 71968 498968
rect 706000 479968 780000 499032
rect -2000 457968 72000 477032
rect 11097 436032 71968 457968
rect 706032 456032 766903 479968
rect 706000 436968 780000 456032
rect -2000 416968 72000 436032
rect 11097 395032 71968 416968
rect 706032 413032 766903 436968
rect -2000 375968 72000 395032
rect 706000 393968 780000 413032
rect 11097 354032 71968 375968
rect 706032 370032 766903 393968
rect -2000 334968 72000 354032
rect 706000 350968 780000 370032
rect 11097 313032 71968 334968
rect 706032 327032 766903 350968
rect -2000 293968 72000 313032
rect 706000 307968 780000 327032
rect 11097 272032 71968 293968
rect 706032 284032 766903 307968
rect -2000 252968 72000 272032
rect 706000 264968 780000 284032
rect 11097 231032 71968 252968
rect 706032 241032 766903 264968
rect -2000 211968 72000 231032
rect 706000 221968 780000 241032
rect 11097 190032 71968 211968
rect 706032 198032 766903 221968
rect -2000 170968 72000 190032
rect 706000 178968 780000 198032
rect 11097 149032 71968 170968
rect 706032 155032 766903 178968
rect 706000 154330 780000 155032
rect 705730 149690 780000 154330
rect -2000 129968 72000 149032
rect 706000 142390 780000 149690
rect 705770 136600 780000 142390
rect 706000 135968 780000 136600
rect 11097 108032 71968 129968
rect 706032 112032 766903 135968
rect -2000 88968 72000 108032
rect 706000 92968 780000 112032
rect 11097 73000 71968 88968
rect 706032 73000 766903 92968
rect -2000 71968 73000 73000
rect 104968 71968 124032 72000
rect 159968 71968 179032 72000
rect 214968 71968 234032 72000
rect 269968 71968 289032 72000
rect 324968 71968 344032 72000
rect 379968 71968 399032 72000
rect 434968 71968 454032 72000
rect 489968 71968 509032 72000
rect 544968 71968 564032 72000
rect 599968 71968 619032 72000
rect 654968 71968 674032 72000
rect 705000 71968 780000 73000
rect -2000 11097 780000 71968
rect -2000 -2000 73000 11097
rect 104968 -2000 124032 11097
rect 159968 -2000 179032 11097
rect 214968 -2000 234032 11097
rect 269968 -2000 289032 11097
rect 324968 -2000 344032 11097
rect 379968 -2000 399032 11097
rect 434968 -2000 454032 11097
rect 489968 -2000 509032 11097
rect 544968 -2000 564032 11097
rect 599968 -2000 619032 11097
rect 654968 -2000 674032 11097
rect 705000 -2000 780000 11097
<< metal2 >>
rect 106752 949800 106828 950076
rect 106898 949800 106974 950076
rect 107044 949800 107120 950076
rect 107190 949800 107266 950076
rect 118647 949800 118723 950076
rect 118858 949800 118934 950076
rect 119360 949800 119436 950076
rect 119502 949800 119578 950076
rect 119731 949800 119807 950076
rect 120252 949800 120328 950076
rect 161752 949800 161828 950076
rect 161898 949800 161974 950076
rect 162044 949800 162120 950076
rect 162190 949800 162266 950076
rect 173647 949800 173723 950076
rect 173858 949800 173934 950076
rect 174360 949800 174436 950076
rect 174502 949800 174578 950076
rect 174731 949800 174807 950076
rect 175252 949800 175328 950076
rect 216752 949800 216828 950076
rect 216898 949800 216974 950076
rect 217044 949800 217120 950076
rect 217190 949800 217266 950076
rect 228647 949800 228723 950076
rect 228858 949800 228934 950076
rect 229360 949800 229436 950076
rect 229502 949800 229578 950076
rect 229731 949800 229807 950076
rect 230252 949800 230328 950076
rect 271752 949800 271828 950076
rect 271898 949800 271974 950076
rect 272044 949800 272120 950076
rect 272190 949800 272266 950076
rect 283647 949800 283723 950076
rect 283858 949800 283934 950076
rect 284360 949800 284436 950076
rect 284502 949800 284578 950076
rect 284731 949800 284807 950076
rect 285252 949800 285328 950076
rect 326752 949800 326828 950076
rect 326898 949800 326974 950076
rect 327044 949800 327120 950076
rect 327190 949800 327266 950076
rect 338647 949800 338723 950076
rect 338858 949800 338934 950076
rect 339360 949800 339436 950076
rect 339502 949800 339578 950076
rect 339731 949800 339807 950076
rect 340252 949800 340328 950076
rect 436752 949800 436828 950076
rect 436898 949800 436974 950076
rect 437044 949800 437120 950076
rect 437190 949800 437266 950076
rect 448647 949800 448723 950076
rect 448858 949800 448934 950076
rect 449360 949800 449436 950076
rect 449502 949800 449578 950076
rect 449731 949800 449807 950076
rect 450252 949800 450328 950076
rect 491752 949800 491828 950076
rect 491898 949800 491974 950076
rect 492044 949800 492120 950076
rect 492190 949800 492266 950076
rect 503647 949800 503723 950076
rect 503858 949800 503934 950076
rect 504360 949800 504436 950076
rect 504502 949800 504578 950076
rect 504731 949800 504807 950076
rect 505252 949800 505328 950076
rect 546752 949800 546828 950076
rect 546898 949800 546974 950076
rect 547044 949800 547120 950076
rect 547190 949800 547266 950076
rect 558647 949800 558723 950076
rect 558858 949800 558934 950076
rect 559360 949800 559436 950076
rect 559502 949800 559578 950076
rect 559731 949800 559807 950076
rect 560252 949800 560328 950076
rect 656752 949800 656828 950076
rect 656898 949800 656974 950076
rect 657044 949800 657120 950076
rect 657190 949800 657266 950076
rect 668647 949800 668723 950076
rect 668858 949800 668934 950076
rect 669360 949800 669436 950076
rect 669502 949800 669578 950076
rect 669731 949800 669807 950076
rect 670252 949800 670328 950076
rect 707800 926172 708076 926248
rect 707800 926026 708076 926102
rect 707800 925880 708076 925956
rect 707800 925734 708076 925810
rect 69924 925252 70200 925328
rect 69924 924731 70200 924807
rect 69924 924502 70200 924578
rect 69924 924360 70200 924436
rect 69924 923858 70200 923934
rect 69924 923647 70200 923723
rect 707800 914277 708076 914353
rect 707800 914066 708076 914142
rect 707800 913564 708076 913640
rect 707800 913422 708076 913498
rect 707800 913193 708076 913269
rect 707800 912672 708076 912748
rect 69924 912190 70200 912266
rect 69924 912044 70200 912120
rect 69924 911898 70200 911974
rect 69924 911752 70200 911828
rect 707800 840172 708076 840248
rect 707800 840026 708076 840102
rect 707800 839880 708076 839956
rect 707800 839734 708076 839810
rect 707800 828277 708076 828353
rect 707800 828066 708076 828142
rect 707800 827564 708076 827640
rect 707800 827422 708076 827498
rect 707800 827193 708076 827269
rect 707800 826672 708076 826748
rect 69924 761252 70200 761328
rect 69924 760731 70200 760807
rect 69924 760502 70200 760578
rect 69924 760360 70200 760436
rect 69924 759858 70200 759934
rect 69924 759647 70200 759723
rect 707800 754172 708076 754248
rect 707800 754026 708076 754102
rect 707800 753880 708076 753956
rect 707800 753734 708076 753810
rect 69924 748190 70200 748266
rect 69924 748044 70200 748120
rect 69924 747898 70200 747974
rect 69924 747752 70200 747828
rect 707800 742277 708076 742353
rect 707800 742066 708076 742142
rect 707800 741564 708076 741640
rect 707800 741422 708076 741498
rect 707800 741193 708076 741269
rect 707800 740672 708076 740748
rect 69924 720252 70200 720328
rect 69924 719731 70200 719807
rect 69924 719502 70200 719578
rect 69924 719360 70200 719436
rect 69924 718858 70200 718934
rect 69924 718647 70200 718723
rect 707800 711172 708076 711248
rect 707800 711026 708076 711102
rect 707800 710880 708076 710956
rect 707800 710734 708076 710810
rect 69924 707190 70200 707266
rect 69924 707044 70200 707120
rect 69924 706898 70200 706974
rect 69924 706752 70200 706828
rect 707800 699277 708076 699353
rect 707800 699066 708076 699142
rect 707800 698564 708076 698640
rect 707800 698422 708076 698498
rect 707800 698193 708076 698269
rect 707800 697672 708076 697748
rect 69924 679252 70200 679328
rect 69924 678731 70200 678807
rect 69924 678502 70200 678578
rect 69924 678360 70200 678436
rect 69924 677858 70200 677934
rect 69924 677647 70200 677723
rect 707800 668172 708076 668248
rect 707800 668026 708076 668102
rect 707800 667880 708076 667956
rect 707800 667734 708076 667810
rect 69924 666190 70200 666266
rect 69924 666044 70200 666120
rect 69924 665898 70200 665974
rect 69924 665752 70200 665828
rect 707800 656277 708076 656353
rect 707800 656066 708076 656142
rect 707800 655564 708076 655640
rect 707800 655422 708076 655498
rect 707800 655193 708076 655269
rect 707800 654672 708076 654748
rect 69924 638252 70200 638328
rect 69924 637731 70200 637807
rect 69924 637502 70200 637578
rect 69924 637360 70200 637436
rect 69924 636858 70200 636934
rect 69924 636647 70200 636723
rect 69924 625190 70200 625266
rect 707800 625172 708076 625248
rect 69924 625044 70200 625120
rect 707800 625026 708076 625102
rect 69924 624898 70200 624974
rect 707800 624880 708076 624956
rect 69924 624752 70200 624828
rect 707800 624734 708076 624810
rect 707800 613277 708076 613353
rect 707800 613066 708076 613142
rect 707800 612564 708076 612640
rect 707800 612422 708076 612498
rect 707800 612193 708076 612269
rect 707800 611672 708076 611748
rect 69924 597252 70200 597328
rect 69924 596731 70200 596807
rect 69924 596502 70200 596578
rect 69924 596360 70200 596436
rect 69924 595858 70200 595934
rect 69924 595647 70200 595723
rect 69924 584190 70200 584266
rect 69924 584044 70200 584120
rect 69924 583898 70200 583974
rect 69924 583752 70200 583828
rect 707800 582172 708076 582248
rect 707800 582026 708076 582102
rect 707800 581880 708076 581956
rect 707800 581734 708076 581810
rect 707800 570277 708076 570353
rect 707800 570066 708076 570142
rect 707800 569564 708076 569640
rect 707800 569422 708076 569498
rect 707800 569193 708076 569269
rect 707800 568672 708076 568748
rect 69924 556252 70200 556328
rect 69924 555731 70200 555807
rect 69924 555502 70200 555578
rect 69924 555360 70200 555436
rect 69924 554858 70200 554934
rect 69924 554647 70200 554723
rect 69924 543190 70200 543266
rect 69924 543044 70200 543120
rect 69924 542898 70200 542974
rect 69924 542752 70200 542828
rect 707800 539172 708076 539248
rect 707800 539026 708076 539102
rect 707800 538880 708076 538956
rect 707800 538734 708076 538810
rect 707800 527277 708076 527353
rect 707800 527066 708076 527142
rect 707800 526564 708076 526640
rect 707800 526422 708076 526498
rect 707800 526193 708076 526269
rect 707800 525672 708076 525748
rect 69924 515252 70200 515328
rect 69924 514731 70200 514807
rect 69924 514502 70200 514578
rect 69924 514360 70200 514436
rect 69924 513858 70200 513934
rect 69924 513647 70200 513723
rect 69924 502190 70200 502266
rect 69924 502044 70200 502120
rect 69924 501898 70200 501974
rect 69924 501752 70200 501828
rect 69924 392252 70200 392328
rect 69924 391731 70200 391807
rect 69924 391502 70200 391578
rect 69924 391360 70200 391436
rect 69924 390858 70200 390934
rect 69924 390647 70200 390723
rect 69924 379190 70200 379266
rect 69924 379044 70200 379120
rect 69924 378898 70200 378974
rect 69924 378752 70200 378828
rect 707800 367172 708076 367248
rect 707800 367026 708076 367102
rect 707800 366880 708076 366956
rect 707800 366734 708076 366810
rect 707800 355277 708076 355353
rect 707800 355066 708076 355142
rect 707800 354564 708076 354640
rect 707800 354422 708076 354498
rect 707800 354193 708076 354269
rect 707800 353672 708076 353748
rect 69924 351252 70200 351328
rect 69924 350731 70200 350807
rect 69924 350502 70200 350578
rect 69924 350360 70200 350436
rect 69924 349858 70200 349934
rect 69924 349647 70200 349723
rect 69924 338190 70200 338266
rect 69924 338044 70200 338120
rect 69924 337898 70200 337974
rect 69924 337752 70200 337828
rect 707800 324172 708076 324248
rect 707800 324026 708076 324102
rect 707800 323880 708076 323956
rect 707800 323734 708076 323810
rect 707800 312277 708076 312353
rect 707800 312066 708076 312142
rect 707800 311564 708076 311640
rect 707800 311422 708076 311498
rect 707800 311193 708076 311269
rect 707800 310672 708076 310748
rect 69924 310252 70200 310328
rect 69924 309731 70200 309807
rect 69924 309502 70200 309578
rect 69924 309360 70200 309436
rect 69924 308858 70200 308934
rect 69924 308647 70200 308723
rect 69924 297190 70200 297266
rect 69924 297044 70200 297120
rect 69924 296898 70200 296974
rect 69924 296752 70200 296828
rect 707800 281172 708076 281248
rect 707800 281026 708076 281102
rect 707800 280880 708076 280956
rect 707800 280734 708076 280810
rect 69924 269252 70200 269328
rect 707800 269277 708076 269353
rect 707800 269066 708076 269142
rect 69924 268731 70200 268807
rect 69924 268502 70200 268578
rect 707800 268564 708076 268640
rect 69924 268360 70200 268436
rect 707800 268422 708076 268498
rect 707800 268193 708076 268269
rect 69924 267858 70200 267934
rect 69924 267647 70200 267723
rect 707800 267672 708076 267748
rect 69924 256190 70200 256266
rect 69924 256044 70200 256120
rect 69924 255898 70200 255974
rect 69924 255752 70200 255828
rect 707800 238172 708076 238248
rect 707800 238026 708076 238102
rect 707800 237880 708076 237956
rect 707800 237734 708076 237810
rect 69924 228252 70200 228328
rect 69924 227731 70200 227807
rect 69924 227502 70200 227578
rect 69924 227360 70200 227436
rect 69924 226858 70200 226934
rect 69924 226647 70200 226723
rect 707800 226277 708076 226353
rect 707800 226066 708076 226142
rect 707800 225564 708076 225640
rect 707800 225422 708076 225498
rect 707800 225193 708076 225269
rect 707800 224672 708076 224748
rect 69924 215190 70200 215266
rect 69924 215044 70200 215120
rect 69924 214898 70200 214974
rect 69924 214752 70200 214828
rect 707800 195172 708076 195248
rect 707800 195026 708076 195102
rect 707800 194880 708076 194956
rect 707800 194734 708076 194810
rect 69924 187252 70200 187328
rect 69924 186731 70200 186807
rect 69924 186502 70200 186578
rect 69924 186360 70200 186436
rect 69924 185858 70200 185934
rect 69924 185647 70200 185723
rect 707800 183277 708076 183353
rect 707800 183066 708076 183142
rect 707800 182564 708076 182640
rect 707800 182422 708076 182498
rect 707800 182193 708076 182269
rect 707800 181672 708076 181748
rect 69924 174190 70200 174266
rect 69924 174044 70200 174120
rect 69924 173898 70200 173974
rect 69924 173752 70200 173828
rect 707621 152172 708010 152248
rect 707621 152026 708010 152102
rect 707621 151880 708010 151956
rect 707621 151734 708010 151810
rect 707621 140277 708020 140353
rect 707621 140066 708020 140142
rect 707621 139564 708020 139640
rect 707621 139422 708020 139498
rect 707621 139193 708020 139269
rect 707621 138672 708020 138748
rect 707800 109172 708076 109248
rect 707800 109026 708076 109102
rect 707800 108880 708076 108956
rect 707800 108734 708076 108810
rect 707800 97277 708076 97353
rect 707800 97066 708076 97142
rect 707800 96564 708076 96640
rect 707800 96422 708076 96498
rect 707800 96193 708076 96269
rect 707800 95672 708076 95748
rect 176172 69924 176248 70200
rect 231172 69924 231248 70200
rect 340880 69924 340956 70200
rect 341026 69924 341102 70200
rect 395880 69924 395956 70200
rect 396026 69924 396102 70200
rect 439277 69924 439353 70200
rect 450880 69924 450956 70200
rect 451026 69924 451102 70200
rect 451171 69924 451247 70200
rect 494277 69924 494353 70200
rect 505880 69924 505956 70200
rect 506026 69924 506102 70200
rect 506172 69924 506248 70200
rect 547672 69924 547748 70200
rect 548193 69924 548269 70200
rect 548422 69924 548498 70200
rect 548564 69923 548640 70199
rect 549066 69924 549142 70200
rect 549277 69924 549353 70200
rect 560734 69924 560810 70200
rect 560880 69924 560956 70200
rect 561026 69924 561102 70200
rect 561172 69924 561248 70200
<< metal5 >>
rect 107500 1007600 119500 1019600
rect 162500 1007600 174500 1019600
rect 217500 1007600 229500 1019600
rect 272500 1007600 284500 1019600
rect 327500 1007600 339500 1019600
rect 382500 1007600 394500 1019600
rect 437500 1007600 449500 1019600
rect 492500 1007600 504500 1019600
rect 547500 1007600 559500 1019600
rect 602500 1007600 614500 1019600
rect 657500 1007600 669500 1019600
rect 400 912500 12400 924500
rect 765600 913500 777600 925500
rect 400 871500 12400 883500
rect 765600 870500 777600 882500
rect 400 830500 12400 842500
rect 765600 827500 777600 839500
rect 400 789500 12400 801500
rect 765600 784500 777600 796500
rect 400 748500 12400 760500
rect 765600 741500 777600 753500
rect 400 707500 12400 719500
rect 765600 698500 777600 710500
rect 400 666500 12400 678500
rect 765600 655500 777600 667500
rect 400 625500 12400 637500
rect 765600 612500 777600 624500
rect 400 584500 12400 596500
rect 765600 569500 777600 581500
rect 400 543500 12400 555500
rect 765600 526500 777600 538500
rect 400 502500 12400 514500
rect 765600 483500 777600 495500
rect 400 461500 12400 473500
rect 765600 440500 777600 452500
rect 400 420500 12400 432500
rect 765600 397500 777600 409500
rect 400 379500 12400 391500
rect 765600 354500 777600 366500
rect 400 338500 12400 350500
rect 765600 311500 777600 323500
rect 400 297500 12400 309500
rect 765600 268500 777600 280500
rect 400 256500 12400 268500
rect 400 215500 12400 227500
rect 765600 225500 777600 237500
rect 400 174500 12400 186500
rect 765600 182500 777600 194500
rect 400 133500 12400 145500
rect 765600 139500 777600 151500
rect 400 92500 12400 104500
rect 765600 96500 777600 108500
rect 108500 400 120500 12400
rect 163500 400 175500 12400
rect 218500 400 230500 12400
rect 273500 400 285500 12400
rect 328500 400 340500 12400
rect 383500 400 395500 12400
rect 438500 400 450500 12400
rect 493500 400 505500 12400
rect 548500 400 560500 12400
rect 603500 400 615500 12400
rect 658500 400 670500 12400
use GF_NI_BI_T  GF_NI_BI_T_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 327000 0 1 0
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_1
timestamp 1654889802
transform 1 0 382000 0 1 0
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_2
timestamp 1654889802
transform 1 0 437000 0 1 0
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_3
timestamp 1654889802
transform 1 0 492000 0 1 0
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_4
timestamp 1654889802
transform 1 0 547000 0 1 0
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_5
timestamp 1654889802
transform 0 -1 778000 1 0 95000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_6
timestamp 1654889802
transform 0 -1 778000 1 0 138000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_7
timestamp 1654889802
transform 0 -1 778000 1 0 181000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_8
timestamp 1654889802
transform 0 -1 778000 1 0 224000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_9
timestamp 1654889802
transform 0 -1 778000 1 0 267000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_10
timestamp 1654889802
transform 0 -1 778000 1 0 310000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_11
timestamp 1654889802
transform 0 -1 778000 1 0 353000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_12
timestamp 1654889802
transform -1 0 451000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_13
timestamp 1654889802
transform -1 0 176000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_14
timestamp 1654889802
transform -1 0 341000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_15
timestamp 1654889802
transform 0 -1 778000 1 0 525000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_16
timestamp 1654889802
transform 0 -1 778000 1 0 568000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_17
timestamp 1654889802
transform 0 -1 778000 1 0 611000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_18
timestamp 1654889802
transform 0 -1 778000 1 0 654000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_19
timestamp 1654889802
transform 0 -1 778000 1 0 697000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_20
timestamp 1654889802
transform 0 -1 778000 1 0 740000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_21
timestamp 1654889802
transform -1 0 286000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_22
timestamp 1654889802
transform 0 -1 778000 1 0 826000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_23
timestamp 1654889802
transform -1 0 231000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_24
timestamp 1654889802
transform 0 -1 778000 1 0 912000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_25
timestamp 1654889802
transform -1 0 671000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_26
timestamp 1654889802
transform -1 0 561000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_27
timestamp 1654889802
transform -1 0 506000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_28
timestamp 1654889802
transform -1 0 121000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_29
timestamp 1654889802
transform 0 1 0 -1 0 926000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_30
timestamp 1654889802
transform 0 1 0 -1 0 639000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_31
timestamp 1654889802
transform 0 1 0 -1 0 598000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_32
timestamp 1654889802
transform 0 1 0 -1 0 557000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_33
timestamp 1654889802
transform 0 1 0 -1 0 762000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_34
timestamp 1654889802
transform 0 1 0 -1 0 721000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_35
timestamp 1654889802
transform 0 1 0 -1 0 680000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_36
timestamp 1654889802
transform 0 1 0 -1 0 516000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_37
timestamp 1654889802
transform 0 1 0 -1 0 188000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_38
timestamp 1654889802
transform 0 1 0 -1 0 270000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_39
timestamp 1654889802
transform 0 1 0 -1 0 393000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_40
timestamp 1654889802
transform 0 1 0 -1 0 352000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_41
timestamp 1654889802
transform 0 1 0 -1 0 311000
box -32 0 15032 70000
use GF_NI_BI_T  GF_NI_BI_T_42
timestamp 1654889802
transform 0 1 0 -1 0 229000
box -32 0 15032 70000
use GF_NI_COR  GF_NI_COR_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 0 0 1 0
box 0 0 71000 71000
use GF_NI_COR  GF_NI_COR_1
timestamp 1654889802
transform -1 0 778000 0 1 0
box 0 0 71000 71000
use GF_NI_COR  GF_NI_COR_2
timestamp 1654889802
transform -1 0 778000 0 -1 1020000
box 0 0 71000 71000
use GF_NI_COR  GF_NI_COR_3
timestamp 1654889802
transform 1 0 0 0 -1 1020000
box 0 0 71000 71000
use GF_NI_DVDD  GF_NI_DVDD_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 657000 0 1 0
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_1
timestamp 1654889802
transform 0 -1 778000 1 0 482000
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_2
timestamp 1654889802
transform 0 -1 778000 1 0 783000
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_3
timestamp 1654889802
transform 0 -1 778000 1 0 869000
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_4
timestamp 1654889802
transform 0 1 0 -1 0 475000
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_5
timestamp 1654889802
transform 0 1 0 -1 0 106000
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_7
timestamp 1654889802
transform 0 1 0 -1 0 885000
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_8
timestamp 1654889802
transform 0 1 0 -1 0 844000
box -32 0 15032 70000
use GF_NI_DVDD  GF_NI_DVDD_9
timestamp 1654889802
transform 0 1 0 -1 0 147000
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 107000 0 1 0
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_1
timestamp 1654889802
transform 1 0 272000 0 1 0
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_2
timestamp 1654889802
transform 1 0 602000 0 1 0
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_3
timestamp 1654889802
transform 0 -1 778000 1 0 396000
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_4
timestamp 1654889802
transform 0 -1 778000 1 0 439000
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_5
timestamp 1654889802
transform -1 0 396000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_6
timestamp 1654889802
transform 0 1 0 -1 0 434000
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_8
timestamp 1654889802
transform -1 0 616000 0 -1 1020000
box -32 0 15032 70000
use GF_NI_DVSS  GF_NI_DVSS_9
timestamp 1654889802
transform 0 1 0 -1 0 803000
box -32 0 15032 70000
use GF_NI_FILL5  GF_NI_FILL5_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 706000 0 1 0
box -32 13097 1032 69968
use GF_NI_FILL5  GF_NI_FILL5_1
timestamp 1654889802
transform -1 0 72000 0 -1 1020000
box -32 13097 1032 69968
use GF_NI_FILL5  GF_NI_FILL5_2
timestamp 1654889802
transform 0 1 0 -1 0 949000
box -32 13097 1032 69968
use GF_NI_FILL10  GF_NI_FILL10_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 71000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1
timestamp 1654889802
transform 1 0 73000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_2
timestamp 1654889802
transform 1 0 75000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_3
timestamp 1654889802
transform 1 0 77000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_4
timestamp 1654889802
transform 1 0 79000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_5
timestamp 1654889802
transform 1 0 81000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_6
timestamp 1654889802
transform 1 0 83000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_7
timestamp 1654889802
transform 1 0 85000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_8
timestamp 1654889802
transform 1 0 87000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_9
timestamp 1654889802
transform 1 0 89000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_10
timestamp 1654889802
transform 1 0 91000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_11
timestamp 1654889802
transform 1 0 93000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_12
timestamp 1654889802
transform 1 0 95000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_13
timestamp 1654889802
transform 1 0 97000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_14
timestamp 1654889802
transform 1 0 99000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_15
timestamp 1654889802
transform 1 0 101000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_16
timestamp 1654889802
transform 1 0 103000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_17
timestamp 1654889802
transform 1 0 105000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_18
timestamp 1654889802
transform 1 0 122000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_19
timestamp 1654889802
transform 1 0 124000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_20
timestamp 1654889802
transform 1 0 126000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_21
timestamp 1654889802
transform 1 0 128000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_22
timestamp 1654889802
transform 1 0 130000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_23
timestamp 1654889802
transform 1 0 132000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_24
timestamp 1654889802
transform 1 0 134000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_25
timestamp 1654889802
transform 1 0 136000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_26
timestamp 1654889802
transform 1 0 138000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_27
timestamp 1654889802
transform 1 0 140000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_28
timestamp 1654889802
transform 1 0 142000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_29
timestamp 1654889802
transform 1 0 144000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_30
timestamp 1654889802
transform 1 0 146000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_31
timestamp 1654889802
transform 1 0 148000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_32
timestamp 1654889802
transform 1 0 150000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_33
timestamp 1654889802
transform 1 0 152000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_34
timestamp 1654889802
transform 1 0 154000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_35
timestamp 1654889802
transform 1 0 156000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_36
timestamp 1654889802
transform 1 0 158000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_37
timestamp 1654889802
transform 1 0 160000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_38
timestamp 1654889802
transform 1 0 177000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_39
timestamp 1654889802
transform 1 0 179000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_40
timestamp 1654889802
transform 1 0 181000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_41
timestamp 1654889802
transform 1 0 183000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_42
timestamp 1654889802
transform 1 0 185000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_43
timestamp 1654889802
transform 1 0 187000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_44
timestamp 1654889802
transform 1 0 189000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_45
timestamp 1654889802
transform 1 0 191000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_46
timestamp 1654889802
transform 1 0 215000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_47
timestamp 1654889802
transform 1 0 213000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_48
timestamp 1654889802
transform 1 0 211000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_49
timestamp 1654889802
transform 1 0 209000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_50
timestamp 1654889802
transform 1 0 207000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_51
timestamp 1654889802
transform 1 0 205000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_52
timestamp 1654889802
transform 1 0 203000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_53
timestamp 1654889802
transform 1 0 201000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_54
timestamp 1654889802
transform 1 0 199000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_55
timestamp 1654889802
transform 1 0 197000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_56
timestamp 1654889802
transform 1 0 195000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_57
timestamp 1654889802
transform 1 0 193000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_58
timestamp 1654889802
transform 1 0 248000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_59
timestamp 1654889802
transform 1 0 232000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_60
timestamp 1654889802
transform 1 0 234000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_61
timestamp 1654889802
transform 1 0 236000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_62
timestamp 1654889802
transform 1 0 238000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_63
timestamp 1654889802
transform 1 0 240000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_64
timestamp 1654889802
transform 1 0 242000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_65
timestamp 1654889802
transform 1 0 244000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_66
timestamp 1654889802
transform 1 0 246000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_67
timestamp 1654889802
transform 1 0 270000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_68
timestamp 1654889802
transform 1 0 268000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_69
timestamp 1654889802
transform 1 0 266000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_70
timestamp 1654889802
transform 1 0 264000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_71
timestamp 1654889802
transform 1 0 262000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_72
timestamp 1654889802
transform 1 0 260000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_73
timestamp 1654889802
transform 1 0 258000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_74
timestamp 1654889802
transform 1 0 256000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_75
timestamp 1654889802
transform 1 0 254000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_76
timestamp 1654889802
transform 1 0 252000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_77
timestamp 1654889802
transform 1 0 250000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_78
timestamp 1654889802
transform 1 0 305000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_79
timestamp 1654889802
transform 1 0 303000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_80
timestamp 1654889802
transform 1 0 287000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_81
timestamp 1654889802
transform 1 0 289000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_82
timestamp 1654889802
transform 1 0 291000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_83
timestamp 1654889802
transform 1 0 293000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_84
timestamp 1654889802
transform 1 0 295000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_85
timestamp 1654889802
transform 1 0 297000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_86
timestamp 1654889802
transform 1 0 299000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_87
timestamp 1654889802
transform 1 0 301000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_88
timestamp 1654889802
transform 1 0 325000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_89
timestamp 1654889802
transform 1 0 323000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_90
timestamp 1654889802
transform 1 0 321000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_91
timestamp 1654889802
transform 1 0 319000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_92
timestamp 1654889802
transform 1 0 317000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_93
timestamp 1654889802
transform 1 0 315000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_94
timestamp 1654889802
transform 1 0 313000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_95
timestamp 1654889802
transform 1 0 311000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_96
timestamp 1654889802
transform 1 0 309000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_97
timestamp 1654889802
transform 1 0 307000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_98
timestamp 1654889802
transform 1 0 362000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_99
timestamp 1654889802
transform 1 0 360000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_100
timestamp 1654889802
transform 1 0 358000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_101
timestamp 1654889802
transform 1 0 342000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_102
timestamp 1654889802
transform 1 0 344000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_103
timestamp 1654889802
transform 1 0 346000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_104
timestamp 1654889802
transform 1 0 348000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_105
timestamp 1654889802
transform 1 0 350000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_106
timestamp 1654889802
transform 1 0 352000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_107
timestamp 1654889802
transform 1 0 354000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_108
timestamp 1654889802
transform 1 0 356000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_109
timestamp 1654889802
transform 1 0 380000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_110
timestamp 1654889802
transform 1 0 378000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_111
timestamp 1654889802
transform 1 0 376000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_112
timestamp 1654889802
transform 1 0 374000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_113
timestamp 1654889802
transform 1 0 372000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_114
timestamp 1654889802
transform 1 0 370000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_115
timestamp 1654889802
transform 1 0 368000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_116
timestamp 1654889802
transform 1 0 366000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_117
timestamp 1654889802
transform 1 0 364000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_118
timestamp 1654889802
transform 1 0 417000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_119
timestamp 1654889802
transform 1 0 415000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_120
timestamp 1654889802
transform 1 0 413000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_121
timestamp 1654889802
transform 1 0 397000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_122
timestamp 1654889802
transform 1 0 399000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_123
timestamp 1654889802
transform 1 0 401000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_124
timestamp 1654889802
transform 1 0 403000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_125
timestamp 1654889802
transform 1 0 405000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_126
timestamp 1654889802
transform 1 0 407000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_127
timestamp 1654889802
transform 1 0 409000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_128
timestamp 1654889802
transform 1 0 411000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_129
timestamp 1654889802
transform 1 0 435000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_130
timestamp 1654889802
transform 1 0 433000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_131
timestamp 1654889802
transform 1 0 431000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_132
timestamp 1654889802
transform 1 0 429000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_133
timestamp 1654889802
transform 1 0 427000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_134
timestamp 1654889802
transform 1 0 425000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_135
timestamp 1654889802
transform 1 0 423000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_136
timestamp 1654889802
transform 1 0 421000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_137
timestamp 1654889802
transform 1 0 419000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_138
timestamp 1654889802
transform 1 0 452000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_139
timestamp 1654889802
transform 1 0 454000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_140
timestamp 1654889802
transform 1 0 456000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_141
timestamp 1654889802
transform 1 0 458000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_142
timestamp 1654889802
transform 1 0 460000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_143
timestamp 1654889802
transform 1 0 462000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_144
timestamp 1654889802
transform 1 0 464000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_145
timestamp 1654889802
transform 1 0 468000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_146
timestamp 1654889802
transform 1 0 466000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_147
timestamp 1654889802
transform 1 0 472000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_148
timestamp 1654889802
transform 1 0 470000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_149
timestamp 1654889802
transform 1 0 476000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_150
timestamp 1654889802
transform 1 0 474000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_151
timestamp 1654889802
transform 1 0 480000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_152
timestamp 1654889802
transform 1 0 478000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_153
timestamp 1654889802
transform 1 0 484000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_154
timestamp 1654889802
transform 1 0 482000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_155
timestamp 1654889802
transform 1 0 488000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_156
timestamp 1654889802
transform 1 0 486000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_157
timestamp 1654889802
transform 1 0 490000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_158
timestamp 1654889802
transform 1 0 507000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_159
timestamp 1654889802
transform 1 0 509000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_160
timestamp 1654889802
transform 1 0 511000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_161
timestamp 1654889802
transform 1 0 513000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_162
timestamp 1654889802
transform 1 0 515000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_163
timestamp 1654889802
transform 1 0 517000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_164
timestamp 1654889802
transform 1 0 519000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_165
timestamp 1654889802
transform 1 0 523000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_166
timestamp 1654889802
transform 1 0 521000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_167
timestamp 1654889802
transform 1 0 527000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_168
timestamp 1654889802
transform 1 0 525000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_169
timestamp 1654889802
transform 1 0 531000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_170
timestamp 1654889802
transform 1 0 529000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_171
timestamp 1654889802
transform 1 0 535000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_172
timestamp 1654889802
transform 1 0 533000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_173
timestamp 1654889802
transform 1 0 539000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_174
timestamp 1654889802
transform 1 0 537000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_175
timestamp 1654889802
transform 1 0 543000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_176
timestamp 1654889802
transform 1 0 541000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_177
timestamp 1654889802
transform 1 0 545000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_178
timestamp 1654889802
transform 1 0 562000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_179
timestamp 1654889802
transform 1 0 564000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_180
timestamp 1654889802
transform 1 0 566000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_181
timestamp 1654889802
transform 1 0 568000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_182
timestamp 1654889802
transform 1 0 570000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_183
timestamp 1654889802
transform 1 0 572000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_184
timestamp 1654889802
transform 1 0 574000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_185
timestamp 1654889802
transform 1 0 578000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_186
timestamp 1654889802
transform 1 0 576000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_187
timestamp 1654889802
transform 1 0 582000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_188
timestamp 1654889802
transform 1 0 580000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_189
timestamp 1654889802
transform 1 0 586000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_190
timestamp 1654889802
transform 1 0 584000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_191
timestamp 1654889802
transform 1 0 590000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_192
timestamp 1654889802
transform 1 0 588000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_193
timestamp 1654889802
transform 1 0 594000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_194
timestamp 1654889802
transform 1 0 592000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_195
timestamp 1654889802
transform 1 0 598000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_196
timestamp 1654889802
transform 1 0 596000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_197
timestamp 1654889802
transform 1 0 600000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_198
timestamp 1654889802
transform 1 0 617000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_199
timestamp 1654889802
transform 1 0 619000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_200
timestamp 1654889802
transform 1 0 621000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_201
timestamp 1654889802
transform 1 0 623000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_202
timestamp 1654889802
transform 1 0 625000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_203
timestamp 1654889802
transform 1 0 627000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_204
timestamp 1654889802
transform 1 0 629000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_205
timestamp 1654889802
transform 1 0 633000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_206
timestamp 1654889802
transform 1 0 631000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_207
timestamp 1654889802
transform 1 0 637000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_208
timestamp 1654889802
transform 1 0 635000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_209
timestamp 1654889802
transform 1 0 641000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_210
timestamp 1654889802
transform 1 0 639000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_211
timestamp 1654889802
transform 1 0 645000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_212
timestamp 1654889802
transform 1 0 643000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_213
timestamp 1654889802
transform 1 0 649000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_214
timestamp 1654889802
transform 1 0 647000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_215
timestamp 1654889802
transform 1 0 653000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_216
timestamp 1654889802
transform 1 0 651000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_217
timestamp 1654889802
transform 1 0 655000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_218
timestamp 1654889802
transform 1 0 672000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_219
timestamp 1654889802
transform 1 0 674000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_220
timestamp 1654889802
transform 1 0 676000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_221
timestamp 1654889802
transform 1 0 678000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_222
timestamp 1654889802
transform 1 0 680000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_223
timestamp 1654889802
transform 1 0 682000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_224
timestamp 1654889802
transform 1 0 684000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_225
timestamp 1654889802
transform 1 0 688000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_226
timestamp 1654889802
transform 1 0 686000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_227
timestamp 1654889802
transform 1 0 692000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_228
timestamp 1654889802
transform 1 0 690000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_229
timestamp 1654889802
transform 1 0 696000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_230
timestamp 1654889802
transform 1 0 694000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_231
timestamp 1654889802
transform 1 0 700000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_232
timestamp 1654889802
transform 1 0 698000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_233
timestamp 1654889802
transform 1 0 704000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_234
timestamp 1654889802
transform 1 0 702000 0 1 0
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_235
timestamp 1654889802
transform 0 -1 778000 1 0 71000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_236
timestamp 1654889802
transform 0 -1 778000 1 0 73000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_237
timestamp 1654889802
transform 0 -1 778000 1 0 75000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_238
timestamp 1654889802
transform 0 -1 778000 1 0 77000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_239
timestamp 1654889802
transform 0 -1 778000 1 0 79000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_240
timestamp 1654889802
transform 0 -1 778000 1 0 81000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_241
timestamp 1654889802
transform 0 -1 778000 1 0 83000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_242
timestamp 1654889802
transform 0 -1 778000 1 0 85000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_243
timestamp 1654889802
transform 0 -1 778000 1 0 87000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_244
timestamp 1654889802
transform 0 -1 778000 1 0 89000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_245
timestamp 1654889802
transform 0 -1 778000 1 0 91000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_246
timestamp 1654889802
transform 0 -1 778000 1 0 93000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_247
timestamp 1654889802
transform 0 -1 778000 1 0 118000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_248
timestamp 1654889802
transform 0 -1 778000 1 0 114000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_249
timestamp 1654889802
transform 0 -1 778000 1 0 116000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_250
timestamp 1654889802
transform 0 -1 778000 1 0 122000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_251
timestamp 1654889802
transform 0 -1 778000 1 0 120000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_252
timestamp 1654889802
transform 0 -1 778000 1 0 126000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_253
timestamp 1654889802
transform 0 -1 778000 1 0 124000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_254
timestamp 1654889802
transform 0 -1 778000 1 0 130000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_255
timestamp 1654889802
transform 0 -1 778000 1 0 128000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_256
timestamp 1654889802
transform 0 -1 778000 1 0 134000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_257
timestamp 1654889802
transform 0 -1 778000 1 0 132000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_258
timestamp 1654889802
transform 0 -1 778000 1 0 136000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_259
timestamp 1654889802
transform 0 -1 778000 1 0 112000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_260
timestamp 1654889802
transform 0 -1 778000 1 0 110000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_261
timestamp 1654889802
transform 0 -1 778000 1 0 153000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_262
timestamp 1654889802
transform 0 -1 778000 1 0 155000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_263
timestamp 1654889802
transform 0 -1 778000 1 0 157000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_264
timestamp 1654889802
transform 0 -1 778000 1 0 159000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_265
timestamp 1654889802
transform 0 -1 778000 1 0 163000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_266
timestamp 1654889802
transform 0 -1 778000 1 0 161000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_267
timestamp 1654889802
transform 0 -1 778000 1 0 167000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_268
timestamp 1654889802
transform 0 -1 778000 1 0 165000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_269
timestamp 1654889802
transform 0 -1 778000 1 0 171000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_270
timestamp 1654889802
transform 0 -1 778000 1 0 169000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_271
timestamp 1654889802
transform 0 -1 778000 1 0 175000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_272
timestamp 1654889802
transform 0 -1 778000 1 0 173000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_273
timestamp 1654889802
transform 0 -1 778000 1 0 179000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_274
timestamp 1654889802
transform 0 -1 778000 1 0 177000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_275
timestamp 1654889802
transform 0 -1 778000 1 0 196000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_276
timestamp 1654889802
transform 0 -1 778000 1 0 198000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_277
timestamp 1654889802
transform 0 -1 778000 1 0 200000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_278
timestamp 1654889802
transform 0 -1 778000 1 0 202000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_279
timestamp 1654889802
transform 0 -1 778000 1 0 206000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_280
timestamp 1654889802
transform 0 -1 778000 1 0 204000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_281
timestamp 1654889802
transform 0 -1 778000 1 0 210000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_282
timestamp 1654889802
transform 0 -1 778000 1 0 208000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_283
timestamp 1654889802
transform 0 -1 778000 1 0 214000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_284
timestamp 1654889802
transform 0 -1 778000 1 0 212000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_285
timestamp 1654889802
transform 0 -1 778000 1 0 218000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_286
timestamp 1654889802
transform 0 -1 778000 1 0 216000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_287
timestamp 1654889802
transform 0 -1 778000 1 0 222000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_288
timestamp 1654889802
transform 0 -1 778000 1 0 220000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_289
timestamp 1654889802
transform 0 -1 778000 1 0 239000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_290
timestamp 1654889802
transform 0 -1 778000 1 0 241000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_291
timestamp 1654889802
transform 0 -1 778000 1 0 243000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_292
timestamp 1654889802
transform 0 -1 778000 1 0 245000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_293
timestamp 1654889802
transform 0 -1 778000 1 0 249000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_294
timestamp 1654889802
transform 0 -1 778000 1 0 247000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_295
timestamp 1654889802
transform 0 -1 778000 1 0 253000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_296
timestamp 1654889802
transform 0 -1 778000 1 0 251000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_297
timestamp 1654889802
transform 0 -1 778000 1 0 257000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_298
timestamp 1654889802
transform 0 -1 778000 1 0 255000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_299
timestamp 1654889802
transform 0 -1 778000 1 0 261000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_300
timestamp 1654889802
transform 0 -1 778000 1 0 259000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_301
timestamp 1654889802
transform 0 -1 778000 1 0 265000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_302
timestamp 1654889802
transform 0 -1 778000 1 0 263000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_303
timestamp 1654889802
transform 0 -1 778000 1 0 282000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_304
timestamp 1654889802
transform 0 -1 778000 1 0 284000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_305
timestamp 1654889802
transform 0 -1 778000 1 0 286000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_306
timestamp 1654889802
transform 0 -1 778000 1 0 288000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_307
timestamp 1654889802
transform 0 -1 778000 1 0 292000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_308
timestamp 1654889802
transform 0 -1 778000 1 0 290000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_309
timestamp 1654889802
transform 0 -1 778000 1 0 296000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_310
timestamp 1654889802
transform 0 -1 778000 1 0 294000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_311
timestamp 1654889802
transform 0 -1 778000 1 0 300000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_312
timestamp 1654889802
transform 0 -1 778000 1 0 298000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_313
timestamp 1654889802
transform 0 -1 778000 1 0 304000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_314
timestamp 1654889802
transform 0 -1 778000 1 0 302000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_315
timestamp 1654889802
transform 0 -1 778000 1 0 308000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_316
timestamp 1654889802
transform 0 -1 778000 1 0 306000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_317
timestamp 1654889802
transform 0 -1 778000 1 0 325000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_318
timestamp 1654889802
transform 0 -1 778000 1 0 327000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_319
timestamp 1654889802
transform 0 -1 778000 1 0 329000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_320
timestamp 1654889802
transform 0 -1 778000 1 0 331000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_321
timestamp 1654889802
transform 0 -1 778000 1 0 335000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_322
timestamp 1654889802
transform 0 -1 778000 1 0 333000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_323
timestamp 1654889802
transform 0 -1 778000 1 0 339000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_324
timestamp 1654889802
transform 0 -1 778000 1 0 337000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_325
timestamp 1654889802
transform 0 -1 778000 1 0 343000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_326
timestamp 1654889802
transform 0 -1 778000 1 0 341000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_327
timestamp 1654889802
transform 0 -1 778000 1 0 347000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_328
timestamp 1654889802
transform 0 -1 778000 1 0 345000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_329
timestamp 1654889802
transform 0 -1 778000 1 0 351000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_330
timestamp 1654889802
transform 0 -1 778000 1 0 349000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_331
timestamp 1654889802
transform 0 -1 778000 1 0 368000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_332
timestamp 1654889802
transform 0 -1 778000 1 0 370000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_333
timestamp 1654889802
transform 0 -1 778000 1 0 372000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_334
timestamp 1654889802
transform 0 -1 778000 1 0 374000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_335
timestamp 1654889802
transform 0 -1 778000 1 0 378000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_336
timestamp 1654889802
transform 0 -1 778000 1 0 376000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_337
timestamp 1654889802
transform 0 -1 778000 1 0 382000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_338
timestamp 1654889802
transform 0 -1 778000 1 0 380000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_339
timestamp 1654889802
transform 0 -1 778000 1 0 386000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_340
timestamp 1654889802
transform 0 -1 778000 1 0 384000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_341
timestamp 1654889802
transform 0 -1 778000 1 0 390000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_342
timestamp 1654889802
transform 0 -1 778000 1 0 388000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_343
timestamp 1654889802
transform 0 -1 778000 1 0 394000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_344
timestamp 1654889802
transform 0 -1 778000 1 0 392000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_345
timestamp 1654889802
transform 0 -1 778000 1 0 411000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_346
timestamp 1654889802
transform 0 -1 778000 1 0 413000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_347
timestamp 1654889802
transform 0 -1 778000 1 0 415000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_348
timestamp 1654889802
transform 0 -1 778000 1 0 417000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_349
timestamp 1654889802
transform 0 -1 778000 1 0 421000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_350
timestamp 1654889802
transform 0 -1 778000 1 0 419000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_351
timestamp 1654889802
transform 0 -1 778000 1 0 425000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_352
timestamp 1654889802
transform 0 -1 778000 1 0 423000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_353
timestamp 1654889802
transform 0 -1 778000 1 0 429000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_354
timestamp 1654889802
transform 0 -1 778000 1 0 427000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_355
timestamp 1654889802
transform 0 -1 778000 1 0 433000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_356
timestamp 1654889802
transform 0 -1 778000 1 0 431000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_357
timestamp 1654889802
transform 0 -1 778000 1 0 437000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_358
timestamp 1654889802
transform 0 -1 778000 1 0 435000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_359
timestamp 1654889802
transform 0 -1 778000 1 0 454000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_360
timestamp 1654889802
transform 0 -1 778000 1 0 456000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_361
timestamp 1654889802
transform 0 -1 778000 1 0 458000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_362
timestamp 1654889802
transform 0 -1 778000 1 0 460000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_363
timestamp 1654889802
transform 0 -1 778000 1 0 464000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_364
timestamp 1654889802
transform 0 -1 778000 1 0 462000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_365
timestamp 1654889802
transform 0 -1 778000 1 0 468000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_366
timestamp 1654889802
transform 0 -1 778000 1 0 466000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_367
timestamp 1654889802
transform 0 -1 778000 1 0 472000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_368
timestamp 1654889802
transform 0 -1 778000 1 0 470000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_369
timestamp 1654889802
transform 0 -1 778000 1 0 476000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_370
timestamp 1654889802
transform 0 -1 778000 1 0 474000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_371
timestamp 1654889802
transform 0 -1 778000 1 0 480000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_372
timestamp 1654889802
transform 0 -1 778000 1 0 478000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_373
timestamp 1654889802
transform 0 -1 778000 1 0 497000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_374
timestamp 1654889802
transform 0 -1 778000 1 0 499000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_375
timestamp 1654889802
transform 0 -1 778000 1 0 501000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_376
timestamp 1654889802
transform 0 -1 778000 1 0 503000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_377
timestamp 1654889802
transform 0 -1 778000 1 0 507000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_378
timestamp 1654889802
transform 0 -1 778000 1 0 505000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_379
timestamp 1654889802
transform 0 -1 778000 1 0 511000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_380
timestamp 1654889802
transform 0 -1 778000 1 0 509000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_381
timestamp 1654889802
transform 0 -1 778000 1 0 515000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_382
timestamp 1654889802
transform 0 -1 778000 1 0 513000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_383
timestamp 1654889802
transform 0 -1 778000 1 0 519000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_384
timestamp 1654889802
transform 0 -1 778000 1 0 517000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_385
timestamp 1654889802
transform 0 -1 778000 1 0 523000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_386
timestamp 1654889802
transform 0 -1 778000 1 0 521000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_387
timestamp 1654889802
transform 0 -1 778000 1 0 540000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_388
timestamp 1654889802
transform 0 -1 778000 1 0 542000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_389
timestamp 1654889802
transform 0 -1 778000 1 0 544000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_390
timestamp 1654889802
transform 0 -1 778000 1 0 546000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_391
timestamp 1654889802
transform 0 -1 778000 1 0 550000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_392
timestamp 1654889802
transform 0 -1 778000 1 0 548000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_393
timestamp 1654889802
transform 0 -1 778000 1 0 554000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_394
timestamp 1654889802
transform 0 -1 778000 1 0 552000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_395
timestamp 1654889802
transform 0 -1 778000 1 0 558000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_396
timestamp 1654889802
transform 0 -1 778000 1 0 556000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_397
timestamp 1654889802
transform 0 -1 778000 1 0 562000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_398
timestamp 1654889802
transform 0 -1 778000 1 0 560000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_399
timestamp 1654889802
transform 0 -1 778000 1 0 566000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_400
timestamp 1654889802
transform 0 -1 778000 1 0 564000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_401
timestamp 1654889802
transform 0 -1 778000 1 0 583000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_402
timestamp 1654889802
transform 0 -1 778000 1 0 585000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_403
timestamp 1654889802
transform 0 -1 778000 1 0 587000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_404
timestamp 1654889802
transform 0 -1 778000 1 0 589000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_405
timestamp 1654889802
transform 0 -1 778000 1 0 593000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_406
timestamp 1654889802
transform 0 -1 778000 1 0 591000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_407
timestamp 1654889802
transform 0 -1 778000 1 0 597000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_408
timestamp 1654889802
transform 0 -1 778000 1 0 595000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_409
timestamp 1654889802
transform 0 -1 778000 1 0 601000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_410
timestamp 1654889802
transform 0 -1 778000 1 0 599000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_411
timestamp 1654889802
transform 0 -1 778000 1 0 605000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_412
timestamp 1654889802
transform 0 -1 778000 1 0 603000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_413
timestamp 1654889802
transform 0 -1 778000 1 0 609000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_414
timestamp 1654889802
transform 0 -1 778000 1 0 607000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_415
timestamp 1654889802
transform 0 -1 778000 1 0 626000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_416
timestamp 1654889802
transform 0 -1 778000 1 0 628000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_417
timestamp 1654889802
transform 0 -1 778000 1 0 630000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_418
timestamp 1654889802
transform 0 -1 778000 1 0 632000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_419
timestamp 1654889802
transform 0 -1 778000 1 0 636000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_420
timestamp 1654889802
transform 0 -1 778000 1 0 634000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_421
timestamp 1654889802
transform 0 -1 778000 1 0 640000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_422
timestamp 1654889802
transform 0 -1 778000 1 0 638000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_423
timestamp 1654889802
transform 0 -1 778000 1 0 644000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_424
timestamp 1654889802
transform 0 -1 778000 1 0 642000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_425
timestamp 1654889802
transform 0 -1 778000 1 0 648000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_426
timestamp 1654889802
transform 0 -1 778000 1 0 646000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_427
timestamp 1654889802
transform 0 -1 778000 1 0 652000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_428
timestamp 1654889802
transform 0 -1 778000 1 0 650000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_429
timestamp 1654889802
transform 0 -1 778000 1 0 669000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_430
timestamp 1654889802
transform 0 -1 778000 1 0 671000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_431
timestamp 1654889802
transform 0 -1 778000 1 0 673000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_432
timestamp 1654889802
transform 0 -1 778000 1 0 675000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_433
timestamp 1654889802
transform 0 -1 778000 1 0 679000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_434
timestamp 1654889802
transform 0 -1 778000 1 0 677000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_435
timestamp 1654889802
transform 0 -1 778000 1 0 683000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_436
timestamp 1654889802
transform 0 -1 778000 1 0 681000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_437
timestamp 1654889802
transform 0 -1 778000 1 0 687000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_438
timestamp 1654889802
transform 0 -1 778000 1 0 685000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_439
timestamp 1654889802
transform 0 -1 778000 1 0 691000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_440
timestamp 1654889802
transform 0 -1 778000 1 0 689000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_441
timestamp 1654889802
transform 0 -1 778000 1 0 695000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_442
timestamp 1654889802
transform 0 -1 778000 1 0 693000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_443
timestamp 1654889802
transform 0 -1 778000 1 0 712000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_444
timestamp 1654889802
transform 0 -1 778000 1 0 714000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_445
timestamp 1654889802
transform 0 -1 778000 1 0 716000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_446
timestamp 1654889802
transform 0 -1 778000 1 0 718000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_447
timestamp 1654889802
transform 0 -1 778000 1 0 722000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_448
timestamp 1654889802
transform 0 -1 778000 1 0 720000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_449
timestamp 1654889802
transform 0 -1 778000 1 0 726000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_450
timestamp 1654889802
transform 0 -1 778000 1 0 724000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_451
timestamp 1654889802
transform 0 -1 778000 1 0 730000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_452
timestamp 1654889802
transform 0 -1 778000 1 0 728000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_453
timestamp 1654889802
transform 0 -1 778000 1 0 734000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_454
timestamp 1654889802
transform 0 -1 778000 1 0 732000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_455
timestamp 1654889802
transform 0 -1 778000 1 0 738000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_456
timestamp 1654889802
transform 0 -1 778000 1 0 736000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_457
timestamp 1654889802
transform 0 -1 778000 1 0 755000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_458
timestamp 1654889802
transform 0 -1 778000 1 0 757000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_459
timestamp 1654889802
transform 0 -1 778000 1 0 759000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_460
timestamp 1654889802
transform 0 -1 778000 1 0 761000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_461
timestamp 1654889802
transform 0 -1 778000 1 0 765000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_462
timestamp 1654889802
transform 0 -1 778000 1 0 763000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_463
timestamp 1654889802
transform 0 -1 778000 1 0 769000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_464
timestamp 1654889802
transform 0 -1 778000 1 0 767000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_465
timestamp 1654889802
transform 0 -1 778000 1 0 773000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_466
timestamp 1654889802
transform 0 -1 778000 1 0 771000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_467
timestamp 1654889802
transform 0 -1 778000 1 0 777000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_468
timestamp 1654889802
transform 0 -1 778000 1 0 775000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_469
timestamp 1654889802
transform 0 -1 778000 1 0 781000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_470
timestamp 1654889802
transform 0 -1 778000 1 0 779000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_471
timestamp 1654889802
transform 0 -1 778000 1 0 798000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_472
timestamp 1654889802
transform 0 -1 778000 1 0 800000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_473
timestamp 1654889802
transform 0 -1 778000 1 0 802000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_474
timestamp 1654889802
transform 0 -1 778000 1 0 804000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_475
timestamp 1654889802
transform 0 -1 778000 1 0 808000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_476
timestamp 1654889802
transform 0 -1 778000 1 0 806000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_477
timestamp 1654889802
transform 0 -1 778000 1 0 812000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_478
timestamp 1654889802
transform 0 -1 778000 1 0 810000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_479
timestamp 1654889802
transform 0 -1 778000 1 0 816000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_480
timestamp 1654889802
transform 0 -1 778000 1 0 814000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_481
timestamp 1654889802
transform 0 -1 778000 1 0 820000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_482
timestamp 1654889802
transform 0 -1 778000 1 0 818000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_483
timestamp 1654889802
transform 0 -1 778000 1 0 824000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_484
timestamp 1654889802
transform 0 -1 778000 1 0 822000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_485
timestamp 1654889802
transform 0 -1 778000 1 0 841000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_486
timestamp 1654889802
transform 0 -1 778000 1 0 843000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_487
timestamp 1654889802
transform 0 -1 778000 1 0 845000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_488
timestamp 1654889802
transform 0 -1 778000 1 0 847000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_489
timestamp 1654889802
transform 0 -1 778000 1 0 851000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_490
timestamp 1654889802
transform 0 -1 778000 1 0 849000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_491
timestamp 1654889802
transform 0 -1 778000 1 0 855000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_492
timestamp 1654889802
transform 0 -1 778000 1 0 853000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_493
timestamp 1654889802
transform 0 -1 778000 1 0 859000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_494
timestamp 1654889802
transform 0 -1 778000 1 0 857000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_495
timestamp 1654889802
transform 0 -1 778000 1 0 863000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_496
timestamp 1654889802
transform 0 -1 778000 1 0 861000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_497
timestamp 1654889802
transform 0 -1 778000 1 0 867000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_498
timestamp 1654889802
transform 0 -1 778000 1 0 865000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_499
timestamp 1654889802
transform 0 -1 778000 1 0 884000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_500
timestamp 1654889802
transform 0 -1 778000 1 0 886000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_501
timestamp 1654889802
transform 0 -1 778000 1 0 888000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_502
timestamp 1654889802
transform 0 -1 778000 1 0 890000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_503
timestamp 1654889802
transform 0 -1 778000 1 0 894000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_504
timestamp 1654889802
transform 0 -1 778000 1 0 892000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_505
timestamp 1654889802
transform 0 -1 778000 1 0 898000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_506
timestamp 1654889802
transform 0 -1 778000 1 0 896000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_507
timestamp 1654889802
transform 0 -1 778000 1 0 902000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_508
timestamp 1654889802
transform 0 -1 778000 1 0 900000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_509
timestamp 1654889802
transform 0 -1 778000 1 0 906000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_510
timestamp 1654889802
transform 0 -1 778000 1 0 904000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_511
timestamp 1654889802
transform 0 -1 778000 1 0 910000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_512
timestamp 1654889802
transform 0 -1 778000 1 0 908000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_513
timestamp 1654889802
transform 0 -1 778000 1 0 931000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_514
timestamp 1654889802
transform 0 -1 778000 1 0 927000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_515
timestamp 1654889802
transform 0 -1 778000 1 0 929000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_516
timestamp 1654889802
transform 0 -1 778000 1 0 935000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_517
timestamp 1654889802
transform 0 -1 778000 1 0 933000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_518
timestamp 1654889802
transform 0 -1 778000 1 0 939000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_519
timestamp 1654889802
transform 0 -1 778000 1 0 937000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_520
timestamp 1654889802
transform 0 -1 778000 1 0 943000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_521
timestamp 1654889802
transform 0 -1 778000 1 0 941000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_522
timestamp 1654889802
transform 0 -1 778000 1 0 947000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_523
timestamp 1654889802
transform 0 -1 778000 1 0 945000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_524
timestamp 1654889802
transform -1 0 695000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_525
timestamp 1654889802
transform -1 0 697000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_526
timestamp 1654889802
transform -1 0 707000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_527
timestamp 1654889802
transform -1 0 705000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_528
timestamp 1654889802
transform -1 0 703000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_529
timestamp 1654889802
transform -1 0 701000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_530
timestamp 1654889802
transform -1 0 699000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_531
timestamp 1654889802
transform -1 0 679000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_532
timestamp 1654889802
transform -1 0 681000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_533
timestamp 1654889802
transform -1 0 683000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_534
timestamp 1654889802
transform -1 0 685000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_535
timestamp 1654889802
transform -1 0 687000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_536
timestamp 1654889802
transform -1 0 689000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_537
timestamp 1654889802
transform -1 0 693000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_538
timestamp 1654889802
transform -1 0 691000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_539
timestamp 1654889802
transform -1 0 677000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_540
timestamp 1654889802
transform -1 0 675000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_541
timestamp 1654889802
transform -1 0 673000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_542
timestamp 1654889802
transform -1 0 654000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_543
timestamp 1654889802
transform -1 0 652000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_544
timestamp 1654889802
transform -1 0 650000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_545
timestamp 1654889802
transform -1 0 656000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_546
timestamp 1654889802
transform -1 0 638000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_547
timestamp 1654889802
transform -1 0 636000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_548
timestamp 1654889802
transform -1 0 634000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_549
timestamp 1654889802
transform -1 0 646000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_550
timestamp 1654889802
transform -1 0 644000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_551
timestamp 1654889802
transform -1 0 642000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_552
timestamp 1654889802
transform -1 0 640000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_553
timestamp 1654889802
transform -1 0 648000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_554
timestamp 1654889802
transform -1 0 624000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_555
timestamp 1654889802
transform -1 0 622000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_556
timestamp 1654889802
transform -1 0 620000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_557
timestamp 1654889802
transform -1 0 632000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_558
timestamp 1654889802
transform -1 0 630000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_559
timestamp 1654889802
transform -1 0 628000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_560
timestamp 1654889802
transform -1 0 626000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_561
timestamp 1654889802
transform -1 0 618000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_562
timestamp 1654889802
transform -1 0 589000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_563
timestamp 1654889802
transform -1 0 591000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_564
timestamp 1654889802
transform -1 0 593000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_565
timestamp 1654889802
transform -1 0 595000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_566
timestamp 1654889802
transform -1 0 597000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_567
timestamp 1654889802
transform -1 0 599000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_568
timestamp 1654889802
transform -1 0 601000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_569
timestamp 1654889802
transform -1 0 577000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_570
timestamp 1654889802
transform -1 0 575000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_571
timestamp 1654889802
transform -1 0 583000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_572
timestamp 1654889802
transform -1 0 581000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_573
timestamp 1654889802
transform -1 0 579000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_574
timestamp 1654889802
transform -1 0 585000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_575
timestamp 1654889802
transform -1 0 587000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_576
timestamp 1654889802
transform -1 0 567000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_577
timestamp 1654889802
transform -1 0 565000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_578
timestamp 1654889802
transform -1 0 563000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_579
timestamp 1654889802
transform -1 0 573000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_580
timestamp 1654889802
transform -1 0 571000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_581
timestamp 1654889802
transform -1 0 569000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_582
timestamp 1654889802
transform -1 0 546000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_583
timestamp 1654889802
transform -1 0 544000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_584
timestamp 1654889802
transform -1 0 530000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_585
timestamp 1654889802
transform -1 0 532000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_586
timestamp 1654889802
transform -1 0 528000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_587
timestamp 1654889802
transform -1 0 538000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_588
timestamp 1654889802
transform -1 0 536000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_589
timestamp 1654889802
transform -1 0 534000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_590
timestamp 1654889802
transform -1 0 542000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_591
timestamp 1654889802
transform -1 0 540000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_592
timestamp 1654889802
transform -1 0 514000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_593
timestamp 1654889802
transform -1 0 516000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_594
timestamp 1654889802
transform -1 0 518000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_595
timestamp 1654889802
transform -1 0 520000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_596
timestamp 1654889802
transform -1 0 522000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_597
timestamp 1654889802
transform -1 0 524000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_598
timestamp 1654889802
transform -1 0 526000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_599
timestamp 1654889802
transform -1 0 508000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_600
timestamp 1654889802
transform -1 0 510000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_601
timestamp 1654889802
transform -1 0 512000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_602
timestamp 1654889802
transform -1 0 485000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_603
timestamp 1654889802
transform -1 0 483000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_604
timestamp 1654889802
transform -1 0 487000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_605
timestamp 1654889802
transform -1 0 489000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_606
timestamp 1654889802
transform -1 0 491000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_607
timestamp 1654889802
transform -1 0 469000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_608
timestamp 1654889802
transform -1 0 471000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_609
timestamp 1654889802
transform -1 0 473000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_610
timestamp 1654889802
transform -1 0 475000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_611
timestamp 1654889802
transform -1 0 477000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_612
timestamp 1654889802
transform -1 0 479000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_613
timestamp 1654889802
transform -1 0 481000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_614
timestamp 1654889802
transform -1 0 455000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_615
timestamp 1654889802
transform -1 0 453000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_616
timestamp 1654889802
transform -1 0 463000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_617
timestamp 1654889802
transform -1 0 461000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_618
timestamp 1654889802
transform -1 0 459000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_619
timestamp 1654889802
transform -1 0 457000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_620
timestamp 1654889802
transform -1 0 465000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_621
timestamp 1654889802
transform -1 0 467000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_622
timestamp 1654889802
transform -1 0 424000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_623
timestamp 1654889802
transform -1 0 426000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_624
timestamp 1654889802
transform -1 0 428000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_625
timestamp 1654889802
transform -1 0 430000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_626
timestamp 1654889802
transform -1 0 432000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_627
timestamp 1654889802
transform -1 0 434000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_628
timestamp 1654889802
transform -1 0 436000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_629
timestamp 1654889802
transform -1 0 408000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_630
timestamp 1654889802
transform -1 0 410000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_631
timestamp 1654889802
transform -1 0 412000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_632
timestamp 1654889802
transform -1 0 414000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_633
timestamp 1654889802
transform -1 0 416000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_634
timestamp 1654889802
transform -1 0 418000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_635
timestamp 1654889802
transform -1 0 420000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_636
timestamp 1654889802
transform -1 0 422000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_637
timestamp 1654889802
transform -1 0 402000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_638
timestamp 1654889802
transform -1 0 400000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_639
timestamp 1654889802
transform -1 0 398000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_640
timestamp 1654889802
transform -1 0 404000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_641
timestamp 1654889802
transform -1 0 406000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_642
timestamp 1654889802
transform -1 0 381000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_643
timestamp 1654889802
transform -1 0 379000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_644
timestamp 1654889802
transform -1 0 367000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_645
timestamp 1654889802
transform -1 0 369000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_646
timestamp 1654889802
transform -1 0 365000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_647
timestamp 1654889802
transform -1 0 363000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_648
timestamp 1654889802
transform -1 0 371000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_649
timestamp 1654889802
transform -1 0 377000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_650
timestamp 1654889802
transform -1 0 375000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_651
timestamp 1654889802
transform -1 0 373000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_652
timestamp 1654889802
transform -1 0 355000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_653
timestamp 1654889802
transform -1 0 353000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_654
timestamp 1654889802
transform -1 0 351000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_655
timestamp 1654889802
transform -1 0 349000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_656
timestamp 1654889802
transform -1 0 359000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_657
timestamp 1654889802
transform -1 0 357000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_658
timestamp 1654889802
transform -1 0 361000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_659
timestamp 1654889802
transform -1 0 347000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_660
timestamp 1654889802
transform -1 0 345000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_661
timestamp 1654889802
transform -1 0 343000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_662
timestamp 1654889802
transform -1 0 324000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_663
timestamp 1654889802
transform -1 0 322000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_664
timestamp 1654889802
transform -1 0 320000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_665
timestamp 1654889802
transform -1 0 318000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_666
timestamp 1654889802
transform -1 0 326000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_667
timestamp 1654889802
transform -1 0 304000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_668
timestamp 1654889802
transform -1 0 302000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_669
timestamp 1654889802
transform -1 0 308000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_670
timestamp 1654889802
transform -1 0 306000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_671
timestamp 1654889802
transform -1 0 314000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_672
timestamp 1654889802
transform -1 0 310000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_673
timestamp 1654889802
transform -1 0 312000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_674
timestamp 1654889802
transform -1 0 316000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_675
timestamp 1654889802
transform -1 0 288000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_676
timestamp 1654889802
transform -1 0 292000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_677
timestamp 1654889802
transform -1 0 290000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_678
timestamp 1654889802
transform -1 0 296000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_679
timestamp 1654889802
transform -1 0 294000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_680
timestamp 1654889802
transform -1 0 298000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_681
timestamp 1654889802
transform -1 0 300000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_682
timestamp 1654889802
transform -1 0 257000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_683
timestamp 1654889802
transform -1 0 259000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_684
timestamp 1654889802
transform -1 0 261000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_685
timestamp 1654889802
transform -1 0 263000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_686
timestamp 1654889802
transform -1 0 265000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_687
timestamp 1654889802
transform -1 0 267000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_688
timestamp 1654889802
transform -1 0 269000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_689
timestamp 1654889802
transform -1 0 271000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_690
timestamp 1654889802
transform -1 0 243000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_691
timestamp 1654889802
transform -1 0 245000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_692
timestamp 1654889802
transform -1 0 247000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_693
timestamp 1654889802
transform -1 0 249000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_694
timestamp 1654889802
transform -1 0 253000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_695
timestamp 1654889802
transform -1 0 251000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_696
timestamp 1654889802
transform -1 0 255000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_697
timestamp 1654889802
transform -1 0 239000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_698
timestamp 1654889802
transform -1 0 241000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_699
timestamp 1654889802
transform -1 0 235000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_700
timestamp 1654889802
transform -1 0 237000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_701
timestamp 1654889802
transform -1 0 233000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_702
timestamp 1654889802
transform -1 0 212000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_703
timestamp 1654889802
transform -1 0 214000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_704
timestamp 1654889802
transform -1 0 216000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_705
timestamp 1654889802
transform -1 0 198000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_706
timestamp 1654889802
transform -1 0 210000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_707
timestamp 1654889802
transform -1 0 208000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_708
timestamp 1654889802
transform -1 0 206000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_709
timestamp 1654889802
transform -1 0 204000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_710
timestamp 1654889802
transform -1 0 200000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_711
timestamp 1654889802
transform -1 0 202000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_712
timestamp 1654889802
transform -1 0 182000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_713
timestamp 1654889802
transform -1 0 184000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_714
timestamp 1654889802
transform -1 0 196000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_715
timestamp 1654889802
transform -1 0 192000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_716
timestamp 1654889802
transform -1 0 194000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_717
timestamp 1654889802
transform -1 0 188000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_718
timestamp 1654889802
transform -1 0 190000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_719
timestamp 1654889802
transform -1 0 186000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_720
timestamp 1654889802
transform -1 0 180000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_721
timestamp 1654889802
transform -1 0 178000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_722
timestamp 1654889802
transform -1 0 153000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_723
timestamp 1654889802
transform -1 0 157000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_724
timestamp 1654889802
transform -1 0 155000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_725
timestamp 1654889802
transform -1 0 161000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_726
timestamp 1654889802
transform -1 0 159000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_727
timestamp 1654889802
transform -1 0 141000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_728
timestamp 1654889802
transform -1 0 137000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_729
timestamp 1654889802
transform -1 0 139000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_730
timestamp 1654889802
transform -1 0 143000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_731
timestamp 1654889802
transform -1 0 151000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_732
timestamp 1654889802
transform -1 0 149000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_733
timestamp 1654889802
transform -1 0 145000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_734
timestamp 1654889802
transform -1 0 147000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_735
timestamp 1654889802
transform -1 0 125000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_736
timestamp 1654889802
transform -1 0 127000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_737
timestamp 1654889802
transform -1 0 123000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_738
timestamp 1654889802
transform -1 0 133000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_739
timestamp 1654889802
transform -1 0 135000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_740
timestamp 1654889802
transform -1 0 129000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_741
timestamp 1654889802
transform -1 0 131000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_742
timestamp 1654889802
transform -1 0 92000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_743
timestamp 1654889802
transform -1 0 94000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_744
timestamp 1654889802
transform -1 0 96000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_745
timestamp 1654889802
transform -1 0 98000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_746
timestamp 1654889802
transform -1 0 100000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_747
timestamp 1654889802
transform -1 0 106000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_748
timestamp 1654889802
transform -1 0 104000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_749
timestamp 1654889802
transform -1 0 102000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_750
timestamp 1654889802
transform -1 0 76000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_751
timestamp 1654889802
transform -1 0 78000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_752
timestamp 1654889802
transform -1 0 80000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_753
timestamp 1654889802
transform -1 0 82000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_754
timestamp 1654889802
transform -1 0 84000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_755
timestamp 1654889802
transform -1 0 86000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_756
timestamp 1654889802
transform -1 0 88000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_757
timestamp 1654889802
transform -1 0 90000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_758
timestamp 1654889802
transform -1 0 74000 0 -1 1020000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_759
timestamp 1654889802
transform 0 1 0 -1 0 946000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_760
timestamp 1654889802
transform 0 1 0 -1 0 948000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_761
timestamp 1654889802
transform 0 1 0 -1 0 108000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_762
timestamp 1654889802
transform 0 1 0 -1 0 940000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_763
timestamp 1654889802
transform 0 1 0 -1 0 942000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_764
timestamp 1654889802
transform 0 1 0 -1 0 944000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_765
timestamp 1654889802
transform 0 1 0 -1 0 938000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_766
timestamp 1654889802
transform 0 1 0 -1 0 934000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_767
timestamp 1654889802
transform 0 1 0 -1 0 936000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_768
timestamp 1654889802
transform 0 1 0 -1 0 928000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_769
timestamp 1654889802
transform 0 1 0 -1 0 932000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_770
timestamp 1654889802
transform 0 1 0 -1 0 930000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_771
timestamp 1654889802
transform 0 1 0 -1 0 909000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_772
timestamp 1654889802
transform 0 1 0 -1 0 911000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_773
timestamp 1654889802
transform 0 1 0 -1 0 110000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_774
timestamp 1654889802
transform 0 1 0 -1 0 901000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_775
timestamp 1654889802
transform 0 1 0 -1 0 899000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_776
timestamp 1654889802
transform 0 1 0 -1 0 905000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_777
timestamp 1654889802
transform 0 1 0 -1 0 907000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_778
timestamp 1654889802
transform 0 1 0 -1 0 903000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_779
timestamp 1654889802
transform 0 1 0 -1 0 895000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_780
timestamp 1654889802
transform 0 1 0 -1 0 897000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_781
timestamp 1654889802
transform 0 1 0 -1 0 887000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_782
timestamp 1654889802
transform 0 1 0 -1 0 893000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_783
timestamp 1654889802
transform 0 1 0 -1 0 889000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_784
timestamp 1654889802
transform 0 1 0 -1 0 891000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_785
timestamp 1654889802
transform 0 1 0 -1 0 112000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_786
timestamp 1654889802
transform 0 1 0 -1 0 866000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_787
timestamp 1654889802
transform 0 1 0 -1 0 868000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_788
timestamp 1654889802
transform 0 1 0 -1 0 870000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_789
timestamp 1654889802
transform 0 1 0 -1 0 860000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_790
timestamp 1654889802
transform 0 1 0 -1 0 864000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_791
timestamp 1654889802
transform 0 1 0 -1 0 862000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_792
timestamp 1654889802
transform 0 1 0 -1 0 852000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_793
timestamp 1654889802
transform 0 1 0 -1 0 856000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_794
timestamp 1654889802
transform 0 1 0 -1 0 854000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_795
timestamp 1654889802
transform 0 1 0 -1 0 858000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_796
timestamp 1654889802
transform 0 1 0 -1 0 848000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_797
timestamp 1654889802
transform 0 1 0 -1 0 846000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_798
timestamp 1654889802
transform 0 1 0 -1 0 850000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_799
timestamp 1654889802
transform 0 1 0 -1 0 823000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_800
timestamp 1654889802
transform 0 1 0 -1 0 114000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_801
timestamp 1654889802
transform 0 1 0 -1 0 829000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_802
timestamp 1654889802
transform 0 1 0 -1 0 827000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_803
timestamp 1654889802
transform 0 1 0 -1 0 825000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_804
timestamp 1654889802
transform 0 1 0 -1 0 821000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_805
timestamp 1654889802
transform 0 1 0 -1 0 817000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_806
timestamp 1654889802
transform 0 1 0 -1 0 819000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_807
timestamp 1654889802
transform 0 1 0 -1 0 815000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_808
timestamp 1654889802
transform 0 1 0 -1 0 811000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_809
timestamp 1654889802
transform 0 1 0 -1 0 809000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_810
timestamp 1654889802
transform 0 1 0 -1 0 813000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_811
timestamp 1654889802
transform 0 1 0 -1 0 807000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_812
timestamp 1654889802
transform 0 1 0 -1 0 805000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_813
timestamp 1654889802
transform 0 1 0 -1 0 782000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_814
timestamp 1654889802
transform 0 1 0 -1 0 780000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_815
timestamp 1654889802
transform 0 1 0 -1 0 784000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_816
timestamp 1654889802
transform 0 1 0 -1 0 786000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_817
timestamp 1654889802
transform 0 1 0 -1 0 788000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_818
timestamp 1654889802
transform 0 1 0 -1 0 116000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_819
timestamp 1654889802
transform 0 1 0 -1 0 778000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_820
timestamp 1654889802
transform 0 1 0 -1 0 766000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_821
timestamp 1654889802
transform 0 1 0 -1 0 770000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_822
timestamp 1654889802
transform 0 1 0 -1 0 768000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_823
timestamp 1654889802
transform 0 1 0 -1 0 774000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_824
timestamp 1654889802
transform 0 1 0 -1 0 772000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_825
timestamp 1654889802
transform 0 1 0 -1 0 776000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_826
timestamp 1654889802
transform 0 1 0 -1 0 764000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_827
timestamp 1654889802
transform 0 1 0 -1 0 118000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_828
timestamp 1654889802
transform 0 1 0 -1 0 747000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_829
timestamp 1654889802
transform 0 1 0 -1 0 745000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_830
timestamp 1654889802
transform 0 1 0 -1 0 743000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_831
timestamp 1654889802
transform 0 1 0 -1 0 739000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_832
timestamp 1654889802
transform 0 1 0 -1 0 741000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_833
timestamp 1654889802
transform 0 1 0 -1 0 737000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_834
timestamp 1654889802
transform 0 1 0 -1 0 735000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_835
timestamp 1654889802
transform 0 1 0 -1 0 731000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_836
timestamp 1654889802
transform 0 1 0 -1 0 733000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_837
timestamp 1654889802
transform 0 1 0 -1 0 727000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_838
timestamp 1654889802
transform 0 1 0 -1 0 729000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_839
timestamp 1654889802
transform 0 1 0 -1 0 725000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_840
timestamp 1654889802
transform 0 1 0 -1 0 723000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_841
timestamp 1654889802
transform 0 1 0 -1 0 706000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_842
timestamp 1654889802
transform 0 1 0 -1 0 704000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_843
timestamp 1654889802
transform 0 1 0 -1 0 702000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_844
timestamp 1654889802
transform 0 1 0 -1 0 698000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_845
timestamp 1654889802
transform 0 1 0 -1 0 700000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_846
timestamp 1654889802
transform 0 1 0 -1 0 696000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_847
timestamp 1654889802
transform 0 1 0 -1 0 120000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_848
timestamp 1654889802
transform 0 1 0 -1 0 694000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_849
timestamp 1654889802
transform 0 1 0 -1 0 690000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_850
timestamp 1654889802
transform 0 1 0 -1 0 686000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_851
timestamp 1654889802
transform 0 1 0 -1 0 688000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_852
timestamp 1654889802
transform 0 1 0 -1 0 682000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_853
timestamp 1654889802
transform 0 1 0 -1 0 684000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_854
timestamp 1654889802
transform 0 1 0 -1 0 692000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_855
timestamp 1654889802
transform 0 1 0 -1 0 665000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_856
timestamp 1654889802
transform 0 1 0 -1 0 122000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_857
timestamp 1654889802
transform 0 1 0 -1 0 659000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_858
timestamp 1654889802
transform 0 1 0 -1 0 657000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_859
timestamp 1654889802
transform 0 1 0 -1 0 661000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_860
timestamp 1654889802
transform 0 1 0 -1 0 663000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_861
timestamp 1654889802
transform 0 1 0 -1 0 651000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_862
timestamp 1654889802
transform 0 1 0 -1 0 655000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_863
timestamp 1654889802
transform 0 1 0 -1 0 653000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_864
timestamp 1654889802
transform 0 1 0 -1 0 643000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_865
timestamp 1654889802
transform 0 1 0 -1 0 647000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_866
timestamp 1654889802
transform 0 1 0 -1 0 645000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_867
timestamp 1654889802
transform 0 1 0 -1 0 649000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_868
timestamp 1654889802
transform 0 1 0 -1 0 641000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_869
timestamp 1654889802
transform 0 1 0 -1 0 622000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_870
timestamp 1654889802
transform 0 1 0 -1 0 624000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_871
timestamp 1654889802
transform 0 1 0 -1 0 124000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_872
timestamp 1654889802
transform 0 1 0 -1 0 618000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_873
timestamp 1654889802
transform 0 1 0 -1 0 616000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_874
timestamp 1654889802
transform 0 1 0 -1 0 620000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_875
timestamp 1654889802
transform 0 1 0 -1 0 614000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_876
timestamp 1654889802
transform 0 1 0 -1 0 610000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_877
timestamp 1654889802
transform 0 1 0 -1 0 608000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_878
timestamp 1654889802
transform 0 1 0 -1 0 612000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_879
timestamp 1654889802
transform 0 1 0 -1 0 602000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_880
timestamp 1654889802
transform 0 1 0 -1 0 600000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_881
timestamp 1654889802
transform 0 1 0 -1 0 606000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_882
timestamp 1654889802
transform 0 1 0 -1 0 604000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_883
timestamp 1654889802
transform 0 1 0 -1 0 579000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_884
timestamp 1654889802
transform 0 1 0 -1 0 581000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_885
timestamp 1654889802
transform 0 1 0 -1 0 583000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_886
timestamp 1654889802
transform 0 1 0 -1 0 126000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_887
timestamp 1654889802
transform 0 1 0 -1 0 577000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_888
timestamp 1654889802
transform 0 1 0 -1 0 575000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_889
timestamp 1654889802
transform 0 1 0 -1 0 565000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_890
timestamp 1654889802
transform 0 1 0 -1 0 569000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_891
timestamp 1654889802
transform 0 1 0 -1 0 567000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_892
timestamp 1654889802
transform 0 1 0 -1 0 571000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_893
timestamp 1654889802
transform 0 1 0 -1 0 573000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_894
timestamp 1654889802
transform 0 1 0 -1 0 561000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_895
timestamp 1654889802
transform 0 1 0 -1 0 563000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_896
timestamp 1654889802
transform 0 1 0 -1 0 559000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_897
timestamp 1654889802
transform 0 1 0 -1 0 536000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_898
timestamp 1654889802
transform 0 1 0 -1 0 538000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_899
timestamp 1654889802
transform 0 1 0 -1 0 540000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_900
timestamp 1654889802
transform 0 1 0 -1 0 542000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_901
timestamp 1654889802
transform 0 1 0 -1 0 128000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_902
timestamp 1654889802
transform 0 1 0 -1 0 532000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_903
timestamp 1654889802
transform 0 1 0 -1 0 534000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_904
timestamp 1654889802
transform 0 1 0 -1 0 524000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_905
timestamp 1654889802
transform 0 1 0 -1 0 522000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_906
timestamp 1654889802
transform 0 1 0 -1 0 528000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_907
timestamp 1654889802
transform 0 1 0 -1 0 526000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_908
timestamp 1654889802
transform 0 1 0 -1 0 530000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_909
timestamp 1654889802
transform 0 1 0 -1 0 518000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_910
timestamp 1654889802
transform 0 1 0 -1 0 520000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_911
timestamp 1654889802
transform 0 1 0 -1 0 495000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_912
timestamp 1654889802
transform 0 1 0 -1 0 493000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_913
timestamp 1654889802
transform 0 1 0 -1 0 497000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_914
timestamp 1654889802
transform 0 1 0 -1 0 499000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_915
timestamp 1654889802
transform 0 1 0 -1 0 501000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_916
timestamp 1654889802
transform 0 1 0 -1 0 130000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_917
timestamp 1654889802
transform 0 1 0 -1 0 479000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_918
timestamp 1654889802
transform 0 1 0 -1 0 483000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_919
timestamp 1654889802
transform 0 1 0 -1 0 481000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_920
timestamp 1654889802
transform 0 1 0 -1 0 487000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_921
timestamp 1654889802
transform 0 1 0 -1 0 485000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_922
timestamp 1654889802
transform 0 1 0 -1 0 489000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_923
timestamp 1654889802
transform 0 1 0 -1 0 491000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_924
timestamp 1654889802
transform 0 1 0 -1 0 477000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_925
timestamp 1654889802
transform 0 1 0 -1 0 132000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_926
timestamp 1654889802
transform 0 1 0 -1 0 460000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_927
timestamp 1654889802
transform 0 1 0 -1 0 458000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_928
timestamp 1654889802
transform 0 1 0 -1 0 456000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_929
timestamp 1654889802
transform 0 1 0 -1 0 454000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_930
timestamp 1654889802
transform 0 1 0 -1 0 450000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_931
timestamp 1654889802
transform 0 1 0 -1 0 452000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_932
timestamp 1654889802
transform 0 1 0 -1 0 448000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_933
timestamp 1654889802
transform 0 1 0 -1 0 444000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_934
timestamp 1654889802
transform 0 1 0 -1 0 446000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_935
timestamp 1654889802
transform 0 1 0 -1 0 442000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_936
timestamp 1654889802
transform 0 1 0 -1 0 440000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_937
timestamp 1654889802
transform 0 1 0 -1 0 436000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_938
timestamp 1654889802
transform 0 1 0 -1 0 438000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_940
timestamp 1654889802
transform 0 1 0 -1 0 411000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_941
timestamp 1654889802
transform 0 1 0 -1 0 413000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_942
timestamp 1654889802
transform 0 1 0 -1 0 419000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_943
timestamp 1654889802
transform 0 1 0 -1 0 417000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_944
timestamp 1654889802
transform 0 1 0 -1 0 415000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_945
timestamp 1654889802
transform 0 1 0 -1 0 407000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_946
timestamp 1654889802
transform 0 1 0 -1 0 409000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_947
timestamp 1654889802
transform 0 1 0 -1 0 405000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_948
timestamp 1654889802
transform 0 1 0 -1 0 403000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_949
timestamp 1654889802
transform 0 1 0 -1 0 399000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_950
timestamp 1654889802
transform 0 1 0 -1 0 401000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_951
timestamp 1654889802
transform 0 1 0 -1 0 397000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_952
timestamp 1654889802
transform 0 1 0 -1 0 395000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_953
timestamp 1654889802
transform 0 1 0 -1 0 378000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_955
timestamp 1654889802
transform 0 1 0 -1 0 372000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_956
timestamp 1654889802
transform 0 1 0 -1 0 374000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_957
timestamp 1654889802
transform 0 1 0 -1 0 376000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_958
timestamp 1654889802
transform 0 1 0 -1 0 368000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_959
timestamp 1654889802
transform 0 1 0 -1 0 366000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_960
timestamp 1654889802
transform 0 1 0 -1 0 370000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_961
timestamp 1654889802
transform 0 1 0 -1 0 364000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_962
timestamp 1654889802
transform 0 1 0 -1 0 360000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_963
timestamp 1654889802
transform 0 1 0 -1 0 358000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_964
timestamp 1654889802
transform 0 1 0 -1 0 362000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_965
timestamp 1654889802
transform 0 1 0 -1 0 356000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_966
timestamp 1654889802
transform 0 1 0 -1 0 354000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_967
timestamp 1654889802
transform 0 1 0 -1 0 335000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_968
timestamp 1654889802
transform 0 1 0 -1 0 337000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_970
timestamp 1654889802
transform 0 1 0 -1 0 331000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_971
timestamp 1654889802
transform 0 1 0 -1 0 329000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_972
timestamp 1654889802
transform 0 1 0 -1 0 333000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_973
timestamp 1654889802
transform 0 1 0 -1 0 327000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_974
timestamp 1654889802
transform 0 1 0 -1 0 323000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_975
timestamp 1654889802
transform 0 1 0 -1 0 321000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_976
timestamp 1654889802
transform 0 1 0 -1 0 325000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_977
timestamp 1654889802
transform 0 1 0 -1 0 319000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_978
timestamp 1654889802
transform 0 1 0 -1 0 315000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_979
timestamp 1654889802
transform 0 1 0 -1 0 313000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_980
timestamp 1654889802
transform 0 1 0 -1 0 317000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_981
timestamp 1654889802
transform 0 1 0 -1 0 292000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_982
timestamp 1654889802
transform 0 1 0 -1 0 294000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_983
timestamp 1654889802
transform 0 1 0 -1 0 296000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_985
timestamp 1654889802
transform 0 1 0 -1 0 290000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_986
timestamp 1654889802
transform 0 1 0 -1 0 278000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_987
timestamp 1654889802
transform 0 1 0 -1 0 282000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_988
timestamp 1654889802
transform 0 1 0 -1 0 280000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_989
timestamp 1654889802
transform 0 1 0 -1 0 286000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_990
timestamp 1654889802
transform 0 1 0 -1 0 284000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_991
timestamp 1654889802
transform 0 1 0 -1 0 288000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_992
timestamp 1654889802
transform 0 1 0 -1 0 276000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_993
timestamp 1654889802
transform 0 1 0 -1 0 272000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_994
timestamp 1654889802
transform 0 1 0 -1 0 274000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_995
timestamp 1654889802
transform 0 1 0 -1 0 251000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_996
timestamp 1654889802
transform 0 1 0 -1 0 253000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_997
timestamp 1654889802
transform 0 1 0 -1 0 255000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_999
timestamp 1654889802
transform 0 1 0 -1 0 249000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1000
timestamp 1654889802
transform 0 1 0 -1 0 237000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1001
timestamp 1654889802
transform 0 1 0 -1 0 241000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1002
timestamp 1654889802
transform 0 1 0 -1 0 239000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1003
timestamp 1654889802
transform 0 1 0 -1 0 245000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1004
timestamp 1654889802
transform 0 1 0 -1 0 243000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1005
timestamp 1654889802
transform 0 1 0 -1 0 247000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1006
timestamp 1654889802
transform 0 1 0 -1 0 233000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1007
timestamp 1654889802
transform 0 1 0 -1 0 235000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1008
timestamp 1654889802
transform 0 1 0 -1 0 231000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1009
timestamp 1654889802
transform 0 1 0 -1 0 212000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1010
timestamp 1654889802
transform 0 1 0 -1 0 210000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1011
timestamp 1654889802
transform 0 1 0 -1 0 208000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1013
timestamp 1654889802
transform 0 1 0 -1 0 214000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1014
timestamp 1654889802
transform 0 1 0 -1 0 206000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1015
timestamp 1654889802
transform 0 1 0 -1 0 194000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1016
timestamp 1654889802
transform 0 1 0 -1 0 196000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1017
timestamp 1654889802
transform 0 1 0 -1 0 202000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1018
timestamp 1654889802
transform 0 1 0 -1 0 204000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1019
timestamp 1654889802
transform 0 1 0 -1 0 198000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1020
timestamp 1654889802
transform 0 1 0 -1 0 200000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1021
timestamp 1654889802
transform 0 1 0 -1 0 190000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1022
timestamp 1654889802
transform 0 1 0 -1 0 192000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1024
timestamp 1654889802
transform 0 1 0 -1 0 173000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1025
timestamp 1654889802
transform 0 1 0 -1 0 171000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1026
timestamp 1654889802
transform 0 1 0 -1 0 169000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1027
timestamp 1654889802
transform 0 1 0 -1 0 165000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1028
timestamp 1654889802
transform 0 1 0 -1 0 167000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1029
timestamp 1654889802
transform 0 1 0 -1 0 163000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1030
timestamp 1654889802
transform 0 1 0 -1 0 161000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1031
timestamp 1654889802
transform 0 1 0 -1 0 157000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1032
timestamp 1654889802
transform 0 1 0 -1 0 159000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1033
timestamp 1654889802
transform 0 1 0 -1 0 155000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1034
timestamp 1654889802
transform 0 1 0 -1 0 153000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1035
timestamp 1654889802
transform 0 1 0 -1 0 149000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1036
timestamp 1654889802
transform 0 1 0 -1 0 151000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1038
timestamp 1654889802
transform 0 1 0 -1 0 91000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1039
timestamp 1654889802
transform 0 1 0 -1 0 89000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1040
timestamp 1654889802
transform 0 1 0 -1 0 87000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1041
timestamp 1654889802
transform 0 1 0 -1 0 85000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1042
timestamp 1654889802
transform 0 1 0 -1 0 83000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1043
timestamp 1654889802
transform 0 1 0 -1 0 79000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1044
timestamp 1654889802
transform 0 1 0 -1 0 81000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1045
timestamp 1654889802
transform 0 1 0 -1 0 75000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1046
timestamp 1654889802
transform 0 1 0 -1 0 77000
box -32 13097 2032 69968
use GF_NI_FILL10  GF_NI_FILL10_1047
timestamp 1654889802
transform 0 1 0 -1 0 73000
box -32 13097 2032 69968
use GF_NI_IN_C  GF_NI_IN_C_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 217000 0 1 0
box -32 0 15032 70000
use GF_NI_IN_S  GF_NI_IN_S_0 $PDKPATH/libs.ref/gf180mcu_io/mag
timestamp 1654889802
transform 1 0 162000 0 1 0
box -32 0 15032 70000
<< labels >>
flabel metal5 108500 400 120500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 163500 400 175500 12400 0 FreeSans 24000 0 0 0 resetb
port 446 nsew
flabel metal5 273500 400 285500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 328500 400 340500 12400 0 FreeSans 24000 0 0 0 flash_csb
port 5 nsew
flabel metal5 383500 400 395500 12400 0 FreeSans 24000 0 0 0 flash_clk
port 2 nsew
flabel metal5 438500 400 450500 12400 0 FreeSans 24000 0 0 0 flash_io0
port 8 nsew
flabel metal5 493500 400 505500 12400 0 FreeSans 24000 0 0 0 flash_io1
port 13 nsew
flabel metal5 548500 400 560500 12400 0 FreeSans 24000 0 0 0 gpio
port 18 nsew
flabel metal5 603500 400 615500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 658500 400 670500 12400 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 96500 777600 108500 0 FreeSans 24000 0 0 0 mprj_io[0]
port 29 nsew
flabel metal5 765600 139500 777600 151500 0 FreeSans 24000 0 0 0 mprj_io[1]
port 40 nsew
flabel metal5 765600 182500 777600 194500 0 FreeSans 24000 0 0 0 mprj_io[2]
port 51 nsew
flabel metal5 765600 225500 777600 237500 0 FreeSans 24000 0 0 0 mprj_io[3]
port 60 nsew
flabel metal5 765600 268500 777600 280500 0 FreeSans 24000 0 0 0 mprj_io[4]
port 61 nsew
flabel metal5 765600 311500 777600 323500 0 FreeSans 24000 0 0 0 mprj_io[5]
port 62 nsew
flabel metal5 765600 354500 777600 366500 0 FreeSans 24000 0 0 0 mprj_io[6]
port 63 nsew
flabel metal5 765600 397500 777600 409500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 765600 440500 777600 452500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 765600 483500 777600 495500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 526500 777600 538500 0 FreeSans 24000 0 0 0 mprj_io[7]
port 64 nsew
flabel metal5 765600 569500 777600 581500 0 FreeSans 24000 0 0 0 mprj_io[8]
port 65 nsew
flabel metal5 765600 612500 777600 624500 0 FreeSans 24000 0 0 0 mprj_io[9]
port 66 nsew
flabel metal5 765600 655500 777600 667500 0 FreeSans 24000 0 0 0 mprj_io[10]
port 30 nsew
flabel metal5 765600 698500 777600 710500 0 FreeSans 24000 0 0 0 mprj_io[11]
port 31 nsew
flabel metal5 765600 741500 777600 753500 0 FreeSans 24000 0 0 0 mprj_io[12]
port 32 nsew
flabel metal5 765600 784500 777600 796500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 827500 777600 839500 0 FreeSans 24000 0 0 0 mprj_io[13]
port 33 nsew
flabel metal5 765600 870500 777600 882500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 913500 777600 925500 0 FreeSans 24000 0 0 0 mprj_io[14]
port 34 nsew
flabel metal5 657500 1007600 669500 1019600 0 FreeSans 24000 0 0 0 mprj_io[15]
port 35 nsew
flabel metal5 602500 1007600 614500 1019600 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 547500 1007600 559500 1019600 0 FreeSans 24000 0 0 0 mprj_io[16]
port 36 nsew
flabel metal5 492500 1007600 504500 1019600 0 FreeSans 24000 0 0 0 mprj_io[17]
port 37 nsew
flabel metal5 437500 1007600 449500 1019600 0 FreeSans 24000 0 0 0 mprj_io[18]
port 38 nsew
flabel metal5 382500 1007600 394500 1019600 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 327500 1007600 339500 1019600 0 FreeSans 24000 0 0 0 mprj_io[19]
port 39 nsew
flabel metal5 272500 1007600 284500 1019600 0 FreeSans 24000 0 0 0 mprj_io[20]
port 41 nsew
flabel metal5 217500 1007600 229500 1019600 0 FreeSans 24000 0 0 0 mprj_io[21]
port 42 nsew
flabel metal5 162500 1007600 174500 1019600 0 FreeSans 24000 0 0 0 mprj_io[22]
port 43 nsew
flabel metal5 107500 1007600 119500 1019600 0 FreeSans 24000 0 0 0 mprj_io[23]
port 44 nsew
flabel metal5 400 912500 12400 924500 0 FreeSans 24000 0 0 0 mprj_io[24]
port 45 nsew
flabel metal5 400 871500 12400 883500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 830500 12400 842500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 789500 12400 801500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 400 748500 12400 760500 0 FreeSans 24000 0 0 0 mprj_io[25]
port 46 nsew
flabel metal5 400 707500 12400 719500 0 FreeSans 24000 0 0 0 mprj_io[26]
port 47 nsew
flabel metal5 400 666500 12400 678500 0 FreeSans 24000 0 0 0 mprj_io[27]
port 48 nsew
flabel metal5 400 625500 12400 637500 0 FreeSans 24000 0 0 0 mprj_io[28]
port 49 nsew
flabel metal5 400 584500 12400 596500 0 FreeSans 24000 0 0 0 mprj_io[29]
port 50 nsew
flabel metal5 400 543500 12400 555500 0 FreeSans 24000 0 0 0 mprj_io[30]
port 52 nsew
flabel metal5 400 502500 12400 514500 0 FreeSans 24000 0 0 0 mprj_io[31]
port 53 nsew
flabel metal5 400 461500 12400 473500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 420500 12400 432500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 400 379500 12400 391500 0 FreeSans 24000 0 0 0 mprj_io[32]
port 54 nsew
flabel metal5 400 338500 12400 350500 0 FreeSans 24000 0 0 0 mprj_io[33]
port 55 nsew
flabel metal5 400 297500 12400 309500 0 FreeSans 24000 0 0 0 mprj_io[34]
port 56 nsew
flabel metal5 400 256500 12400 268500 0 FreeSans 24000 0 0 0 mprj_io[35]
port 57 nsew
flabel metal5 400 215500 12400 227500 0 FreeSans 24000 0 0 0 mprj_io[36]
port 58 nsew
flabel metal5 400 174500 12400 186500 0 FreeSans 24000 0 0 0 mprj_io[37]
port 59 nsew
flabel metal5 400 133500 12400 145500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 92500 12400 104500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 218500 400 230500 12400 0 FreeSans 24000 0 0 0 clock
port 0 nsew
flabel metal2 176172 69924 176248 70200 0 FreeSans 480 90 0 0 resetb_core
port 447 nsew
flabel metal2 231172 69924 231248 70200 0 FreeSans 480 90 0 0 clock_core
port 1 nsew
flabel metal2 395880 69924 395956 70200 0 FreeSans 480 90 0 0 flash_clk_core
port 3 nsew
flabel metal2 396026 69924 396102 70200 0 FreeSans 480 90 0 0 flash_clk_oe_core
port 4 nsew
flabel metal2 340880 69924 340956 70200 0 FreeSans 480 90 0 0 flash_csb_core
port 6 nsew
flabel metal2 341026 69924 341102 70200 0 FreeSans 480 90 0 0 flash_csb_oe_core
port 7 nsew
flabel metal2 439277 69924 439353 70200 0 FreeSans 480 90 0 0 flash_io0_ie_core
port 11 nsew
flabel metal2 450880 69924 450956 70200 0 FreeSans 480 90 0 0 flash_io0_do_core
port 10 nsew
flabel metal2 451026 69924 451102 70200 0 FreeSans 480 90 0 0 flash_io0_oe_core
port 12 nsew
flabel metal2 451171 69924 451247 70200 0 FreeSans 480 90 0 0 flash_io0_di_core
port 9 nsew
flabel metal2 494277 69924 494353 70200 0 FreeSans 480 90 0 0 flash_io1_ie_core
port 16 nsew
flabel metal2 505880 69924 505956 70200 0 FreeSans 480 90 0 0 flash_io1_do_core
port 15 nsew
flabel metal2 506026 69924 506102 70200 0 FreeSans 480 90 0 0 flash_io1_oe_core
port 17 nsew
flabel metal2 506172 69924 506248 70200 0 FreeSans 480 90 0 0 flash_io1_di_core
port 14 nsew
flabel metal2 547672 69924 547748 70200 0 FreeSans 480 90 0 0 gpio_schmitt_select
port 27 nsew
flabel metal2 548193 69924 548269 70200 0 FreeSans 480 90 0 0 gpio_pu_select
port 26 nsew
flabel metal2 548422 69924 548498 70200 0 FreeSans 480 90 0 0 gpio_drive_select_core[0]
port 19 nsew
flabel metal2 548564 69923 548640 70199 0 FreeSans 480 90 0 0 gpio_drive_select_core[1]
port 20 nsew
flabel metal2 549066 69924 549142 70200 0 FreeSans 480 90 0 0 gpio_pd_select
port 25 nsew
flabel metal2 549277 69924 549353 70200 0 FreeSans 480 90 0 0 gpio_inen_core
port 22 nsew
flabel metal2 560734 69924 560810 70200 0 FreeSans 480 90 0 0 gpio_slew_select
port 28 nsew
flabel metal2 560880 69924 560956 70200 0 FreeSans 480 90 0 0 gpio_out_core
port 23 nsew
flabel metal2 561172 69924 561248 70200 0 FreeSans 480 90 0 0 gpio_in_core
port 21 nsew
flabel metal2 561026 69924 561102 70200 0 FreeSans 480 90 0 0 gpio_outen_core
port 24 nsew
flabel metal2 707800 95672 708076 95748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[0]
port 370 nsew
flabel metal2 707800 96193 708076 96269 0 FreeSans 480 0 0 0 mprj_io_pu_select[0]
port 332 nsew
flabel metal2 707800 96422 708076 96498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[0]
port 67 nsew
flabel metal2 707800 96564 708076 96640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[1]
port 78 nsew
flabel metal2 707800 97066 708076 97142 0 FreeSans 480 0 0 0 mprj_io_pd_select[0]
port 294 nsew
flabel metal2 707800 97277 708076 97353 0 FreeSans 480 0 0 0 mprj_io_inen[0]
port 180 nsew
flabel metal2 707800 108734 708076 108810 0 FreeSans 480 0 0 0 mprj_io_slew_select[0]
port 408 nsew
flabel metal2 707800 108880 708076 108956 0 FreeSans 480 0 0 0 mprj_io_out[0]
port 218 nsew
flabel metal2 707800 109026 708076 109102 0 FreeSans 480 0 0 0 mprj_io_outen[0]
port 256 nsew
flabel metal2 707800 109172 708076 109248 0 FreeSans 480 0 0 0 mprj_io_in[0]
port 142 nsew
flabel metal2 707621 138672 707897 138748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[1]
port 381 nsew
flabel metal2 707621 139193 707897 139269 0 FreeSans 480 0 0 0 mprj_io_pu_select[1]
port 343 nsew
flabel metal2 707621 139422 707897 139498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[2]
port 89 nsew
flabel metal2 707621 139564 707897 139640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[3]
port 100 nsew
flabel metal2 707621 140066 707897 140142 0 FreeSans 480 0 0 0 mprj_io_pd_select[1]
port 305 nsew
flabel metal2 707621 140277 707897 140353 0 FreeSans 480 0 0 0 mprj_io_inen[1]
port 191 nsew
flabel metal2 707621 151734 707897 151810 0 FreeSans 480 0 0 0 mprj_io_slew_select[1]
port 419 nsew
flabel metal2 707621 151880 707897 151956 0 FreeSans 480 0 0 0 mprj_io_out[1]
port 229 nsew
flabel metal2 707621 152026 707897 152102 0 FreeSans 480 0 0 0 mprj_io_outen[1]
port 267 nsew
flabel metal2 707621 152172 707897 152248 0 FreeSans 480 0 0 0 mprj_io_in[1]
port 153 nsew
flabel metal2 707800 195172 708076 195248 0 FreeSans 480 0 0 0 mprj_io_in[2]
port 164 nsew
flabel metal2 707800 195026 708076 195102 0 FreeSans 480 0 0 0 mprj_io_outen[2]
port 278 nsew
flabel metal2 707800 194880 708076 194956 0 FreeSans 480 0 0 0 mprj_io_out[2]
port 240 nsew
flabel metal2 707800 194734 708076 194810 0 FreeSans 480 0 0 0 mprj_io_slew_select[2]
port 430 nsew
flabel metal2 707800 183277 708076 183353 0 FreeSans 480 0 0 0 mprj_io_inen[2]
port 202 nsew
flabel metal2 707800 183066 708076 183142 0 FreeSans 480 0 0 0 mprj_io_pd_select[2]
port 316 nsew
flabel metal2 707800 182564 708076 182640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[4]
port 111 nsew
flabel metal2 707800 182422 708076 182498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[5]
port 122 nsew
flabel metal2 707800 182193 708076 182269 0 FreeSans 480 0 0 0 mprj_io_pu_select[2]
port 354 nsew
flabel metal2 707800 181672 708076 181748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[2]
port 392 nsew
flabel metal2 707800 238172 708076 238248 0 FreeSans 480 0 0 0 mprj_io_in[3]
port 173 nsew
flabel metal2 707800 238026 708076 238102 0 FreeSans 480 0 0 0 mprj_io_outen[3]
port 287 nsew
flabel metal2 707800 237880 708076 237956 0 FreeSans 480 0 0 0 mprj_io_out[3]
port 249 nsew
flabel metal2 707800 237734 708076 237810 0 FreeSans 480 0 0 0 mprj_io_slew_select[3]
port 439 nsew
flabel metal2 707800 226277 708076 226353 0 FreeSans 480 0 0 0 mprj_io_inen[3]
port 211 nsew
flabel metal2 707800 226066 708076 226142 0 FreeSans 480 0 0 0 mprj_io_pd_select[3]
port 325 nsew
flabel metal2 707800 225564 708076 225640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[6]
port 132 nsew
flabel metal2 707800 225422 708076 225498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[7]
port 139 nsew
flabel metal2 707800 225193 708076 225269 0 FreeSans 480 0 0 0 mprj_io_pu_select[3]
port 363 nsew
flabel metal2 707800 224672 708076 224748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[3]
port 401 nsew
flabel metal2 707800 281172 708076 281248 0 FreeSans 480 0 0 0 mprj_io_in[4]
port 174 nsew
flabel metal2 707800 281026 708076 281102 0 FreeSans 480 0 0 0 mprj_io_outen[4]
port 288 nsew
flabel metal2 707800 280880 708076 280956 0 FreeSans 480 0 0 0 mprj_io_out[4]
port 250 nsew
flabel metal2 707800 280734 708076 280810 0 FreeSans 480 0 0 0 mprj_io_slew_select[4]
port 440 nsew
flabel metal2 707800 269277 708076 269353 0 FreeSans 480 0 0 0 mprj_io_inen[4]
port 212 nsew
flabel metal2 707800 269066 708076 269142 0 FreeSans 480 0 0 0 mprj_io_pd_select[4]
port 326 nsew
flabel metal2 707800 268564 708076 268640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[8]
port 140 nsew
flabel metal2 707800 268422 708076 268498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[9]
port 141 nsew
flabel metal2 707800 268193 708076 268269 0 FreeSans 480 0 0 0 mprj_io_pu_select[4]
port 364 nsew
flabel metal2 707800 267672 708076 267748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[4]
port 402 nsew
flabel metal2 707800 324172 708076 324248 0 FreeSans 480 0 0 0 mprj_io_in[5]
port 175 nsew
flabel metal2 707800 324026 708076 324102 0 FreeSans 480 0 0 0 mprj_io_outen[5]
port 289 nsew
flabel metal2 707800 323880 708076 323956 0 FreeSans 480 0 0 0 mprj_io_out[5]
port 251 nsew
flabel metal2 707800 323734 708076 323810 0 FreeSans 480 0 0 0 mprj_io_slew_select[5]
port 441 nsew
flabel metal2 707800 312277 708076 312353 0 FreeSans 480 0 0 0 mprj_io_inen[5]
port 213 nsew
flabel metal2 707800 312066 708076 312142 0 FreeSans 480 0 0 0 mprj_io_pd_select[5]
port 327 nsew
flabel metal2 707800 311564 708076 311640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[10]
port 68 nsew
flabel metal2 707800 311422 708076 311498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[11]
port 69 nsew
flabel metal2 707800 311193 708076 311269 0 FreeSans 480 0 0 0 mprj_io_pu_select[5]
port 365 nsew
flabel metal2 707800 310672 708076 310748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[5]
port 403 nsew
flabel metal2 707800 367172 708076 367248 0 FreeSans 480 0 0 0 mprj_io_in[6]
port 176 nsew
flabel metal2 707800 367026 708076 367102 0 FreeSans 480 0 0 0 mprj_io_outen[6]
port 290 nsew
flabel metal2 707800 366880 708076 366956 0 FreeSans 480 0 0 0 mprj_io_out[6]
port 252 nsew
flabel metal2 707800 366734 708076 366810 0 FreeSans 480 0 0 0 mprj_io_slew_select[6]
port 442 nsew
flabel metal2 707800 355277 708076 355353 0 FreeSans 480 0 0 0 mprj_io_inen[6]
port 214 nsew
flabel metal2 707800 355066 708076 355142 0 FreeSans 480 0 0 0 mprj_io_pd_select[6]
port 328 nsew
flabel metal2 707800 354564 708076 354640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[12]
port 70 nsew
flabel metal2 707800 354422 708076 354498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[13]
port 71 nsew
flabel metal2 707800 354193 708076 354269 0 FreeSans 480 0 0 0 mprj_io_pu_select[6]
port 366 nsew
flabel metal2 707800 353672 708076 353748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[6]
port 404 nsew
flabel metal2 707800 539172 708076 539248 0 FreeSans 480 0 0 0 mprj_io_in[7]
port 177 nsew
flabel metal2 707800 539026 708076 539102 0 FreeSans 480 0 0 0 mprj_io_outen[7]
port 291 nsew
flabel metal2 707800 538880 708076 538956 0 FreeSans 480 0 0 0 mprj_io_out[7]
port 253 nsew
flabel metal2 707800 538734 708076 538810 0 FreeSans 480 0 0 0 mprj_io_slew_select[7]
port 443 nsew
flabel metal2 707800 527277 708076 527353 0 FreeSans 480 0 0 0 mprj_io_inen[7]
port 215 nsew
flabel metal2 707800 527066 708076 527142 0 FreeSans 480 0 0 0 mprj_io_pd_select[7]
port 329 nsew
flabel metal2 707800 526564 708076 526640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[14]
port 72 nsew
flabel metal2 707800 526422 708076 526498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[15]
port 73 nsew
flabel metal2 707800 526193 708076 526269 0 FreeSans 480 0 0 0 mprj_io_pu_select[7]
port 367 nsew
flabel metal2 707800 525672 708076 525748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[7]
port 405 nsew
flabel metal2 707800 582172 708076 582248 0 FreeSans 480 0 0 0 mprj_io_in[8]
port 178 nsew
flabel metal2 707800 582026 708076 582102 0 FreeSans 480 0 0 0 mprj_io_outen[8]
port 292 nsew
flabel metal2 707800 581880 708076 581956 0 FreeSans 480 0 0 0 mprj_io_out[8]
port 254 nsew
flabel metal2 707800 581734 708076 581810 0 FreeSans 480 0 0 0 mprj_io_slew_select[8]
port 444 nsew
flabel metal2 707800 570277 708076 570353 0 FreeSans 480 0 0 0 mprj_io_inen[8]
port 216 nsew
flabel metal2 707800 570066 708076 570142 0 FreeSans 480 0 0 0 mprj_io_pd_select[8]
port 330 nsew
flabel metal2 707800 569564 708076 569640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[16]
port 74 nsew
flabel metal2 707800 569422 708076 569498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[17]
port 75 nsew
flabel metal2 707800 569193 708076 569269 0 FreeSans 480 0 0 0 mprj_io_pu_select[8]
port 368 nsew
flabel metal2 707800 568672 708076 568748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[8]
port 406 nsew
flabel metal2 707800 625172 708076 625248 0 FreeSans 480 0 0 0 mprj_io_in[9]
port 179 nsew
flabel metal2 707800 625026 708076 625102 0 FreeSans 480 0 0 0 mprj_io_outen[9]
port 293 nsew
flabel metal2 707800 624880 708076 624956 0 FreeSans 480 0 0 0 mprj_io_out[9]
port 255 nsew
flabel metal2 707800 624734 708076 624810 0 FreeSans 480 0 0 0 mprj_io_slew_select[9]
port 445 nsew
flabel metal2 707800 613277 708076 613353 0 FreeSans 480 0 0 0 mprj_io_inen[9]
port 217 nsew
flabel metal2 707800 613066 708076 613142 0 FreeSans 480 0 0 0 mprj_io_pd_select[9]
port 331 nsew
flabel metal2 707800 612564 708076 612640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[18]
port 76 nsew
flabel metal2 707800 612422 708076 612498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[19]
port 77 nsew
flabel metal2 707800 612193 708076 612269 0 FreeSans 480 0 0 0 mprj_io_pu_select[9]
port 369 nsew
flabel metal2 707800 611672 708076 611748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[9]
port 407 nsew
flabel metal2 707800 668172 708076 668248 0 FreeSans 480 0 0 0 mprj_io_in[10]
port 143 nsew
flabel metal2 707800 668026 708076 668102 0 FreeSans 480 0 0 0 mprj_io_outen[10]
port 257 nsew
flabel metal2 707800 667880 708076 667956 0 FreeSans 480 0 0 0 mprj_io_out[10]
port 219 nsew
flabel metal2 707800 667734 708076 667810 0 FreeSans 480 0 0 0 mprj_io_slew_select[10]
port 409 nsew
flabel metal2 707800 656277 708076 656353 0 FreeSans 480 0 0 0 mprj_io_inen[10]
port 181 nsew
flabel metal2 707800 656066 708076 656142 0 FreeSans 480 0 0 0 mprj_io_pd_select[10]
port 295 nsew
flabel metal2 707800 655564 708076 655640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[20]
port 79 nsew
flabel metal2 707800 655422 708076 655498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[21]
port 80 nsew
flabel metal2 707800 655193 708076 655269 0 FreeSans 480 0 0 0 mprj_io_pu_select[10]
port 333 nsew
flabel metal2 707800 654672 708076 654748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[10]
port 371 nsew
flabel metal2 707800 711172 708076 711248 0 FreeSans 480 0 0 0 mprj_io_in[11]
port 144 nsew
flabel metal2 707800 711026 708076 711102 0 FreeSans 480 0 0 0 mprj_io_outen[11]
port 258 nsew
flabel metal2 707800 710880 708076 710956 0 FreeSans 480 0 0 0 mprj_io_out[11]
port 220 nsew
flabel metal2 707800 710734 708076 710810 0 FreeSans 480 0 0 0 mprj_io_slew_select[11]
port 410 nsew
flabel metal2 707800 699277 708076 699353 0 FreeSans 480 0 0 0 mprj_io_inen[11]
port 182 nsew
flabel metal2 707800 699066 708076 699142 0 FreeSans 480 0 0 0 mprj_io_pd_select[11]
port 296 nsew
flabel metal2 707800 698564 708076 698640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[22]
port 81 nsew
flabel metal2 707800 698422 708076 698498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[23]
port 82 nsew
flabel metal2 707800 698193 708076 698269 0 FreeSans 480 0 0 0 mprj_io_pu_select[11]
port 334 nsew
flabel metal2 707800 697672 708076 697748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[11]
port 372 nsew
flabel metal2 707800 840172 708076 840248 0 FreeSans 480 0 0 0 mprj_io_in[12]
port 145 nsew
flabel metal2 707800 840026 708076 840102 0 FreeSans 480 0 0 0 mprj_io_outen[12]
port 259 nsew
flabel metal2 707800 839880 708076 839956 0 FreeSans 480 0 0 0 mprj_io_out[12]
port 221 nsew
flabel metal2 707800 839734 708076 839810 0 FreeSans 480 0 0 0 mprj_io_slew_select[12]
port 411 nsew
flabel metal2 707800 828277 708076 828353 0 FreeSans 480 0 0 0 mprj_io_inen[12]
port 183 nsew
flabel metal2 707800 828066 708076 828142 0 FreeSans 480 0 0 0 mprj_io_pd_select[12]
port 297 nsew
flabel metal2 707800 827564 708076 827640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[24]
port 83 nsew
flabel metal2 707800 827422 708076 827498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[25]
port 84 nsew
flabel metal2 707800 827193 708076 827269 0 FreeSans 480 0 0 0 mprj_io_pu_select[12]
port 335 nsew
flabel metal2 707800 826672 708076 826748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[12]
port 373 nsew
flabel metal2 707800 740672 708076 740748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[13]
port 374 nsew
flabel metal2 707800 741193 708076 741269 0 FreeSans 480 0 0 0 mprj_io_pu_select[13]
port 336 nsew
flabel metal2 707800 741422 708076 741498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[26]
port 85 nsew
flabel metal2 707800 741564 708076 741640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[27]
port 86 nsew
flabel metal2 707800 742066 708076 742142 0 FreeSans 480 0 0 0 mprj_io_pd_select[13]
port 298 nsew
flabel metal2 707800 742277 708076 742353 0 FreeSans 480 0 0 0 mprj_io_inen[13]
port 184 nsew
flabel metal2 707800 753734 708076 753810 0 FreeSans 480 0 0 0 mprj_io_slew_select[13]
port 412 nsew
flabel metal2 707800 753880 708076 753956 0 FreeSans 480 0 0 0 mprj_io_out[13]
port 222 nsew
flabel metal2 707800 754026 708076 754102 0 FreeSans 480 0 0 0 mprj_io_outen[13]
port 260 nsew
flabel metal2 707800 754172 708076 754248 0 FreeSans 480 0 0 0 mprj_io_in[13]
port 146 nsew
flabel metal2 707800 912672 708076 912748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[14]
port 375 nsew
flabel metal2 707800 913193 708076 913269 0 FreeSans 480 0 0 0 mprj_io_pu_select[14]
port 337 nsew
flabel metal2 707800 913422 708076 913498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[28]
port 87 nsew
flabel metal2 707800 913564 708076 913640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[29]
port 88 nsew
flabel metal2 707800 914066 708076 914142 0 FreeSans 480 0 0 0 mprj_io_pd_select[14]
port 299 nsew
flabel metal2 707800 914277 708076 914353 0 FreeSans 480 0 0 0 mprj_io_inen[14]
port 185 nsew
flabel metal2 707800 925734 708076 925810 0 FreeSans 480 0 0 0 mprj_io_slew_select[14]
port 413 nsew
flabel metal2 707800 925880 708076 925956 0 FreeSans 480 0 0 0 mprj_io_out[14]
port 223 nsew
flabel metal2 707800 926026 708076 926102 0 FreeSans 480 0 0 0 mprj_io_outen[14]
port 261 nsew
flabel metal2 707800 926172 708076 926248 0 FreeSans 480 0 0 0 mprj_io_in[14]
port 147 nsew
flabel metal2 670252 949800 670328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[15]
port 376 nsew
flabel metal2 669731 949800 669807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[15]
port 338 nsew
flabel metal2 669502 949800 669578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[30]
port 90 nsew
flabel metal2 669360 949800 669436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[31]
port 91 nsew
flabel metal2 668858 949800 668934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[15]
port 300 nsew
flabel metal2 668647 949800 668723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[15]
port 186 nsew
flabel metal2 657190 949800 657266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[15]
port 414 nsew
flabel metal2 657044 949800 657120 950076 0 FreeSans 480 270 0 0 mprj_io_out[15]
port 224 nsew
flabel metal2 656898 949800 656974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[15]
port 262 nsew
flabel metal2 656752 949800 656828 950076 0 FreeSans 480 270 0 0 mprj_io_in[15]
port 148 nsew
flabel metal2 560252 949800 560328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[16]
port 377 nsew
flabel metal2 559731 949800 559807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[16]
port 339 nsew
flabel metal2 559502 949800 559578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[32]
port 92 nsew
flabel metal2 559360 949800 559436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[33]
port 93 nsew
flabel metal2 558858 949800 558934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[16]
port 301 nsew
flabel metal2 558647 949800 558723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[16]
port 187 nsew
flabel metal2 547190 949800 547266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[16]
port 415 nsew
flabel metal2 547044 949800 547120 950076 0 FreeSans 480 270 0 0 mprj_io_out[16]
port 225 nsew
flabel metal2 546898 949800 546974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[16]
port 263 nsew
flabel metal2 546752 949800 546828 950076 0 FreeSans 480 270 0 0 mprj_io_in[16]
port 149 nsew
flabel metal2 505252 949800 505328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[17]
port 378 nsew
flabel metal2 504731 949800 504807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[17]
port 340 nsew
flabel metal2 504502 949800 504578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[34]
port 94 nsew
flabel metal2 504360 949800 504436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[35]
port 95 nsew
flabel metal2 503858 949800 503934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[17]
port 302 nsew
flabel metal2 503647 949800 503723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[17]
port 188 nsew
flabel metal2 492190 949800 492266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[17]
port 416 nsew
flabel metal2 492044 949800 492120 950076 0 FreeSans 480 270 0 0 mprj_io_out[17]
port 226 nsew
flabel metal2 491898 949800 491974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[17]
port 264 nsew
flabel metal2 491752 949800 491828 950076 0 FreeSans 480 270 0 0 mprj_io_in[17]
port 150 nsew
flabel metal2 450252 949800 450328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[18]
port 379 nsew
flabel metal2 449731 949800 449807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[18]
port 341 nsew
flabel metal2 449502 949800 449578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[36]
port 96 nsew
flabel metal2 449360 949800 449436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[37]
port 97 nsew
flabel metal2 448858 949800 448934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[18]
port 303 nsew
flabel metal2 448647 949800 448723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[18]
port 189 nsew
flabel metal2 437190 949800 437266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[18]
port 417 nsew
flabel metal2 437044 949800 437120 950076 0 FreeSans 480 270 0 0 mprj_io_out[18]
port 227 nsew
flabel metal2 436898 949800 436974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[18]
port 265 nsew
flabel metal2 436752 949800 436828 950076 0 FreeSans 480 270 0 0 mprj_io_in[18]
port 151 nsew
flabel metal2 340252 949800 340328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[19]
port 380 nsew
flabel metal2 339731 949800 339807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[19]
port 342 nsew
flabel metal2 339502 949800 339578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[38]
port 98 nsew
flabel metal2 339360 949800 339436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[39]
port 99 nsew
flabel metal2 338858 949800 338934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[19]
port 304 nsew
flabel metal2 338647 949800 338723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[19]
port 190 nsew
flabel metal2 327190 949800 327266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[19]
port 418 nsew
flabel metal2 327044 949800 327120 950076 0 FreeSans 480 270 0 0 mprj_io_out[19]
port 228 nsew
flabel metal2 326898 949800 326974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[19]
port 266 nsew
flabel metal2 326752 949800 326828 950076 0 FreeSans 480 270 0 0 mprj_io_in[19]
port 152 nsew
flabel metal2 285252 949800 285328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[20]
port 382 nsew
flabel metal2 284731 949800 284807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[20]
port 344 nsew
flabel metal2 284502 949800 284578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[40]
port 101 nsew
flabel metal2 284360 949800 284436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[41]
port 102 nsew
flabel metal2 283858 949800 283934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[20]
port 306 nsew
flabel metal2 283647 949800 283723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[20]
port 192 nsew
flabel metal2 272190 949800 272266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[20]
port 420 nsew
flabel metal2 272044 949800 272120 950076 0 FreeSans 480 270 0 0 mprj_io_out[20]
port 230 nsew
flabel metal2 271898 949800 271974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[20]
port 268 nsew
flabel metal2 271752 949800 271828 950076 0 FreeSans 480 270 0 0 mprj_io_in[20]
port 154 nsew
flabel metal2 230252 949800 230328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[21]
port 383 nsew
flabel metal2 229731 949800 229807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[21]
port 345 nsew
flabel metal2 229502 949800 229578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[42]
port 103 nsew
flabel metal2 229360 949800 229436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[43]
port 104 nsew
flabel metal2 228858 949800 228934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[21]
port 307 nsew
flabel metal2 228647 949800 228723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[21]
port 193 nsew
flabel metal2 217190 949800 217266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[21]
port 421 nsew
flabel metal2 217044 949800 217120 950076 0 FreeSans 480 270 0 0 mprj_io_out[21]
port 231 nsew
flabel metal2 216898 949800 216974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[21]
port 269 nsew
flabel metal2 216752 949800 216828 950076 0 FreeSans 480 270 0 0 mprj_io_in[21]
port 155 nsew
flabel metal2 175252 949800 175328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[22]
port 384 nsew
flabel metal2 174731 949800 174807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[22]
port 346 nsew
flabel metal2 174502 949800 174578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[44]
port 105 nsew
flabel metal2 174360 949800 174436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[45]
port 106 nsew
flabel metal2 173858 949800 173934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[22]
port 308 nsew
flabel metal2 173647 949800 173723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[22]
port 194 nsew
flabel metal2 162190 949800 162266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[22]
port 422 nsew
flabel metal2 162044 949800 162120 950076 0 FreeSans 480 270 0 0 mprj_io_out[22]
port 232 nsew
flabel metal2 161898 949800 161974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[22]
port 270 nsew
flabel metal2 161752 949800 161828 950076 0 FreeSans 480 270 0 0 mprj_io_in[22]
port 156 nsew
flabel metal2 120252 949800 120328 950076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[23]
port 385 nsew
flabel metal2 119731 949800 119807 950076 0 FreeSans 480 270 0 0 mprj_io_pu_select[23]
port 347 nsew
flabel metal2 119502 949800 119578 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[46]
port 107 nsew
flabel metal2 119360 949800 119436 950076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[47]
port 108 nsew
flabel metal2 118858 949800 118934 950076 0 FreeSans 480 270 0 0 mprj_io_pd_select[23]
port 309 nsew
flabel metal2 118647 949800 118723 950076 0 FreeSans 480 270 0 0 mprj_io_inen[23]
port 195 nsew
flabel metal2 107190 949800 107266 950076 0 FreeSans 480 270 0 0 mprj_io_slew_select[23]
port 423 nsew
flabel metal2 107044 949800 107120 950076 0 FreeSans 480 270 0 0 mprj_io_out[23]
port 233 nsew
flabel metal2 106898 949800 106974 950076 0 FreeSans 480 270 0 0 mprj_io_outen[23]
port 271 nsew
flabel metal2 106752 949800 106828 950076 0 FreeSans 480 270 0 0 mprj_io_in[23]
port 157 nsew
flabel metal2 69924 173752 70200 173828 0 FreeSans 480 180 0 0 mprj_io_in[37]
port 172 nsew
flabel metal2 69924 173898 70200 173974 0 FreeSans 480 180 0 0 mprj_io_outen[37]
port 286 nsew
flabel metal2 69924 174044 70200 174120 0 FreeSans 480 180 0 0 mprj_io_out[37]
port 248 nsew
flabel metal2 69924 174190 70200 174266 0 FreeSans 480 180 0 0 mprj_io_slew_select[37]
port 438 nsew
flabel metal2 69924 185647 70200 185723 0 FreeSans 480 180 0 0 mprj_io_inen[37]
port 210 nsew
flabel metal2 69924 185858 70200 185934 0 FreeSans 480 180 0 0 mprj_io_pd_select[37]
port 324 nsew
flabel metal2 69924 186360 70200 186436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[75]
port 138 nsew
flabel metal2 69924 186502 70200 186578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[74]
port 137 nsew
flabel metal2 69924 186731 70200 186807 0 FreeSans 480 180 0 0 mprj_io_pu_select[37]
port 362 nsew
flabel metal2 69924 187252 70200 187328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[37]
port 400 nsew
flabel metal2 69924 214752 70200 214828 0 FreeSans 480 180 0 0 mprj_io_in[36]
port 171 nsew
flabel metal2 69924 214898 70200 214974 0 FreeSans 480 180 0 0 mprj_io_outen[36]
port 285 nsew
flabel metal2 69924 215044 70200 215120 0 FreeSans 480 180 0 0 mprj_io_out[36]
port 247 nsew
flabel metal2 69924 215190 70200 215266 0 FreeSans 480 180 0 0 mprj_io_slew_select[36]
port 437 nsew
flabel metal2 69924 226647 70200 226723 0 FreeSans 480 180 0 0 mprj_io_inen[36]
port 209 nsew
flabel metal2 69924 226858 70200 226934 0 FreeSans 480 180 0 0 mprj_io_pd_select[36]
port 323 nsew
flabel metal2 69924 227360 70200 227436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[73]
port 136 nsew
flabel metal2 69924 227502 70200 227578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[72]
port 135 nsew
flabel metal2 69924 227731 70200 227807 0 FreeSans 480 180 0 0 mprj_io_pu_select[36]
port 361 nsew
flabel metal2 69924 228252 70200 228328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[36]
port 399 nsew
flabel metal2 69924 255752 70200 255828 0 FreeSans 480 180 0 0 mprj_io_in[35]
port 170 nsew
flabel metal2 69924 255898 70200 255974 0 FreeSans 480 180 0 0 mprj_io_outen[35]
port 284 nsew
flabel metal2 69924 256044 70200 256120 0 FreeSans 480 180 0 0 mprj_io_out[35]
port 246 nsew
flabel metal2 69924 256190 70200 256266 0 FreeSans 480 180 0 0 mprj_io_slew_select[35]
port 436 nsew
flabel metal2 69924 267647 70200 267723 0 FreeSans 480 180 0 0 mprj_io_inen[35]
port 208 nsew
flabel metal2 69924 267858 70200 267934 0 FreeSans 480 180 0 0 mprj_io_pd_select[35]
port 322 nsew
flabel metal2 69924 268360 70200 268436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[71]
port 134 nsew
flabel metal2 69924 268502 70200 268578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[70]
port 133 nsew
flabel metal2 69924 268731 70200 268807 0 FreeSans 480 180 0 0 mprj_io_pu_select[35]
port 360 nsew
flabel metal2 69924 269252 70200 269328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[35]
port 398 nsew
flabel metal2 69924 296752 70200 296828 0 FreeSans 480 180 0 0 mprj_io_in[34]
port 169 nsew
flabel metal2 69924 296898 70200 296974 0 FreeSans 480 180 0 0 mprj_io_outen[34]
port 283 nsew
flabel metal2 69924 297044 70200 297120 0 FreeSans 480 180 0 0 mprj_io_out[34]
port 245 nsew
flabel metal2 69924 297190 70200 297266 0 FreeSans 480 180 0 0 mprj_io_slew_select[34]
port 435 nsew
flabel metal2 69924 308647 70200 308723 0 FreeSans 480 180 0 0 mprj_io_inen[34]
port 207 nsew
flabel metal2 69924 308858 70200 308934 0 FreeSans 480 180 0 0 mprj_io_pd_select[34]
port 321 nsew
flabel metal2 69924 309360 70200 309436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[69]
port 131 nsew
flabel metal2 69924 309502 70200 309578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[68]
port 130 nsew
flabel metal2 69924 309731 70200 309807 0 FreeSans 480 180 0 0 mprj_io_pu_select[34]
port 359 nsew
flabel metal2 69924 310252 70200 310328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[34]
port 397 nsew
flabel metal2 69924 337752 70200 337828 0 FreeSans 480 180 0 0 mprj_io_in[33]
port 168 nsew
flabel metal2 69924 337898 70200 337974 0 FreeSans 480 180 0 0 mprj_io_outen[33]
port 282 nsew
flabel metal2 69924 338044 70200 338120 0 FreeSans 480 180 0 0 mprj_io_out[33]
port 244 nsew
flabel metal2 69924 338190 70200 338266 0 FreeSans 480 180 0 0 mprj_io_slew_select[33]
port 434 nsew
flabel metal2 69924 349647 70200 349723 0 FreeSans 480 180 0 0 mprj_io_inen[33]
port 206 nsew
flabel metal2 69924 349858 70200 349934 0 FreeSans 480 180 0 0 mprj_io_pd_select[33]
port 320 nsew
flabel metal2 69924 350360 70200 350436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[67]
port 129 nsew
flabel metal2 69924 350502 70200 350578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[66]
port 128 nsew
flabel metal2 69924 350731 70200 350807 0 FreeSans 480 180 0 0 mprj_io_pu_select[33]
port 358 nsew
flabel metal2 69924 351252 70200 351328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[33]
port 396 nsew
flabel metal2 69924 378752 70200 378828 0 FreeSans 480 180 0 0 mprj_io_in[32]
port 167 nsew
flabel metal2 69924 378898 70200 378974 0 FreeSans 480 180 0 0 mprj_io_outen[32]
port 281 nsew
flabel metal2 69924 379044 70200 379120 0 FreeSans 480 180 0 0 mprj_io_out[32]
port 243 nsew
flabel metal2 69924 379190 70200 379266 0 FreeSans 480 180 0 0 mprj_io_slew_select[32]
port 433 nsew
flabel metal2 69924 390647 70200 390723 0 FreeSans 480 180 0 0 mprj_io_inen[32]
port 205 nsew
flabel metal2 69924 390858 70200 390934 0 FreeSans 480 180 0 0 mprj_io_pd_select[32]
port 319 nsew
flabel metal2 69924 391360 70200 391436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[65]
port 127 nsew
flabel metal2 69924 391502 70200 391578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[64]
port 126 nsew
flabel metal2 69924 391731 70200 391807 0 FreeSans 480 180 0 0 mprj_io_pu_select[32]
port 357 nsew
flabel metal2 69924 392252 70200 392328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[32]
port 395 nsew
flabel metal2 69924 501752 70200 501828 0 FreeSans 480 180 0 0 mprj_io_in[31]
port 166 nsew
flabel metal2 69924 501898 70200 501974 0 FreeSans 480 180 0 0 mprj_io_outen[31]
port 280 nsew
flabel metal2 69924 502044 70200 502120 0 FreeSans 480 180 0 0 mprj_io_out[31]
port 242 nsew
flabel metal2 69924 502190 70200 502266 0 FreeSans 480 180 0 0 mprj_io_slew_select[31]
port 432 nsew
flabel metal2 69924 513647 70200 513723 0 FreeSans 480 180 0 0 mprj_io_inen[31]
port 204 nsew
flabel metal2 69924 513858 70200 513934 0 FreeSans 480 180 0 0 mprj_io_pd_select[31]
port 318 nsew
flabel metal2 69924 514360 70200 514436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[63]
port 125 nsew
flabel metal2 69924 514502 70200 514578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[62]
port 124 nsew
flabel metal2 69924 514731 70200 514807 0 FreeSans 480 180 0 0 mprj_io_pu_select[31]
port 356 nsew
flabel metal2 69924 515252 70200 515328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[31]
port 394 nsew
flabel metal2 69924 542752 70200 542828 0 FreeSans 480 180 0 0 mprj_io_in[30]
port 165 nsew
flabel metal2 69924 542898 70200 542974 0 FreeSans 480 180 0 0 mprj_io_outen[30]
port 279 nsew
flabel metal2 69924 543044 70200 543120 0 FreeSans 480 180 0 0 mprj_io_out[30]
port 241 nsew
flabel metal2 69924 543190 70200 543266 0 FreeSans 480 180 0 0 mprj_io_slew_select[30]
port 431 nsew
flabel metal2 69924 554647 70200 554723 0 FreeSans 480 180 0 0 mprj_io_inen[30]
port 203 nsew
flabel metal2 69924 554858 70200 554934 0 FreeSans 480 180 0 0 mprj_io_pd_select[30]
port 317 nsew
flabel metal2 69924 555360 70200 555436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[61]
port 123 nsew
flabel metal2 69924 555502 70200 555578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[63]
port 125 nsew
flabel metal2 69924 555731 70200 555807 0 FreeSans 480 180 0 0 mprj_io_pu_select[30]
port 355 nsew
flabel metal2 69924 556252 70200 556328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[30]
port 393 nsew
flabel metal2 69924 583752 70200 583828 0 FreeSans 480 180 0 0 mprj_io_in[29]
port 163 nsew
flabel metal2 69924 583898 70200 583974 0 FreeSans 480 180 0 0 mprj_io_outen[29]
port 277 nsew
flabel metal2 69924 584044 70200 584120 0 FreeSans 480 180 0 0 mprj_io_out[29]
port 239 nsew
flabel metal2 69924 584190 70200 584266 0 FreeSans 480 180 0 0 mprj_io_slew_select[29]
port 429 nsew
flabel metal2 69924 595647 70200 595723 0 FreeSans 480 180 0 0 mprj_io_inen[29]
port 201 nsew
flabel metal2 69924 595858 70200 595934 0 FreeSans 480 180 0 0 mprj_io_pd_select[29]
port 315 nsew
flabel metal2 69924 596360 70200 596436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[59]
port 121 nsew
flabel metal2 69924 596502 70200 596578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[58]
port 120 nsew
flabel metal2 69924 596731 70200 596807 0 FreeSans 480 180 0 0 mprj_io_pu_select[29]
port 353 nsew
flabel metal2 69924 597252 70200 597328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[29]
port 391 nsew
flabel metal2 69924 624752 70200 624828 0 FreeSans 480 180 0 0 mprj_io_in[28]
port 162 nsew
flabel metal2 69924 624898 70200 624974 0 FreeSans 480 180 0 0 mprj_io_outen[28]
port 276 nsew
flabel metal2 69924 625044 70200 625120 0 FreeSans 480 180 0 0 mprj_io_out[28]
port 238 nsew
flabel metal2 69924 625190 70200 625266 0 FreeSans 480 180 0 0 mprj_io_slew_select[28]
port 428 nsew
flabel metal2 69924 636647 70200 636723 0 FreeSans 480 180 0 0 mprj_io_inen[28]
port 200 nsew
flabel metal2 69924 636858 70200 636934 0 FreeSans 480 180 0 0 mprj_io_pd_select[28]
port 314 nsew
flabel metal2 69924 637360 70200 637436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[57]
port 119 nsew
flabel metal2 69924 637502 70200 637578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[56]
port 118 nsew
flabel metal2 69924 637731 70200 637807 0 FreeSans 480 180 0 0 mprj_io_pu_select[28]
port 352 nsew
flabel metal2 69924 638252 70200 638328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[28]
port 390 nsew
flabel metal2 69924 665752 70200 665828 0 FreeSans 480 180 0 0 mprj_io_in[27]
port 161 nsew
flabel metal2 69924 665898 70200 665974 0 FreeSans 480 180 0 0 mprj_io_outen[27]
port 275 nsew
flabel metal2 69924 666044 70200 666120 0 FreeSans 480 180 0 0 mprj_io_out[27]
port 237 nsew
flabel metal2 69924 666190 70200 666266 0 FreeSans 480 180 0 0 mprj_io_slew_select[27]
port 427 nsew
flabel metal2 69924 677647 70200 677723 0 FreeSans 480 180 0 0 mprj_io_inen[27]
port 199 nsew
flabel metal2 69924 677858 70200 677934 0 FreeSans 480 180 0 0 mprj_io_pd_select[27]
port 313 nsew
flabel metal2 69924 678360 70200 678436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[55]
port 117 nsew
flabel metal2 69924 678502 70200 678578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[54]
port 116 nsew
flabel metal2 69924 678731 70200 678807 0 FreeSans 480 180 0 0 mprj_io_pu_select[27]
port 351 nsew
flabel metal2 69924 679252 70200 679328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[27]
port 389 nsew
flabel metal2 69924 706752 70200 706828 0 FreeSans 480 180 0 0 mprj_io_in[26]
port 160 nsew
flabel metal2 69924 706898 70200 706974 0 FreeSans 480 180 0 0 mprj_io_outen[26]
port 274 nsew
flabel metal2 69924 707044 70200 707120 0 FreeSans 480 180 0 0 mprj_io_out[26]
port 236 nsew
flabel metal2 69924 707190 70200 707266 0 FreeSans 480 180 0 0 mprj_io_slew_select[26]
port 426 nsew
flabel metal2 69924 718647 70200 718723 0 FreeSans 480 180 0 0 mprj_io_inen[26]
port 198 nsew
flabel metal2 69924 718858 70200 718934 0 FreeSans 480 180 0 0 mprj_io_pd_select[26]
port 312 nsew
flabel metal2 69924 719360 70200 719436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[53]
port 115 nsew
flabel metal2 69924 719502 70200 719578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[52]
port 114 nsew
flabel metal2 69924 719731 70200 719807 0 FreeSans 480 180 0 0 mprj_io_pu_select[26]
port 350 nsew
flabel metal2 69924 720252 70200 720328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[26]
port 388 nsew
flabel metal2 69924 747752 70200 747828 0 FreeSans 480 180 0 0 mprj_io_in[25]
port 159 nsew
flabel metal2 69924 747898 70200 747974 0 FreeSans 480 180 0 0 mprj_io_outen[25]
port 273 nsew
flabel metal2 69924 748044 70200 748120 0 FreeSans 480 180 0 0 mprj_io_out[25]
port 235 nsew
flabel metal2 69924 748190 70200 748266 0 FreeSans 480 180 0 0 mprj_io_slew_select[25]
port 425 nsew
flabel metal2 69924 759647 70200 759723 0 FreeSans 480 180 0 0 mprj_io_inen[25]
port 197 nsew
flabel metal2 69924 759858 70200 759934 0 FreeSans 480 180 0 0 mprj_io_pd_select[25]
port 311 nsew
flabel metal2 69924 760360 70200 760436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[51]
port 112 nsew
flabel metal2 69924 760502 70200 760578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[525]
port 113 nsew
flabel metal2 69924 760731 70200 760807 0 FreeSans 480 180 0 0 mprj_io_pu_select[25]
port 349 nsew
flabel metal2 69924 761252 70200 761328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[25]
port 387 nsew
flabel metal2 69924 911752 70200 911828 0 FreeSans 480 180 0 0 mprj_io_in[24]
port 158 nsew
flabel metal2 69924 911898 70200 911974 0 FreeSans 480 180 0 0 mprj_io_outen[24]
port 272 nsew
flabel metal2 69924 912044 70200 912120 0 FreeSans 480 180 0 0 mprj_io_out[24]
port 234 nsew
flabel metal2 69924 912190 70200 912266 0 FreeSans 480 180 0 0 mprj_io_slew_select[24]
port 424 nsew
flabel metal2 69924 923647 70200 923723 0 FreeSans 480 180 0 0 mprj_io_inen[24]
port 196 nsew
flabel metal2 69924 923858 70200 923934 0 FreeSans 480 180 0 0 mprj_io_pd_select[24]
port 310 nsew
flabel metal2 69924 924360 70200 924436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[49]
port 110 nsew
flabel metal2 69924 924502 70200 924578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[48]
port 109 nsew
flabel metal2 69924 924731 70200 924807 0 FreeSans 480 180 0 0 mprj_io_pu_select[24]
port 348 nsew
flabel metal2 69924 925252 70200 925328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[24]
port 386 nsew
<< end >>
