VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_id_textblock
  CLASS BLOCK ;
  FOREIGN user_id_textblock ;
  ORIGIN 0.000 0.000 ;
  SIZE 126.650 BY 30.225 ;
  OBS
      LAYER Metal5 ;
        RECT 3.650 9.980 6.890 11.060 ;
        RECT 3.650 4.580 4.730 9.980 ;
        RECT 5.810 4.580 6.890 9.980 ;
        RECT 3.650 3.500 6.890 4.580 ;
        RECT 19.275 9.980 22.515 11.060 ;
        RECT 19.275 4.580 20.355 9.980 ;
        RECT 21.435 4.580 22.515 9.980 ;
        RECT 19.275 3.500 22.515 4.580 ;
        RECT 34.900 9.980 38.140 11.060 ;
        RECT 34.900 4.580 35.980 9.980 ;
        RECT 37.060 4.580 38.140 9.980 ;
        RECT 34.900 3.500 38.140 4.580 ;
        RECT 50.525 9.980 53.765 11.060 ;
        RECT 50.525 4.580 51.605 9.980 ;
        RECT 52.685 4.580 53.765 9.980 ;
        RECT 50.525 3.500 53.765 4.580 ;
        RECT 66.150 9.980 69.390 11.060 ;
        RECT 66.150 4.580 67.230 9.980 ;
        RECT 68.310 4.580 69.390 9.980 ;
        RECT 66.150 3.500 69.390 4.580 ;
        RECT 81.775 9.980 85.015 11.060 ;
        RECT 81.775 4.580 82.855 9.980 ;
        RECT 83.935 4.580 85.015 9.980 ;
        RECT 81.775 3.500 85.015 4.580 ;
        RECT 97.400 9.980 100.640 11.060 ;
        RECT 97.400 4.580 98.480 9.980 ;
        RECT 99.560 4.580 100.640 9.980 ;
        RECT 97.400 3.500 100.640 4.580 ;
        RECT 113.325 9.980 116.565 11.060 ;
        RECT 113.325 4.580 114.405 9.980 ;
        RECT 115.485 4.580 116.565 9.980 ;
        RECT 113.325 3.500 116.565 4.580 ;
  END
END user_id_textblock
END LIBRARY

