magic
tech gf180mcuC
magscale 1 5
timestamp 1655473080
<< obsm1 >>
rect 336 211 17416 6302
<< metal2 >>
rect 1260 6600 1316 7000
rect 3836 6600 3892 7000
rect 6412 6600 6468 7000
rect 8988 6600 9044 7000
rect 11564 6600 11620 7000
rect 14140 6600 14196 7000
rect 16716 6600 16772 7000
<< obsm2 >>
rect 490 6570 1230 6600
rect 1346 6570 3806 6600
rect 3922 6570 6382 6600
rect 6498 6570 8958 6600
rect 9074 6570 11534 6600
rect 11650 6570 14110 6600
rect 14226 6570 16686 6600
rect 16802 6570 17374 6600
rect 490 205 17374 6570
<< metal3 >>
rect 17600 6524 18000 6580
rect 17600 5628 18000 5684
rect 17600 4788 18000 4844
rect 17600 3892 18000 3948
rect 17600 2996 18000 3052
rect 17600 2156 18000 2212
rect 17600 1260 18000 1316
rect 17600 420 18000 476
<< obsm3 >>
rect 485 6494 17570 6566
rect 485 5714 17600 6494
rect 485 5598 17570 5714
rect 485 4874 17600 5598
rect 485 4758 17570 4874
rect 485 3978 17600 4758
rect 485 3862 17570 3978
rect 485 3082 17600 3862
rect 485 2966 17570 3082
rect 485 2242 17600 2966
rect 485 2126 17570 2242
rect 485 1346 17600 2126
rect 485 1230 17570 1346
rect 485 506 17600 1230
rect 485 390 17570 506
rect 485 266 17600 390
<< metal4 >>
rect 2394 362 2554 6302
rect 4532 362 4692 6302
rect 6670 362 6830 6302
rect 8808 362 8968 6302
rect 10946 362 11106 6302
rect 13084 362 13244 6302
rect 15222 362 15382 6302
<< obsm4 >>
rect 1666 6332 17206 6571
rect 1666 485 2364 6332
rect 2584 485 4502 6332
rect 4722 485 6640 6332
rect 6860 485 8778 6332
rect 8998 485 10916 6332
rect 11136 485 13054 6332
rect 13274 485 15192 6332
rect 15412 485 17206 6332
<< metal5 >>
rect 306 5751 17446 5911
rect 306 4974 17446 5134
rect 306 4197 17446 4357
rect 306 3420 17446 3580
rect 306 2643 17446 2803
rect 306 1866 17446 2026
rect 306 1089 17446 1249
<< obsm5 >>
rect 3282 4407 17214 4882
rect 3282 3630 17214 4147
rect 3282 2853 17214 3370
rect 3282 2076 17214 2593
rect 3282 1299 17214 1816
rect 3282 518 17214 1039
<< labels >>
rlabel metal4 s 2394 362 2554 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 6670 362 6830 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 10946 362 11106 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 15222 362 15382 6302 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 306 1089 17446 1249 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 306 2643 17446 2803 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 306 4197 17446 4357 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 306 5751 17446 5911 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 4532 362 4692 6302 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 8808 362 8968 6302 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 13084 362 13244 6302 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 306 1866 17446 2026 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 306 3420 17446 3580 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 306 4974 17446 5134 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 6412 6600 6468 7000 6 core_clk
port 3 nsew signal output
rlabel metal2 s 3836 6600 3892 7000 6 ext_clk
port 4 nsew signal input
rlabel metal3 s 17600 420 18000 476 6 ext_clk_sel
port 5 nsew signal input
rlabel metal3 s 17600 6524 18000 6580 6 ext_reset
port 6 nsew signal input
rlabel metal2 s 14140 6600 14196 7000 6 pll_clk
port 7 nsew signal input
rlabel metal2 s 16716 6600 16772 7000 6 pll_clk90
port 8 nsew signal input
rlabel metal2 s 1260 6600 1316 7000 6 resetb
port 9 nsew signal input
rlabel metal2 s 11564 6600 11620 7000 6 resetb_sync
port 10 nsew signal output
rlabel metal3 s 17600 3892 18000 3948 6 sel2[0]
port 11 nsew signal input
rlabel metal3 s 17600 4788 18000 4844 6 sel2[1]
port 12 nsew signal input
rlabel metal3 s 17600 5628 18000 5684 6 sel2[2]
port 13 nsew signal input
rlabel metal3 s 17600 1260 18000 1316 6 sel[0]
port 14 nsew signal input
rlabel metal3 s 17600 2156 18000 2212 6 sel[1]
port 15 nsew signal input
rlabel metal3 s 17600 2996 18000 3052 6 sel[2]
port 16 nsew signal input
rlabel metal2 s 8988 6600 9044 7000 6 user_clk
port 17 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 18000 7000
string GDS_END 695170
string GDS_FILE ../gds/caravel_clocking.gds.gz
string GDS_START 171610
string LEFclass BLOCK
string LEFview TRUE
<< end >>
