VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_id_programming
  CLASS BLOCK ;
  FOREIGN user_id_programming ;
  ORIGIN 0.430 2.100 ;
  SIZE 109.500 BY 10.760 ;
  PIN mask_rev[0]
    PORT
      LAYER Metal1 ;
        RECT 9.060 6.190 9.435 7.310 ;
      LAYER Via1 ;
        RECT 9.090 6.290 9.390 6.590 ;
      LAYER Metal2 ;
        RECT 5.290 6.280 9.500 6.600 ;
        RECT 5.290 2.440 5.570 6.280 ;
        RECT 0.140 2.160 5.570 2.440 ;
        RECT 0.140 -2.100 0.420 2.160 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    PORT
      LAYER Metal1 ;
        RECT 40.420 6.190 40.795 7.310 ;
      LAYER Via1 ;
        RECT 40.450 6.290 40.750 6.590 ;
      LAYER Metal2 ;
        RECT 34.860 6.280 40.860 6.600 ;
        RECT 34.860 -2.100 35.140 6.280 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    PORT
      LAYER Metal1 ;
        RECT 40.420 0.530 40.795 1.650 ;
      LAYER Via1 ;
        RECT 40.450 1.250 40.750 1.550 ;
      LAYER Metal2 ;
        RECT 38.780 1.240 40.860 1.560 ;
        RECT 38.780 -2.100 39.060 1.240 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    PORT
      LAYER Metal1 ;
        RECT 46.020 6.190 46.395 7.310 ;
      LAYER Via1 ;
        RECT 46.050 6.290 46.350 6.590 ;
      LAYER Metal2 ;
        RECT 42.140 6.280 46.470 6.600 ;
        RECT 42.140 -2.100 42.420 6.280 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    PORT
      LAYER Metal1 ;
        RECT 46.020 0.530 46.395 1.650 ;
      LAYER Via1 ;
        RECT 46.050 1.250 46.350 1.550 ;
      LAYER Metal2 ;
        RECT 44.365 1.240 46.500 1.560 ;
        RECT 45.500 -2.100 45.780 1.240 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    PORT
      LAYER Metal1 ;
        RECT 52.740 6.190 53.115 7.310 ;
      LAYER Via1 ;
        RECT 52.770 6.290 53.070 6.590 ;
      LAYER Metal2 ;
        RECT 48.860 6.280 53.170 6.600 ;
        RECT 48.860 -2.100 49.140 6.280 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    PORT
      LAYER Metal1 ;
        RECT 52.740 0.530 53.115 1.650 ;
      LAYER Via1 ;
        RECT 52.770 1.250 53.070 1.550 ;
      LAYER Metal2 ;
        RECT 51.085 1.240 53.175 1.560 ;
        RECT 52.220 -2.100 52.500 1.240 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    PORT
      LAYER Metal1 ;
        RECT 58.340 6.190 58.715 7.310 ;
      LAYER Via1 ;
        RECT 58.370 6.290 58.670 6.590 ;
      LAYER Metal2 ;
        RECT 56.140 6.280 58.770 6.600 ;
        RECT 56.140 3.030 56.420 6.280 ;
        RECT 56.115 2.725 56.420 3.030 ;
        RECT 56.115 0.395 56.395 2.725 ;
        RECT 56.115 0.115 56.420 0.395 ;
        RECT 56.140 -2.100 56.420 0.115 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    PORT
      LAYER Metal1 ;
        RECT 58.340 0.530 58.715 1.650 ;
      LAYER Via1 ;
        RECT 58.370 1.250 58.670 1.550 ;
      LAYER Metal2 ;
        RECT 56.685 1.240 59.780 1.560 ;
        RECT 59.500 -2.100 59.780 1.240 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    PORT
      LAYER Metal1 ;
        RECT 65.060 6.190 65.435 7.310 ;
      LAYER Via1 ;
        RECT 65.090 6.290 65.390 6.590 ;
      LAYER Metal2 ;
        RECT 62.860 6.280 65.490 6.600 ;
        RECT 62.860 3.160 63.140 6.280 ;
        RECT 62.835 2.860 63.140 3.160 ;
        RECT 62.835 0.075 63.115 2.860 ;
        RECT 62.835 -0.210 63.140 0.075 ;
        RECT 62.860 -2.100 63.140 -0.210 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    PORT
      LAYER Metal1 ;
        RECT 65.060 0.530 65.435 1.650 ;
      LAYER Via1 ;
        RECT 65.090 1.250 65.390 1.550 ;
      LAYER Metal2 ;
        RECT 63.405 1.240 66.500 1.560 ;
        RECT 66.220 -2.100 66.500 1.240 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    PORT
      LAYER Metal1 ;
        RECT 9.060 0.530 9.435 1.650 ;
      LAYER Via1 ;
        RECT 9.090 1.250 9.390 1.550 ;
      LAYER Metal2 ;
        RECT 3.500 1.240 9.500 1.560 ;
        RECT 3.500 -2.100 3.780 1.240 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    PORT
      LAYER Metal1 ;
        RECT 70.660 6.190 71.035 7.310 ;
      LAYER Via1 ;
        RECT 70.690 6.290 70.990 6.590 ;
      LAYER Metal2 ;
        RECT 68.160 6.280 71.090 6.600 ;
        RECT 68.160 0.195 68.440 6.280 ;
        RECT 68.160 -0.085 70.420 0.195 ;
        RECT 70.140 -2.100 70.420 -0.085 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    PORT
      LAYER Metal1 ;
        RECT 70.660 0.530 71.035 1.650 ;
      LAYER Via1 ;
        RECT 70.690 1.250 70.990 1.550 ;
      LAYER Metal2 ;
        RECT 69.005 1.240 73.780 1.560 ;
        RECT 73.500 -2.100 73.780 1.240 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    PORT
      LAYER Metal1 ;
        RECT 77.380 6.190 77.755 7.310 ;
      LAYER Via1 ;
        RECT 77.410 6.290 77.710 6.590 ;
      LAYER Metal2 ;
        RECT 74.925 6.280 77.800 6.600 ;
        RECT 74.925 0.605 75.205 6.280 ;
        RECT 74.925 0.325 77.140 0.605 ;
        RECT 76.860 -2.100 77.140 0.325 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    PORT
      LAYER Metal1 ;
        RECT 77.380 0.530 77.755 1.650 ;
      LAYER Via1 ;
        RECT 77.410 1.250 77.710 1.550 ;
      LAYER Metal2 ;
        RECT 75.725 1.240 80.500 1.560 ;
        RECT 80.220 -2.100 80.500 1.240 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    PORT
      LAYER Metal1 ;
        RECT 82.980 6.190 83.355 7.310 ;
        RECT 83.590 1.885 83.890 2.305 ;
        RECT 83.610 1.005 83.875 1.885 ;
        RECT 83.590 0.585 83.890 1.005 ;
      LAYER Via1 ;
        RECT 83.010 6.290 83.310 6.590 ;
        RECT 83.590 1.945 83.890 2.245 ;
        RECT 83.590 0.645 83.890 0.945 ;
      LAYER Metal2 ;
        RECT 81.320 6.280 83.890 6.600 ;
        RECT 83.610 2.255 83.890 6.280 ;
        RECT 83.520 1.935 83.985 2.255 ;
        RECT 83.475 0.645 83.985 0.955 ;
        RECT 83.580 0.635 83.985 0.645 ;
        RECT 83.580 -2.100 83.860 0.635 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    PORT
      LAYER Metal1 ;
        RECT 82.980 0.530 83.355 1.650 ;
      LAYER Via1 ;
        RECT 83.010 1.250 83.310 1.550 ;
      LAYER Metal2 ;
        RECT 81.325 1.240 87.755 1.560 ;
        RECT 87.475 -0.040 87.755 1.240 ;
        RECT 87.475 -0.515 87.780 -0.040 ;
        RECT 87.500 -2.100 87.780 -0.515 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    PORT
      LAYER Metal1 ;
        RECT 89.700 6.190 90.075 7.310 ;
        RECT 90.375 1.860 90.675 2.280 ;
        RECT 90.395 0.980 90.660 1.860 ;
        RECT 90.375 0.560 90.675 0.980 ;
      LAYER Via1 ;
        RECT 89.730 6.290 90.030 6.590 ;
        RECT 90.375 1.920 90.675 2.220 ;
        RECT 90.375 0.620 90.675 0.920 ;
      LAYER Metal2 ;
        RECT 88.045 6.280 90.665 6.600 ;
        RECT 90.385 2.230 90.665 6.280 ;
        RECT 90.315 1.910 90.735 2.230 ;
        RECT 90.315 0.610 91.140 0.930 ;
        RECT 90.860 -2.100 91.140 0.610 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    PORT
      LAYER Metal1 ;
        RECT 89.700 0.530 90.075 1.650 ;
      LAYER Via1 ;
        RECT 89.730 1.250 90.030 1.550 ;
      LAYER Metal2 ;
        RECT 88.045 1.240 92.035 1.560 ;
        RECT 91.755 0.715 92.035 1.240 ;
        RECT 91.755 0.435 94.500 0.715 ;
        RECT 94.220 -2.100 94.500 0.435 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    PORT
      LAYER Metal1 ;
        RECT 95.300 6.190 95.675 7.310 ;
        RECT 95.950 1.885 96.250 2.305 ;
        RECT 95.970 1.005 96.235 1.885 ;
        RECT 95.950 0.585 96.250 1.005 ;
      LAYER Via1 ;
        RECT 95.330 6.290 95.630 6.590 ;
        RECT 95.950 1.945 96.250 2.245 ;
        RECT 95.950 0.645 96.250 0.945 ;
      LAYER Metal2 ;
        RECT 93.650 6.280 96.240 6.600 ;
        RECT 95.960 2.255 96.240 6.280 ;
        RECT 95.890 1.930 96.310 2.255 ;
        RECT 95.890 0.675 97.860 0.955 ;
        RECT 95.890 0.630 96.310 0.675 ;
        RECT 97.580 -2.100 97.860 0.675 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    PORT
      LAYER Metal1 ;
        RECT 95.300 0.530 95.675 1.650 ;
      LAYER Via1 ;
        RECT 95.330 1.250 95.630 1.550 ;
      LAYER Metal2 ;
        RECT 93.635 1.240 98.995 1.560 ;
        RECT 98.715 0.895 98.995 1.240 ;
        RECT 98.715 0.615 101.780 0.895 ;
        RECT 101.500 -2.100 101.780 0.615 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    PORT
      LAYER Metal1 ;
        RECT 15.780 6.190 16.155 7.310 ;
      LAYER Via1 ;
        RECT 15.810 6.290 16.110 6.590 ;
      LAYER Metal2 ;
        RECT 11.725 6.280 16.220 6.600 ;
        RECT 11.725 0.890 12.005 6.280 ;
        RECT 7.420 0.610 12.005 0.890 ;
        RECT 7.420 -2.100 7.700 0.610 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    PORT
      LAYER Metal1 ;
        RECT 102.020 6.190 102.395 7.310 ;
        RECT 102.655 1.860 102.955 2.280 ;
        RECT 102.680 0.980 102.945 1.860 ;
        RECT 102.655 0.560 102.955 0.980 ;
      LAYER Via1 ;
        RECT 102.050 6.290 102.350 6.590 ;
        RECT 102.655 1.920 102.955 2.220 ;
        RECT 102.655 0.620 102.955 0.920 ;
      LAYER Metal2 ;
        RECT 100.365 6.280 102.945 6.600 ;
        RECT 102.665 2.230 102.945 6.280 ;
        RECT 102.595 1.910 103.015 2.230 ;
        RECT 102.595 0.905 103.015 0.930 ;
        RECT 102.595 0.625 105.140 0.905 ;
        RECT 102.595 0.610 103.015 0.625 ;
        RECT 104.860 -2.100 105.140 0.625 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    PORT
      LAYER Metal1 ;
        RECT 102.020 0.530 102.395 1.650 ;
      LAYER Via1 ;
        RECT 102.050 1.250 102.350 1.550 ;
      LAYER Metal2 ;
        RECT 100.365 1.240 108.500 1.560 ;
        RECT 108.220 -2.100 108.500 1.240 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    PORT
      LAYER Metal1 ;
        RECT 15.780 0.530 16.155 1.650 ;
      LAYER Via1 ;
        RECT 15.810 1.250 16.110 1.550 ;
      LAYER Metal2 ;
        RECT 12.745 1.240 16.220 1.560 ;
        RECT 12.745 0.190 13.025 1.240 ;
        RECT 10.780 -0.090 13.025 0.190 ;
        RECT 10.780 -2.100 11.060 -0.090 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    PORT
      LAYER Metal1 ;
        RECT 21.380 6.190 21.755 7.310 ;
      LAYER Via1 ;
        RECT 21.410 6.290 21.710 6.590 ;
      LAYER Metal2 ;
        RECT 16.600 6.280 21.820 6.600 ;
        RECT 16.600 0.240 16.880 6.280 ;
        RECT 14.140 -0.040 16.880 0.240 ;
        RECT 14.140 -2.100 14.420 -0.040 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    PORT
      LAYER Metal1 ;
        RECT 21.380 0.530 21.755 1.650 ;
      LAYER Via1 ;
        RECT 21.410 1.250 21.710 1.550 ;
      LAYER Metal2 ;
        RECT 17.390 1.240 21.820 1.560 ;
        RECT 17.500 -2.100 17.780 1.240 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    PORT
      LAYER Metal1 ;
        RECT 28.100 6.190 28.475 7.310 ;
      LAYER Via1 ;
        RECT 28.130 6.290 28.430 6.590 ;
      LAYER Metal2 ;
        RECT 23.735 6.280 28.540 6.600 ;
        RECT 23.735 0.670 24.015 6.280 ;
        RECT 20.860 0.390 24.015 0.670 ;
        RECT 20.860 -2.100 21.140 0.390 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    PORT
      LAYER Metal1 ;
        RECT 28.100 0.530 28.475 1.650 ;
      LAYER Via1 ;
        RECT 28.130 1.250 28.430 1.550 ;
      LAYER Metal2 ;
        RECT 24.670 1.240 28.540 1.560 ;
        RECT 24.780 -2.100 25.060 1.240 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    PORT
      LAYER Metal1 ;
        RECT 33.700 6.190 34.075 7.310 ;
      LAYER Via1 ;
        RECT 33.730 6.290 34.030 6.590 ;
      LAYER Metal2 ;
        RECT 30.370 6.280 34.140 6.600 ;
        RECT 30.370 0.445 30.650 6.280 ;
        RECT 28.140 0.165 30.650 0.445 ;
        RECT 28.140 -2.100 28.420 0.165 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    PORT
      LAYER Metal1 ;
        RECT 33.700 0.530 34.075 1.650 ;
      LAYER Via1 ;
        RECT 33.730 1.250 34.030 1.550 ;
      LAYER Metal2 ;
        RECT 31.500 1.240 34.140 1.560 ;
        RECT 31.500 -2.100 31.780 1.240 ;
    END
  END mask_rev[9]
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 4.220 1.995 5.350 ;
        RECT 4.005 4.220 4.235 5.350 ;
        RECT 4.850 4.220 5.190 5.920 ;
        RECT 5.850 4.220 6.080 5.480 ;
        RECT 8.185 4.220 8.415 5.495 ;
        RECT 11.845 4.220 12.075 5.350 ;
        RECT 12.570 4.220 12.800 5.480 ;
        RECT 14.905 4.220 15.135 5.495 ;
        RECT 17.190 4.220 17.530 5.910 ;
        RECT 18.170 4.220 18.400 5.480 ;
        RECT 20.505 4.220 20.735 5.495 ;
        RECT 24.165 4.220 24.395 5.350 ;
        RECT 24.890 4.220 25.120 5.480 ;
        RECT 27.225 4.220 27.455 5.495 ;
        RECT 29.510 4.220 29.850 5.910 ;
        RECT 30.490 4.220 30.720 5.480 ;
        RECT 32.825 4.220 33.055 5.495 ;
        RECT 36.485 4.220 36.715 5.350 ;
        RECT 37.210 4.220 37.440 5.480 ;
        RECT 39.545 4.220 39.775 5.495 ;
        RECT 41.830 4.220 42.170 5.910 ;
        RECT 42.810 4.220 43.040 5.480 ;
        RECT 45.145 4.220 45.375 5.495 ;
        RECT 48.805 4.220 49.035 5.350 ;
        RECT 49.530 4.220 49.760 5.480 ;
        RECT 51.865 4.220 52.095 5.495 ;
        RECT 54.150 4.220 54.490 5.910 ;
        RECT 55.130 4.220 55.360 5.480 ;
        RECT 57.465 4.220 57.695 5.495 ;
        RECT 61.125 4.220 61.355 5.350 ;
        RECT 61.850 4.220 62.080 5.480 ;
        RECT 64.185 4.220 64.415 5.495 ;
        RECT 66.470 4.220 66.810 5.910 ;
        RECT 67.450 4.220 67.680 5.480 ;
        RECT 69.785 4.220 70.015 5.495 ;
        RECT 73.445 4.220 73.675 5.350 ;
        RECT 74.170 4.220 74.400 5.480 ;
        RECT 76.505 4.220 76.735 5.495 ;
        RECT 78.790 4.220 79.130 5.910 ;
        RECT 79.770 4.220 80.000 5.480 ;
        RECT 82.105 4.220 82.335 5.495 ;
        RECT 85.765 4.220 85.995 5.350 ;
        RECT 86.490 4.220 86.720 5.480 ;
        RECT 88.825 4.220 89.055 5.495 ;
        RECT 91.110 4.220 91.450 5.910 ;
        RECT 92.090 4.220 92.320 5.480 ;
        RECT 94.425 4.220 94.655 5.495 ;
        RECT 98.085 4.220 98.315 5.350 ;
        RECT 98.810 4.220 99.040 5.480 ;
        RECT 101.145 4.220 101.375 5.495 ;
        RECT 103.410 4.220 103.750 5.920 ;
        RECT 105.925 4.220 106.155 5.350 ;
        RECT 108.165 4.220 108.395 5.350 ;
        RECT 0.000 3.620 108.640 4.220 ;
        RECT 1.765 2.490 1.995 3.620 ;
        RECT 4.005 2.490 4.235 3.620 ;
        RECT 4.850 1.920 5.190 3.620 ;
        RECT 5.850 2.360 6.080 3.620 ;
        RECT 8.185 2.345 8.415 3.620 ;
        RECT 11.845 2.490 12.075 3.620 ;
        RECT 12.570 2.360 12.800 3.620 ;
        RECT 14.905 2.345 15.135 3.620 ;
        RECT 17.190 1.930 17.530 3.620 ;
        RECT 18.170 2.360 18.400 3.620 ;
        RECT 20.505 2.345 20.735 3.620 ;
        RECT 24.165 2.490 24.395 3.620 ;
        RECT 24.890 2.360 25.120 3.620 ;
        RECT 27.225 2.345 27.455 3.620 ;
        RECT 29.510 1.930 29.850 3.620 ;
        RECT 30.490 2.360 30.720 3.620 ;
        RECT 32.825 2.345 33.055 3.620 ;
        RECT 36.485 2.490 36.715 3.620 ;
        RECT 37.210 2.360 37.440 3.620 ;
        RECT 39.545 2.345 39.775 3.620 ;
        RECT 41.830 1.930 42.170 3.620 ;
        RECT 42.810 2.360 43.040 3.620 ;
        RECT 45.145 2.345 45.375 3.620 ;
        RECT 48.805 2.490 49.035 3.620 ;
        RECT 49.530 2.360 49.760 3.620 ;
        RECT 51.865 2.345 52.095 3.620 ;
        RECT 54.150 1.930 54.490 3.620 ;
        RECT 55.130 2.360 55.360 3.620 ;
        RECT 57.465 2.345 57.695 3.620 ;
        RECT 61.125 2.490 61.355 3.620 ;
        RECT 61.850 2.360 62.080 3.620 ;
        RECT 64.185 2.345 64.415 3.620 ;
        RECT 66.470 1.930 66.810 3.620 ;
        RECT 67.450 2.360 67.680 3.620 ;
        RECT 69.785 2.345 70.015 3.620 ;
        RECT 73.445 2.490 73.675 3.620 ;
        RECT 74.170 2.360 74.400 3.620 ;
        RECT 76.505 2.345 76.735 3.620 ;
        RECT 78.790 1.930 79.130 3.620 ;
        RECT 79.770 2.360 80.000 3.620 ;
        RECT 82.105 2.345 82.335 3.620 ;
        RECT 85.765 2.490 85.995 3.620 ;
        RECT 86.490 2.360 86.720 3.620 ;
        RECT 88.825 2.345 89.055 3.620 ;
        RECT 91.110 1.930 91.450 3.620 ;
        RECT 92.090 2.360 92.320 3.620 ;
        RECT 94.425 2.345 94.655 3.620 ;
        RECT 98.085 2.490 98.315 3.620 ;
        RECT 98.810 2.360 99.040 3.620 ;
        RECT 101.145 2.345 101.375 3.620 ;
        RECT 103.410 1.920 103.750 3.620 ;
        RECT 105.925 2.490 106.155 3.620 ;
        RECT 108.165 2.490 108.395 3.620 ;
      LAYER Via1 ;
        RECT 31.080 3.620 32.530 4.220 ;
        RECT 76.080 3.620 77.530 4.220 ;
      LAYER Metal2 ;
        RECT 31.015 3.185 32.600 4.785 ;
        RECT 76.015 3.185 77.600 4.785 ;
      LAYER Via2 ;
        RECT 31.080 3.260 32.530 4.710 ;
        RECT 76.080 3.260 77.530 4.710 ;
      LAYER Metal3 ;
        RECT 30.985 -0.840 32.635 8.660 ;
        RECT 75.985 -0.840 77.635 8.660 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.540 108.640 8.140 ;
        RECT 0.245 6.745 0.475 7.540 ;
        RECT 2.485 6.745 2.715 7.540 ;
        RECT 4.850 6.650 5.190 7.540 ;
        RECT 5.850 6.680 6.080 7.540 ;
        RECT 8.085 6.680 8.315 7.540 ;
        RECT 10.325 6.745 10.555 7.540 ;
        RECT 12.570 6.680 12.800 7.540 ;
        RECT 14.805 6.680 15.035 7.540 ;
        RECT 17.190 6.655 17.530 7.540 ;
        RECT 18.170 6.680 18.400 7.540 ;
        RECT 20.405 6.680 20.635 7.540 ;
        RECT 22.645 6.745 22.875 7.540 ;
        RECT 24.890 6.680 25.120 7.540 ;
        RECT 27.125 6.680 27.355 7.540 ;
        RECT 29.510 6.655 29.850 7.540 ;
        RECT 30.490 6.680 30.720 7.540 ;
        RECT 32.725 6.680 32.955 7.540 ;
        RECT 34.965 6.745 35.195 7.540 ;
        RECT 37.210 6.680 37.440 7.540 ;
        RECT 39.445 6.680 39.675 7.540 ;
        RECT 41.830 6.655 42.170 7.540 ;
        RECT 42.810 6.680 43.040 7.540 ;
        RECT 45.045 6.680 45.275 7.540 ;
        RECT 47.285 6.745 47.515 7.540 ;
        RECT 49.530 6.680 49.760 7.540 ;
        RECT 51.765 6.680 51.995 7.540 ;
        RECT 54.150 6.655 54.490 7.540 ;
        RECT 55.130 6.680 55.360 7.540 ;
        RECT 57.365 6.680 57.595 7.540 ;
        RECT 59.605 6.745 59.835 7.540 ;
        RECT 61.850 6.680 62.080 7.540 ;
        RECT 64.085 6.680 64.315 7.540 ;
        RECT 66.470 6.655 66.810 7.540 ;
        RECT 67.450 6.680 67.680 7.540 ;
        RECT 69.685 6.680 69.915 7.540 ;
        RECT 71.925 6.745 72.155 7.540 ;
        RECT 74.170 6.680 74.400 7.540 ;
        RECT 76.405 6.680 76.635 7.540 ;
        RECT 78.790 6.655 79.130 7.540 ;
        RECT 79.770 6.680 80.000 7.540 ;
        RECT 82.005 6.680 82.235 7.540 ;
        RECT 84.245 6.745 84.475 7.540 ;
        RECT 86.490 6.680 86.720 7.540 ;
        RECT 88.725 6.680 88.955 7.540 ;
        RECT 91.110 6.655 91.450 7.540 ;
        RECT 92.090 6.680 92.320 7.540 ;
        RECT 94.325 6.680 94.555 7.540 ;
        RECT 96.565 6.745 96.795 7.540 ;
        RECT 98.810 6.680 99.040 7.540 ;
        RECT 101.045 6.680 101.275 7.540 ;
        RECT 103.410 6.650 103.750 7.540 ;
        RECT 104.405 6.745 104.635 7.540 ;
        RECT 106.645 6.745 106.875 7.540 ;
        RECT 0.245 0.300 0.475 1.095 ;
        RECT 2.485 0.300 2.715 1.095 ;
        RECT 4.850 0.300 5.190 1.190 ;
        RECT 5.850 0.300 6.080 1.160 ;
        RECT 8.085 0.300 8.315 1.160 ;
        RECT 10.325 0.300 10.555 1.095 ;
        RECT 12.570 0.300 12.800 1.160 ;
        RECT 14.805 0.300 15.035 1.160 ;
        RECT 17.190 0.300 17.530 1.185 ;
        RECT 18.170 0.300 18.400 1.160 ;
        RECT 20.405 0.300 20.635 1.160 ;
        RECT 22.645 0.300 22.875 1.095 ;
        RECT 24.890 0.300 25.120 1.160 ;
        RECT 27.125 0.300 27.355 1.160 ;
        RECT 29.510 0.300 29.850 1.185 ;
        RECT 30.490 0.300 30.720 1.160 ;
        RECT 32.725 0.300 32.955 1.160 ;
        RECT 34.965 0.300 35.195 1.095 ;
        RECT 37.210 0.300 37.440 1.160 ;
        RECT 39.445 0.300 39.675 1.160 ;
        RECT 41.830 0.300 42.170 1.185 ;
        RECT 42.810 0.300 43.040 1.160 ;
        RECT 45.045 0.300 45.275 1.160 ;
        RECT 47.285 0.300 47.515 1.095 ;
        RECT 49.530 0.300 49.760 1.160 ;
        RECT 51.765 0.300 51.995 1.160 ;
        RECT 54.150 0.300 54.490 1.185 ;
        RECT 55.130 0.300 55.360 1.160 ;
        RECT 57.365 0.300 57.595 1.160 ;
        RECT 59.605 0.300 59.835 1.095 ;
        RECT 61.850 0.300 62.080 1.160 ;
        RECT 64.085 0.300 64.315 1.160 ;
        RECT 66.470 0.300 66.810 1.185 ;
        RECT 67.450 0.300 67.680 1.160 ;
        RECT 69.685 0.300 69.915 1.160 ;
        RECT 71.925 0.300 72.155 1.095 ;
        RECT 74.170 0.300 74.400 1.160 ;
        RECT 76.405 0.300 76.635 1.160 ;
        RECT 78.790 0.300 79.130 1.185 ;
        RECT 79.770 0.300 80.000 1.160 ;
        RECT 82.005 0.300 82.235 1.160 ;
        RECT 84.245 0.300 84.475 1.095 ;
        RECT 86.490 0.300 86.720 1.160 ;
        RECT 88.725 0.300 88.955 1.160 ;
        RECT 91.110 0.300 91.450 1.185 ;
        RECT 92.090 0.300 92.320 1.160 ;
        RECT 94.325 0.300 94.555 1.160 ;
        RECT 96.565 0.300 96.795 1.095 ;
        RECT 98.810 0.300 99.040 1.160 ;
        RECT 101.045 0.300 101.275 1.160 ;
        RECT 103.410 0.300 103.750 1.190 ;
        RECT 104.405 0.300 104.635 1.095 ;
        RECT 106.645 0.300 106.875 1.095 ;
        RECT 0.000 -0.300 108.640 0.300 ;
      LAYER Via1 ;
        RECT 8.570 7.550 10.035 8.120 ;
        RECT 53.570 7.550 55.035 8.120 ;
        RECT 98.570 7.550 100.035 8.120 ;
        RECT 8.580 -0.285 10.020 0.285 ;
        RECT 53.580 -0.285 55.020 0.285 ;
        RECT 98.580 -0.285 100.020 0.285 ;
      LAYER Metal2 ;
        RECT 8.505 7.535 10.105 8.625 ;
        RECT 53.515 8.140 55.105 8.625 ;
        RECT 98.515 8.140 100.105 8.625 ;
        RECT 53.505 7.535 55.105 8.140 ;
        RECT 98.505 7.535 100.105 8.140 ;
        RECT 8.515 7.025 10.105 7.535 ;
        RECT 53.515 7.025 55.105 7.535 ;
        RECT 98.515 7.025 100.105 7.535 ;
        RECT 8.515 -0.815 10.100 0.300 ;
        RECT 53.515 -0.815 55.100 0.300 ;
        RECT 98.515 -0.815 100.100 0.300 ;
      LAYER Via2 ;
        RECT 8.570 7.070 10.035 8.570 ;
        RECT 53.570 7.070 55.035 8.570 ;
        RECT 98.570 7.070 100.035 8.570 ;
        RECT 8.630 -0.720 10.000 0.255 ;
        RECT 53.630 -0.720 55.000 0.255 ;
        RECT 98.630 -0.720 100.000 0.255 ;
      LAYER Metal3 ;
        RECT 8.485 -0.840 10.135 8.660 ;
        RECT 53.485 -0.840 55.135 8.660 ;
        RECT 98.485 -0.840 100.135 8.660 ;
    END
  END VSS
  OBS
      LAYER Pwell ;
        RECT -0.430 6.080 109.070 8.270 ;
      LAYER Nwell ;
        RECT -0.430 1.760 109.070 6.080 ;
      LAYER Pwell ;
        RECT -0.430 -0.430 109.070 1.760 ;
      LAYER Metal1 ;
        RECT 0.245 6.285 1.520 6.515 ;
        RECT 0.245 4.450 0.475 6.285 ;
        RECT 1.765 5.880 1.995 7.310 ;
        RECT 0.730 5.650 1.995 5.880 ;
        RECT 2.485 6.285 3.760 6.515 ;
        RECT 2.485 4.450 2.715 6.285 ;
        RECT 4.005 5.880 4.235 7.310 ;
        RECT 6.970 6.505 7.200 7.310 ;
        RECT 6.475 6.270 7.200 6.505 ;
      LAYER Metal1 ;
        RECT 7.470 5.990 7.845 7.260 ;
      LAYER Metal1 ;
        RECT 2.970 5.650 4.235 5.880 ;
      LAYER Metal1 ;
        RECT 6.820 5.630 7.845 5.990 ;
      LAYER Metal1 ;
        RECT 10.325 6.285 11.600 6.515 ;
        RECT 8.710 5.655 9.435 5.890 ;
      LAYER Metal1 ;
        RECT 6.820 4.450 7.180 5.630 ;
      LAYER Metal1 ;
        RECT 9.205 4.450 9.435 5.655 ;
        RECT 10.325 4.450 10.555 6.285 ;
        RECT 11.845 5.880 12.075 7.310 ;
        RECT 13.690 6.505 13.920 7.310 ;
        RECT 13.195 6.270 13.920 6.505 ;
      LAYER Metal1 ;
        RECT 14.190 5.990 14.565 7.260 ;
      LAYER Metal1 ;
        RECT 19.290 6.505 19.520 7.310 ;
        RECT 18.795 6.270 19.520 6.505 ;
      LAYER Metal1 ;
        RECT 19.790 5.990 20.165 7.260 ;
      LAYER Metal1 ;
        RECT 10.810 5.650 12.075 5.880 ;
      LAYER Metal1 ;
        RECT 13.540 5.630 14.565 5.990 ;
      LAYER Metal1 ;
        RECT 15.430 5.655 16.155 5.890 ;
      LAYER Metal1 ;
        RECT 13.540 4.450 13.900 5.630 ;
      LAYER Metal1 ;
        RECT 15.925 4.450 16.155 5.655 ;
      LAYER Metal1 ;
        RECT 19.140 5.630 20.165 5.990 ;
      LAYER Metal1 ;
        RECT 22.645 6.285 23.920 6.515 ;
        RECT 21.030 5.655 21.755 5.890 ;
      LAYER Metal1 ;
        RECT 19.140 4.450 19.500 5.630 ;
      LAYER Metal1 ;
        RECT 21.525 4.450 21.755 5.655 ;
        RECT 22.645 4.450 22.875 6.285 ;
        RECT 24.165 5.880 24.395 7.310 ;
        RECT 26.010 6.505 26.240 7.310 ;
        RECT 25.515 6.270 26.240 6.505 ;
      LAYER Metal1 ;
        RECT 26.510 5.990 26.885 7.260 ;
      LAYER Metal1 ;
        RECT 31.610 6.505 31.840 7.310 ;
        RECT 31.115 6.270 31.840 6.505 ;
      LAYER Metal1 ;
        RECT 32.110 5.990 32.485 7.260 ;
      LAYER Metal1 ;
        RECT 23.130 5.650 24.395 5.880 ;
      LAYER Metal1 ;
        RECT 25.860 5.630 26.885 5.990 ;
      LAYER Metal1 ;
        RECT 27.750 5.655 28.475 5.890 ;
      LAYER Metal1 ;
        RECT 25.860 4.450 26.220 5.630 ;
      LAYER Metal1 ;
        RECT 28.245 4.450 28.475 5.655 ;
      LAYER Metal1 ;
        RECT 31.460 5.630 32.485 5.990 ;
      LAYER Metal1 ;
        RECT 34.965 6.285 36.240 6.515 ;
        RECT 33.350 5.655 34.075 5.890 ;
      LAYER Metal1 ;
        RECT 31.460 4.450 31.820 5.630 ;
      LAYER Metal1 ;
        RECT 33.845 4.450 34.075 5.655 ;
        RECT 34.965 4.450 35.195 6.285 ;
        RECT 36.485 5.880 36.715 7.310 ;
        RECT 38.330 6.505 38.560 7.310 ;
        RECT 37.835 6.270 38.560 6.505 ;
      LAYER Metal1 ;
        RECT 38.830 5.990 39.205 7.260 ;
      LAYER Metal1 ;
        RECT 43.930 6.505 44.160 7.310 ;
        RECT 43.435 6.270 44.160 6.505 ;
      LAYER Metal1 ;
        RECT 44.430 5.990 44.805 7.260 ;
      LAYER Metal1 ;
        RECT 35.450 5.650 36.715 5.880 ;
      LAYER Metal1 ;
        RECT 38.180 5.630 39.205 5.990 ;
      LAYER Metal1 ;
        RECT 40.070 5.655 40.795 5.890 ;
      LAYER Metal1 ;
        RECT 38.180 4.450 38.540 5.630 ;
      LAYER Metal1 ;
        RECT 40.565 4.450 40.795 5.655 ;
      LAYER Metal1 ;
        RECT 43.780 5.630 44.805 5.990 ;
      LAYER Metal1 ;
        RECT 47.285 6.285 48.560 6.515 ;
        RECT 45.670 5.655 46.395 5.890 ;
      LAYER Metal1 ;
        RECT 43.780 4.450 44.140 5.630 ;
      LAYER Metal1 ;
        RECT 46.165 4.450 46.395 5.655 ;
        RECT 47.285 4.450 47.515 6.285 ;
        RECT 48.805 5.880 49.035 7.310 ;
        RECT 50.650 6.505 50.880 7.310 ;
        RECT 50.155 6.270 50.880 6.505 ;
      LAYER Metal1 ;
        RECT 51.150 5.990 51.525 7.260 ;
      LAYER Metal1 ;
        RECT 56.250 6.505 56.480 7.310 ;
        RECT 55.755 6.270 56.480 6.505 ;
      LAYER Metal1 ;
        RECT 56.750 5.990 57.125 7.260 ;
      LAYER Metal1 ;
        RECT 47.770 5.650 49.035 5.880 ;
      LAYER Metal1 ;
        RECT 50.500 5.630 51.525 5.990 ;
      LAYER Metal1 ;
        RECT 52.390 5.655 53.115 5.890 ;
      LAYER Metal1 ;
        RECT 50.500 4.450 50.860 5.630 ;
      LAYER Metal1 ;
        RECT 52.885 4.450 53.115 5.655 ;
      LAYER Metal1 ;
        RECT 56.100 5.630 57.125 5.990 ;
      LAYER Metal1 ;
        RECT 59.605 6.285 60.880 6.515 ;
        RECT 57.990 5.655 58.715 5.890 ;
      LAYER Metal1 ;
        RECT 56.100 4.450 56.460 5.630 ;
      LAYER Metal1 ;
        RECT 58.485 4.450 58.715 5.655 ;
        RECT 59.605 4.450 59.835 6.285 ;
        RECT 61.125 5.880 61.355 7.310 ;
        RECT 62.970 6.505 63.200 7.310 ;
        RECT 62.475 6.270 63.200 6.505 ;
      LAYER Metal1 ;
        RECT 63.470 5.990 63.845 7.260 ;
      LAYER Metal1 ;
        RECT 68.570 6.505 68.800 7.310 ;
        RECT 68.075 6.270 68.800 6.505 ;
      LAYER Metal1 ;
        RECT 69.070 5.990 69.445 7.260 ;
      LAYER Metal1 ;
        RECT 60.090 5.650 61.355 5.880 ;
      LAYER Metal1 ;
        RECT 62.820 5.630 63.845 5.990 ;
      LAYER Metal1 ;
        RECT 64.710 5.655 65.435 5.890 ;
      LAYER Metal1 ;
        RECT 62.820 4.450 63.180 5.630 ;
      LAYER Metal1 ;
        RECT 65.205 4.450 65.435 5.655 ;
      LAYER Metal1 ;
        RECT 68.420 5.630 69.445 5.990 ;
      LAYER Metal1 ;
        RECT 71.925 6.285 73.200 6.515 ;
        RECT 70.310 5.655 71.035 5.890 ;
      LAYER Metal1 ;
        RECT 68.420 4.450 68.780 5.630 ;
      LAYER Metal1 ;
        RECT 70.805 4.450 71.035 5.655 ;
        RECT 71.925 4.450 72.155 6.285 ;
        RECT 73.445 5.880 73.675 7.310 ;
        RECT 75.290 6.505 75.520 7.310 ;
        RECT 74.795 6.270 75.520 6.505 ;
      LAYER Metal1 ;
        RECT 75.790 5.990 76.165 7.260 ;
      LAYER Metal1 ;
        RECT 80.890 6.505 81.120 7.310 ;
        RECT 80.395 6.270 81.120 6.505 ;
      LAYER Metal1 ;
        RECT 81.390 5.990 81.765 7.260 ;
      LAYER Metal1 ;
        RECT 72.410 5.650 73.675 5.880 ;
      LAYER Metal1 ;
        RECT 75.140 5.630 76.165 5.990 ;
      LAYER Metal1 ;
        RECT 77.030 5.655 77.755 5.890 ;
      LAYER Metal1 ;
        RECT 75.140 4.450 75.500 5.630 ;
      LAYER Metal1 ;
        RECT 77.525 4.450 77.755 5.655 ;
      LAYER Metal1 ;
        RECT 80.740 5.630 81.765 5.990 ;
      LAYER Metal1 ;
        RECT 84.245 6.285 85.520 6.515 ;
        RECT 82.630 5.655 83.355 5.890 ;
      LAYER Metal1 ;
        RECT 80.740 4.450 81.100 5.630 ;
      LAYER Metal1 ;
        RECT 83.125 4.450 83.355 5.655 ;
        RECT 84.245 4.450 84.475 6.285 ;
        RECT 85.765 5.880 85.995 7.310 ;
        RECT 87.610 6.505 87.840 7.310 ;
        RECT 87.115 6.270 87.840 6.505 ;
      LAYER Metal1 ;
        RECT 88.110 5.990 88.485 7.260 ;
      LAYER Metal1 ;
        RECT 93.210 6.505 93.440 7.310 ;
        RECT 92.715 6.270 93.440 6.505 ;
      LAYER Metal1 ;
        RECT 93.710 5.990 94.085 7.260 ;
      LAYER Metal1 ;
        RECT 84.730 5.650 85.995 5.880 ;
      LAYER Metal1 ;
        RECT 87.460 5.630 88.485 5.990 ;
      LAYER Metal1 ;
        RECT 89.350 5.655 90.075 5.890 ;
      LAYER Metal1 ;
        RECT 87.460 4.450 87.820 5.630 ;
      LAYER Metal1 ;
        RECT 89.845 4.450 90.075 5.655 ;
      LAYER Metal1 ;
        RECT 93.060 5.630 94.085 5.990 ;
      LAYER Metal1 ;
        RECT 96.565 6.285 97.840 6.515 ;
        RECT 94.950 5.655 95.675 5.890 ;
      LAYER Metal1 ;
        RECT 93.060 4.450 93.420 5.630 ;
      LAYER Metal1 ;
        RECT 95.445 4.450 95.675 5.655 ;
        RECT 96.565 4.450 96.795 6.285 ;
        RECT 98.085 5.880 98.315 7.310 ;
        RECT 99.930 6.505 100.160 7.310 ;
        RECT 99.435 6.270 100.160 6.505 ;
      LAYER Metal1 ;
        RECT 100.430 5.990 100.805 7.260 ;
      LAYER Metal1 ;
        RECT 97.050 5.650 98.315 5.880 ;
      LAYER Metal1 ;
        RECT 99.780 5.630 100.805 5.990 ;
      LAYER Metal1 ;
        RECT 104.405 6.285 105.680 6.515 ;
        RECT 101.670 5.655 102.395 5.890 ;
      LAYER Metal1 ;
        RECT 99.780 4.450 100.140 5.630 ;
      LAYER Metal1 ;
        RECT 102.165 4.450 102.395 5.655 ;
        RECT 104.405 4.450 104.635 6.285 ;
        RECT 105.925 5.880 106.155 7.310 ;
        RECT 104.890 5.650 106.155 5.880 ;
        RECT 106.645 6.285 107.920 6.515 ;
        RECT 106.645 4.450 106.875 6.285 ;
        RECT 108.165 5.880 108.395 7.310 ;
        RECT 107.130 5.650 108.395 5.880 ;
        RECT 0.245 1.555 0.475 3.390 ;
        RECT 0.730 1.960 1.995 2.190 ;
        RECT 0.245 1.325 1.520 1.555 ;
        RECT 1.765 0.530 1.995 1.960 ;
        RECT 2.485 1.555 2.715 3.390 ;
      LAYER Metal1 ;
        RECT 6.820 2.210 7.180 3.390 ;
      LAYER Metal1 ;
        RECT 2.970 1.960 4.235 2.190 ;
        RECT 2.485 1.325 3.760 1.555 ;
        RECT 4.005 0.530 4.235 1.960 ;
      LAYER Metal1 ;
        RECT 6.820 1.850 7.845 2.210 ;
      LAYER Metal1 ;
        RECT 9.205 2.185 9.435 3.390 ;
        RECT 8.710 1.950 9.435 2.185 ;
        RECT 6.475 1.335 7.200 1.570 ;
        RECT 6.970 0.530 7.200 1.335 ;
      LAYER Metal1 ;
        RECT 7.470 0.580 7.845 1.850 ;
      LAYER Metal1 ;
        RECT 10.325 1.555 10.555 3.390 ;
      LAYER Metal1 ;
        RECT 13.540 2.210 13.900 3.390 ;
      LAYER Metal1 ;
        RECT 10.810 1.960 12.075 2.190 ;
        RECT 10.325 1.325 11.600 1.555 ;
        RECT 11.845 0.530 12.075 1.960 ;
      LAYER Metal1 ;
        RECT 13.540 1.850 14.565 2.210 ;
      LAYER Metal1 ;
        RECT 15.925 2.185 16.155 3.390 ;
        RECT 15.430 1.950 16.155 2.185 ;
      LAYER Metal1 ;
        RECT 19.140 2.210 19.500 3.390 ;
        RECT 19.140 1.850 20.165 2.210 ;
      LAYER Metal1 ;
        RECT 21.525 2.185 21.755 3.390 ;
        RECT 21.030 1.950 21.755 2.185 ;
        RECT 13.195 1.335 13.920 1.570 ;
        RECT 13.690 0.530 13.920 1.335 ;
      LAYER Metal1 ;
        RECT 14.190 0.580 14.565 1.850 ;
      LAYER Metal1 ;
        RECT 18.795 1.335 19.520 1.570 ;
        RECT 19.290 0.530 19.520 1.335 ;
      LAYER Metal1 ;
        RECT 19.790 0.580 20.165 1.850 ;
      LAYER Metal1 ;
        RECT 22.645 1.555 22.875 3.390 ;
      LAYER Metal1 ;
        RECT 25.860 2.210 26.220 3.390 ;
      LAYER Metal1 ;
        RECT 23.130 1.960 24.395 2.190 ;
        RECT 22.645 1.325 23.920 1.555 ;
        RECT 24.165 0.530 24.395 1.960 ;
      LAYER Metal1 ;
        RECT 25.860 1.850 26.885 2.210 ;
      LAYER Metal1 ;
        RECT 28.245 2.185 28.475 3.390 ;
        RECT 27.750 1.950 28.475 2.185 ;
      LAYER Metal1 ;
        RECT 31.460 2.210 31.820 3.390 ;
        RECT 31.460 1.850 32.485 2.210 ;
      LAYER Metal1 ;
        RECT 33.845 2.185 34.075 3.390 ;
        RECT 33.350 1.950 34.075 2.185 ;
        RECT 25.515 1.335 26.240 1.570 ;
        RECT 26.010 0.530 26.240 1.335 ;
      LAYER Metal1 ;
        RECT 26.510 0.580 26.885 1.850 ;
      LAYER Metal1 ;
        RECT 31.115 1.335 31.840 1.570 ;
        RECT 31.610 0.530 31.840 1.335 ;
      LAYER Metal1 ;
        RECT 32.110 0.580 32.485 1.850 ;
      LAYER Metal1 ;
        RECT 34.965 1.555 35.195 3.390 ;
      LAYER Metal1 ;
        RECT 38.180 2.210 38.540 3.390 ;
      LAYER Metal1 ;
        RECT 35.450 1.960 36.715 2.190 ;
        RECT 34.965 1.325 36.240 1.555 ;
        RECT 36.485 0.530 36.715 1.960 ;
      LAYER Metal1 ;
        RECT 38.180 1.850 39.205 2.210 ;
      LAYER Metal1 ;
        RECT 40.565 2.185 40.795 3.390 ;
        RECT 40.070 1.950 40.795 2.185 ;
      LAYER Metal1 ;
        RECT 43.780 2.210 44.140 3.390 ;
        RECT 43.780 1.850 44.805 2.210 ;
      LAYER Metal1 ;
        RECT 46.165 2.185 46.395 3.390 ;
        RECT 45.670 1.950 46.395 2.185 ;
        RECT 37.835 1.335 38.560 1.570 ;
        RECT 38.330 0.530 38.560 1.335 ;
      LAYER Metal1 ;
        RECT 38.830 0.580 39.205 1.850 ;
      LAYER Metal1 ;
        RECT 43.435 1.335 44.160 1.570 ;
        RECT 43.930 0.530 44.160 1.335 ;
      LAYER Metal1 ;
        RECT 44.430 0.580 44.805 1.850 ;
      LAYER Metal1 ;
        RECT 47.285 1.555 47.515 3.390 ;
      LAYER Metal1 ;
        RECT 50.500 2.210 50.860 3.390 ;
      LAYER Metal1 ;
        RECT 47.770 1.960 49.035 2.190 ;
        RECT 47.285 1.325 48.560 1.555 ;
        RECT 48.805 0.530 49.035 1.960 ;
      LAYER Metal1 ;
        RECT 50.500 1.850 51.525 2.210 ;
      LAYER Metal1 ;
        RECT 52.885 2.185 53.115 3.390 ;
        RECT 52.390 1.950 53.115 2.185 ;
      LAYER Metal1 ;
        RECT 56.100 2.210 56.460 3.390 ;
        RECT 56.100 1.850 57.125 2.210 ;
      LAYER Metal1 ;
        RECT 58.485 2.185 58.715 3.390 ;
        RECT 57.990 1.950 58.715 2.185 ;
        RECT 50.155 1.335 50.880 1.570 ;
        RECT 50.650 0.530 50.880 1.335 ;
      LAYER Metal1 ;
        RECT 51.150 0.580 51.525 1.850 ;
      LAYER Metal1 ;
        RECT 55.755 1.335 56.480 1.570 ;
        RECT 56.250 0.530 56.480 1.335 ;
      LAYER Metal1 ;
        RECT 56.750 0.580 57.125 1.850 ;
      LAYER Metal1 ;
        RECT 59.605 1.555 59.835 3.390 ;
      LAYER Metal1 ;
        RECT 62.820 2.210 63.180 3.390 ;
      LAYER Metal1 ;
        RECT 60.090 1.960 61.355 2.190 ;
        RECT 59.605 1.325 60.880 1.555 ;
        RECT 61.125 0.530 61.355 1.960 ;
      LAYER Metal1 ;
        RECT 62.820 1.850 63.845 2.210 ;
      LAYER Metal1 ;
        RECT 65.205 2.185 65.435 3.390 ;
        RECT 64.710 1.950 65.435 2.185 ;
      LAYER Metal1 ;
        RECT 68.420 2.210 68.780 3.390 ;
        RECT 68.420 1.850 69.445 2.210 ;
      LAYER Metal1 ;
        RECT 70.805 2.185 71.035 3.390 ;
        RECT 70.310 1.950 71.035 2.185 ;
        RECT 62.475 1.335 63.200 1.570 ;
        RECT 62.970 0.530 63.200 1.335 ;
      LAYER Metal1 ;
        RECT 63.470 0.580 63.845 1.850 ;
      LAYER Metal1 ;
        RECT 68.075 1.335 68.800 1.570 ;
        RECT 68.570 0.530 68.800 1.335 ;
      LAYER Metal1 ;
        RECT 69.070 0.580 69.445 1.850 ;
      LAYER Metal1 ;
        RECT 71.925 1.555 72.155 3.390 ;
      LAYER Metal1 ;
        RECT 75.140 2.210 75.500 3.390 ;
      LAYER Metal1 ;
        RECT 72.410 1.960 73.675 2.190 ;
        RECT 71.925 1.325 73.200 1.555 ;
        RECT 73.445 0.530 73.675 1.960 ;
      LAYER Metal1 ;
        RECT 75.140 1.850 76.165 2.210 ;
      LAYER Metal1 ;
        RECT 77.525 2.185 77.755 3.390 ;
        RECT 77.030 1.950 77.755 2.185 ;
      LAYER Metal1 ;
        RECT 80.740 2.210 81.100 3.390 ;
        RECT 80.740 1.850 81.765 2.210 ;
      LAYER Metal1 ;
        RECT 83.125 2.185 83.355 3.390 ;
        RECT 82.630 1.950 83.355 2.185 ;
        RECT 74.795 1.335 75.520 1.570 ;
        RECT 75.290 0.530 75.520 1.335 ;
      LAYER Metal1 ;
        RECT 75.790 0.580 76.165 1.850 ;
      LAYER Metal1 ;
        RECT 80.395 1.335 81.120 1.570 ;
        RECT 80.890 0.530 81.120 1.335 ;
      LAYER Metal1 ;
        RECT 81.390 0.580 81.765 1.850 ;
      LAYER Metal1 ;
        RECT 84.245 1.555 84.475 3.390 ;
      LAYER Metal1 ;
        RECT 87.460 2.210 87.820 3.390 ;
      LAYER Metal1 ;
        RECT 84.730 1.960 85.995 2.190 ;
        RECT 84.245 1.325 85.520 1.555 ;
        RECT 85.765 0.530 85.995 1.960 ;
      LAYER Metal1 ;
        RECT 87.460 1.850 88.485 2.210 ;
      LAYER Metal1 ;
        RECT 89.845 2.185 90.075 3.390 ;
        RECT 89.350 1.950 90.075 2.185 ;
      LAYER Metal1 ;
        RECT 93.060 2.210 93.420 3.390 ;
        RECT 93.060 1.850 94.085 2.210 ;
      LAYER Metal1 ;
        RECT 95.445 2.185 95.675 3.390 ;
        RECT 94.950 1.950 95.675 2.185 ;
        RECT 87.115 1.335 87.840 1.570 ;
        RECT 87.610 0.530 87.840 1.335 ;
      LAYER Metal1 ;
        RECT 88.110 0.580 88.485 1.850 ;
      LAYER Metal1 ;
        RECT 92.715 1.335 93.440 1.570 ;
        RECT 93.210 0.530 93.440 1.335 ;
      LAYER Metal1 ;
        RECT 93.710 0.580 94.085 1.850 ;
      LAYER Metal1 ;
        RECT 96.565 1.555 96.795 3.390 ;
      LAYER Metal1 ;
        RECT 99.780 2.210 100.140 3.390 ;
      LAYER Metal1 ;
        RECT 97.050 1.960 98.315 2.190 ;
        RECT 96.565 1.325 97.840 1.555 ;
        RECT 98.085 0.530 98.315 1.960 ;
      LAYER Metal1 ;
        RECT 99.780 1.850 100.805 2.210 ;
      LAYER Metal1 ;
        RECT 102.165 2.185 102.395 3.390 ;
        RECT 101.670 1.950 102.395 2.185 ;
        RECT 99.435 1.335 100.160 1.570 ;
        RECT 99.930 0.530 100.160 1.335 ;
      LAYER Metal1 ;
        RECT 100.430 0.580 100.805 1.850 ;
      LAYER Metal1 ;
        RECT 104.405 1.555 104.635 3.390 ;
        RECT 104.890 1.960 106.155 2.190 ;
        RECT 104.405 1.325 105.680 1.555 ;
        RECT 105.925 0.530 106.155 1.960 ;
        RECT 106.645 1.555 106.875 3.390 ;
        RECT 107.130 1.960 108.395 2.190 ;
        RECT 106.645 1.325 107.920 1.555 ;
        RECT 108.165 0.530 108.395 1.960 ;
  END
END user_id_programming
END LIBRARY

