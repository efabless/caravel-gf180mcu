magic
tech gf180mcuC
magscale 1 10
timestamp 1655473235
<< checkpaint >>
rect -2056 -2056 17000 16000
<< obsm1 >>
rect 1120 1318 14822 12906
<< metal2 >>
rect -56 13200 56 14000
rect 1288 13200 1400 14000
rect 2632 13200 2744 14000
rect 3976 13200 4088 14000
rect 5320 13200 5432 14000
rect 6664 13200 6776 14000
rect 8008 13200 8120 14000
rect 9352 13200 9464 14000
rect 10696 13200 10808 14000
rect 12040 13200 12152 14000
rect 13384 13200 13496 14000
rect 14728 13200 14840 14000
rect 0 -56 800 56
rect 1288 0 1400 800
rect 2632 0 2744 800
rect 3976 0 4088 800
rect 5320 0 5432 800
rect 6664 0 6776 800
rect 8008 0 8120 800
rect 9352 0 9464 800
rect 10696 0 10808 800
rect 12040 0 12152 800
rect 13384 0 13496 800
rect 14728 0 14840 800
<< obsm2 >>
rect -28 13140 28 13200
rect 116 13140 1228 13356
rect 1460 13140 2572 13356
rect 2804 13140 3916 13356
rect 4148 13140 5260 13356
rect 5492 13140 6604 13356
rect 6836 13140 7948 13356
rect 8180 13140 9292 13356
rect 9524 13140 10636 13356
rect 10868 13140 11980 13356
rect 12212 13140 13324 13356
rect 13556 13140 14668 13356
rect -28 12740 14812 13140
rect 0 860 14812 12740
rect 0 116 1228 860
rect 860 28 1228 116
rect 800 0 1228 28
rect 1460 0 2572 860
rect 2804 0 3916 860
rect 4148 0 5260 860
rect 5492 0 6604 860
rect 6836 0 7948 860
rect 8180 0 9292 860
rect 9524 0 10636 860
rect 10868 0 11980 860
rect 12212 0 13324 860
rect 13556 0 14668 860
rect 800 -28 1148 0
<< metal3 >>
rect 0 12824 800 12936
rect 14200 12824 15000 12936
rect 0 11480 800 11592
rect 14200 11480 15000 11592
rect 0 10136 800 10248
rect 14200 10136 15000 10248
rect 0 8792 800 8904
rect 14200 8792 15000 8904
rect 0 7448 800 7560
rect 14200 7448 15000 7560
rect 0 6104 800 6216
rect 14200 6104 15000 6216
rect 0 4760 800 4872
rect 14200 4760 15000 4872
rect 0 3416 800 3528
rect 14200 3416 15000 3528
rect 0 2072 800 2184
rect 14200 2072 15000 2184
rect 0 728 800 840
rect 14200 728 15000 840
<< obsm3 >>
rect 860 12764 14140 12908
rect 74 11652 14364 12764
rect 860 11420 14140 11652
rect 74 10308 14364 11420
rect 860 10076 14140 10308
rect 74 8964 14364 10076
rect 860 8732 14140 8964
rect 74 7620 14364 8732
rect 860 7388 14140 7620
rect 74 6276 14364 7388
rect 860 6044 14140 6276
rect 74 4932 14364 6044
rect 860 4700 14140 4932
rect 74 3588 14364 4700
rect 860 3356 14140 3588
rect 74 2244 14364 3356
rect 860 2012 14140 2244
rect 74 900 14364 2012
rect 860 756 14140 900
<< metal4 >>
rect 2555 1508 2875 11820
rect 4150 1508 4470 11820
rect 5745 1508 6065 11820
rect 7340 1508 7660 11820
rect 8935 1508 9255 11820
rect 10530 1508 10850 11820
rect 12125 1508 12445 11820
<< metal5 >>
rect 1060 10914 13836 11234
rect 1060 9556 13836 9876
rect 1060 8198 13836 8518
rect 1060 6840 13836 7160
rect 1060 5482 13836 5802
rect 1060 4124 13836 4444
rect 1060 2766 13836 3086
<< labels >>
rlabel metal4 s 2555 1508 2875 11820 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 5745 1508 6065 11820 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 8935 1508 9255 11820 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 12125 1508 12445 11820 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1060 2766 13836 3086 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1060 5482 13836 5802 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1060 8198 13836 8518 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1060 10914 13836 11234 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 4150 1508 4470 11820 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 7340 1508 7660 11820 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 10530 1508 10850 11820 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 1060 4124 13836 4444 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 1060 6840 13836 7160 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 1060 9556 13836 9876 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 4760 800 4872 6 spare_xfq[0]
port 3 nsew signal output
rlabel metal2 s 13384 0 13496 800 6 spare_xfq[1]
port 4 nsew signal output
rlabel metal2 s 6664 13200 6776 14000 6 spare_xi[0]
port 5 nsew signal output
rlabel metal2 s 5320 0 5432 800 6 spare_xi[1]
port 6 nsew signal output
rlabel metal3 s 14200 2072 15000 2184 6 spare_xi[2]
port 7 nsew signal output
rlabel metal3 s 0 10136 800 10248 6 spare_xi[3]
port 8 nsew signal output
rlabel metal3 s 14200 728 15000 840 6 spare_xib
port 9 nsew signal output
rlabel metal2 s 14728 0 14840 800 6 spare_xmx[0]
port 10 nsew signal output
rlabel metal3 s 14200 10136 15000 10248 6 spare_xmx[1]
port 11 nsew signal output
rlabel metal2 s -56 13200 56 14000 4 spare_xna[0]
port 12 nsew signal output
rlabel metal2 s 8008 0 8120 800 6 spare_xna[1]
port 13 nsew signal output
rlabel metal3 s 0 3416 800 3528 6 spare_xno[0]
port 14 nsew signal output
rlabel metal2 s 10696 0 10808 800 6 spare_xno[1]
port 15 nsew signal output
rlabel metal3 s 14200 11480 15000 11592 6 spare_xz[0]
port 16 nsew signal output
rlabel metal3 s 0 7448 800 7560 6 spare_xz[10]
port 17 nsew signal output
rlabel metal2 s 2632 0 2744 800 6 spare_xz[11]
port 18 nsew signal output
rlabel metal2 s 13384 13200 13496 14000 6 spare_xz[12]
port 19 nsew signal output
rlabel metal2 s 9352 13200 9464 14000 6 spare_xz[13]
port 20 nsew signal output
rlabel metal3 s 14200 7448 15000 7560 6 spare_xz[14]
port 21 nsew signal output
rlabel metal2 s 12040 13200 12152 14000 6 spare_xz[15]
port 22 nsew signal output
rlabel metal3 s 0 2072 800 2184 6 spare_xz[16]
port 23 nsew signal output
rlabel metal3 s 14200 12824 15000 12936 6 spare_xz[17]
port 24 nsew signal output
rlabel metal2 s 2632 13200 2744 14000 6 spare_xz[18]
port 25 nsew signal output
rlabel metal2 s 0 -56 800 56 8 spare_xz[19]
port 26 nsew signal output
rlabel metal2 s 8008 13200 8120 14000 6 spare_xz[1]
port 27 nsew signal output
rlabel metal3 s 14200 8792 15000 8904 6 spare_xz[20]
port 28 nsew signal output
rlabel metal2 s 1288 13200 1400 14000 6 spare_xz[21]
port 29 nsew signal output
rlabel metal3 s 0 728 800 840 6 spare_xz[22]
port 30 nsew signal output
rlabel metal2 s 12040 0 12152 800 6 spare_xz[23]
port 31 nsew signal output
rlabel metal2 s 10696 13200 10808 14000 6 spare_xz[24]
port 32 nsew signal output
rlabel metal3 s 14200 3416 15000 3528 6 spare_xz[25]
port 33 nsew signal output
rlabel metal2 s 1288 0 1400 800 6 spare_xz[26]
port 34 nsew signal output
rlabel metal2 s 3976 0 4088 800 6 spare_xz[27]
port 35 nsew signal output
rlabel metal3 s 0 11480 800 11592 6 spare_xz[28]
port 36 nsew signal output
rlabel metal3 s 14200 4760 15000 4872 6 spare_xz[29]
port 37 nsew signal output
rlabel metal2 s 6664 0 6776 800 6 spare_xz[2]
port 38 nsew signal output
rlabel metal3 s 0 8792 800 8904 6 spare_xz[30]
port 39 nsew signal output
rlabel metal2 s 14728 13200 14840 14000 6 spare_xz[3]
port 40 nsew signal output
rlabel metal2 s 3976 13200 4088 14000 6 spare_xz[4]
port 41 nsew signal output
rlabel metal2 s 5320 13200 5432 14000 6 spare_xz[5]
port 42 nsew signal output
rlabel metal2 s 9352 0 9464 800 6 spare_xz[6]
port 43 nsew signal output
rlabel metal3 s 0 6104 800 6216 6 spare_xz[7]
port 44 nsew signal output
rlabel metal3 s 0 12824 800 12936 6 spare_xz[8]
port 45 nsew signal output
rlabel metal3 s 14200 6104 15000 6216 6 spare_xz[9]
port 46 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 15000 14000
string GDS_END 193670
string GDS_FILE ../gds/spare_logic_block.gds.gz
string GDS_START 78910
string LEFclass BLOCK
string LEFview TRUE
<< end >>
