* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_20 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_12 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_20 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_16 I ZN VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_95_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6914_ _6914_/D _7315_/RN _6914_/CLK _6914_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ hold41/Z _7300_/RN _6845_/CLK hold40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3988_ _6899_/Q _5891_/A4 _5560_/A1 _4408_/A1 _4016_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6776_ _6776_/D _7359_/RN _6776_/CLK _6776_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5727_ hold79/Z hold407/Z _5731_/S _7093_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5658_ hold38/Z _7032_/Q hold8/Z hold39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ _4773_/C _4702_/B _5306_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_124_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ hold363/Z hold836/Z _5596_/S _5589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold362 _7332_/Q hold362/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold351 _5895_/Z _7239_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold340 _7263_/Q hold340/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7328_ _7328_/D _7331_/CLK _7328_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7259_ _7259_/D _7286_/RN _7259_/CLK _7259_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold395 _7104_/Q hold395/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold384 _6829_/Q hold384/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold373 _7020_/Q hold373/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _4960_/A1 _4960_/A2 _4483_/B _4711_/B _4964_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4891_ _4691_/C _5490_/B _5308_/B _5353_/A4 _5361_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3911_ _4402_/A4 _5872_/A4 _5581_/A3 _4402_/A3 _4015_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6630_ _6632_/A2 _6894_/Q _6675_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3842_ _7246_/Q _4019_/A2 _4320_/S input37/Z _3914_/A2 _7222_/Q _3845_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_32_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6561_ _6561_/A1 _6561_/A2 _6561_/A3 _6561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5512_ _5512_/A1 _5512_/A2 _5514_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3773_ _7110_/Q _4009_/B1 _3855_/B1 _6944_/Q _3776_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6492_ _7023_/Q _6321_/Z _6342_/Z _7249_/Q _6493_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5443_ _5515_/A1 _5482_/A2 _5443_/B _5444_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5374_ _5515_/A1 _5482_/A2 _5374_/B _5375_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ hold99/Z hold238/Z _4328_/S _6827_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7113_ hold95/Z _7322_/RN _7113_/CLK hold94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _7044_/D _7286_/RN _7044_/CLK _7044_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_101_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ hold825/Z hold323/Z _4256_/S _4256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4187_ hold59/Z hold369/Z _4193_/S _4187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6828_ _6828_/D input75/Z _6828_/CLK _6828_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _6759_/D _7359_/RN _6759_/CLK _6759_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold170 _7176_/Q hold170/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold181 _5600_/Z _6980_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold192 _7126_/Q hold192/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet679_320 net429_90/I _6967_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet679_331 net779_438/I _6956_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_342 net429_96/I _6945_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5090_ _5085_/Z _5251_/A1 _5483_/A2 _5253_/A1 _5092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4110_ _6727_/Q _6726_/Q _6792_/Q _3496_/Z _4110_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4041_ _7018_/Q _4041_/A2 _4041_/B1 input34/Z _4044_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _6387_/A2 _6337_/A4 _6593_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4943_ _5407_/B _5224_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4874_ _5516_/A1 _4874_/A2 _5463_/A1 _4874_/A4 _4876_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_138_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6613_ _6848_/Q _6613_/A2 _6613_/B _6613_/C _6615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3825_ _6996_/Q _5669_/A1 _5827_/A1 _5863_/A3 _3854_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6544_ _7147_/Q _6323_/Z _6334_/Z _7033_/Q _6352_/Z _7155_/Q _6547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3756_ _3752_/Z _3756_/A2 _3756_/A3 _3756_/A4 _3756_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_134_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6475_ _7168_/Q _6604_/A2 _6337_/Z _7070_/Q _6476_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5426_ _5508_/A4 _5508_/A2 _5507_/A2 _5470_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3687_ _7226_/Q _3914_/A2 _4033_/A2 _7234_/Q _3688_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput242 _7377_/Z mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput253 _4156_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput220 _4137_/ZN mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput231 _7374_/Z mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5357_ _5417_/C _5359_/A1 _5359_/A2 _5405_/A1 _4775_/Z _5358_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xoutput264 _6942_/Q pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput275 _6741_/Q pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput286 _6735_/Q pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4308_ hold630/Z hold323/Z _4320_/S _4308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5288_ _5216_/C _4518_/Z _5319_/A1 _5138_/B _5364_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput297 _6954_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4239_ _5564_/A1 _5882_/A2 _6677_/A3 _4241_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7027_ _7027_/D _7300_/RN _7027_/CLK _7027_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_28_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_261 net729_396/I _7026_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_294 net629_296/I _6993_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_272 net629_272/I _7015_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_283 net779_427/I _7004_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4590_ _4590_/A1 _4590_/A2 _4590_/A3 _4598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3610_ _3906_/A1 _5872_/A2 _3509_/Z _5872_/A3 _4037_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _4395_/A2 hold67/Z _3541_/B hold68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_127_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold906 _4290_/Z _6809_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_155_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6260_ _6915_/Q _6294_/A2 _6289_/B1 _6871_/Q _6262_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3472_ _4063_/A2 _3472_/A2 _6795_/Q _3472_/B _3473_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_170_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5211_ _5421_/A2 _5406_/A1 _5218_/B _5213_/B _5314_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6191_ _7039_/Q _6295_/A2 _6294_/B1 _7103_/Q _6192_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5142_ _5324_/A3 _5324_/A4 _5142_/B _5142_/C _5387_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_24__1403_ clkbuf_4_9_0__1403_/Z _4150__9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104__1403_ clkbuf_4_1_0__1403_/Z net429_99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5073_ _5073_/A1 _5375_/A1 _5074_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_87__1403_ clkbuf_4_4_0__1403_/Z net429_97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ _7172_/Q _4024_/A2 _4024_/B1 _6951_/Q _4024_/C _4025_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5975_ _5975_/I _7290_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4926_ _4926_/A1 _4926_/A2 _5320_/A1 _5320_/A2 _5320_/C _5052_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _4483_/B _4097_/B _4711_/B _5313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_138_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3808_ input14/Z _4031_/A2 _3914_/A2 _7223_/Q _3809_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4788_ _4787_/B _5040_/A4 _4788_/B _5342_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6527_ _7258_/Q _6319_/Z _6321_/Z _7024_/Q _6530_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3739_ _6733_/Q _3914_/B1 _5777_/A2 _5566_/A1 _3742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ _6458_/A1 _6458_/A2 _6989_/Q _6613_/A2 _6613_/C _6460_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_107_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ _5440_/C _5409_/A2 _5409_/B _5429_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6389_ _7181_/Q _6320_/Z _6325_/Z _7083_/Q _6337_/Z _7067_/Q _6392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_55 net429_55/I _7232_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_77 net429_89/I _7210_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_88 net429_90/I _7199_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_66 net429_83/I _7221_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet429_99 net429_99/I _7188_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ hold363/Z hold887/Z _5767_/S _5760_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _4959_/A1 _4730_/C _4711_/B _4718_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5691_ hold79/Z hold400/Z _5695_/S _5691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _4505_/Z _5534_/A1 _5380_/B _5061_/A3 _4643_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_175_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ _5295_/B2 _3402_/I _5475_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold703 _6941_/Q hold703/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7361_ _7361_/D _6713_/Z _4152_/I1 _7361_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6312_ _6543_/A2 _6355_/A4 _7296_/Q _6540_/A4 _6312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7292_ _7292_/D _7322_/RN _7322_/CLK _7292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3524_ _3884_/A1 _3554_/B _4405_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold714 _5707_/Z _7075_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold736 _5725_/Z _7091_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold725 _7074_/Q hold725/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold747 _7268_/Q hold747/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold769 _6955_/Q hold769/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3455_ _3421_/B _4160_/B _3472_/B _4058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xhold758 _7181_/Q hold758/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6243_ _7105_/Q _6294_/B1 _6292_/B1 _7073_/Q _6244_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet829_467 _4150__40/I _6760_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6174_ _6174_/I0 _7307_/Q _6434_/S _7307_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet829_478 net829_498/I _6749_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_456 net429_99/I _6771_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3386_ _7013_/Q _3386_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5125_ _5406_/A1 _5280_/B _5130_/B1 _5309_/B _5431_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet829_489 net829_498/I _6738_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5056_ _5384_/A1 _5059_/A2 _5261_/A2 _5482_/C _5487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4007_ _4007_/A1 _4007_/A2 _4007_/A3 _4007_/A4 _4008_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ _7287_/Q _5965_/A1 _5952_/B _6017_/A3 _5960_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_111_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _4691_/C _5421_/C _5206_/B _5353_/A4 _5313_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5889_ hold38/Z hold444/Z _5890_/S _5889_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold41 hold41/I hold41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold30 hold30/I hold30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_70__1403_ clkbuf_4_7_0__1403_/Z net629_298/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold63 hold63/I hold63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold52 hold52/I hold52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold74 hold74/I hold74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold96 hold96/I hold96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold85 hold85/I hold85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_16_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7319_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6930_ _6930_/D _6688_/Z _4152_/I1 _6930_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_35_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _6861_/D input75/Z _6861_/CLK _6861_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5812_ _5812_/A1 _5812_/A2 hold310/Z hold79/Z _5813_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6792_ _6792_/D _6683_/Z _4152_/I1 _6792_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_50_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ hold323/Z hold811/Z _5749_/S _7107_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5674_ hold59/Z hold293/Z _5677_/S _5674_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4625_ _5099_/C _4499_/B _4634_/A1 _4787_/B _5377_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold500 _5939_/Z _7278_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4556_ _4702_/B _5305_/B _4694_/B _5425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7344_ _7344_/D _6698_/Z _4152_/I1 _7344_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold511 _4418_/Z _6907_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold522 _5894_/Z _7238_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold544 _7393_/I hold544/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3507_ _3436_/B _3507_/A2 _4178_/S _3556_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold533 _6777_/Q hold533/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7275_ _7275_/D _7286_/RN _7275_/CLK _7275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4487_ _4483_/B _4523_/A2 _4488_/B _5441_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_143_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold566 _7158_/Q hold566/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold555 _7076_/Q hold555/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold577 _7376_/I hold577/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold588 _7375_/I hold588/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3438_ hold182/Z _6795_/Q _3440_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6226_ _6434_/S _6226_/A2 _6226_/B _7309_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold599 _4340_/Z _6840_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3369_ _7143_/Q _3369_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6157_ _7094_/Q _6290_/A2 _6293_/A2 _7078_/Q _6157_/C _6160_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _5406_/A1 _5108_/A2 _5130_/B1 _5353_/A3 _5354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ _6302_/A1 _6302_/A2 _6987_/Q _7293_/Q _6089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _4788_/B _5450_/A2 _5401_/A2 _5040_/A4 _5039_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_122_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput120 wb_adr_i[3] _4751_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_0_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput142 wb_dat_i[22] _6662_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput153 wb_dat_i[3] _6650_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput131 wb_dat_i[12] _6653_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput164 wb_sel_i[3] _6672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_91_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_400 net429_72/I _6836_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_4_0__1403_ clkbuf_0__1403_/Z clkbuf_4_9_0__1403_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4410_ hold323/Z hold695/Z _4410_/S _4410_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5390_ _5529_/B1 _5005_/Z _5390_/B _5390_/C _5454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ hold99/Z _6841_/Q _4346_/S _4341_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4272_ _4271_/Z hold903/Z _4286_/S _4272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7060_ _7060_/D _7315_/RN _7060_/CLK _7060_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_98_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6011_ _6805_/Q _6807_/Q _6007_/B _6011_/B _7299_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_39_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6913_ _6913_/D _7315_/RN _6913_/CLK _6913_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6844_ hold62/Z _7300_/RN _6844_/CLK hold61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3987_ _6756_/Q _5560_/A1 _5827_/A1 _6677_/A1 _4029_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6775_ _6775_/D _7359_/RN _6775_/CLK _6775_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5726_ hold99/Z hold552/Z _5731_/S _7092_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5657_ hold50/Z hold57/Z hold8/Z _7031_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4608_ _4634_/A1 _5252_/A2 _4716_/B _4608_/A4 _5374_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5588_ _5588_/A1 _5863_/A4 hold18/Z _6677_/A3 _5596_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold341 _5922_/Z _7263_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4539_ _3399_/I _5162_/A2 _4751_/B _4691_/C _5320_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold330 _4336_/Z _6837_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7327_ _7327_/D _7331_/CLK _7327_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold352 _6785_/Q hold352/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7258_ _7258_/D _7286_/RN _7258_/CLK _7258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold374 _7256_/Q hold374/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold363 _4178_/Z hold363/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold396 _6748_/Q hold396/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold385 _7190_/Q hold385/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6209_ _6209_/A1 _6209_/A2 _6209_/A3 _6209_/A4 _6210_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7189_ _7189_/D input75/Z _7189_/CLK _7189_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _4890_/A1 _5308_/B _5497_/A1 _4715_/B _4892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3910_ _3910_/A1 _3521_/Z _3523_/B _5872_/A4 _3913_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3841_ _3841_/A1 _3841_/A2 _3841_/A3 _3859_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6560_ _7283_/Q _6610_/A2 _6347_/C hold55/I _6561_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3772_ _5585_/A2 _3509_/Z _3504_/Z _5872_/A3 _3855_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_158_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _5511_/A1 _5511_/A2 _5511_/A3 _5512_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6491_ _7047_/Q _6609_/B1 _6341_/Z _6999_/Q _6493_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5442_ _5442_/A1 _5442_/A2 _5442_/A3 _5442_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5373_ _5373_/A1 _5373_/A2 _5373_/A3 _5373_/A4 _5376_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _7112_/D _7322_/RN _7112_/CLK _7112_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4324_ hold323/Z hold820/Z _4328_/S _6826_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7043_ _7043_/D _7315_/RN _7043_/CLK _7043_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_113_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4255_ hold893/Z hold363/Z _4256_/S _4255_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4186_ hold58/Z _7336_/Q _6881_/Q hold59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_27_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6827_ _6827_/D _7359_/RN _6827_/CLK _7397_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _6758_/D _7359_/RN _6758_/CLK _6758_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5709_ hold79/Z hold411/Z _5713_/S _5709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6689_ input75/Z _7012_/Q _4069_/C _6689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold160 _7133_/Q hold160/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold171 _5823_/Z _7176_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold182 _7366_/Q hold182/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold193 _5764_/Z _7126_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_58_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet679_321 _4150__8/I _6966_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_310 net679_317/I _6977_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet679_332 net779_451/I _6955_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_343 net429_96/I _6944_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4040_ _7034_/Q _4040_/A2 _4040_/B1 _6736_/Q _4040_/C _4044_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5991_ _7294_/Q _6006_/B1 _5991_/B _7294_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _5324_/A4 _5405_/A2 _6896_/Q _5407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_80_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _5490_/B _5111_/B1 _4873_/B _4873_/C _5463_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6612_ _6612_/A1 _6612_/A2 _6612_/A3 _6611_/Z _6613_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_47__1403_ clkbuf_4_15_0__1403_/Z net779_434/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3824_ _6988_/Q _5750_/A2 hold68/I _5750_/A3 _3856_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6543_ _7163_/Q _6543_/A2 _6566_/A2 _6594_/A3 _6551_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3755_ _7280_/Q _4027_/A2 _4040_/A2 _7038_/Q _3756_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6474_ _7144_/Q _6323_/Z _6334_/Z _7030_/Q _6352_/Z _7152_/Q _6476_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3686_ hold52/I _3981_/A2 _4045_/C2 input27/Z _3688_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _5515_/A1 _5425_/A2 _5218_/B _5310_/B _5508_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput210 _4129_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput232 _7395_/Z mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput221 _7385_/Z mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput243 _4132_/Z mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5356_ _5356_/A1 _5356_/A2 _5437_/A1 _5363_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput254 _7398_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput265 _6943_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput276 _6742_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _5287_/A1 _5287_/A2 _5534_/B1 _5421_/B _5287_/C _5494_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4307_ _4306_/Z hold895/Z _4321_/S _4307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput287 _6951_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput298 _3993_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4238_ hold323/Z hold420/Z _4238_/S _4238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7026_ _7026_/D _7300_/RN _7026_/CLK _7026_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_56_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4169_ _7361_/Q input75/Z _4169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_4_7_0__1403_ clkbuf_4_7_0__1403_/I clkbuf_4_7_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_55_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet629_262 net729_396/I _7025_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_273 _4150__22/I _7014_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_295 net629_301/I _6992_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_284 net629_284/I _7003_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3540_ _4178_/S hold82/Z _3540_/B hold83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_128_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold907 _7058_/Q hold907/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _5210_/A1 _5511_/A1 _5313_/B _5466_/B _5210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3471_ _6726_/Q _6725_/Q _6792_/Q _6727_/Q _3473_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6190_ _7095_/Q _6290_/A2 _6293_/A2 _7079_/Q _6192_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5141_ _5162_/A2 _5177_/B1 _4751_/B _5214_/A4 _5406_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_123_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _5320_/A1 _5301_/B _5374_/B _5228_/A2 _5375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4023_ _6861_/Q _4023_/A2 _4023_/B1 _6954_/Q _4025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _6805_/Q _6807_/Q _7290_/Q _5974_/B _5975_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4925_ _5425_/A2 _5413_/A2 _5218_/B _5310_/B _4926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4856_ _5417_/C _5193_/A1 _5359_/A2 _4876_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_176_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3807_ _7101_/Q _4006_/B1 _4008_/A2 _7093_/Q _4009_/B1 _7109_/Q _3809_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4787_ _4694_/B _4456_/Z _4787_/B _4789_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_118_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ hold53/I _6315_/Z _6354_/Z _7218_/Q _6530_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3738_ _3738_/A1 _3738_/A2 _3743_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6457_ _6457_/A1 _6456_/Z _6458_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3669_ _3868_/A1 _5576_/A2 _5750_/A4 _4402_/A3 _4045_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_69_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5408_ _5262_/B _5408_/A2 _5408_/B _5409_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6388_ _6388_/A1 _6388_/A2 _6393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5339_ _5339_/A1 _5473_/B _5473_/C _5142_/C _5142_/B _5405_/A1 _5340_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_133_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7009_ hold30/Z _7300_/RN _7009_/CLK hold29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_28_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7322_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30__1403_ clkbuf_4_14_0__1403_/Z net429_55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_110__1403_ net779_410/I net829_483/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_93__1403_ clkbuf_4_1_0__1403_/Z net679_334/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_166_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet429_78 net429_89/I _7209_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_56 net429_59/I _7231_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_67 net429_67/I _7220_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet429_89 net429_89/I _7198_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ _4832_/A1 _4710_/A2 _4839_/A3 _4839_/A2 _5291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5690_ hold99/Z hold542/Z _5695_/S _5690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _4693_/B _5172_/A1 _5060_/B _4641_/C _5250_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_156_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4572_ _5296_/A3 _4691_/C _4751_/B _4518_/Z _5065_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_116_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7360_ _7360_/D _6712_/Z _7364_/CLK _7360_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_183_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold715 _7269_/Q hold715/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_155_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6311_ _7298_/Q _7299_/Q _6540_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_116_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7291_ _7291_/D _7322_/RN _7319_/CLK _7291_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3523_ _6881_/Q hold31/Z _3523_/B _3523_/C hold185/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xhold737 _7131_/Q hold737/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold704 _6847_/Q hold704/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold726 _5706_/Z _7074_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold748 _5928_/Z _7268_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3454_ _6795_/Q _6794_/Q _6792_/Q _3464_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold759 _5829_/Z _7181_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6242_ hold29/I _6295_/B1 _6292_/A2 _7017_/Q _6244_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ _6806_/Q _6173_/A2 _6173_/A3 _6173_/B _6174_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xnet829_468 _4150__3/I _6759_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_479 net829_482/I _6748_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_457 net829_457/I _6770_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3385_ hold93/I _3385_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5124_ _5440_/A2 _5280_/B _5534_/B1 _5308_/B _5124_/C _5128_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5055_ _5320_/C _6894_/Q hold31/I _5225_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4006_ _7074_/Q _4006_/A2 _4006_/B1 _7098_/Q _4007_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5957_ _6017_/A3 _5957_/A2 _5959_/A2 _5954_/B _7286_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4908_ _5417_/C _5416_/A2 _5475_/A2 _5466_/A2 _4910_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5888_ hold50/Z hold482/Z _5890_/S _5888_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4839_ _5440_/B1 _4839_/A2 _4839_/A3 _4839_/A4 _4842_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_107_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6509_ _6613_/A2 _6503_/Z _6508_/Z _6510_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold31 hold31/I hold31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold20 hold20/I hold20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_188_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold53 hold53/I hold53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold64 hold64/I hold64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold42 hold42/I hold42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold97 hold97/I hold97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_90_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold75 hold75/I hold75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold86 hold86/I hold86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _6860_/D _7325_/CLK _6860_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ hold358/Z hold99/Z _5817_/S _5811_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _6791_/D _7359_/RN _6791_/CLK _6791_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5742_ hold363/Z hold897/Z _5749_/S _7106_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5673_ hold79/Z hold304/Z _5677_/S _5673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4624_ _5421_/C _5461_/A4 _5534_/A2 _5322_/A2 _4630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4555_ _4693_/B _5310_/B _5199_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold501 _7248_/Q hold501/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7343_ _7343_/D _6697_/Z _7364_/CLK _7343_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
Xhold545 _5593_/Z _6974_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3506_ _3421_/B _7368_/Q _3507_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold523 _7015_/Q hold523/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold534 _4247_/Z _6777_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold512 _6908_/Q hold512/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7274_ _7274_/D _7286_/RN _7274_/CLK _7274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold567 _7182_/Q hold567/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4486_ _5382_/A1 _5382_/A2 _5252_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xhold556 _7068_/Q hold556/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold578 _4298_/Z _6813_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6225_ _5951_/B _6614_/B _7309_/Q _6226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3437_ _7368_/Q _3437_/I1 _3448_/S _7368_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold589 _4296_/Z _6812_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3368_ _7151_/Q _3368_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6156_ _6156_/A1 _6156_/A2 _6265_/C _6157_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _5107_/A1 _5492_/A1 _5269_/A1 _5107_/A4 _5109_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_100_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _7293_/Q _6074_/Z _6087_/B _6087_/C _6090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5038_ _5038_/A1 _5038_/A2 _5038_/A3 _5038_/A4 _5038_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_72_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6989_ _6989_/D _7322_/RN _6989_/CLK _6989_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_53_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput110 wb_adr_i[23] _4929_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_150_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput132 wb_dat_i[13] _6657_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput154 wb_dat_i[4] _6654_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput121 wb_adr_i[4] _4694_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput143 wb_dat_i[23] _6666_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput165 wb_stb_i _4103_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_189_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_401 net779_430/I _6835_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ hold323/Z hold598/Z _4346_/S _4340_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4271_ hold711/Z _4178_/Z _4285_/S _4271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6010_ _6010_/A1 _6599_/A2 _6807_/Q _6011_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6912_ _6912_/D input75/Z _6912_/CLK _6912_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6843_ hold66/Z _7300_/RN _6843_/CLK hold65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3986_ _5808_/A4 _4402_/A4 _3986_/A3 _5872_/A3 _4023_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6774_ _6774_/D _7359_/RN _6774_/CLK _6774_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5725_ hold323/Z hold735/Z _5731_/S _5725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5656_ hold59/Z _7030_/Q hold8/Z hold60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _5239_/A3 _4607_/A2 _4607_/A3 _4634_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_163_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold320 _7124_/Q hold320/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5587_ hold812/Z hold323/Z _5587_/S _6969_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4538_ _4751_/B _4691_/C _5180_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold342 _7231_/Q hold342/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold331 _7163_/Q hold331/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7326_ _7326_/D _7331_/CLK _7326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold353 _4259_/Z _6785_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7257_ _7257_/D _7315_/RN _7257_/CLK _7257_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4469_ _4762_/A4 _5162_/A2 _4751_/B _3402_/I _5172_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold375 _6764_/Q hold375/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold386 _5839_/Z _7190_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold364 _4258_/Z _6784_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6208_ _7162_/Q _6295_/A2 _6294_/B1 _7226_/Q _6209_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold397 _4208_/Z _6748_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7188_ _7188_/D _7243_/RN _7188_/CLK _7188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6139_ _7109_/Q _7231_/Q _7293_/Q _6139_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3840_ _7262_/Q _4017_/A2 _4017_/B1 input63/Z _3841_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3771_ _7144_/Q _3771_/A2 _4012_/A2 _7200_/Q _3776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _4787_/B _5510_/A2 _5533_/A3 _4693_/B _5511_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_12_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6490_ _7209_/Q _6316_/Z _6338_/Z _7079_/Q _6493_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5441_ _5384_/B _5450_/A1 _5441_/A3 _5441_/A4 _5480_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5372_ _5373_/A1 _5373_/A2 _5373_/A3 _5373_/A4 _5372_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7111_ hold97/Z _7315_/RN _7111_/CLK hold96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4323_ hold363/Z hold665/Z _4328_/S _6825_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7042_ _7042_/D _7315_/RN _7042_/CLK _7042_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_87_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4254_ _5578_/B _5808_/A2 _5581_/A3 _5872_/A4 _4256_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4185_ hold79/Z hold494/Z _4193_/S _4185_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6826_ _6826_/D input75/Z _6826_/CLK _6826_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _6757_/D input75/Z _6757_/CLK _6757_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ hold99/Z hold555/Z _5713_/S _7076_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3969_ _7373_/I _5732_/A4 _5891_/A3 _5566_/A1 _4046_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6688_ input75/Z _7012_/Q _4069_/C _6688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_136_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5639_ hold50/Z hold523/Z _5639_/S _7015_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold150 _7049_/Q hold150/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold161 _5772_/Z _7133_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7309_ _7309_/D _7322_/RN _7322_/CLK _7309_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_2_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold183 hold183/I hold183/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold194 _7168_/Q hold194/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold172 _7217_/Q hold172/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_160_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet679_322 net429_63/I _6965_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_311 net779_431/I _6976_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_344 net779_451/I _6943_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_333 net679_333/I _6954_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _4083_/B _7294_/Q _5991_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _5450_/A2 _5336_/A2 _5401_/A2 _5405_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_17_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _5417_/C _5294_/C _5199_/A3 _5457_/A1 _4873_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_178_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6611_ _6613_/A2 _6611_/A2 _6611_/A3 _6611_/A4 _6611_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3823_ _3868_/A1 _4402_/A1 _4402_/A3 _5750_/A4 _4037_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_32_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ hold27/I _6566_/A2 _6593_/A3 _6594_/A3 _6547_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3754_ _7030_/Q _4046_/A2 _4045_/A2 hold71/I _3756_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_185_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6473_ _7224_/Q _6317_/Z _6354_/Z _7216_/Q _6387_/Z _7062_/Q _6476_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3685_ _6734_/Q _3914_/B1 _4020_/A2 _7242_/Q _3688_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput200 _4123_/ZN mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5424_ _5439_/A1 _5424_/A2 _5424_/B _5424_/C _5427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_173_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput233 _7396_/Z mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput211 _7379_/Z mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput222 _7386_/Z mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput244 _7378_/Z mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5355_ _5355_/A1 _5355_/A2 _5437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput266 _6944_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput277 _6743_/Q pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput255 _4154_/I pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5286_ _5457_/A1 _5286_/A2 _5268_/B _5286_/A4 _5287_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_160_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4306_ hold708/Z _4178_/Z _4320_/S _4306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput288 _6952_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput299 _4162_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7025_ hold14/Z _7300_/RN _7025_/CLK _7025_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4237_ hold363/Z hold459/Z _4238_/S _4237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7341_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _7362_/Q input75/Z _4168_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4099_ _4099_/A1 _4099_/A2 _4099_/A3 _4103_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _6809_/D _7300_/RN _6809_/CLK _6809_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_252 net429_71/I _7035_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet629_263 net629_296/I _7024_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_285 net779_427/I _7002_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_274 net729_389/I _7013_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_53__1403_ net579_205/I net579_240/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_296 net629_296/I _6991_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold908 _7082_/Q hold908/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_155_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3470_ input58/Z _7356_/Q _3470_/S _7356_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5140_ _5238_/B1 _5497_/A2 _5140_/B _5263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _5445_/B1 _5238_/B1 _5071_/B _5071_/C _5073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4022_ input52/Z _4287_/A1 _4022_/B1 _6913_/Q _4022_/C _4025_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5973_ _6302_/A1 _6807_/Q _6268_/A1 _5974_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4924_ _5525_/A1 _5320_/A2 _4924_/B _4924_/C _4926_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_21_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _5310_/B _5306_/C _5196_/B1 _4694_/B _4889_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_60_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4786_ _4693_/B _5460_/A2 _5040_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_138_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ _7077_/Q _4006_/A2 _3916_/B1 _7069_/Q _4010_/B1 _7117_/Q _3819_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6525_ _6521_/Z _6525_/A2 _6525_/A3 _6525_/A4 _6537_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3737_ _4045_/B1 _3736_/Z input49/Z _4285_/S _3738_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150__2 _4150__3/I _7359_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _6613_/A2 _6456_/A2 _6456_/A3 _6456_/A4 _6456_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3668_ _3548_/B _3521_/Z _3884_/A1 _3556_/B _5576_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5407_ _5407_/A1 _5407_/A2 _5407_/B _5407_/C _5408_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6387_ _6387_/A1 _6387_/A2 _7294_/Q _6540_/A4 _6387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3599_ _3906_/A1 _3910_/A1 _3509_/Z _5808_/A3 _4006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5338_ _5326_/C _5338_/A2 _4953_/Z _5396_/B1 _5474_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_161_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5269_ _5269_/A1 _5269_/A2 _5351_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7008_ hold75/Z _7300_/RN _7008_/CLK hold74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_28_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet429_79 net429_81/I _7208_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_57 net429_57/I _7230_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_68 net429_97/I _7219_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4640_ _5236_/A4 _5320_/A1 _5309_/B _5441_/A3 _4643_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ _5417_/A2 _5296_/A3 _5457_/A1 _5344_/C _4577_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_128_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6310_ _6594_/A3 _6387_/A1 _6387_/A2 _6337_/A4 _6310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xhold716 _5929_/Z _7269_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7290_ _7290_/D _7322_/RN _7322_/CLK _7290_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3522_ _6881_/Q hold31/Z _3523_/C _3554_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold727 _7067_/Q hold727/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold705 _4348_/Z _6847_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold749 _6773_/Q hold749/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6241_ _7097_/Q _6290_/A2 _6289_/A2 hold88/I _6291_/C1 _7001_/Q _6244_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold738 _5770_/Z _7131_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3453_ _3453_/A1 _4095_/A1 _7364_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _6806_/Q _7306_/Q _6173_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5123_ _5123_/A1 _5526_/A1 _5123_/A3 _5361_/A4 _5124_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet829_458 net429_64/I _6769_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_469 net429_74/I _6758_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3384_ hold90/I _3384_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _5054_/A1 _5054_/A2 _5054_/B _6921_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ _4005_/A1 _4005_/A2 _4005_/A3 _4008_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _5952_/B _6017_/A3 _6808_/Q _6806_/Q _5959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5887_ hold59/Z hold315/Z _5890_/S _5887_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4907_ _4698_/C _5417_/C _5416_/A2 _5466_/A2 _4910_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4838_ _4838_/A1 _5498_/B _4838_/A3 _4842_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_166_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4769_ _5283_/A2 _5268_/B _5270_/A2 _5473_/A2 _4770_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_153_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6508_ _6508_/A1 _6508_/A2 _6508_/A3 _6508_/A4 _6508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_162_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6439_ _6439_/A1 _6439_/A2 _6444_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold21 hold21/I hold21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold10 hold10/I hold10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold32 hold32/I hold32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold65 hold65/I hold65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold54 hold54/I hold54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold43 hold43/I hold43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold98 hold98/I hold98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold76 hold76/I hold76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold87 hold87/I hold87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5810_ hold808/Z hold323/Z _5817_/S _7165_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6790_ _6790_/D _7359_/RN _6790_/CLK _6790_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ _5891_/A1 _5741_/A2 _5759_/A3 _5891_/A4 _5749_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_62_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ hold99/Z hold486/Z _5677_/S _5672_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _4623_/A1 _4623_/A2 _4623_/A3 _4630_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4554_ _4694_/B _4787_/B _5184_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_129_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold502 _5905_/Z _7248_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7342_ _7342_/D _6696_/Z _7364_/CLK _7342_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_7273_ _7273_/D _7315_/RN _7273_/CLK _7273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold535 _6964_/Q hold535/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3505_ _4178_/S hold6/Z _3505_/B _3556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold524 _7055_/Q hold524/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold513 _4419_/Z _6908_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4485_ _4482_/Z _4485_/A2 _4447_/Z _4485_/A4 _5382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold568 _5830_/Z _7182_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold546 _7391_/I hold546/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold557 _7084_/Q hold557/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6224_ _6224_/A1 _6224_/A2 _6806_/Q _7308_/Q _6226_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold579 _7377_/I hold579/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3436_ _6795_/Q _3426_/B _3436_/A3 _3436_/B _3437_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3367_ _3367_/I _5803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6155_ _7038_/Q _6295_/A2 _6289_/B1 _7022_/Q _6156_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _5267_/B _5356_/A1 _5107_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6086_ _7293_/Q _6086_/A2 _6086_/B1 _6086_/B2 _6087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5037_ _5406_/A1 _4796_/Z _5336_/A2 _5401_/A2 _5038_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6988_ _6988_/D _7322_/RN _6988_/CLK _6988_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5939_ hold99/Z hold499/Z _5944_/S _5939_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput111 wb_adr_i[24] _4101_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput100 wb_adr_i[14] _4443_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput122 wb_adr_i[5] _4787_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput144 wb_dat_i[24] _6637_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput133 wb_dat_i[14] _6661_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput155 wb_dat_i[5] _6658_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput166 wb_we_i _6673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_64_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _4285_/S _4269_/Z _4305_/B1 _4402_/A1 _4305_/C _4286_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_97_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _6911_/D input75/Z _6911_/CLK _6911_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _6842_/D _7300_/RN _6842_/CLK _6842_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3985_ input43/Z _4285_/S _3985_/B1 _6754_/Q _4018_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6773_ _6773_/D _7359_/RN _6773_/CLK _6773_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5724_ hold363/Z hold778/Z _5731_/S _5724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ hold79/Z hold90/Z hold8/Z _7029_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _5061_/A3 _5196_/A1 _4608_/A4 _5305_/B _4613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xhold310 _4305_/C hold310/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5586_ hold881/Z hold363/Z _5587_/S _6968_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7325_ _7325_/D _7325_/CLK _7325_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold332 _7116_/Q hold332/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold343 _5886_/Z _7231_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold321 _5762_/Z _7124_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4537_ _5214_/A4 _5460_/A1 _5295_/B2 _5416_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_2_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold387 _7247_/Q hold387/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4468_ _5214_/A4 _5460_/A1 _5295_/B2 _5322_/A2 _5395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold376 _4229_/Z _6764_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7256_ _7256_/D _7286_/RN _7256_/CLK _7256_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold354 _7064_/Q hold354/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold365 _7132_/Q hold365/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet479_150 net429_89/I _7137_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6207_ hold48/I _6289_/B1 _6291_/C1 _7128_/Q _6209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3419_ _7370_/Q hold81/I _7368_/Q _3416_/Z _3419_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7187_ _7187_/D _7243_/RN _7187_/CLK _7187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold398 _6747_/Q hold398/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6138_ _6138_/A1 _7293_/Q _6142_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4399_ _5891_/A1 _4408_/A1 _5732_/A4 _5550_/A1 _4401_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_58_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6069_ _7051_/Q _6291_/A2 _6289_/B1 _7019_/Q _6294_/A2 _7107_/Q _6074_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ _3770_/A1 _3770_/A2 _3770_/A3 _3770_/A4 _3784_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_158_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _5497_/A2 _5440_/A2 _5440_/B1 _5228_/B _5440_/C _5459_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_145_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _5515_/A1 _5482_/A2 _5482_/C _5371_/C _5373_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _5588_/A1 _6677_/A3 _5863_/A4 hold185/Z hold186/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7110_ _7110_/D _7322_/RN _7110_/CLK _7110_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7041_ hold3/Z _7300_/RN _7041_/CLK _7041_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4253_ hold323/Z hold701/Z _4253_/S _4253_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4184_ hold78/Z _7335_/Q _6881_/Q hold79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_95_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _4144_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _6825_/D input75/Z _6825_/CLK _6825_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6756_ _6756_/D input75/Z _6756_/CLK _6756_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3968_ _6780_/Q _5891_/A2 _4426_/A3 _4024_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5707_ hold323/Z hold713/Z _5713_/S _5707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3899_ _4405_/A3 _4402_/A4 _3986_/A3 _3830_/B _3985_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6687_ input75/Z _7012_/Q _4069_/C _6687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_163_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5638_ hold59/Z hold302/Z _5641_/S _5638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5569_ _5578_/B _5585_/A2 _3830_/B _5581_/A3 _5571_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold151 _5677_/Z _7049_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold162 _7267_/Q hold162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold140 _5881_/Z _7227_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7308_ _7308_/D _7322_/RN _7322_/CLK _7308_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold184 _3565_/C _3523_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold195 _5814_/Z _7168_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold173 _5869_/Z _7217_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7239_ _7239_/D _7315_/RN _7239_/CLK _7239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_13__1403_ net479_128/I net679_317/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_312 net679_317/I _6975_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76__1403_ clkbuf_4_7_0__1403_/Z net679_330/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet679_323 net729_359/I _6964_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_334 net679_334/I _6953_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_345 net679_347/I _6942_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4940_ _5336_/A2 _4991_/B _4963_/A2 _4963_/A3 _5142_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_64_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _5416_/B _5359_/A2 _5417_/C _5417_/B _4873_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6610_ _6914_/Q _6610_/A2 _6610_/B1 _6918_/Q _6787_/Q _6310_/Z _6611_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3822_ _3821_/Z _6933_/Q _3961_/S _6933_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ _7267_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6550_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3753_ _3753_/A1 _4303_/S _4287_/A1 input56/Z _4038_/B1 _7014_/Q _3756_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _6472_/A1 _6472_/A2 _6472_/A3 _6472_/A4 _6472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3684_ _7218_/Q _4028_/A2 _3919_/B1 _6750_/Q _3688_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput201 _4121_/ZN mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ _5423_/A1 _5423_/A2 _5509_/A1 _5512_/A1 _5424_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5354_ _5354_/A1 _5354_/A2 _5354_/A3 _5355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput234 _4126_/Z mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput212 _7380_/Z mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput223 _7387_/Z mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _4320_/S _4269_/Z _4305_/B1 _4305_/B2 _4305_/C _4321_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
Xoutput245 _4131_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput256 _4154_/ZN pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput267 _6938_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5285_ _5279_/Z _5281_/Z _5362_/A1 _5285_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_142_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput289 _6746_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput278 _6728_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7024_ _7024_/D _7322_/RN _7024_/CLK _7024_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4236_ _5550_/A1 _5780_/A3 _5818_/A2 _5891_/A1 _4238_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4167_ _4172_/A1 _6898_/Q _6889_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4098_ _4098_/A1 _4098_/A2 _4099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _6808_/D _7315_/RN _4144_/I1 _6808_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _6739_/D _7243_/RN _6739_/CLK _6739_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_149_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_253 net629_269/I _7034_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet629_275 net779_418/I _7012_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_264 net629_264/I _7023_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_286 net629_286/I _7001_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_297 net629_297/I _6990_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0__1403_ clkbuf_4_2_0__1403_/Z net729_357/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold909 _7196_/Q hold909/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _5070_/A1 _5446_/A1 _5071_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ _4021_/A1 _4021_/A2 _4021_/A3 _4021_/A4 _4035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5972_ _6043_/A1 _6231_/A1 _6302_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_80_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _4751_/B _5228_/B _5322_/A2 _5462_/A2 _5098_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_178_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4854_ _5490_/B _5214_/A4 _5162_/A2 _5180_/B2 _5196_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_60_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4785_ _4694_/B _4456_/Z _4787_/B _4788_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3805_ hold93/I _4041_/A2 _3805_/B _3805_/C _3820_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_119_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6524_ _7096_/Q _6331_/Z _6608_/B1 _7112_/Q _6525_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3736_ _7312_/Q _6960_/Q _6962_/Q _3736_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _7109_/Q _6608_/B1 _6347_/C _7239_/Q _6456_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150__3 _4150__3/I _7358_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3667_ _3554_/B _3523_/B _3509_/Z _3504_/Z _5777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5406_ _5406_/A1 _5039_/Z _5406_/B _5406_/C _5407_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3598_ _4402_/A4 _4402_/A3 _3830_/B _5808_/A3 _3963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6386_ _7123_/Q _6308_/Z _6336_/Z _7099_/Q _6388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5337_ _5337_/A1 _5396_/B1 _5337_/B _5337_/C _5340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5268_ _5416_/B _5405_/A1 _5268_/B _5344_/C _5269_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4219_ hold363/Z hold774/Z _4220_/S _4219_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7007_ _7007_/D _7300_/RN _7007_/CLK _7007_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5199_ _5439_/A1 _5417_/C _5199_/A3 _5306_/C _5464_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_56_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet429_58 _4150__9/I _7229_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_69 net429_93/I _7218_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4570_ _5214_/A4 _5162_/A2 _4751_/B _4691_/C _5457_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3521_ _3519_/Z _3523_/C _3521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_183_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold706 _7083_/Q hold706/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold728 _7059_/Q hold728/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold717 _7099_/Q hold717/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6240_ _6240_/A1 _6240_/A2 _6240_/A3 _6240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xhold739 _6952_/Q hold739/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3452_ _7344_/Q _6792_/Q _3409_/Z _4095_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3383_ _7037_/Q _3383_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6171_ _6302_/A1 _6302_/A2 _6990_/Q _7293_/Q _6173_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _5406_/A1 _5525_/A2 _5130_/B1 _5308_/B _5361_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet829_459 net829_473/I _6768_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5053_ _5053_/A1 _5224_/A1 _5053_/B _5053_/C _5054_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4004_ _7122_/Q _5836_/A3 _5863_/A3 _6677_/A1 _4034_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5955_ _7285_/Q _7286_/Q _6012_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5886_ hold79/Z hold342/Z _5890_/S _5886_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4906_ _4906_/A1 _5196_/B1 _4906_/B _4906_/C _4910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_40_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4837_ _5295_/B2 _5439_/A2 _4691_/C _4995_/A4 _4838_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_21_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ _5283_/A2 _5268_/B _5270_/A2 _5405_/A1 _4770_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_147_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4699_ _4747_/A2 _5462_/A2 _5310_/B _4741_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_107_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6507_ _7119_/Q _6322_/Z _6334_/Z hold57/I _6508_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3719_ _7153_/Q _3981_/A2 _4012_/A2 _7201_/Q _3720_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6438_ _7125_/Q _6308_/Z _6336_/Z _7101_/Q _6439_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6369_ _6760_/Q _6328_/Z _6338_/Z _7074_/Q _6370_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold22 hold22/I hold22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold11 hold11/I hold11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold44 hold44/I hold44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold33 hold33/I hold33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold55 hold55/I hold55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold99 hold99/I hold99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold77 hold77/I hold77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold88 hold88/I hold88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold66 hold66/I hold66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_56_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5740_ hold2/Z hold135/Z _5740_/S _5740_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ hold323/Z hold793/Z _5677_/S _5671_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ _5322_/A2 _5417_/C _5416_/C _5196_/B2 _4623_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7341_ _7341_/D _7341_/RN _7341_/CLK _7341_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_175_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4553_ _4702_/B _5305_/B _5510_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_129_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold514 _7206_/Q hold514/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4484_ _4482_/Z _4485_/A2 _4447_/Z _4485_/A4 _4488_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xhold503 _7160_/Q hold503/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7272_ _7272_/D _7286_/RN _7272_/CLK _7272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold525 _6914_/Q hold525/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold536 _5580_/Z _6964_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3504_ _3505_/B _3503_/Z _3504_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_143_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold547 _5591_/Z _6972_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold569 _7167_/Q _3366_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6223_ _6806_/Q _6223_/A2 _6224_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3435_ _7368_/Q _3416_/Z _3436_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold558 _6815_/Q hold558/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3366_ _3366_/I _5813_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6154_ _7070_/Q _6292_/B1 _6291_/B1 _7030_/Q _7006_/Q _6295_/B1 _6160_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _5515_/A1 _5228_/A2 _5216_/B _5105_/C _5356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_112_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6085_ _6085_/A1 _6085_/A2 _6085_/A3 _6085_/A4 _6086_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _5324_/A4 _5326_/C _5220_/A3 _5338_/A2 _5450_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6987_ _6987_/D _7315_/RN _6987_/CLK _6987_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5938_ hold323/Z hold600/Z _5944_/S _5938_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5869_ hold50/Z hold172/Z _5871_/S _5869_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 wb_adr_i[15] _4443_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput134 wb_dat_i[15] _6665_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput123 wb_adr_i[6] _4702_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xinput145 wb_dat_i[25] _6641_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput112 wb_adr_i[25] _3350_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput156 wb_dat_i[6] _6662_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _6926_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _6910_/D _7359_/RN _6910_/CLK _6910_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _6841_/D _7300_/RN _6841_/CLK _6841_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ input36/Z _4303_/S _4320_/S input71/Z _4018_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6772_ _6772_/D _7359_/RN _6772_/CLK _6772_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ _5891_/A1 _5741_/A2 _5759_/A3 _5732_/A4 _5731_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_176_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ hold99/Z hold300/Z hold8/Z _7028_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _5061_/A3 _4608_/A4 _5305_/B _5241_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xhold311 _5641_/S _5639_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5585_ _5578_/B _5585_/A2 _5808_/A3 _5808_/A4 _5587_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7324_ _7324_/D _7325_/CLK _7324_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold300 _7028_/Q hold300/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold333 _5753_/Z _7116_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold322 _7346_/Q hold322/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4536_ _3399_/I _5162_/A2 _4751_/B _5461_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold344 _6836_/Q hold344/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold377 _7207_/Q hold377/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7255_ _7255_/D _7315_/RN _7255_/CLK _7255_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4467_ _4762_/A4 _5162_/A2 _4995_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xhold355 _5694_/Z _7064_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold366 _5771_/Z _7132_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold388 _5904_/Z _7247_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7186_ _7186_/D _7286_/RN _7186_/CLK _7186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6206_ _6766_/Q _6292_/A2 _6290_/B1 _7170_/Q _6209_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3418_ hold81/I _7368_/Q _3416_/Z _3418_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xhold399 _4207_/Z _6747_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet479_140 net479_145/I _7147_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_151 net479_151/I _7136_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4398_ hold323/Z hold733/Z _4398_/S _4398_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3349_ _4792_/B _4711_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_6137_ _6137_/A1 _6137_/A2 _6137_/A3 _6141_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ _7091_/Q _6290_/A2 _6293_/B1 _7059_/Q _6074_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _5238_/B1 _4796_/Z _5336_/A2 _5336_/A3 _5020_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_73_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36__1403_ clkbuf_4_10_0__1403_/Z net429_81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116__1403_ net779_410/I net679_347/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_99__1403_ net629_288/I net429_86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5370_ _5487_/A1 _5487_/A4 _5487_/A3 _5376_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4321_ _4320_/Z hold550/Z _4321_/S _4321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7040_ _7040_/D _7315_/RN _7040_/CLK _7040_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4252_ hold363/Z hold776/Z _4253_/S _4252_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4183_ hold99/Z hold334/Z _4193_/S _4183_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _6824_/D _7286_/RN _6824_/CLK _6824_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6755_ _6755_/D _7315_/RN _6755_/CLK _6755_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3967_ _7188_/Q _5891_/A3 _5836_/A3 _5891_/A2 _4007_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5706_ hold363/Z hold725/Z _5713_/S _5706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6686_ _7359_/RN _7012_/Q _4069_/C _6686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3898_ _4402_/A4 _3986_/A3 _5581_/A3 _3830_/B _3926_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_164_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5637_ hold79/Z hold259/Z _5641_/S _5637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5568_ _5578_/B hold693/Z _5568_/A3 hold694/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold152 _7211_/Q hold152/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4519_ _5295_/B2 _5322_/A2 _3399_/I _5162_/A2 _5515_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7307_ _7307_/D _7322_/RN _7322_/CLK _7307_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold130 _5843_/Z _7194_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold141 _7242_/Q hold141/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7238_ _7238_/D _7315_/RN _7238_/CLK _7238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5499_ _5499_/A1 _5499_/A2 _5499_/A3 _5499_/A4 _5500_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold163 _5926_/Z _7267_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold185 hold185/I hold185/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold174 _7192_/Q hold174/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold196 _7072_/Q hold196/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7169_ hold73/Z _7243_/RN _7169_/CLK hold72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_302 net779_414/I _6985_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_313 net679_315/I _6974_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0__1403_ clkbuf_3_6_0__1403_/Z net429_73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet679_324 net429_91/I _6963_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_335 net429_95/I _6952_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_346 net679_347/I _6941_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ _5417_/B _4751_/B _5416_/A2 _4691_/C _5111_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_33_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3821_ _6932_/Q _6624_/I0 _3960_/S _3821_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6540_ _7049_/Q _6566_/A2 _6593_/A3 _6540_/A4 _6562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3752_ _3752_/A1 _3752_/A2 _3752_/A3 _3752_/A4 _3752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_173_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3683_ _7000_/Q _3963_/A2 _3683_/B _3703_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6471_ _7200_/Q _6313_/Z _6331_/Z _7094_/Q _6335_/Z _7006_/Q _6472_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_127_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5422_ _5422_/A1 _5422_/A2 _5422_/A3 _5422_/A4 _5512_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput235 _4127_/Z mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ _4691_/C _5490_/B _5353_/A3 _5353_/A4 _5354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput213 _4145_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput224 _7388_/Z mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput202 _3386_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput246 _4130_/Z mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xoutput257 _6948_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput268 _6945_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4304_ hold540/Z _4303_/Z _4304_/S _4304_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5284_ _5287_/A1 _5284_/A2 _5534_/B1 _5309_/B _5284_/C _5362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_141_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput279 _6729_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4235_ hold802/Z hold323/Z _4235_/S _4235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7023_ _7023_/D _7322_/RN _7023_/CLK _7023_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ _6969_/Q input39/Z _4166_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4097_ _4715_/B _4711_/B _4097_/B _5414_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_83_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_82__1403_ clkbuf_4_5_0__1403_/Z net629_281/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _6807_/D _7315_/RN _4144_/I1 _6807_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4999_ _5395_/A1 _5529_/A1 _5529_/B2 _5138_/A2 _5000_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6738_ _6738_/D _7243_/RN _6738_/CLK _6738_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6669_ _4392_/Z _6895_/Q _6888_/Q _6669_/A4 _6670_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_152_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_265 net629_288/I _7022_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_254 net779_427/I _7033_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_276 net729_389/I _7011_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_287 net429_57/I _7000_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_298 net629_298/I _6989_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4020_ _7236_/Q _4020_/A2 _4020_/B1 _7156_/Q _4021_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5971_ _7290_/Q _7289_/Q _6299_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_64_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4922_ _5417_/A2 _5473_/A2 _5217_/B _5344_/C _4924_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_92_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _5417_/C _5416_/A2 _4751_/B _4691_/C _5534_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4784_ _5324_/A3 _5268_/B _5134_/A3 _5283_/A4 _5278_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3804_ _3804_/A1 _3804_/A2 _3804_/A3 _3805_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6523_ _7016_/Q _6329_/Z _6604_/A2 _7170_/Q _6525_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3735_ hold57/I _4046_/A2 _4038_/B1 _7015_/Q _3738_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _7191_/Q _6318_/Z _6325_/Z _7085_/Q _7037_/Q _6312_/Z _6456_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5405_ _5405_/A1 _5405_/A2 _5405_/B _5406_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4150__4 _4150__5/I _7283_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3666_ _7282_/Q _4027_/A2 _4017_/A2 _7266_/Q _3673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6385_ _7043_/Q _6566_/A2 _6593_/A3 _6540_/A4 _6405_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3597_ _3910_/A1 _3509_/Z _3504_/Z _5808_/A3 _4009_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5336_ _4796_/Z _5336_/A2 _5336_/A3 _5529_/A2 _5337_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_142_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _5267_/A1 _5270_/A4 _5267_/B _5355_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7006_ _7006_/D _7300_/RN _7006_/CLK _7006_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4218_ _5550_/A1 _5836_/A3 _5818_/A2 _6677_/A3 _4220_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5198_ _5198_/A1 _5306_/A1 _5198_/B _5200_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4149_ _6881_/Q _4149_/A2 _4149_/B1 _4149_/B2 _4149_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet429_59 net429_59/I _7228_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3520_ hold183/Z _3520_/A2 _6881_/Q _3565_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold707 _5716_/Z _7083_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold718 _5734_/Z _7099_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_3_7_0__1403_ clkbuf_0__1403_/Z clkbuf_3_7_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_115_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold729 _5689_/Z _7059_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3451_ _4112_/A1 _7364_/Q _3453_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3382_ _7045_/Q _6121_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6170_ _6170_/A1 _6170_/A2 _6294_/A2 _6151_/Z _6170_/C _6173_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5121_ _5196_/B2 _5196_/B1 _5121_/B _5278_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _4395_/C _5052_/A2 _5053_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ _7066_/Q _5750_/A4 _5909_/A3 _5750_/A3 _4011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_93_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5954_ _6808_/Q _5964_/A2 _5954_/B _7285_/Q _5957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5885_ hold99/Z hold336/Z _5890_/S _5885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4905_ _4691_/C _5490_/B _5421_/B _5353_/A4 _4906_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_52_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _5359_/A2 _5286_/A2 _5291_/C _5134_/A3 _5498_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_178_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4767_ _5283_/A2 _5268_/B _5270_/A2 _5274_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_146_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _7225_/Q _6317_/Z _6347_/C _7241_/Q _6508_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4698_ _5214_/A4 _5460_/A1 _5294_/B _4698_/C _4773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_107_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3718_ _7185_/Q _4014_/A2 _4040_/B1 _6741_/Q _3720_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6437_ _7117_/Q _6594_/A2 _6594_/A3 _6594_/A4 _6439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3649_ _7081_/Q _4006_/A2 _4006_/B1 _7105_/Q _3658_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6368_ _7252_/Q _6319_/Z _6608_/B1 _7106_/Q _6372_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ _5319_/A1 _5320_/A2 _5319_/B _5319_/C _5347_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6299_ _6920_/Q _6265_/C _6299_/B _6299_/C _6300_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xhold12 hold12/I hold12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold23 hold23/I hold23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold34 hold34/I hold34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold45 hold45/I hold45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold56 hold56/I hold56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold78 hold78/I hold78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold67 hold67/I hold67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold89 hold89/I hold89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_72_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_0_0__1403_ clkbuf_4_1_0__1403_/I net779_410/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_105_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7331_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_187_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ hold363/Z hold867/Z _5677_/S _5670_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4621_ _5417_/C _5417_/A2 _5306_/B _5306_/C _4623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_176_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _7340_/D _7341_/RN _7341_/CLK _7340_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4552_ _5395_/A1 _5252_/A2 _5236_/A4 _5095_/A2 _4582_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold515 _5857_/Z _7206_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4483_ _4959_/A1 _4483_/A2 _4483_/B _5382_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7271_ _7271_/D _7315_/RN _7271_/CLK _7271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_144_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold504 _6996_/Q hold504/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold526 _4428_/Z _6914_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3503_ _4178_/S hold6/Z _3503_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold548 _7279_/Q hold548/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6222_ _6302_/A1 _6302_/A2 _6992_/Q _7293_/Q _6223_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3434_ hold638/Z _6795_/Q _3436_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold559 _4302_/Z _6815_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold537 _7201_/Q hold537/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3365_ _7175_/Q _3365_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6153_ _6152_/Z _6265_/B1 _7289_/Q _7290_/Q _6169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _5291_/B _5268_/B _5134_/A4 _5104_/B1 _5104_/B2 _5269_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_98_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6084_ _7229_/Q _6294_/A2 _6293_/A2 _7197_/Q _6085_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ _5327_/A4 _4927_/Z _4794_/Z _5441_/A4 _5038_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6986_ _6986_/D _7286_/RN _6986_/CLK _6986_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_81_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _4178_/Z _7276_/Q _5944_/S _5937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5868_ hold59/Z hold190/Z _5871_/S _5868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4819_ _4819_/A1 _4819_/A2 _4819_/A3 _4819_/A4 _4823_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5799_ hold910/Z _4178_/Z _5807_/S _7156_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput102 wb_adr_i[16] _4448_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput135 wb_dat_i[16] _6638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput124 wb_adr_i[7] _5305_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput113 wb_adr_i[26] _4098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput157 wb_dat_i[7] _6666_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput146 wb_dat_i[26] _6645_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_59__1403_ net579_205/I net629_299/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6840_ _6840_/D _7300_/RN _6840_/CLK _6840_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _6771_/D _7243_/RN _6771_/CLK _6771_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3983_ _7268_/Q _5936_/A1 hold18/I _5927_/A3 _4022_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5722_ hold2/Z hold88/Z _5722_/S hold89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5653_ hold323/Z hold672/Z hold8/Z _7027_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5584_ hold843/Z hold363/Z _5584_/S _6967_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4604_ _5061_/A3 _5305_/B _5239_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4535_ _4500_/B _5305_/B _4694_/B _4787_/B _5102_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7323_ _7323_/D _7341_/RN _7341_/CLK _7323_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold301 _7142_/Q hold301/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold312 _5636_/Z _7012_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold323 _4180_/Z hold323/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold334 _6730_/Q hold334/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold378 _5858_/Z _7207_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold356 _7208_/Q hold356/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7254_ _7254_/D _7315_/RN _7254_/CLK _7254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4466_ _5305_/B _4452_/Z _4456_/Z _4792_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_132_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold345 _4335_/Z _6836_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold367 _7174_/Q hold367/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet479_130 net829_452/I _7157_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6205_ _7218_/Q _6290_/A2 _6291_/B1 hold52/I _6209_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold389 _7215_/Q hold389/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3417_ _7368_/Q _7367_/Q _7366_/Q _7365_/Q _3426_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xnet479_141 net479_145/I _7146_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4397_ hold363/Z hold817/Z _4398_/S _4397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7185_ _7185_/D _7243_/RN _7185_/CLK _7185_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3348_ _4483_/B _4715_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_112_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6136_ _7199_/Q _6293_/A2 _6292_/B1 _7191_/Q _7175_/Q _6291_/A2 _6137_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6067_ _7075_/Q _6293_/A2 _6291_/B1 _7027_/Q _6074_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5018_ _5482_/A2 _4796_/Z _5336_/A2 _5336_/A3 _5020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_26_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6969_ _6969_/D _7359_/RN _6969_/CLK _6969_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold890 _6758_/Q hold890/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ hold35/Z hold2/Z _4320_/S _4320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4251_ _5891_/A2 _4426_/A3 _6677_/A3 _4253_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_101_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4182_ hold98/Z _7334_/Q _6881_/Q hold99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_68_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6823_ _6823_/D _7322_/RN _6823_/CLK _6823_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6754_ _6754_/D _7315_/RN _6754_/CLK _6754_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3966_ _6907_/Q _5560_/A1 _5780_/A3 _5741_/A2 _4005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5705_ _5891_/A1 _5741_/A2 _5759_/A3 _5780_/A3 _5713_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6685_ _7359_/RN _7012_/Q _4069_/C _6685_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_176_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5636_ hold99/Z _7012_/Q _5639_/S _5636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3897_ _5808_/A4 _4402_/A4 _5581_/A3 _4402_/A3 _3953_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_163_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5567_ _5872_/A4 _5872_/A3 _3830_/C _4178_/Z _5568_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xhold153 _5862_/Z _7211_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4518_ _3399_/I _5162_/A2 _4518_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_5498_ _5515_/A1 _5498_/A2 _5498_/B _5498_/C _5499_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7306_ _7306_/D _7322_/RN _7322_/CLK _7306_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_2_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold120 _5628_/Z _7005_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold131 _7218_/Q hold131/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold142 _5898_/Z _7242_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4449_ _4463_/A1 _4463_/A2 _4463_/A3 _4960_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xclkbuf_leaf_42__1403_ clkbuf_4_15_0__1403_/Z net429_57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold186 hold186/I _4328_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold175 _5841_/Z _7192_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold164 _7193_/Q hold164/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7237_ _7237_/D _7243_/RN _7237_/CLK _7237_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_160_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold197 _7096_/Q hold197/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7168_ _7168_/D _7243_/RN _7168_/CLK _7168_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6119_ _6434_/S _6119_/A2 _6119_/B _7305_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7099_ _7099_/D _7322_/RN _7099_/CLK _7099_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_303 net779_418/I _6984_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_314 net679_315/I _6973_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet679_336 net829_495/I _6951_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_347 net679_347/I _6940_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_325 net679_330/I _6962_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3820_ _3795_/Z _3820_/A2 _3820_/A3 _3819_/Z _6624_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3751_ _7272_/Q _3921_/A2 _4031_/A2 input16/Z _3752_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3682_ _3682_/A1 _3682_/A2 _3682_/A3 _3682_/A4 _3683_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6470_ _7232_/Q _6599_/A2 _6329_/Z _7014_/Q _6338_/Z _7078_/Q _6472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_127_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _5517_/A1 _5421_/A2 _5421_/B _5421_/C _5422_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5352_ _5356_/A1 _5356_/A2 _5492_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput225 _7389_/Z mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput214 _4144_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_99_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput203 _3385_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput236 _7397_/Z mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput258 _6949_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4303_ hold4/Z hold2/Z _4303_/S _4303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput247 _4152_/Z pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_5283_ _5457_/A1 _5283_/A2 _5268_/B _5283_/A4 _5284_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_142_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ _7022_/D _7359_/RN _7022_/CLK _7022_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xoutput269 _6946_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4234_ hold877/Z hold363/Z _4235_/S _4234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _6968_/Q input70/Z _4165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4096_ _4929_/A3 _4929_/A2 _4097_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_82_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6806_ _6806_/D _7322_/RN _7319_/CLK _6806_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_51_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ _4794_/Z _5171_/A2 _5336_/A3 _5342_/A2 _5333_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_11_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _6737_/D _7243_/RN _6737_/CLK _6737_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3949_ input35/Z _4041_/B1 _3949_/B _3949_/C _3950_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_176_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _6668_/I0 _7339_/Q _6668_/S _7339_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5619_ hold79/Z hold325/Z _5623_/S _5619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6599_ _6773_/Q _6599_/A2 _6329_/Z _6862_/Q _6338_/Z _6906_/Q _6601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_277 net429_89/I _7010_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet629_255 net729_396/I _7032_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_266 net629_266/I _7021_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_299 net629_299/I _6988_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet629_288 net629_288/I _6999_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _7290_/Q _7289_/Q _6268_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _4691_/C _5228_/B _5287_/A1 _5218_/B _5469_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_80_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _5417_/C _5475_/A1 _5416_/A2 _5466_/A2 _4910_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_61_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3803_ hold90/I _4046_/A2 _4043_/A2 input29/Z _4047_/B1 _7143_/Q _3804_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4783_ _4691_/C _5287_/A1 _5525_/A2 _5121_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _7234_/Q _6599_/A2 _6324_/Z _7056_/Q _6328_/Z _6766_/Q _6525_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3734_ _3734_/A1 _3734_/A2 _3734_/A3 _3734_/A4 _3743_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6453_ _7255_/Q _6319_/Z _6328_/Z _6763_/Q _6610_/B1 _7271_/Q _6456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3665_ _7024_/Q _4041_/A2 _4045_/A2 _7056_/Q _3673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _5525_/A1 _5039_/Z _5404_/B _5404_/C _5407_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4150__5 _4150__5/I _7282_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _7115_/Q _6594_/A2 _6594_/A3 _6594_/A4 _6388_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3596_ _5750_/A4 _5750_/A3 _3910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5335_ _5323_/C _5323_/B _5406_/A1 _5335_/B _5400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5266_ _5287_/A1 _5322_/A2 _4454_/Z _5133_/B _5270_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4217_ hold323/Z hold659/Z _4217_/S _4217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7005_ _7005_/D _7300_/RN _7005_/CLK _7005_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5197_ _5534_/A2 _5310_/A1 _5197_/B _5419_/C _5198_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_141_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ _4148_/A1 _6964_/Q input67/Z _6881_/Q _4149_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_29_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4079_ _5999_/I0 _6963_/Q _5945_/B _6805_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7325_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold708 _6978_/Q hold708/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold719 _7098_/Q hold719/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_155_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _6727_/Q _6726_/Q _6725_/Q _6792_/Q _4112_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_130_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3381_ _7053_/Q _3381_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _5440_/A2 _5525_/A2 _5534_/B1 _5534_/A2 _5123_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _5051_/A1 _5051_/A2 _5053_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4002_ _6849_/Q _6677_/A2 hold68/I _5557_/A2 _4036_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_77_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5953_ _5952_/B _5965_/A1 _5953_/B _7285_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5884_ hold323/Z hold854/Z _5890_/S _7229_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4904_ _4904_/A1 _4904_/A2 _5312_/C _4906_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_33_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _4835_/A1 _4716_/B _4483_/B _5359_/A2 _5440_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_139_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4766_ _5283_/A2 _5268_/B _5270_/A2 _5433_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_21_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6505_ _7193_/Q _6318_/Z _6610_/B1 _7273_/Q _6508_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3717_ hold96/I _4009_/B1 _4010_/B1 _7119_/Q _3720_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4697_ _4751_/B _4691_/C _4694_/B _4787_/B _4697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_174_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ _7263_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6447_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3648_ _7065_/Q _4009_/A2 _4008_/A2 _7097_/Q hold94/I _4009_/B1 _3658_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6367_ _7090_/Q _6331_/Z _6342_/Z _7244_/Q _6372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3579_ _3554_/B _3523_/B _3509_/Z _3504_/Z _4305_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5318_ _4518_/Z _5475_/A1 _5466_/A2 _5217_/B _5319_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_96_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6298_ _6245_/C _7291_/Q _6771_/Q _7293_/Q _6300_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold13 hold13/I hold13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold35 hold35/I hold35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5249_ _5244_/Z _5246_/Z _5248_/Z _5255_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold46 hold46/I hold46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold24 hold24/I hold24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold79 hold79/I hold79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold68 hold68/I hold68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold57 hold57/I hold57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_19__1403_ clkbuf_4_11_0__1403_/Z net429_90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _4620_/A1 _5240_/A1 _4620_/A3 _5195_/A3 _4623_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_184_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4551_ _5441_/A3 _4523_/C _5368_/A3 _4716_/B _5059_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4482_ _4483_/B _4792_/B _4482_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7270_ _7270_/D _7315_/RN _7270_/CLK _7270_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold505 _5618_/Z _6996_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold516 _7394_/I hold516/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold527 _6913_/Q hold527/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3502_ _3440_/B hold639/Z _4178_/S _3548_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold549 _5940_/Z _7279_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold538 _7392_/I hold538/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6221_ _7293_/Q _6220_/Z _6221_/B _6221_/C _6224_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3433_ hold81/I _3433_/I1 _3448_/S _7369_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6152_ _7046_/Q _7168_/Q _7293_/Q _6152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _5108_/A2 _5440_/A2 _5216_/A2 _5517_/A2 _5267_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3364_ _7183_/Q _3364_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6083_ _7157_/Q _6295_/A2 _6289_/B1 _7141_/Q _6085_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _5220_/A1 _5338_/A2 _5220_/A3 _5162_/A2 _5327_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ hold36/Z _7286_/RN _6985_/CLK hold35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5936_ _5936_/A1 hold7/Z hold32/Z _4305_/C _5944_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_178_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ hold79/Z hold389/Z _5871_/S _5867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4818_ _3399_/I _5287_/A2 _5460_/A1 _4454_/Z _4819_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5798_ _5578_/B _5808_/A2 _5872_/A3 _5872_/A4 _5807_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_182_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4749_ _4829_/A4 _4750_/A3 _4835_/A1 _5102_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_135_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6419_ _7182_/Q _6320_/Z _6325_/Z _7084_/Q _6337_/Z _7068_/Q _6423_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_162_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7399_ _7399_/I _7399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput136 wb_dat_i[17] _6642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput114 wb_adr_i[27] _4099_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput125 wb_adr_i[8] _4105_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput103 wb_adr_i[17] _4448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput147 wb_dat_i[27] _6649_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput158 wb_dat_i[8] _6637_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_6__1403_ clkbuf_4_3_0__1403_/Z net779_438/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_180_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3982_ _6968_/Q _5812_/A1 _5750_/A3 hold68/I _4039_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6770_ _6770_/D _7243_/RN _6770_/CLK _6770_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_94_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5721_ hold38/Z hold203/Z _5722_/S _5721_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5652_ hold363/Z hold724/Z hold8/Z _7026_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5583_ hold762/Z hold323/Z _5584_/S _6966_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4603_ _4603_/A1 _4603_/A2 _4787_/B _4608_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_117_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold302 _7014_/Q hold302/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4534_ _4773_/C _4693_/B _5310_/B _4702_/B _5300_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7322_ _7322_/D _7322_/RN _7322_/CLK _7322_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold313 _7108_/Q hold313/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold324 _5540_/Z _6929_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold335 _4183_/Z _6730_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold357 _5859_/Z _7208_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4465_ _4773_/C _5305_/C _5460_/A2 _4793_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7253_ _7253_/D _7315_/RN _7253_/CLK _7253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_144_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet479_120 net429_64/I _7167_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold368 _5821_/Z _7174_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold346 _6750_/Q hold346/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold379 _7240_/Q hold379/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7184_ _7184_/D _7286_/RN _7184_/CLK _7184_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet479_131 net779_445/I _7156_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6204_ _6204_/A1 _6204_/A2 _6204_/A3 _6204_/A4 _6210_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3416_ _7367_/Q _7366_/Q _7365_/Q _3416_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xnet479_142 net479_151/I _7145_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4396_ _4408_/A1 _4426_/A3 _6677_/A3 _4398_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_131_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3347_ _7299_/Q _6007_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_6135_ _7159_/Q _6295_/A2 _6291_/C1 _7125_/Q _6137_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6066_ _7115_/Q _6265_/C _6299_/B _6299_/C _6087_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _5017_/A1 _5017_/A2 _5020_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6968_ _6968_/D _7359_/RN _6968_/CLK _6968_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_65__1403_ clkbuf_4_7_0__1403_/Z net629_296/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5919_ hold363/Z hold869/Z _5926_/S _5919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6899_ _6899_/D _7359_/RN _6899_/CLK _6899_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold880 _4264_/Z _6788_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold891 _4222_/Z _6758_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_3_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4250_ hold323/Z hold596/Z _4250_/S _4250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4181_ hold323/Z hold797/Z _4193_/S _4181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6822_ _6822_/D _7286_/RN _6822_/CLK _6822_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6753_ _6753_/D _7359_/RN _6753_/CLK _6753_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3965_ _6903_/Q hold83/I _5557_/A2 _4411_/A2 _4011_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3896_ _3523_/B _5808_/A2 _3521_/Z _5808_/A4 _4012_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5704_ hold2/Z _7073_/Q hold84/Z hold85/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6684_ input75/Z _7012_/Q _4069_/C _6684_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5635_ hold323/Z hold730/Z _5639_/S _7011_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5566_ _5566_/A1 hold574/Z _5566_/B hold693/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold110 _4342_/Z _6842_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4517_ _3399_/I _5162_/A2 _5462_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5497_ _5497_/A1 _5497_/A2 _5497_/B1 _5216_/C _5497_/C _5499_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7305_ _7305_/D _7322_/RN _7322_/CLK _7305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold132 _5870_/Z _7218_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold143 _7185_/Q hold143/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold121 _7097_/Q hold121/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4448_ _4448_/A1 _4448_/A2 _4448_/A3 _4448_/A4 _4463_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7236_ _7236_/D _7315_/RN _7236_/CLK _7236_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold154 _7109_/Q hold154/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold176 _7144_/Q hold176/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold165 _5842_/Z _7193_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold187 _4328_/Z _6830_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold198 _5730_/Z _7096_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4379_ hold323/Z hold673/Z _4379_/S _4379_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7167_ _7167_/D _7315_/RN _7167_/CLK _7167_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_58_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _5951_/B _6614_/B _7305_/Q _6119_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _7098_/D _7322_/RN _7098_/CLK _7098_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6049_ _7140_/Q _6289_/B1 _6291_/C1 _7122_/Q _6052_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet679_304 net779_404/I _6983_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet679_315 net679_315/I _6972_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_337 net429_96/I _6950_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_326 net679_330/I _6961_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_348 net829_475/I _6939_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3750_ input30/Z _4043_/A2 _4041_/B1 input7/Z _3752_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3681_ _7064_/Q _4009_/A2 _4037_/A2 _7210_/Q _3682_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5420_ _5412_/Z _5518_/A2 _5463_/A2 _5514_/A2 _5423_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _5105_/C _5497_/B1 _5351_/B _5351_/C _5356_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xoutput226 _7390_/Z mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput215 _4143_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xoutput204 _3384_/ZN mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_57_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput237 _4128_/Z mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5282_ _5282_/A1 _5282_/A2 _5282_/A3 _5432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput259 _6950_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput248 _4169_/Z pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4302_ hold558/Z _4301_/Z _4304_/S _4302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4233_ _5578_/B _5872_/A2 _4405_/A3 _5808_/A4 _4235_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_4_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _7021_/D _7300_/RN _7021_/CLK hold93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4164_ input1/Z input36/Z _4164_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4095_ _4095_/A1 _7345_/Q _4095_/B _6793_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6805_ _6805_/D _7315_/RN _7319_/CLK _6805_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_63_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4997_ _5326_/C _5305_/B _5473_/B _4991_/B _5529_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6736_ _6736_/D _7300_/RN _6736_/CLK _6736_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_176_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3948_ _3948_/A1 _3948_/A2 _3948_/A3 _3948_/A4 _3949_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6667_ _6667_/A1 _6667_/A2 _6668_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ _3556_/B _5808_/A2 _3509_/Z _5581_/A3 _3981_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5618_ hold99/Z hold504/Z _5623_/S _5618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6598_ _6598_/A1 _6598_/A2 _6598_/A3 _6598_/A4 _6607_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5549_ hold265/Z hold59/Z _5549_/S _5549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _6880_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7219_ hold43/Z _7243_/RN _7219_/CLK hold42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet629_256 net729_396/I _7031_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_267 net829_493/I _7020_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_289 net429_63/I _6998_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_278 net629_284/I _7009_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4920_ _3399_/I _5319_/A1 _5228_/B _5218_/B _5508_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_92_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _5417_/C _3399_/I _5460_/A1 _5475_/A1 _5130_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3802_ _7215_/Q _4028_/A2 _4019_/B1 _6948_/Q _4038_/A2 _6989_/Q _3804_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_60_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4782_ _4782_/A1 _4782_/A2 _4782_/A3 _4798_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6521_ _6521_/A1 _6521_/A2 _6521_/A3 _6520_/Z _6521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3733_ _7135_/Q _4046_/B1 _4047_/A2 hold72/I _3734_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _7279_/Q _6610_/A2 _6321_/Z hold93/I _6337_/Z _7069_/Q _6457_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3664_ _3663_/Z _6937_/Q _3961_/S _6937_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5403_ _5503_/A1 _5400_/Z _5404_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4150__6 _4150__6/I _7281_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6383_ _7261_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6396_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3595_ _3868_/A1 hold68/Z _3624_/A2 hold227/Z _4423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5334_ _5529_/A1 _5529_/A2 _5334_/B _5390_/C _5337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5265_ _5501_/A1 _5501_/A2 _5265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5196_ _5196_/A1 _5198_/A1 _5196_/B1 _5196_/B2 _5419_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4216_ hold363/Z hold663/Z _4217_/S _4216_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7004_ _7004_/D _7300_/RN _7004_/CLK _7004_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_56_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4147_ _7302_/Q _6958_/Q _6962_/Q _4147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _7286_/Q _6808_/Q _6017_/A2 _5952_/B _5945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6719_ _7359_/RN _7012_/Q _4069_/C _6719_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold709 _5598_/Z _6978_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3380_ _7061_/Q _3380_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5050_ _5450_/A2 _5327_/A4 _5407_/C _5051_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _6752_/Q hold83/I _5557_/A2 _6677_/A2 _4036_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_77_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _4062_/Z _6806_/Q _5952_/B _5952_/C _5953_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_1_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _5417_/C _5475_/A1 _5416_/A2 _4906_/A1 _5312_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_18_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ hold363/Z hold860/Z _5890_/S _7228_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4834_ _5416_/B _5439_/A2 _4834_/B _5498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xnet529_200 net629_298/I _7087_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4765_ _5214_/A4 _5272_/B _5162_/A2 _4698_/C _4770_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_159_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _7039_/Q _6312_/Z _6610_/A2 _7281_/Q _6508_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3716_ _7225_/Q _3914_/A2 _3919_/B1 _6749_/Q _3720_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4696_ _5462_/A2 _4747_/A2 _4747_/B _4832_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_134_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6435_ _7045_/Q _6566_/A2 _6593_/A3 _6540_/A4 _6443_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3647_ _7073_/Q _3916_/B1 _4010_/A2 hold88/I _7121_/Q _4010_/B1 _3658_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6366_ _7228_/Q _6599_/A2 _6310_/Z _7172_/Q _6372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3578_ _3548_/B _3521_/Z _3884_/A1 _3556_/B _5812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5317_ _5462_/A2 _5319_/A1 _5206_/B _5218_/B _5469_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6297_ _6297_/A1 _6297_/A2 _6297_/A3 _6296_/Z _6297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xhold14 hold14/I hold14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold36 hold36/I hold36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5248_ _5381_/A1 _5381_/A3 _5248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold47 hold47/I hold47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold25 hold25/I hold25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold58 hold58/I hold58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5179_ _5344_/C _5473_/A2 _5344_/B _5405_/A2 _5368_/A2 _5345_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xhold69 hold69/I hold69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4550_ _4641_/C _4787_/B _4694_/B _5172_/A1 _5384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4481_ _4483_/B _4792_/B _4945_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xhold506 _7271_/Q hold506/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold517 _5594_/Z _6975_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3501_ _3421_/B hold638/Z hold639/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold539 _5592_/Z _6973_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold528 _4427_/Z _6913_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6220_ _6220_/A1 _6220_/A2 _6220_/A3 _6219_/Z _6220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3432_ _6795_/Q _3418_/Z _3432_/A3 _3432_/B _3433_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3363_ _7191_/Q _3363_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6151_ _7110_/Q _7232_/Q _7293_/Q _6151_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _5102_/A1 _5268_/B _5134_/A4 _5473_/A2 _5102_/B2 _5492_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_112_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ _6245_/B _6299_/B _7173_/Q _7292_/Q _6085_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _5238_/B1 _5342_/A2 _4796_/Z _5401_/A2 _5038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6984_ hold92/Z _7286_/RN _6984_/CLK hold91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ hold2/Z hold166/Z _5935_/S _5935_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5866_ hold99/Z hold721/Z _5871_/S _7214_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4817_ _3399_/I _5287_/A2 _5460_/A1 _5180_/B2 _4819_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5797_ hold2/Z _7155_/Q hold33/Z hold34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4748_ _5270_/A2 _5286_/A4 _4750_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ _5214_/A4 _5322_/A2 _4751_/B _5162_/A2 _5416_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_162_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6418_ _6415_/Z _6418_/A2 _6418_/A3 _6418_/A4 _6430_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7398_ _7398_/I _7398_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_25__1403_ clkbuf_4_11_0__1403_/Z _4150__15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6349_ _6348_/Z _6342_/Z _6335_/Z _6608_/B1 _6349_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_115_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_105__1403_ clkbuf_4_1_0__1403_/Z net829_457/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput115 wb_adr_i[28] _4099_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput104 wb_adr_i[18] _4448_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput126 wb_adr_i[9] _4105_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_88__1403_ clkbuf_4_5_0__1403_/Z net479_151/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput137 wb_dat_i[18] _6646_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput159 wb_dat_i[9] _6641_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput148 wb_dat_i[28] _6653_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_69_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _7148_/Q _3981_/A2 _3981_/B1 _6774_/Q _4021_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5720_ hold50/Z hold217/Z _5722_/S _5720_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5651_ _5678_/A2 _5891_/A1 _5759_/A3 _5732_/A4 hold8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_30_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5582_ hold473/Z hold99/Z _5584_/S _5582_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4602_ _4693_/B _5172_/A1 _5060_/B _5380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _4500_/B _5305_/B _4787_/B _5350_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7321_ _7321_/D _7322_/RN _7322_/CLK _7321_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _7252_/D _7315_/RN _7252_/CLK _7252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold303 _5638_/Z _7014_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold314 _5744_/Z _7108_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold325 _6997_/Q hold325/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4464_ _4442_/Z _4444_/Z _4447_/Z _4792_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_172_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold336 _7230_/Q hold336/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6203_ hold53/I _6295_/B1 _6293_/B1 _7186_/Q _6204_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet479_110 net479_145/I _7177_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold347 _4210_/Z _6750_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold369 _6732_/Q hold369/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold358 _7166_/Q hold358/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet479_121 net429_93/I _7166_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7183_ _7183_/D _7286_/RN _7183_/CLK _7183_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4395_ _6888_/Q _4395_/A2 _4395_/B _4395_/C _6881_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3415_ _6792_/Q _3415_/A2 _3448_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet479_143 net429_95/I _7144_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_132 net629_279/I _7155_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3346_ _7298_/Q _6343_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_112_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6134_ _6231_/A1 _6299_/C _7133_/Q _7290_/Q _6137_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _6063_/Z _6065_/A2 _6614_/B _6065_/B _7303_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_85_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _5326_/C _5220_/A3 _4991_/B _5305_/B _5169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_85_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6967_ _6967_/D _7315_/RN _6967_/CLK _6967_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ _5936_/A1 _5927_/A3 hold32/Z _4305_/C _5926_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_41_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6898_ _6898_/D _7341_/RN _6926_/CLK _6898_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_167_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5849_ hold79/Z hold426/Z _5853_/S _5849_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold870 _5919_/Z _7260_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold881 _6968_/Q hold881/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_107_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold892 _7157_/Q hold892/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_107_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4180_ hold322/Z _7333_/Q _6881_/Q _4180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_122_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_71__1403_ net629_288/I net629_272/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6821_ _6821_/D _7322_/RN _6821_/CLK _7380_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3964_ _6905_/Q _5750_/A4 _5750_/A3 _5777_/A2 _4009_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6752_ _6752_/D _7359_/RN _6752_/CLK _6752_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ hold38/Z hold196/Z hold84/Z _7072_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3895_ _4402_/A4 _5581_/A3 _4402_/A3 _3830_/B _4023_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6683_ input75/Z _7012_/Q _4069_/C _6683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5634_ hold363/Z hold831/Z _5639_/S _7010_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7304_ _7304_/D _7322_/RN _7322_/CLK _7304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5565_ hold363/Z hold769/Z _5565_/S _5565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold100 _4341_/Z _6841_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5496_ _5496_/A1 _5528_/A1 _5496_/A3 _5502_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold133 _7125_/Q hold133/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4516_ _5214_/A4 _4751_/B _4691_/C _5417_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold111 _7006_/Q hold111/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold144 _5833_/Z _7185_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold122 _5731_/Z _7097_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4447_ _4448_/A1 _4448_/A2 _4448_/A3 _4448_/A4 _4447_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7235_ _7235_/D _7286_/RN _7235_/CLK _7235_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold166 _7275_/Q hold166/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold155 _5745_/Z _7109_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold177 _7161_/Q hold177/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold188 _6833_/Q hold188/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold199 _7112_/Q hold199/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7166_ _7166_/D _7243_/RN _7166_/CLK _7166_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4378_ hold363/Z hold675/Z _4379_/S _4378_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _6117_/A1 _6117_/A2 _6806_/Q _7304_/Q _6119_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ _6881_/Q _4395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_7097_ _7097_/D _7322_/RN _7097_/CLK _7097_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _6048_/A1 _6048_/A2 _6048_/A3 _6048_/A4 _6058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_74_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet679_305 net779_415/I _6982_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_316 net679_317/I _6971_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_338 net829_483/I _6949_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_327 net679_327/I _6960_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_349 net779_451/I _6938_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ _7104_/Q _4006_/B1 _4012_/A2 _7202_/Q _3682_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput216 _7381_/Z mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5350_ _4693_/B _5350_/A2 _5359_/A2 _5268_/B _5351_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xoutput205 _3383_/ZN mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput238 _4119_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5281_ _5282_/A1 _5282_/A2 _5282_/A3 _5281_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_142_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput227 _7391_/Z mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4301_ hold40/Z hold38/Z _4303_/S _4301_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput249 _4151_/Z pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4232_ hold2/Z hold113/Z _4232_/S _4232_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7020_ _7020_/D _7243_/RN _7020_/CLK _7020_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_114_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ _4128_/S input63/Z _4163_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4094_ _4094_/A1 _4094_/A2 _6808_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ _4996_/A1 _4996_/A2 _4996_/A3 _5000_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6804_ _6804_/D _7359_/RN _6804_/CLK _7388_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6735_ _6735_/D _7300_/RN _6735_/CLK _6735_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3947_ _7173_/Q _4024_/A2 _3947_/B1 _7003_/Q _3947_/C1 _6883_/Q _3948_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_51_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6666_ _6896_/Q _6666_/A2 _6666_/B1 _6666_/B2 _6667_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3878_ _6777_/Q _5560_/A1 _5732_/A4 _5891_/A2 _3952_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6597_ _6757_/Q _6315_/Z _6316_/Z _6785_/Q _6598_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5617_ hold323/Z hold690/Z _5623_/S _6995_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ hold257/Z hold79/Z _5549_/S _5548_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _5478_/Z _5479_/A2 _5479_/A3 _5479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_3_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7218_ _7218_/D _7243_/RN _7218_/CLK _7218_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_257 net779_427/I _7030_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_268 net679_334/I _7019_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7149_ _7149_/D input75/Z _7149_/CLK _7149_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_171_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_279 net629_279/I _7008_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _5461_/A1 _5517_/A1 _5510_/A2 _5218_/B _4918_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3801_ _7247_/Q _4019_/A2 _4015_/A2 _7045_/Q input46/Z _4285_/S _3804_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4781_ _3399_/I _5525_/A2 _5460_/A1 _5319_/A1 _4782_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _6520_/A1 _6520_/A2 _6520_/A3 _6520_/A4 _6520_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_174_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3732_ _7217_/Q _4028_/A2 _4042_/A2 _6765_/Q _3734_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6451_ _6447_/Z _6451_/A2 _6451_/A3 _6451_/A4 _6458_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _6936_/Q _6628_/I0 _3960_/S _3663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5402_ _5402_/A1 _5337_/C _5402_/A3 _5402_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4150__7 _4150__9/I _7280_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6382_ _7173_/Q _6310_/Z _6321_/Z _7019_/Q _6404_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5333_ _5333_/A1 _5333_/A2 _5333_/B _5390_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3594_ hold227/Z _3624_/A2 _3868_/A1 _5750_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_126_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5264_ _5323_/B _5493_/B _5133_/C _5497_/A1 _5501_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _5195_/A1 _5195_/A2 _5195_/A3 _5197_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4215_ _5936_/A1 _4305_/C hold641/Z hold185/Z _4217_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_68_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7003_ _7003_/D _7300_/RN _7003_/CLK _7003_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_84_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4146_ _7300_/Q _6959_/Q _6962_/Q _4146_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _7287_/Q _7288_/Q _6017_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4979_ _5326_/C _4691_/C _4751_/B _4995_/A4 _5241_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6718_ _7359_/RN _7012_/Q _4069_/C _6718_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_20_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _6898_/Q _6649_/A2 _6649_/B1 _6897_/Q _6651_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4000_ _6928_/Q _3561_/B _5909_/A2 _5777_/A2 _4025_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_120_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _6808_/Q _6806_/Q _6807_/Q _5951_/B _5961_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_65_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _4698_/C _5417_/C _5416_/A2 _4906_/A1 _4904_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_80_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5882_ _4305_/C _5882_/A2 hold32/Z _5891_/A4 _5890_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_34_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _5216_/C _5138_/B _5439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xnet529_201 net579_217/I _7086_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4764_ _4764_/A1 _4764_/A2 _4764_/A3 _5354_/A3 _4770_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6503_ _6503_/A1 _6503_/A2 _6503_/A3 _6503_/A4 _6503_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3715_ _3715_/A1 _3715_/A2 _3715_/A3 _3745_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4695_ _4693_/B _4773_/B1 _4747_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6434_ _6434_/I0 _7315_/Q _6434_/S _7315_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3646_ _7211_/Q _4037_/A2 _4287_/A1 input60/Z _3646_/C _3659_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6365_ _6365_/A1 _6365_/A2 _6364_/Z _6365_/A4 _6365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3577_ _4402_/A4 _5872_/A4 _5872_/A3 _4402_/A3 _4040_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_142_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _5311_/Z _5511_/A2 _5316_/A3 _5319_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6296_ _6296_/A1 _6296_/A2 _6296_/A3 _6296_/A4 _6296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_170_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5247_ _5395_/A1 _5443_/B _5309_/B _5250_/A1 _5381_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold37 hold37/I hold37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_57_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold26 hold26/I hold26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold15 hold15/I hold15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5178_ _5178_/A1 _5406_/B _5144_/Z _5404_/B _5178_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
Xhold59 hold59/I hold59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_69_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold48 hold48/I hold48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _6819_/Q input58/Z _7364_/Q _4129_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_48__1403_ clkbuf_4_15_0__1403_/Z net779_435/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ _3500_/A1 _4114_/B2 _4160_/B _7342_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold518 _7254_/Q hold518/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold507 _5931_/Z _7271_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4480_ _4715_/B _4792_/B _4795_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3431_ _7368_/Q _6795_/Q _3432_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold529 _7079_/Q hold529/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3362_ _7199_/Q _3362_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6150_ _7144_/Q _7293_/Q _6299_/B _6265_/B1 _6169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _5417_/C _5296_/A3 _5416_/B _5324_/A4 _5102_/B2 _5107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6081_ _7131_/Q _6295_/B1 _6291_/C1 _7123_/Q _6292_/B1 _7189_/Q _6085_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5032_ _5032_/A1 _5032_/A2 _5032_/A3 _5032_/A4 _5038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_57_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _6983_/D _7286_/RN _6983_/CLK _6983_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ hold38/Z hold250/Z _5935_/S _5934_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5865_ hold323/Z hold884/Z _5871_/S _7213_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _4691_/C _5287_/A1 _5287_/A2 _4819_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5796_ hold38/Z hold52/Z hold33/Z _7154_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4747_ _5462_/A2 _4747_/A2 _4747_/B _4787_/B _5286_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_135_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _5460_/A1 _5295_/B2 _4691_/C _3399_/I _5497_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6417_ _7198_/Q _6313_/Z _6331_/Z _7092_/Q _6335_/Z _7004_/Q _6418_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7397_ _7397_/I _7397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3629_ _3906_/A1 _5808_/A2 _3509_/Z _5808_/A3 _4042_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_162_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6348_ _6312_/Z _6610_/B1 _6341_/Z _6348_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
Xinput127 wb_cyc_i _4103_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput116 wb_adr_i[29] _4098_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput105 wb_adr_i[19] _4448_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6279_ _6279_/A1 _6279_/A2 _6806_/Q _7310_/Q _6280_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_76_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput149 wb_dat_i[29] _6657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput138 wb_dat_i[19] _6650_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_15_0__1403_ clkbuf_3_7_0__1403_/Z clkbuf_4_15_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_153_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ _6847_/Q _4435_/A1 hold68/I _5557_/A2 _4049_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5650_ _7025_/Q hold2/Z hold13/Z hold14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31__1403_ clkbuf_4_11_0__1403_/Z net429_63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4601_ _4601_/A1 _5237_/A1 _4601_/A3 _4613_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5581_ _5578_/B _5585_/A2 _5581_/A3 _5872_/A4 _5584_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_111__1403_ net779_410/I net429_98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_94__1403_ clkbuf_4_4_0__1403_/Z net429_71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4532_ _4500_/B _5305_/B _5294_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7320_ _7320_/D _7322_/RN _7322_/CLK _7320_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7251_ _7251_/D _7286_/RN _7251_/CLK _7251_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4463_ _4463_/A1 _4463_/A2 _4463_/A3 _4793_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold304 _7045_/Q hold304/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold315 _7232_/Q hold315/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold326 _5619_/Z _6997_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold337 _5885_/Z _7230_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold348 _7048_/Q hold348/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _6245_/B _6299_/B hold46/I _7292_/Q _6204_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3414_ _6792_/Q _3415_/A2 _3423_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xnet479_111 net429_95/I _7176_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold359 _5811_/Z _7166_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4394_ _4393_/Z _6895_/Q _6890_/Q _4395_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7182_ _7182_/D _7286_/RN _7182_/CLK _7182_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_125_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet479_144 net829_498/I _7143_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_133 net479_151/I _7154_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_122 net829_496/I _7165_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3345_ _7296_/Q _6328_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_6133_ _7053_/Q _6291_/A2 _6133_/B _6133_/C _6143_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_98_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6064_ _6302_/A1 _6302_/A2 _6986_/Q _7293_/Q _6065_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _4796_/Z _5336_/A2 _5024_/A4 _5336_/A3 _5017_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_73_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0_0__1403_ clkbuf_0__1403_/Z clkbuf_4_1_0__1403_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6966_ _6966_/D _7286_/RN _6966_/CLK _6966_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ hold2/Z _7259_/Q _5917_/S _5917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6897_ _6897_/D _7341_/RN _7341_/CLK _6897_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_179_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ hold99/Z hold461/Z _5853_/S _5848_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5779_ hold323/Z hold809/Z _5779_/S _5779_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold871 _7236_/Q hold871/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold860 _7228_/Q hold860/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold882 _6772_/Q hold882/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold893 _6782_/Q hold893/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _6820_/D _7322_/RN _6820_/CLK _7379_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3963_ _6994_/Q _3963_/A2 _3963_/B1 _6851_/Q _4013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6751_ _6751_/D _7300_/RN _6751_/CLK _6751_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_50_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3894_ _4405_/A3 _4402_/A4 _5642_/A3 _4402_/A3 _4037_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5702_ hold50/Z hold216/Z hold84/Z _7071_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6682_ input75/Z _7012_/Q _4069_/C _6682_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_176_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5633_ _5669_/A1 _4305_/C hold32/Z _5927_/A3 _5641_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_31_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5564_ _5564_/A1 _5566_/A1 _6677_/A3 _5565_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold101 _7341_/Q hold101/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4515_ _5060_/C _4787_/B _4499_/B _4515_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7303_ _7303_/D _7322_/RN _7322_/CLK _7303_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold123 _7137_/Q hold123/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5495_ _5495_/A1 _5495_/A2 _5496_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold134 _5763_/Z _7125_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold112 _5629_/Z _7006_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4446_ _4463_/A1 _4463_/A2 _4485_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold156 _7121_/Q hold156/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold167 _5935_/Z _7275_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7234_ _7234_/D _7286_/RN _7234_/CLK _7234_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold145 _7153_/Q hold145/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold189 _4332_/Z _6833_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold178 _7117_/Q hold178/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_160_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4377_ _4305_/C _5669_/A1 _5927_/A3 hold185/Z _4379_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_101_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7165_ _7165_/D _7243_/RN _7165_/CLK _7165_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_113_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6116_ _6806_/Q _6116_/A2 _6117_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3328_ _7353_/Q _4113_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_100_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7096_ _7096_/D _7322_/RN _7096_/CLK _7096_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6047_ _7026_/Q _6291_/B1 _6291_/C1 _6994_/Q _6048_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6949_ _6949_/D _7300_/RN _6949_/CLK _6949_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_42_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet679_306 net779_435/I _6981_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet679_317 net679_317/I _6970_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_328 net779_426/I _6959_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_339 net829_483/I _6948_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold690 _6995_/Q hold690/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput217 _7382_/Z mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput206 _6121_/A1 mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput239 _4118_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5280_ _5421_/A2 _5323_/B _5280_/B _5282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput228 _7392_/Z mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4300_ hold579/Z _4299_/Z _4304_/S _4300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4231_ hold38/Z hold248/Z _4232_/S _4231_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4162_ _4132_/S input68/Z _4162_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4093_ _4093_/A1 _7288_/Q _7287_/Q _6808_/Q _4094_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_67_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ _5295_/B2 _5161_/B _3402_/I _4995_/A4 _4996_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6803_ _6803_/D _7359_/RN _6803_/CLK _7387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3946_ _6987_/Q _4038_/A2 _4037_/C1 _6966_/Q _3948_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6734_ _6734_/D _7300_/RN _6734_/CLK _6734_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_32_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6665_ _6898_/Q _6665_/A2 _6665_/B1 _6897_/Q _6667_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ _6969_/Q _5812_/A1 _5750_/A3 hold68/I _3940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5616_ hold363/Z hold900/Z _5623_/S _6994_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6596_ _6759_/Q _6342_/Z _6355_/Z _6779_/Q _6598_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5547_ hold418/Z hold99/Z _5549_/S _5547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5478_ _5478_/A1 _5478_/A2 _5478_/A3 _4671_/B _5478_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_2_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4429_ _5564_/A1 _6677_/A3 _5557_/A2 hold83/Z _4431_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7217_ _7217_/D _7243_/RN _7217_/CLK _7217_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_258 net779_427/I _7029_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7148_ _7148_/D _7243_/RN _7148_/CLK _7148_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_171_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7079_ _7079_/D _7322_/RN _7079_/CLK _7079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet629_269 net629_269/I _7018_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_3_0__1403_ clkbuf_4_3_0__1403_/I clkbuf_4_3_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_145_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4780_ _5268_/B _5305_/B _4839_/A3 _5134_/A3 _5525_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_178_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3800_ _3800_/I _3805_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ _7209_/Q _4037_/A2 _4024_/A2 hold63/I _3734_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6450_ _7175_/Q _6310_/Z _6604_/A2 _7167_/Q _6451_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3662_ _7356_/Q _6794_/Q _3961_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5401_ _4796_/Z _5401_/A2 _5401_/A3 _5529_/B1 _5402_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4150__8 _4150__8/I _7279_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6381_ _6381_/A1 _6381_/A2 _7313_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3593_ _5872_/A2 _3509_/Z _3504_/Z _5872_/A3 _3930_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_62_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5332_ _5330_/B _5396_/B1 _5332_/B _5332_/C _5334_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_161_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5263_ _5263_/A1 _5263_/A2 _5440_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5194_ _5250_/A1 _5410_/B _5194_/B _5194_/C _5195_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4214_ hold323/Z hold670/Z _4214_/S _6753_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7002_ _7002_/D _7300_/RN _7002_/CLK _7002_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4145_ _6822_/Q input93/Z _6967_/Q _4145_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ _5952_/B _7286_/Q _4093_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ _4978_/A1 _4978_/A2 _4978_/A3 _4983_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6717_ _7359_/RN _7012_/Q _4069_/C _6717_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3929_ _7213_/Q _4028_/A2 _4015_/B1 _6759_/Q _3929_/C _3931_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6648_ _6648_/I0 _7334_/Q _6668_/S _7334_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6579_ _6579_/A1 _6579_/A2 _6579_/A3 _6579_/A4 _6579_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_117_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5950_ _4062_/Z _6806_/Q _5952_/C _5954_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _4901_/A1 _5431_/A3 _4901_/A3 _4904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_18_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5881_ hold139/Z hold2/Z _5881_/S _5881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _4832_/A1 _5286_/A2 _5291_/C _4787_/B _5498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4763_ _4691_/C _5287_/A1 _5112_/A1 _4764_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4694_ _4518_/Z _4454_/Z _4694_/B _4755_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_174_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ _7273_/Q _3921_/A2 _4027_/A2 _7281_/Q _3715_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6502_ hold76/I _6323_/Z _6352_/Z _7153_/Q _6503_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6433_ _6433_/A1 _6433_/A2 _6433_/B _6434_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3645_ _3645_/I _3646_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6364_ _6364_/A1 _6364_/A2 _6364_/A3 _6364_/A4 _6364_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3576_ _3504_/Z _3548_/B hold573/Z _3554_/B hold574/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5315_ _5509_/A1 _5509_/A2 _5316_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6295_ _6885_/Q _6295_/A2 _6295_/B1 _6852_/Q _6296_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5246_ _5246_/A1 _5246_/A2 _5246_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold38 hold38/I hold38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold27 hold27/I hold27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold16 hold16/I hold16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold49 hold49/I hold49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5177_ _5439_/A1 _5460_/A3 _5344_/B _5177_/B1 _5473_/A1 _5404_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_68_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4128_ _6828_/Q input81/Z _4128_/S _4128_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ _6724_/Q _3423_/S _4061_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold508 _6762_/Q hold508/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3430_ _7368_/Q _3416_/Z hold81/I _3432_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold519 _7063_/Q hold519/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3361_ _7207_/Q _3361_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5100_ _5100_/A1 _5262_/A1 _5100_/A3 _5260_/B _5225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_98_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6080_ _6268_/A1 _6080_/A2 _6080_/B1 _6268_/B2 _6080_/C _6086_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _5368_/A2 _5473_/B _5326_/C _5338_/A2 _5032_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_111_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_54__1403_ net579_205/I net779_415/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _6982_/D _7322_/RN _6982_/CLK _6982_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_65_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5933_ hold50/Z hold416/Z _5935_/S _5933_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5864_ hold363/Z hold791/Z _5871_/S _5864_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4815_ _4815_/A1 _4815_/A2 _4815_/A3 _4815_/A4 _4819_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5795_ hold50/Z hold145/Z hold33/Z _7153_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4746_ _4829_/A4 _5525_/A1 _4746_/A3 _4835_/A1 _5491_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4677_ _5395_/A1 _5095_/A2 _5384_/B _5384_/C _4681_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_162_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _7396_/I _7396_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6416_ _7230_/Q _6599_/A2 _6338_/Z _7076_/Q _6329_/Z _7012_/Q _6418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3628_ _3548_/B _5872_/A3 _5808_/A2 _3504_/Z _4020_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6347_ _7298_/Q _6007_/B _6347_/B _6347_/C _6351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_89_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3559_ _6881_/Q _4060_/I0 hold11/Z _4402_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_1_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput117 wb_adr_i[2] _3402_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xinput106 wb_adr_i[1] _4762_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_103_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6278_ _5951_/B _6614_/B _7311_/Q _6280_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput128 wb_dat_i[0] _6638_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput139 wb_dat_i[1] _6642_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5229_ _5482_/C _5229_/A2 _5250_/B1 _5369_/A1 _5486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ _5421_/C _5461_/A3 _5320_/A1 _5184_/A2 _4601_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_157_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5580_ _4178_/Z hold535/Z _5580_/S _5580_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4531_ _4773_/C _4702_/B _5461_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7250_ _7250_/D _7286_/RN _7250_/CLK _7250_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4462_ _3399_/I _5305_/B _4452_/Z _4454_/Z _4991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold305 _5673_/Z _7045_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold316 _5887_/Z _7232_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold338 _6763_/Q hold338/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold349 _5676_/Z _7048_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6201_ _7234_/Q _6294_/A2 _6289_/A2 _7210_/Q _6204_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold327 _6733_/Q hold327/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet479_112 net429_98/I _7175_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3413_ _4063_/A1 _3411_/Z _6795_/Q _3415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4393_ _6895_/D _6892_/Q _6891_/Q _6893_/Q _4393_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
Xnet479_145 net479_145/I _7142_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_123 net829_498/I _7164_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_134 net429_93/I _7153_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7181_ _7181_/D _7243_/RN _7181_/CLK _7181_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3344_ _7297_/Q _6355_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_6132_ _6132_/A1 _6132_/A2 _6132_/A3 _6133_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6063_ _6063_/A1 _6063_/A2 _6063_/A3 _6063_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _5014_/A1 _5337_/A1 _5014_/B _5014_/C _5017_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6965_ _6965_/D _7286_/RN _6965_/CLK _6965_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ hold38/Z hold215/Z _5917_/S _7258_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6896_ _6896_/D _7341_/RN _7341_/CLK _6896_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_139_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5847_ hold323/Z hold840/Z _5853_/S _7197_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5778_ hold363/Z hold823/Z _5779_/S _5778_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4729_ _4693_/B _4773_/B1 _4741_/C _4839_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold872 _6818_/Q hold872/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7379_ _7379_/I _7379_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold861 _7164_/Q hold861/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold850 _6810_/Q hold850/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold894 _4255_/Z _6782_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold883 _4240_/Z _6772_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6750_ _6750_/D _7300_/RN _6750_/CLK _6750_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ hold59/Z hold237/Z hold84/Z _7070_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3962_ _3961_/S _6930_/Q _4053_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6681_ input75/Z _7012_/Q _4069_/C _6681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3893_ _4405_/A3 _4402_/A4 _5872_/A4 _4402_/A3 _4043_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_148_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ hold2/Z hold29/Z _5632_/S hold30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5563_ hold363/Z hold784/Z _5563_/S _5563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4514_ _5060_/C _4787_/B _4499_/B _5371_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7302_ _7302_/D _7322_/RN _7322_/CLK _7302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold113 _6767_/Q hold113/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold124 _5776_/Z _7137_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5494_ _5494_/A1 _5494_/A2 _5494_/A3 _5495_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold102 hold102/I _5578_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold135 _7105_/Q hold135/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold146 _7251_/Q hold146/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4445_ _4105_/B _4105_/C input97/Z input96/Z _4463_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_171_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold157 _5758_/Z _7121_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7233_ _7233_/D _7286_/RN _7233_/CLK _7233_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold168 _7395_/I hold168/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold179 _5754_/Z _7117_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7164_ _7164_/D _7243_/RN _7164_/CLK _7164_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4376_ _6628_/I0 _6870_/Q _4376_/S _6870_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6115_ _6302_/A1 _6302_/A2 _6988_/Q _7293_/Q _6116_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_86_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3327_ _7362_/Q _4158_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ hold51/Z _7243_/RN _7095_/CLK _7095_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6046_ _6231_/A1 _7292_/Q _7291_/Q _7290_/Q _6291_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_74_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6948_ _6948_/D _7300_/RN _6948_/CLK _6948_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6879_ _6879_/D _6880_/CLK _6879_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_307 net779_418/I _6980_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_318 net829_455/I _6969_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_329 net779_426/I _6958_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold680 _6999_/Q hold680/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold691 _7022_/Q hold691/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput207 _3381_/ZN mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput218 _7383_/Z mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput229 _7393_/Z mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4230_ hold50/Z hold285/Z _4232_/S _4230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _3961_/S _4161_/A2 _7343_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4092_ _6806_/Q _4092_/A2 _4092_/A3 _4094_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6802_ _6802_/D _7359_/RN _6802_/CLK _7386_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4994_ _4794_/Z _5171_/A2 _5401_/A3 _5336_/A3 _5161_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6733_ _6733_/D _7300_/RN _6733_/CLK _6733_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3945_ _3945_/A1 _3945_/A2 _3945_/A3 _3949_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6664_ _6664_/I0 _7338_/Q _6668_/S _7338_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _5678_/A2 _5827_/A1 _5759_/A3 _5891_/A1 _5623_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3876_ _5808_/A4 _5872_/A2 _3523_/B _3554_/B _4015_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_136_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6595_ _6753_/Q _6308_/Z _6324_/Z _6900_/Q _6336_/Z _6912_/Q _6598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_129_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5546_ hold703/Z hold323/Z _5549_/S _6941_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5477_ _5402_/Z _5477_/A2 _5477_/A3 _5530_/A3 _5504_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_145_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4428_ hold323/Z hold525/Z _4428_/S _4428_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7216_ _7216_/D _7243_/RN _7216_/CLK _7216_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4149_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7147_ hold24/Z _7300_/RN _7147_/CLK _7147_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4359_ _3859_/Z _6855_/Q _4364_/S _6855_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet629_259 net779_427/I _7028_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _7078_/D _7322_/RN _7078_/CLK _7078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6029_ _7034_/Q _6295_/A2 _6290_/A2 _7090_/Q _6035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _7233_/Q _4033_/A2 _4020_/A2 _7241_/Q _3734_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3661_ _3661_/A1 _3661_/A2 _3659_/Z _3661_/A4 _6628_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5400_ _5400_/A1 _5400_/A2 _5454_/A1 _5400_/A4 _5400_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6380_ _6986_/Q _6613_/A2 _6380_/B _6380_/C _6381_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3592_ _3884_/A1 _5872_/A2 _3521_/Z _5872_/A4 _4028_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5331_ _4796_/Z _5336_/A2 _5331_/A3 _5529_/A2 _5332_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_142_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150__9 _4150__9/I _7278_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5262_ _5262_/A1 _5262_/A2 _5262_/A3 _5262_/B _5347_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7001_ _7001_/D _7322_/RN _7001_/CLK _7001_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5193_ _5193_/A1 _5306_/A1 _5193_/B _5193_/C _5194_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ hold363/Z hold669/Z _4214_/S _6752_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4144_ _6823_/Q _4144_/I1 _6965_/Q _4144_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4075_ _4075_/I _6898_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _5295_/B2 _5330_/B _3402_/I _4995_/A4 _4978_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6716_ _7359_/RN _7012_/Q _4069_/C _6716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3928_ _7359_/Q _4028_/B1 _4012_/B1 _6787_/Q _3935_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6647_ _6647_/A1 _6647_/A2 _6648_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3859_ _3859_/A1 _3859_/A2 _3859_/A3 _3859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
X_6578_ _6756_/Q _6315_/Z _6316_/Z _6784_/Q _6579_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ _5529_/A1 _5529_/A2 _5529_/B1 _5529_/B2 _5529_/C _5530_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ _5309_/B _5322_/A2 _5490_/B _5353_/A4 _4901_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5880_ hold433/Z hold38/Z _5881_/S _5880_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _5457_/A1 _5286_/A2 _5291_/C _5134_/A3 _4834_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_2490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4762_ _5460_/A1 _5295_/B2 _3402_/I _4762_/A4 _5473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_159_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4693_ _5214_/A4 _5460_/A1 _4693_/B _4698_/C _4741_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xclkbuf_leaf_14__1403_ net479_128/I net679_315/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6501_ _7135_/Q _6315_/Z _6355_/Z _7161_/Q _6503_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3713_ input68/Z _4303_/S _4041_/B1 input8/Z _3715_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ _6806_/Q _7314_/Q _6433_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_77__1403_ clkbuf_4_5_0__1403_/Z net779_426/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3644_ _7155_/Q _3981_/A2 _4045_/C2 input28/Z _4041_/B1 input10/Z _3645_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_174_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6363_ _7018_/Q _6321_/Z _6329_/Z _7010_/Q _6364_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3575_ _4402_/A4 _5872_/A4 _4402_/A3 _5808_/A3 _4046_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_130_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5314_ _5439_/A1 _5460_/A3 _5217_/B _5314_/B _5509_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6294_ _6916_/Q _6294_/A2 _6294_/B1 _6912_/Q _6296_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5245_ _5395_/A1 _5377_/B _5308_/B _5250_/A1 _5246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold17 hold17/I hold17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold28 hold28/I hold28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5176_ _4796_/Z _5176_/A2 _5401_/A2 _5342_/A2 _5343_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold39 hold39/I hold39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _6826_/Q input78/Z _4128_/S _4127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4058_ _6725_/Q _4058_/A2 _6725_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold509 _4227_/Z _6762_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_167_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3360_ _7215_/Q _3360_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5030_ _5326_/C _5030_/A2 _4789_/B _5338_/A2 _5340_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6981_ _6981_/D _7286_/RN _6981_/CLK _6981_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_1__1403_ clkbuf_4_2_0__1403_/Z net779_430/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5932_ hold59/Z hold479/Z _5935_/S _5932_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _6677_/A3 _5891_/A2 _5863_/A3 _5863_/A4 _5871_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4814_ _3399_/I _5287_/A2 _5460_/A1 _5319_/A1 _5362_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5794_ hold59/Z hold201/Z hold33/Z _7152_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4745_ _5268_/B _5270_/A2 _5324_/A4 _5134_/A3 _4760_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_166_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4676_ _5095_/A2 _5384_/B _5384_/C _5482_/A2 _5478_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_135_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7395_ _7395_/I _7395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6415_ _6415_/A1 _6415_/A2 _6415_/A3 _6415_/A4 _6415_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3627_ _3906_/A1 _3830_/C _3509_/Z _5872_/A3 _4041_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6346_ _6319_/Z _6321_/Z _6334_/Z _6336_/Z _6347_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_115_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3558_ _4402_/A4 _3986_/A3 _5872_/A3 _5642_/A3 _3921_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_1_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput118 wb_adr_i[30] _4104_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput107 wb_adr_i[20] _4792_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_3489_ hold78/I hold98/I _3491_/S _7348_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _6806_/Q _6277_/A2 _6279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput129 wb_dat_i[10] _6645_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5228_ _5515_/A1 _5228_/A2 _5228_/B _5482_/C _5487_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_88_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5159_ _5392_/A2 _5176_/A2 _5159_/B _5159_/C _5160_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_57_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_60__1403_ net429_73/I net629_291/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _5060_/C _4787_/B _4499_/B _5196_/A1 _4587_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_129_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _5214_/A4 _4773_/C _5305_/C _4698_/C _4960_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_144_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold317 _6740_/Q hold317/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold306 _6734_/Q hold306/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold339 _4228_/Z _6763_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7180_ _7180_/D _7315_/RN _7180_/CLK _7180_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6200_ _7202_/Q _6293_/A2 _6292_/B1 _7194_/Q _6204_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold328 _4189_/Z _6733_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3412_ _6727_/Q _6726_/Q _6725_/Q _6794_/Q _4063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet479_102 net429_93/I _7185_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4392_ _6896_/Q _6897_/Q _6898_/Q _6894_/Q _4392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
Xnet479_124 _4150__6/I _7163_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6131_ _7037_/Q _6295_/A2 _6289_/A2 _7085_/Q _6132_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet479_113 net829_493/I _7174_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_146 net829_496/I _7141_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_135 net829_493/I _7152_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _7294_/Q _6337_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_112_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6062_ _7114_/Q _6265_/C _6299_/B _6299_/C _6063_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _5395_/A1 _5005_/Z _5335_/B _5138_/A2 _5014_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6964_ _6964_/D _7359_/RN _6964_/CLK _6964_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5915_ hold50/Z hold243/Z _5917_/S _7257_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6895_ _6895_/D _7341_/RN _7341_/CLK _6895_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5846_ _4178_/Z hold909/Z _5853_/S _7196_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5777_ _5812_/A2 _5777_/A2 _4305_/C _5779_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4728_ _4829_/A4 _4835_/A1 _5268_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_148_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _5295_/B2 _5162_/A2 _3399_/I _5014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_107_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold873 _4309_/Z _6818_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_163_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold840 _7197_/Q hold840/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold862 _7172_/Q hold862/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold851 _4292_/Z _6810_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7378_ _7378_/I _7378_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold895 _6817_/Q hold895/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6329_ _7295_/Q _7294_/Q _6594_/A4 _6540_/A4 _6329_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold884 _7213_/Q hold884/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3961_ _3960_/Z _6931_/Q _3961_/S _6931_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ hold79/Z hold435/Z hold84/Z _7069_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3892_ _6918_/Q hold185/I _5936_/A1 _5927_/A3 _3934_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6680_ input75/Z _7012_/Q _4069_/C _6680_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ hold38/Z hold74/Z _5632_/S hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _5588_/A1 _5891_/A1 _5750_/A2 _7243_/RN _5563_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_156_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4513_ _5061_/A3 _5061_/A4 _5060_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7301_ _7301_/D _7322_/RN _7322_/CLK _7301_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold114 _4232_/Z _6767_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7232_ _7232_/D _7286_/RN _7232_/CLK _7232_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5493_ _5493_/A1 _5525_/A1 _5493_/B _5494_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold125 _7235_/Q hold125/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold103 _5571_/S _5575_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold158 _6834_/Q hold158/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold147 _5908_/Z _7251_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4444_ _4105_/B _4105_/C input97/Z input96/Z _4444_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_132_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold136 _5740_/Z _7105_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7163_ _7163_/D _7315_/RN _7163_/CLK _7163_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold169 _5595_/Z _6976_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_98_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4375_ _6627_/I0 _6869_/Q _4376_/S _6869_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6114_ _7293_/Q _6114_/A2 _6114_/B _6117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3326_ _7363_/Q _3456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7094_ _7094_/D _7243_/RN _7094_/CLK _7094_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6045_ _6231_/A1 _6245_/B _7292_/Q _7290_/Q _6291_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _6947_/D _7300_/RN _6947_/CLK _6947_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6878_ _6878_/D _7325_/CLK _6878_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5829_ hold323/Z hold758/Z _5835_/S _5829_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_308 net779_416/I _6979_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet679_319 net829_455/I _6968_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold681 _7386_/I hold681/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold670 _6753_/Q hold670/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold692 _7373_/I _5566_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput208 _3380_/ZN mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput219 _7384_/Z mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_175_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4160_ _6796_/Q _6793_/Q _4160_/B _4161_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _4091_/A1 _4092_/A3 _4091_/B _6807_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _6801_/D _7359_/RN _6801_/CLK _7385_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4993_ _4794_/Z _5171_/A2 _5401_/A3 _5336_/A3 _5391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_63_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6732_ _6732_/D _7300_/RN _6732_/CLK _6732_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3944_ _6737_/Q _4040_/B1 _4042_/A2 _6761_/Q _3945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6663_ _6663_/A1 _6663_/A2 _6664_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3875_ _4402_/A1 _5750_/A4 _3533_/Z _3986_/A3 _4014_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_177_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5614_ hold2/Z hold77/Z hold69/Z _6993_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _6920_/Q _6594_/A2 _6594_/A3 _6594_/A4 _6598_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_145_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5545_ hold783/Z hold363/Z _5549_/S _6940_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _5476_/A1 _5476_/A2 _5476_/A3 _5476_/A4 _5530_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_160_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ hold363/Z hold527/Z _4428_/S _4427_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7215_ _7215_/D _7359_/RN _7215_/CLK _7215_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7146_ _7146_/D _7300_/RN _7146_/CLK hold48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4358_ _6622_/I0 _6854_/Q _4364_/S _6854_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7077_ _7077_/D _7322_/RN _7077_/CLK _7077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4289_ hold684/Z _4178_/Z _4303_/S _4289_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6028_ _6231_/A1 _6245_/C _6245_/B _7290_/Q _6290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_58_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3660_ _3509_/Z _3523_/B _3554_/B _3556_/B _4426_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_127_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3591_ _7235_/Q _5891_/A4 _5863_/A3 _5827_/A3 _3661_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5330_ _5333_/A1 _5333_/A2 _5330_/B _5452_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _5093_/C _5261_/A2 _5261_/B _5262_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7000_ _7000_/D _7286_/RN _7000_/CLK _7000_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4212_ _6677_/A3 _6677_/A2 _5557_/A2 hold83/Z _4214_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5192_ _5534_/A1 _5410_/B _5216_/A2 _5301_/B _5193_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4143_ _6824_/Q user_clock _6966_/Q _4143_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4074_ _6898_/Q _4115_/A2 _6893_/Q _4075_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_37__1403_ clkbuf_4_14_0__1403_/Z _4150__46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_117__1403_ net779_410/I net779_411/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4976_ _4794_/Z _5171_/A2 _5331_/A3 _4974_/Z _5330_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6715_ _7359_/RN _7012_/Q _4069_/C _6715_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_52_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3927_ _7197_/Q _4012_/A2 _4014_/B1 _6783_/Q _4015_/C1 _6887_/Q _3935_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6646_ _6896_/Q _6646_/A2 _6646_/B1 _6666_/B2 _6647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3858_ _3845_/Z _3858_/A2 _3850_/Z _3858_/A4 _3859_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3789_ _7191_/Q hold18/I _5827_/A1 _5882_/A2 _3809_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6577_ _6758_/Q _6342_/Z _6355_/Z _6778_/Q _6579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5528_ _5528_/A1 _5528_/A2 _5528_/B _5531_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5459_ _5459_/A1 _5459_/A2 _5459_/B1 _5503_/A2 _5472_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7129_ hold16/Z _7243_/RN _7129_/CLK hold15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4830_ _4830_/A1 _4830_/A2 _4830_/A3 _5135_/A1 _4838_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4761_ _5214_/A4 _5322_/A2 _4751_/B _5162_/A2 _5440_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4692_ _4751_/B _4691_/C _4694_/B _4747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3712_ _7039_/Q _4040_/A2 _4287_/A1 input57/Z _4017_/A2 _7265_/Q _3715_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6500_ _7185_/Q _6320_/Z _6337_/Z _7071_/Q _6503_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6431_ _6613_/A2 _6988_/Q _6613_/C _6433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3643_ _3643_/A1 _3643_/A2 _3643_/A3 _3643_/A4 _3643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_146_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6362_ _7196_/Q _6313_/Z _6315_/Z _7130_/Q _6364_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5313_ _5313_/A1 _5313_/A2 _5313_/B _5313_/C _5509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3574_ _4402_/A4 _3986_/A3 _5872_/A4 _5808_/A3 _4027_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_142_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6293_ _6906_/Q _6293_/A2 _6293_/B1 _6902_/Q _6296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5244_ _5378_/A1 _5242_/Z _5378_/A3 _5244_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5175_ _5473_/B _5473_/C _5333_/A1 _5175_/B _5178_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold18 hold18/I hold18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold29 hold29/I hold29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4126_ _6825_/Q input80/Z _4128_/S _4126_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _6726_/Q _4057_/A2 _6726_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _4959_/A1 _4991_/A1 _4795_/B _4964_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6629_ _6673_/A2 _6629_/A2 _6632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20__1403_ clkbuf_4_11_0__1403_/Z net429_67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100__1403_ clkbuf_4_2_0__1403_/Z net779_437/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_83__1403_ clkbuf_4_5_0__1403_/Z net629_279/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6980_ _6980_/D _7286_/RN _6980_/CLK _6980_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ hold79/Z hold506/Z _5935_/S _5931_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ hold2/Z hold152/Z _5862_/S _5862_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4813_ _5286_/A2 _5268_/B _5405_/A1 _5286_/A4 _4815_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5793_ hold79/Z hold256/Z hold33/Z _7151_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4744_ _4829_/A4 _4746_/A3 _4835_/A1 _5267_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4675_ _5295_/B2 _3402_/I _3399_/I _5162_/A2 _5368_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_128_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7394_ _7394_/I _7394_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6414_ _7132_/Q _6315_/Z _6316_/Z _7206_/Q _6415_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3626_ _7017_/Q _5780_/A3 _5678_/A2 _5759_/A3 _3657_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_131_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6345_ _6344_/Z _6330_/Z _6329_/Z _6610_/A2 _6351_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3557_ _3504_/Z _3548_/B _5642_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_163_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6276_ _6302_/A1 _6302_/A2 _6847_/Q _7293_/Q _6277_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput108 wb_adr_i[21] _4483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_3488_ hold58/I hold78/I _3491_/S _7349_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5227_ _5490_/C _5250_/A1 _5250_/B1 _5061_/Z _5373_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput119 wb_adr_i[31] _4104_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _5451_/B _5162_/A2 _5396_/A1 _5330_/B _5172_/A1 _5159_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_84_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109_ _4109_/A1 _6617_/B _6888_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5089_ _5241_/A1 _5206_/B _5241_/B1 _5482_/B _5253_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _4452_/Z _4456_/Z _4949_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_129_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold307 _4191_/Z _6734_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet479_103 _4150__25/I _7184_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4391_ _6896_/Q _6897_/Q _6898_/Q _6894_/Q _4395_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold329 _6837_/Q hold329/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold318 _4199_/Z _6740_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3411_ _6727_/Q _6726_/Q _6725_/Q _6794_/Q _3411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xnet479_125 _4150__6/I _7162_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3342_ _7295_/Q _6387_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_113_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _7093_/Q _6290_/A2 _6295_/B1 _7005_/Q _6132_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet479_114 net679_334/I _7173_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_136 net779_451/I _7151_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet479_147 net829_457/I _7140_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6061_ _6245_/B _6060_/Z _6096_/B1 _7292_/Q _6063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _4794_/Z _5171_/A2 _5336_/A2 _5336_/A3 _5153_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_112_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _6963_/D _7315_/RN _6963_/CLK _6963_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6894_ _6894_/D _7341_/RN _7341_/CLK _6894_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5914_ hold59/Z hold374/Z _5917_/S _7256_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5845_ _4305_/C _5882_/A2 hold32/Z _5927_/A3 _5853_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ hold2/Z hold123/Z _5776_/S _5776_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4727_ _4829_/A4 _4835_/A1 _5105_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_148_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ _5214_/A4 _5460_/A1 _4751_/B _5323_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_107_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold830 _4226_/Z _6761_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput90 spimemio_flash_io2_oeb input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3609_ _3910_/A1 _3509_/Z _3504_/Z _5872_/A3 _3916_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold852 _7114_/Q hold852/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4589_ _5461_/A1 _5421_/C _5461_/A3 _5320_/A1 _4590_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_122_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold841 _7358_/Q hold841/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7377_ _7377_/I _7377_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold863 _6736_/Q hold863/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold896 _4307_/Z _6817_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6328_ _6593_/A3 _6594_/A3 _6355_/A4 _6328_/A4 _6328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold885 _6886_/Q hold885/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_107_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold874 _7188_/Q hold874/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ _6905_/Q _6293_/A2 _6291_/B1 _6882_/Q _6289_/A2 _6907_/Q _6262_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ _6930_/Q _6622_/I0 _3960_/S _3960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _4405_/A3 _4402_/A4 _3986_/A3 _5642_/A3 _4017_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5630_ hold50/Z hold105/Z _5632_/S _5630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ hold363/Z hold615/Z _5561_/S _5561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5492_ _5492_/A1 _5492_/A2 _5492_/A3 _5492_/A4 _5528_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4512_ _4512_/A1 _6897_/Q _5260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7300_ _7300_/D _7300_/RN _7322_/CLK _7300_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold126 _5890_/Z _7235_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7231_ _7231_/D _7315_/RN _7231_/CLK _7231_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold115 _6925_/Q hold115/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold104 _5572_/Z _6959_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold159 _4333_/Z _6834_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4443_ input99/Z input98/Z _4443_/A3 _4443_/A4 _4463_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold148 _6981_/Q hold148/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold137 _7283_/Q hold137/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7162_ _7162_/D _7315_/RN _7162_/CLK _7162_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4374_ _3745_/Z _6868_/Q _4376_/S _6868_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7093_ _7093_/D _7322_/RN _7093_/CLK _7093_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6113_ _6113_/A1 _7293_/Q _7116_/Q _6142_/B2 _6113_/C _6114_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3325_ _7370_/Q _3426_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6044_ _7066_/Q _6292_/B1 _6290_/B1 _7042_/Q _6048_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _6946_/D input75/Z _6946_/CLK _6946_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_26_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6877_ _6877_/D _6880_/CLK _6877_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5828_ hold363/Z hold898/Z _5835_/S _5828_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5759_ _5891_/A1 _6677_/A1 _5759_/A3 _5836_/A3 _5767_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_154_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet679_309 net779_419/I _6978_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold660 _4217_/Z _6755_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold671 _6962_/Q hold671/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold682 _4282_/Z _6802_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold693 hold693/I hold693/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput209 _4138_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4090_ _6387_/A2 _6340_/A1 _7294_/Q _4092_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_49_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _6800_/D _7286_/RN _6800_/CLK _7384_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ _5326_/C _4991_/B _4953_/Z _5305_/B _5529_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_177_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _6731_/D _7300_/RN _6731_/CLK _6731_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_32_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3943_ _3943_/A1 _3943_/A2 _3943_/A3 _3943_/A4 _3943_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6662_ _6896_/Q _6662_/A2 _6662_/B1 _6666_/B2 _6663_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3874_ _6789_/Q _5891_/A2 _5777_/A2 _3937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5613_ hold38/Z _6992_/Q hold69/Z hold70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6593_ _6929_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6601_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5544_ _5578_/B _5585_/A2 _3830_/B _5872_/A3 _5549_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5475_ _5475_/A1 _5475_/A2 _5475_/B _5475_/C _5476_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7214_ _7214_/D _7359_/RN _7214_/CLK _7214_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4426_ hold116/Z _5909_/A2 _4426_/A3 _4305_/C _4428_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_113_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7145_ _7145_/D _7300_/RN _7145_/CLK hold76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4357_ _4051_/Z _6853_/Q _4364_/S _6853_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7076_ _7076_/D _7322_/RN _7076_/CLK _7076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4288_ _5597_/A3 _4435_/A1 _4288_/B _5578_/B _4304_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_104_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6027_ _7292_/Q _7291_/Q _6268_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _6929_/D _7359_/RN _6929_/CLK _6929_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold490 _6739_/Q hold490/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3590_ _3868_/A1 _4305_/B2 _5750_/A4 _3986_/A3 _4033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_114_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _5259_/B _5182_/C _5260_/B _5260_/C _5261_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4211_ hold291/Z hold2/Z _4211_/S _4211_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5191_ _5421_/C _5191_/A2 _5310_/A1 _5300_/A2 _5191_/C _5193_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_96_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4142_ input1/Z _6989_/Q _4142_/B _4142_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4073_ _4073_/I _6897_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4975_ _4794_/Z _5171_/A2 _5331_/A3 _4974_/Z _4975_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3926_ _7149_/Q _3981_/A2 _4023_/A2 _6862_/Q _3926_/C1 _6929_/Q _3936_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6714_ input75/Z _7012_/Q _4069_/C _6714_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_177_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6645_ _6898_/Q _6645_/A2 _6645_/B1 _6897_/Q _6647_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3857_ input54/Z _4287_/A1 _3857_/B _3857_/C _3858_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xnet729_390 net729_396/I _6846_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3788_ _7263_/Q _4017_/A2 _4027_/B1 _7255_/Q _3795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6576_ _6752_/Q _6308_/Z _6324_/Z _6899_/Q _6336_/Z _6911_/Q _6579_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5527_ _5527_/A1 _5527_/A2 _5528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _5407_/B _5458_/A2 _5407_/C _5503_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5389_ _5395_/A1 _5335_/B _5389_/B1 _5529_/B1 _5389_/C _5400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4409_ hold363/Z hold781/Z _4410_/S _4409_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _7128_/D _7322_/RN _7128_/CLK _7128_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7059_ _7059_/D _7322_/RN _7059_/CLK _7059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_46_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_43__1403_ clkbuf_4_14_0__1403_/Z net629_271/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _4760_/A1 _4760_/A2 _4760_/A3 _4764_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4691_ _3399_/I _5162_/A2 _4751_/B _4691_/C _4773_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_119_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3711_ _3711_/A1 _3711_/A2 _3711_/A3 _3711_/A4 _3745_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_186_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _6430_/A1 _6430_/A2 _6430_/A3 _6433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3642_ _7025_/Q _4041_/A2 _4043_/A2 input33/Z _3643_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6361_ _7188_/Q _6318_/Z _6320_/Z _7180_/Q _6364_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ _5312_/A1 _5421_/B _5421_/C _5312_/B2 _5312_/C _5511_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3573_ _3830_/C _3521_/Z _3523_/B _5642_/A3 _4031_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _6862_/Q _6292_/A2 _6292_/B1 _6904_/Q _6296_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _5250_/A1 _5534_/A2 _5250_/B1 _5075_/Z _5378_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5174_ _5326_/C _5333_/A1 _5338_/A2 _5473_/B _5387_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xhold19 hold19/I hold19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_111_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4125_ _4125_/I _4125_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _6727_/Q _4056_/A2 _6727_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_169_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3_0__1403_ clkbuf_0__1403_/Z clkbuf_4_7_0__1403_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_52_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _4995_/A4 _5326_/B _5326_/C _4751_/B _4958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_24_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4889_ _4889_/A1 _5525_/B _4889_/A3 _4889_/A4 _4892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_138_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3909_ _6757_/Q _5560_/A1 _5836_/A3 _6677_/A1 _3951_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6628_ _6628_/I0 _7331_/Q _6628_/S _7331_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ hold25/I _6310_/Z _6321_/Z _7025_/Q _6561_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5930_ hold99/Z hold467/Z _5935_/S _5930_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5861_ hold38/Z hold233/Z _5862_/S _5861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4812_ _5310_/B _4832_/A1 _5286_/A2 _5268_/B _5287_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5792_ hold99/Z hold319/Z hold33/Z _7150_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4743_ _5268_/B _5270_/A2 _5134_/A3 _5108_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_175_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4674_ _5214_/A4 _5460_/A1 _5322_/A2 _4751_/B _5482_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6413_ _7246_/Q _6342_/Z _6355_/Z _7158_/Q _6415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7393_ _7393_/I _7393_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3625_ _4402_/A4 _5642_/A3 _4402_/A3 _5808_/A3 _4038_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6344_ _6324_/Z _6325_/Z _6337_/Z _6338_/Z _6344_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_115_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3556_ _6881_/Q hold21/Z _3556_/B _3556_/C hold22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_1_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6275_ _7293_/Q _6262_/Z _6275_/B _6275_/C _6279_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xinput109 wb_adr_i[22] _4929_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3487_ hold49/I hold58/I _3491_/S _7350_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5226_ _5482_/C _5413_/C _5241_/B1 _5369_/A1 _5231_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _5172_/A1 _5475_/C _5157_/B _5157_/C _5159_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4108_ _4108_/A1 _6888_/Q _6617_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5088_ _5380_/C _5238_/B1 _4591_/C _4499_/B _5091_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _4039_/A1 _4039_/A2 _4039_/A3 _4039_/A4 _4050_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold308 _7143_/Q hold308/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4390_ _6896_/Q _6897_/Q _6898_/Q _5320_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
Xhold319 _7150_/Q hold319/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3410_ _6727_/Q _6726_/Q _6725_/Q _4114_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xnet479_104 _4150__8/I _7183_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3341_ _6807_/Q _4083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_124_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet479_115 net829_498/I _7172_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_126 net429_70/I _7161_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet479_148 net829_455/I _7139_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_137 net629_279/I _7150_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6060_ _7058_/Q _7180_/Q _7293_/Q _6060_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5011_ _5326_/C _5220_/A3 _4991_/B _5305_/B _5335_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _6962_/D _7243_/RN _6962_/CLK _6962_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_47_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5913_ hold79/Z hold383/Z _5917_/S _7255_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6893_ _6893_/D _7341_/RN _6926_/CLK _6893_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5844_ hold2/Z hold44/Z _5844_/S hold45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ hold38/Z hold53/Z _5776_/S hold54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4726_ _5460_/A1 _5295_/B2 _5322_/A2 _4762_/A4 _5324_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _4691_/C _5421_/C _5461_/A4 _5206_/B _5253_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput91 spimemio_flash_io3_do input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3608_ _4305_/B2 _5750_/A4 _3533_/Z _3986_/A3 _4047_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7376_ _7376_/I _7376_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput80 spi_sck input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold820 _6826_/Q hold820/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold853 _5751_/Z _7114_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold831 _7010_/Q hold831/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4588_ _5236_/A4 _5413_/A2 _5353_/A3 _5441_/A3 _4590_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6327_ _7260_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6365_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold842 _6678_/Z _7358_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold864 _4195_/Z _6736_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold875 _7382_/I hold875/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold897 _7106_/Q hold897/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold886 _4403_/Z _6886_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3539_ _6881_/Q hold67/Z _3540_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6258_ _6258_/A1 _6258_/A2 _6258_/A3 _6258_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5209_ _5209_/A1 _5228_/B _5209_/B _5466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _7087_/Q _6289_/A2 _6291_/B1 hold57/I _6192_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0__1403_ clkbuf_4_7_0__1403_/I net629_288/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_121_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _4402_/A4 _3986_/A3 _5581_/A3 _5642_/A3 _4022_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_188_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _5560_/A1 _5732_/A4 _5566_/A1 _5891_/A1 _5561_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5491_ _5491_/A1 _5491_/A2 _5491_/A3 _5492_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_156_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ _4694_/B _4787_/B _5395_/A1 _5380_/C _5382_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_8_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4442_ input99/Z input98/Z _4443_/A3 _4443_/A4 _4442_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_7230_ _7230_/D _7286_/RN _7230_/CLK _7230_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold116 _3561_/B hold116/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold105 _7007_/Q hold105/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold149 _5601_/Z _6981_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold127 _6983_/Q hold127/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold138 _5944_/Z _7283_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _7161_/D _7243_/RN _7161_/CLK _7161_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4373_ _4385_/I0 _6867_/Q _4376_/S _6867_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7092_ _7092_/D _7322_/RN _7092_/CLK _7092_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_112_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6112_ _7293_/Q _6302_/A1 _6302_/A2 _6112_/B _6113_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_86_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6043_ _6043_/A1 _6231_/A1 _6245_/B _7292_/Q _6290_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_58_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6945_ _6945_/D _7300_/RN _6945_/CLK _6945_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _6876_/D _6880_/CLK _6876_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ _5827_/A1 _5863_/A3 _5827_/A3 _5891_/A1 _5835_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_10_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5758_ hold2/Z hold156/Z _5758_/S _5758_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _4832_/A1 _4710_/A2 _4839_/A3 _4839_/A2 _5216_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_148_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5689_ hold323/Z hold728/Z _5695_/S _5689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold650 _7252_/Q hold650/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold661 _6917_/Q hold661/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7359_ _7359_/D _7359_/RN _7359_/CLK _7359_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold672 _7027_/Q hold672/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold694 hold694/I _6956_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold683 _7003_/Q hold683/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _4991_/A1 _4991_/A2 _4991_/B _5336_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_91_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _6730_/D _7300_/RN _6730_/CLK _6730_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_189_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3942_ input21/Z _4045_/C2 _4038_/B1 _7011_/Q _6962_/Q _4045_/B1 _3943_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6661_ _6898_/Q _6661_/A2 _6661_/B1 _6897_/Q _6663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3873_ _6791_/Q _5560_/A1 _5836_/A3 _5891_/A2 _3952_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6592_ _7139_/Q _6593_/A3 _6594_/A3 _6594_/A4 _6611_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5612_ hold50/Z hold212/Z hold69/Z _6991_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5543_ hold323/Z hold651/Z _5543_/S _5543_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _5173_/C _5474_/A2 _5474_/A3 _5477_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_160_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7213_ _7213_/D _7359_/RN _7213_/CLK _7213_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xclkbuf_leaf_7__1403_ clkbuf_4_3_0__1403_/Z net829_455/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4425_ hold323/Z hold604/Z _4425_/S _4425_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4356_ _6893_/Q _7341_/RN _4364_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7144_ _7144_/D _7243_/RN _7144_/CLK _7144_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4287_ _4287_/A1 _5597_/A3 _4435_/A1 _5588_/A1 _4288_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7075_ _7075_/D _7322_/RN _7075_/CLK _7075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6026_ _6043_/A1 _6245_/B _7292_/Q _7289_/Q _6295_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_2107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_450 net779_451/I _6777_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _6928_/D _7359_/RN _6928_/CLK _6928_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _6859_/D _7325_/CLK _6859_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold480 _5932_/Z _7272_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold491 _4198_/Z _6739_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4210_ hold346/Z hold38/Z _4211_/S _4210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5190_ _5190_/A1 _5190_/A2 _5191_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ input1/Z input2/Z _4142_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4072_ _6897_/Q _4115_/A2 _6891_/Q _4073_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ _4788_/B _5040_/A4 _4974_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_149_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6713_ input75/Z _7012_/Q _4069_/C _6713_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_51_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3925_ _7027_/Q _4046_/A2 _4047_/C1 _6916_/Q _3925_/C _3936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6644_ _6644_/I0 _7333_/Q _6668_/S _7333_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet729_380 net429_83/I _6872_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3856_ _3856_/A1 _3856_/A2 _3857_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xnet729_391 net779_423/I _6845_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6575_ _6575_/A1 _6575_/A2 _6575_/A3 _6575_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3787_ _3786_/Z _6934_/Q _3961_/S _6934_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5526_ _5526_/A1 _5526_/A2 _5526_/A3 _5526_/A4 _5527_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ _5457_/A1 _5460_/A3 _5344_/B _5457_/B _5459_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_106_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _4408_/A1 _6677_/A2 _6677_/A3 _4410_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5388_ _5473_/A1 _5473_/A2 _5529_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7127_ hold87/Z _7300_/RN _7127_/CLK hold86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4339_ hold363/Z hold684/Z _4346_/S _4339_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7058_ _7058_/D _7315_/RN _7058_/CLK _7058_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_101_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _7299_/Q _6339_/A1 _6355_/A4 _6343_/A4 _6599_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_28_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ input40/Z _4320_/S _4015_/A2 _7047_/Q _3711_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _4690_/A1 _4690_/A2 _4690_/A3 _5260_/B _5054_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3641_ _7041_/Q _4040_/A2 _4045_/A2 _7057_/Q _3643_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6360_ _7276_/Q _6610_/A2 _6322_/Z _7114_/Q _6610_/B1 _7268_/Q _6365_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3572_ _3545_/B _3533_/Z _3624_/A2 hold83/I _3830_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_161_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _5311_/A1 _5514_/A1 _5311_/A3 _5311_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_114_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6291_ _6900_/Q _6291_/A2 _6291_/B1 _6883_/Q _6291_/C1 _6850_/Q _6297_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_130_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ _5242_/A1 _5375_/A2 _5522_/A2 _5242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_102_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ _5340_/A1 _5176_/A2 _5173_/B _5173_/C _5175_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4124_ _7263_/Q input82/Z _4128_/S _4125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4055_ _4058_/A2 _6725_/Q _6726_/Q _4056_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4957_ _5342_/A2 _5401_/A3 _4957_/B _4991_/B _5326_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4888_ _4915_/A3 _5417_/C _5457_/A1 _5306_/C _4889_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3908_ _6904_/Q hold83/I _5557_/A2 _4411_/A2 _3915_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_165_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3839_ _7278_/Q _4027_/A2 _4027_/B1 _7254_/Q _3841_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6627_ _6627_/I0 _7330_/Q _6628_/S _7330_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6558_ _7259_/Q _6319_/Z _6328_/Z _6767_/Q _6610_/B1 _7275_/Q _6561_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_180_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _5509_/A1 _5509_/A2 _5509_/A3 _5509_/A4 _5536_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6489_ _7201_/Q _6313_/Z _6387_/Z _7063_/Q _6493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5860_ hold50/Z hold254/Z _5862_/S _5860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4811_ _5283_/A2 _5268_/B _5324_/A4 _5283_/A4 _4815_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_179_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5791_ hold323/Z hold763/Z hold33/Z _7149_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4742_ _5270_/A2 _5134_/A3 _4746_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4673_ _4673_/A1 _4673_/A2 _4673_/A3 _4673_/A4 _4681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6412_ _7124_/Q _6308_/Z _6324_/Z _7052_/Q _6336_/Z _7100_/Q _6415_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3624_ _4305_/B2 _3624_/A2 _3545_/B _4402_/A4 _4015_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7392_ _7392_/I _7392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ _7299_/Q _6594_/A2 _6594_/A4 _6343_/A4 _6347_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3555_ _3523_/B _3521_/Z _5872_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3486_ hold37/I hold49/I _3491_/S _7351_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6274_ _6274_/A1 _6274_/A2 _6274_/B1 _7293_/Q _6275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _5225_/A1 _5225_/A2 _5225_/B _6922_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5156_ _5395_/A1 _5397_/A2 _5156_/B _5397_/C _5157_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ _4116_/A2 _4106_/Z _4108_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5087_ _5209_/A1 _5421_/B _5482_/B _5087_/B2 _5483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4038_ _6986_/Q _4038_/A2 _4038_/B1 _7010_/Q _4039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5989_ _5989_/A1 _5989_/A2 _7293_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 _3362_/ZN mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold309 _7342_/Q hold309/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet479_105 net429_54/I _7182_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_127 net429_61/I _7160_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3340_ _6806_/Q _6613_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_125_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet479_116 net479_151/I _7171_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_149 net829_455/I _7138_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet479_138 net829_483/I _7149_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5010_ _5010_/A1 _5010_/A2 _5014_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ _6961_/D _7243_/RN _6961_/CLK _6961_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ hold99/Z hold518/Z _5917_/S _7254_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6892_ _6895_/Q _7341_/RN _7341_/CLK _6892_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5843_ hold38/Z hold129/Z _5844_/S _5843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ hold50/Z hold261/Z _5776_/S _5774_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4725_ _5214_/A4 _5162_/A2 _4751_/B _4691_/C _5323_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_147_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4656_ _4656_/A1 _4656_/A2 _4656_/A3 _4656_/A4 _4656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4587_ _4587_/A1 _4587_/A2 _4587_/A3 _4590_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold810 _5779_/Z _7139_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput70 mgmt_gpio_in[7] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3607_ _3906_/A1 _3548_/B _5872_/A3 _3830_/C _4040_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput81 spi_sdo input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold821 _7130_/Q hold821/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7375_ _7375_/I _7375_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold843 _6967_/Q hold843/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold854 _7229_/Q hold854/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ _6593_/A3 _6343_/A4 _7299_/Q _6594_/A4 _6326_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xinput92 spimemio_flash_io3_oeb input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3538_ hold82/I _4395_/A2 _3541_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold832 _6775_/Q hold832/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold876 _4274_/Z _6798_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold898 _7180_/Q hold898/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold865 _6728_/Q hold865/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold887 _7122_/Q hold887/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6257_ _6903_/Q _6292_/B1 _6293_/B1 _6901_/Q _6899_/Q _6291_/A2 _6258_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3469_ _6725_/Q _6792_/Q _3469_/A3 _3470_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5208_ _5234_/A2 _5466_/A2 _5217_/B _5313_/A1 _5416_/C _5344_/C _5209_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_88_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6188_ hold96/I _6294_/A2 _6289_/B1 _7023_/Q _6192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5139_ _5497_/A2 _5440_/A2 _5440_/B1 _5228_/B _5499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _5497_/A1 _5493_/A1 _5490_/B _5490_/C _5491_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_145_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _5395_/A1 _4688_/A1 _5384_/B _5384_/C _4512_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_172_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4441_ _5414_/A1 _4795_/A2 _5441_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold117 hold117/I _5917_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold106 _5630_/Z _7007_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_8_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold128 _5603_/Z _6983_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_160_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold139 _7227_/Q hold139/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7160_ _7160_/D _7315_/RN _7160_/CLK _7160_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6111_ _7142_/Q _7293_/Q _6299_/B _6265_/B1 _6112_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4372_ _6624_/I0 _6866_/Q _4376_/S _6866_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _7091_/D _7243_/RN _7091_/CLK _7091_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6042_ _6043_/A1 _6245_/C _7291_/Q _7289_/Q _6292_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6944_ _6944_/D input75/Z _6944_/CLK _6944_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6875_ _6875_/D _7325_/CLK _6875_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5826_ hold2/Z hold25/Z _5826_/S hold26/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5757_ hold38/Z hold270/Z _5758_/S _5757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4708_ _4839_/A3 _4839_/A2 _5286_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_148_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5688_ _4178_/Z hold907/Z _5695_/S _7058_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _5250_/A1 _5309_/B _4639_/B _4643_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold662 _4433_/Z _6917_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap370 _7315_/RN _7286_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_104_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold640 _3548_/C _3505_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7358_ _7358_/D _7359_/RN _7358_/CLK _7358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold651 _6939_/Q hold651/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold673 _6872_/Q hold673/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6309_ _6355_/A4 _7296_/Q _6387_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7289_ _7289_/D _7322_/RN _7319_/CLK _7289_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_104_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold684 _6839_/Q hold684/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold695 _6902_/Q hold695/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26__1403_ net429_73/I net429_61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_106__1403_ clkbuf_4_1_0__1403_/Z net829_496/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_89__1403_ clkbuf_4_5_0__1403_/Z net479_145/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ _5172_/A1 _5326_/C _5220_/A3 _5325_/A2 _4996_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_64_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ _7141_/Q _4047_/B1 _4042_/B1 _7139_/Q _3941_/C _3943_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6660_ _6660_/I0 _7337_/Q _6668_/S _7337_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3872_ _6785_/Q _5560_/A1 hold22/I _5827_/A3 _3929_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_31_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6591_ _6755_/Q _6319_/Z _6347_/C _6769_/Q _6611_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5611_ hold59/Z hold428/Z hold69/Z _6990_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5542_ hold363/Z hold564/Z _5543_/S _5542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5473_ _5473_/A1 _5473_/A2 _5473_/B _5473_/C _5474_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7212_ _7212_/D _7359_/RN _7212_/CLK _7212_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4424_ hold363/Z hold560/Z _4425_/S _4424_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4355_ hold323/Z _6852_/Q _4355_/S _4355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7143_ _7143_/D _7243_/RN _7143_/CLK _7143_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_98_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7074_ _7074_/D _7243_/RN _7074_/CLK _7074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _4285_/Z hold622/Z _4286_/S _4286_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6025_ _6245_/C _7291_/Q _6121_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_440 net429_74/I _6787_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_451 net779_451/I _6776_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6927_ _6927_/D _7341_/RN _7331_/CLK hold10/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6858_ _6858_/D _7325_/CLK _6858_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5809_ hold861/Z hold363/Z _5817_/S _7164_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6789_ _6789_/D _7359_/RN _6789_/CLK _6789_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_108_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold470 _5942_/Z _7281_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold481 _7080_/Q hold481/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold492 _6738_/Q hold492/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4140_ _6989_/Q _4305_/B1 _4140_/B _4140_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4071_ _4071_/I _6896_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4973_ _5172_/A1 _5473_/B _5326_/C _5325_/A2 _4978_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_51_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _7359_/RN _7012_/Q _4069_/C _6712_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3924_ _3924_/A1 _3924_/A2 _3924_/A3 _3924_/A4 _3924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6643_ _6643_/A1 _6643_/A2 _6644_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet729_381 net429_83/I _6871_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_392 net779_423/I _6844_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_370 net779_451/I _6902_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3855_ _7166_/Q _4047_/A2 _3855_/B1 _6942_/Q _4045_/B1 _6959_/Q _3856_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6574_ _6788_/Q _6313_/Z _6331_/Z _6909_/Q _6335_/Z _6851_/Q _6575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3786_ _6933_/Q _4385_/I0 _3960_/S _3786_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5525_ _5525_/A1 _5525_/A2 _5525_/B _5526_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ _5503_/A1 _5456_/A2 _5530_/A2 _5477_/A2 _5457_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_117_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4407_ hold584/Z hold323/Z _4407_/S _4407_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5387_ _5387_/A1 _5340_/C _5387_/A3 _5503_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4338_ _4435_/A1 _5588_/A1 _5597_/A3 _5891_/A1 _4346_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7126_ _7126_/D _7243_/RN _7126_/CLK _7126_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_72__1403_ clkbuf_4_7_0__1403_/Z net529_184/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4269_ _5936_/A1 hold7/Z hold18/Z _5597_/A3 _4269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_87_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7057_ hold20/Z _7243_/RN _7057_/CLK _7057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6008_ _6343_/A4 _7299_/Q _6594_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_27_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3640_ hold55/I _4020_/A2 _3947_/B1 hold29/I _6743_/Q _4040_/B1 _3643_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_143_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3571_ hold227/Z _3533_/Z _3624_/A2 hold83/I _5566_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_155_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5310_ _5310_/A1 _5312_/A1 _5310_/B _5310_/C _5311_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6290_ _6910_/Q _6290_/A2 _6290_/B1 _6887_/Q _6297_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5241_ _5241_/A1 _5410_/B _5241_/B1 _5241_/B2 _5241_/C _5522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _5172_/A1 _5473_/C _4953_/Z _5172_/B1 _5473_/B _5173_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_114_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ _4119_/S _7271_/Q _4123_/B _4123_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4054_ _4058_/A2 _6725_/Q _4057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _5172_/A1 _5326_/C _4956_/A3 _5475_/C _5473_/A1 _5476_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_178_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _5417_/C _5416_/A2 _5475_/A2 _5196_/B2 _5525_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3907_ _6906_/Q hold83/I _5557_/A2 _5777_/A2 _3912_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_177_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3838_ _7270_/Q _3921_/A2 _4020_/A2 _7238_/Q _4037_/C1 _6965_/Q _3841_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6626_ _3745_/Z _7329_/Q _6628_/S _7329_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ hold44/I _6318_/Z _6608_/B1 hold94/I _6341_/Z _7001_/Q _6562_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_134_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _5507_/Z _5508_/A2 _5508_/A3 _5508_/A4 _5509_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3769_ _7126_/Q _3951_/B1 _4020_/B1 _7160_/Q _3770_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6488_ _6765_/Q _6328_/Z _6604_/A2 hold72/I _6494_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5439_ _5439_/A1 _5439_/A2 _5439_/B _5439_/C _5459_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_79_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7109_ _7109_/D _7286_/RN _7109_/CLK _7109_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _5283_/A2 _5324_/A3 _5268_/B _5283_/A4 _4815_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_178_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ hold363/Z hold807/Z hold33/Z _7148_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4741_ _4741_/A1 _4755_/A3 _5294_/B _4773_/B1 _4741_/C _5134_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4672_ _5099_/B _5099_/C _5457_/A1 _5460_/A3 _4673_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_135_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3623_ _4402_/A4 _3986_/A3 _5872_/A4 _5872_/A3 _4287_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6411_ _7116_/Q _6594_/A2 _6594_/A3 _6594_/A4 _6415_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7391_ _7391_/I _7391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6342_ _6593_/A2 _6387_/A2 _7294_/Q _6594_/A4 _6342_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3554_ _6881_/Q hold17/Z _3554_/B _3554_/C hold18/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_170_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3485_ hold1/I hold37/I _3491_/S _7352_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _6273_/A1 _6273_/A2 _6273_/A3 _6273_/A4 _6274_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5224_ _5224_/A1 _5221_/Z _5224_/B _5224_/C _5225_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_115_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5155_ _5324_/A3 _5220_/A3 _5473_/C _5142_/C _5155_/B2 _5156_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_84_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4106_ _4097_/B _4106_/A2 _4106_/A3 _4106_/A4 _4106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5086_ _5241_/A1 _5421_/B _5241_/B1 _5250_/B2 _5251_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ _7204_/Q _4037_/A2 _4037_/B1 _6871_/Q _4037_/C1 _6967_/Q _4039_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_25_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5988_ _6302_/A1 _6302_/A2 _6006_/B1 _7293_/Q _5989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4939_ _4991_/B _4963_/A2 _4963_/A3 _5338_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_21_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _6872_/Q _6321_/Z _6609_/B1 _6887_/Q _6612_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_166_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput180 _3371_/ZN mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput191 _3361_/ZN mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet479_117 net629_291/I _7170_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_106 net629_269/I _7181_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet479_128 net479_128/I _7159_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet479_139 net829_498/I _7148_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6960_ _6960_/D _7243_/RN _6960_/CLK _6960_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ hold323/Z hold645/Z _5917_/S _7253_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6891_ _6891_/D _7341_/RN _6926_/CLK _6891_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_19_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ hold50/Z hold164/Z _5844_/S _5842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5773_ hold59/Z hold220/Z _5776_/S _5773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4724_ _5214_/A4 _5162_/A2 _4751_/B _5287_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_166_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4655_ _5241_/A1 _4693_/B _4787_/B _5510_/A2 _4656_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold800 _7261_/Q hold800/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4586_ _5099_/B _5441_/A3 _5353_/A3 _5441_/A4 _5067_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput71 mgmt_gpio_in[8] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3606_ _3556_/B _3548_/B hold573/Z _3554_/B _5750_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput82 spi_sdoenb input82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7374_ _7374_/I _7374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold811 _7107_/Q hold811/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold855 _7204_/Q hold855/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6325_ _7297_/Q _7296_/Q _6594_/A2 _6540_/A4 _6325_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3537_ _6881_/Q _4060_/I0 _3624_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold844 _6744_/Q hold844/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput93 trap input93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold822 _5769_/Z _7130_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold833 _4244_/Z _6775_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold877 _6768_/Q hold877/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold866 _4179_/Z _6728_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold888 _5760_/Z _7122_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold899 _5828_/Z _7180_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6256_ _6884_/Q _6295_/A2 _6291_/C1 _6849_/Q _6258_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3468_ input58/Z _7357_/Q _3468_/S _7357_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3399_ _3399_/I _5214_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_20
XFILLER_131_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _4518_/Z _5344_/C _5313_/A1 _4751_/B _5423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6187_ _7055_/Q _6291_/A2 _6295_/B1 _7007_/Q _6291_/C1 _6999_/Q _6193_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5138_ _5353_/A4 _5138_/A2 _5138_/B _5216_/C _5499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _5209_/A1 _5353_/A3 _5445_/A2 _5087_/B2 _5446_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49__1403_ clkbuf_4_15_0__1403_/Z net779_416/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold107 _7000_/Q hold107/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4440_ _5414_/A1 _4795_/A2 _4716_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_145_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold118 _5917_/Z _7259_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold129 _7194_/Q hold129/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ _6106_/Z _6110_/A2 _6110_/A3 _6110_/A4 _6113_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4371_ _3859_/Z _6865_/Q _4376_/S _6865_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _7090_/D _7243_/RN _7090_/CLK _7090_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_112_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6041_ _7098_/Q _6294_/B1 _6289_/B1 _7018_/Q _6048_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ _6943_/D _7359_/RN _6943_/CLK _6943_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_26_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _6874_/D _7325_/CLK _6874_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ hold38/Z hold46/Z _5826_/S hold47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ hold50/Z hold289/Z _5758_/S _5756_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _4730_/B _4730_/C _4839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_147_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ _5891_/A1 _5741_/A2 _5863_/A3 _5827_/A1 _5695_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4638_ _4638_/A1 _4638_/A2 _4638_/A3 _4639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold630 _6979_/Q hold630/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4569_ _5460_/A1 _5295_/B2 _5322_/A2 _3399_/I _5421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold663 _6754_/Q hold663/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap371 _7359_/RN _7315_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_78_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap360 hold32/Z _5863_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold641 hold641/I hold641/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7357_ _7357_/D _6711_/Z _7364_/CLK _7357_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold652 _5543_/Z _6939_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold674 _4379_/Z _6872_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6308_ _6594_/A3 _6387_/A2 _7294_/Q _6594_/A4 _6308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_7288_ _7288_/D _7322_/RN _4144_/I1 _7288_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold685 _4339_/Z _6839_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold696 _4410_/Z _6902_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6239_ _7057_/Q _6291_/A2 _6291_/B1 _7033_/Q _6293_/B1 _7065_/Q _6240_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_85_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3940_ _3940_/A1 _3940_/A2 _3941_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _6769_/Q _5891_/A4 _5560_/A1 _5891_/A2 _3952_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6590_ _6590_/A1 _6590_/A2 _6434_/S _6590_/B2 _7321_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5610_ hold79/Z hold393/Z hold69/Z _6989_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _6677_/A3 _5566_/A1 _5863_/A3 _5863_/A4 _5543_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_8_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7211_ _7211_/D _7286_/RN _7211_/CLK _7211_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ _5472_/A1 _5472_/A2 _5472_/A3 _6925_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4423_ _6677_/A3 _4423_/A2 _5732_/A4 _5550_/A1 _4425_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_141_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ hold363/Z hold644/Z _4355_/S _6851_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7142_ _7142_/D _7300_/RN _7142_/CLK _7142_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_98_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7073_ hold85/Z _7322_/RN _7073_/CLK _7073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6024_ _6245_/B _7292_/Q _6265_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4285_ hold223/Z hold2/Z _4285_/S _4285_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6926_ _6926_/D _7341_/RN _6926_/CLK hold67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet779_430 net779_430/I _6802_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_441 net429_74/I _6786_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6857_ _6857_/D _6880_/CLK _6857_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_32__1403_ clkbuf_4_11_0__1403_/Z _4150__8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6788_ _6788_/D _7359_/RN _6788_/CLK _6788_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5808_ _5578_/B _5808_/A2 _5808_/A3 _5808_/A4 _5817_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_23_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112__1403_ net779_410/I net429_75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5739_ hold38/Z hold395/Z _5740_/S _7104_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_95__1403_ clkbuf_4_4_0__1403_/Z net629_269/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold471 _7225_/Q hold471/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold460 _4237_/Z _6770_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold482 _7233_/Q hold482/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold493 _4197_/Z _6738_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _3753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4070_ _6896_/Q _4115_/A2 _6890_/Q _4071_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _4972_/A1 _4972_/A2 _4958_/Z _4978_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6711_ input75/Z _7012_/Q _4069_/C _6711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3923_ _7131_/Q _4046_/B1 _4045_/A2 _7051_/Q _3924_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6642_ _6896_/Q _6642_/A2 _6642_/B1 _6666_/B2 _6643_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_189_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3854_ _3854_/A1 _3854_/A2 _3854_/A3 _3854_/A4 _3857_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_177_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_393 net779_423/I _6843_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_371 net429_96/I _6901_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_360 net729_387/I _6912_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_382 net429_75/I _6862_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6573_ _6772_/Q _6599_/A2 _6329_/Z _6861_/Q _6338_/Z _6905_/Q _6575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3785_ _3756_/Z _3785_/A2 _3785_/A3 _3785_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_157_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _5481_/Z _5524_/A2 _5531_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5455_ _5455_/I _5477_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4406_ hold586/Z hold363/Z _4407_/S _4406_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7125_ _7125_/D _7315_/RN _7125_/CLK _7125_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5386_ _5386_/A1 _4671_/B _5478_/A1 _5385_/Z _5408_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4337_ hold2/Z hold223/Z _4337_/S _4337_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _7056_/D _7243_/RN _7056_/CLK _7056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4268_ hold834/Z hold323/Z _4268_/S _4268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6007_ _7298_/Q _6007_/A2 _6007_/B _6010_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4199_ hold59/Z hold317/Z _4202_/S _4199_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _6909_/D _7359_/RN _6909_/CLK _6909_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold290 _5756_/Z _7119_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _4402_/A4 _3986_/A3 _5872_/A3 _3830_/B _3778_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_154_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5240_ _5240_/A1 _5240_/A2 _5241_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5171_ _4794_/Z _5171_/A2 _5401_/A2 _5525_/A1 _5172_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4122_ _4119_/S input90/Z _4123_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4053_ _4053_/A1 _4053_/A2 _6930_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4955_ _5326_/C _4956_/A3 _5397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3906_ _3906_/A1 _5872_/A2 _3509_/Z _5581_/A3 _3939_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_178_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4886_ _4886_/A1 _5195_/A2 _4886_/A3 _4886_/A4 _4889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6625_ _6625_/I0 _7328_/Q _6628_/S _7328_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3837_ _3834_/Z _3837_/A2 _3837_/A3 _3859_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6556_ _6556_/A1 _6556_/A2 _6556_/A3 _6556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3768_ _6740_/Q _4040_/B1 _4047_/A2 _7168_/Q _3770_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5507_ _5466_/B _5507_/A2 _5507_/A3 _5507_/A4 _5507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_145_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3699_ hold74/I hold18/I _5669_/A1 _5827_/A1 _3701_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6487_ _7257_/Q _6319_/Z _6354_/Z _7217_/Q _6494_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5438_ _5438_/A1 _5135_/Z _5265_/Z _4834_/B _5439_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xoutput340 _6880_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5369_ _5369_/A1 _5521_/B2 _5369_/B _5369_/C _5487_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_86_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _7108_/D _7286_/RN _7108_/CLK _7108_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_86_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7039_ _7039_/D _7322_/RN _7039_/CLK _7039_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _5460_/A1 _4751_/B _4691_/C _3399_/I _5324_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_1591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4671_ _5172_/A1 _5259_/B _5460_/A3 _4671_/B _4673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7390_ _7390_/I _7390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6410_ _7262_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6418_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3622_ _4402_/A4 _3986_/A3 _5642_/A3 _5808_/A3 _4017_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_174_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _7294_/Q _6594_/A4 _6540_/A4 _6387_/A2 _6341_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_155_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _4402_/A4 _3986_/A3 _5872_/A4 _5581_/A3 _4285_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6272_ _6788_/Q _6293_/A2 _6292_/B1 _6790_/Q _6273_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3484_ _4160_/B _6792_/Q _6795_/Q _3491_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5223_ _5140_/B _5222_/Z _6894_/Q _5320_/C _5224_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _5214_/A4 _5154_/A2 _5162_/A2 _5475_/A1 _5389_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_102_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4105_ _4483_/B _4792_/B _4105_/B _4105_/C _4106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5085_ _5082_/Z _5381_/A1 _5381_/A2 _5085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_84_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _4036_/A1 _4036_/A2 _4036_/A3 _4036_/A4 _4050_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _6805_/Q _6807_/Q _5987_/B _5989_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4938_ _4949_/A1 _4502_/B _4991_/A2 _4991_/A1 _5401_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_178_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4869_ _5490_/C _5534_/B1 _4869_/B1 _5353_/A3 _4869_/C _4874_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6608_ _6791_/Q _6318_/Z _6608_/B1 _6916_/Q _6341_/Z _6850_/Q _6612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_165_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _6539_/A1 _6539_/A2 _6434_/S _6539_/B2 _7319_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput170 _4166_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput181 _3370_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput192 _3360_/ZN mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_102_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet479_107 _4150__8/I _7180_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet479_118 net479_151/I _7169_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet479_129 net429_61/I _7158_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ hold363/Z hold650/Z _5917_/S _7252_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6890_ _6890_/D _7341_/RN _6926_/CLK _6890_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5841_ hold59/Z hold174/Z _5844_/S _5841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5772_ hold79/Z hold160/Z _5776_/S _5772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_11_0__1403_ clkbuf_3_5_0__1403_/Z clkbuf_4_11_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_21_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4723_ _5460_/A1 _3399_/I _5475_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ _4500_/B _4773_/C _4693_/B _4787_/B _5466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold801 _5920_/Z _7261_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4585_ _4518_/Z _5417_/C _5475_/A1 _5417_/B _4587_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput72 mgmt_gpio_in[9] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3605_ _3868_/A1 hold68/I _4402_/A3 _4305_/B2 _4009_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold812 _6969_/Q hold812/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7373_ _7373_/I _7373_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _7297_/Q _6594_/A2 _6540_/A4 _6328_/A4 _6324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xclkbuf_0__1403_ _4149_/ZN clkbuf_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold823 _7138_/Q hold823/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput83 spimemio_flash_clk input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3536_ _7371_/Q _6795_/Q _3536_/B _4060_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold845 _4204_/Z _6744_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput94 uart_enabled _4132_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold834 _6791_/Q hold834/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold856 _6760_/Q hold856/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold867 _7042_/Q hold867/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold878 _4234_/Z _6768_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold889 _7066_/Q hold889/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6255_ _6851_/Q _6295_/B1 _6294_/B1 _6911_/Q _6258_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5206_ _5413_/A2 _5497_/A1 _5206_/B _5421_/C _5313_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3467_ _6792_/Q _3960_/S _3468_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3398_ _7291_/Q _6245_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_6186_ _7071_/Q _6292_/B1 _6290_/B1 _7047_/Q _6193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5137_ _5137_/A1 _5500_/A1 _5222_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5068_ _5068_/A1 _5068_/A2 _5235_/A1 _5070_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_85_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4019_ _7244_/Q _4019_/A2 _4019_/B1 _6945_/Q _4019_/C _4021_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold108 _5622_/Z _7000_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold119 _7005_/Q hold119/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4370_ _6622_/I0 _6864_/Q _4376_/S _6864_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6040_ _6245_/B _7292_/Q _7289_/Q _7290_/Q _6289_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6942_ _6942_/D input75/Z _6942_/CLK _6942_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_19_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6873_ _6873_/D _7325_/CLK _6873_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5824_ hold50/Z hold63/Z _5826_/S hold64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5755_ hold59/Z hold436/Z _5758_/S _5755_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4706_ _4452_/Z _4518_/Z _4454_/Z _5305_/B _4730_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_148_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5686_ hold2/Z _7057_/Q hold19/Z hold20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4637_ _5236_/A4 _5517_/A1 _5309_/B _5441_/A3 _4638_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold620 _4262_/Z _6787_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold631 _5599_/Z _6979_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4568_ _5214_/A4 _5162_/A2 _5416_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold642 hold642/I _4355_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap372 input75/Z _7359_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_2_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7356_ _7356_/D _6710_/Z _7364_/CLK _7356_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold653 _6848_/Q hold653/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold675 _6871_/Q hold675/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4499_ _5172_/A1 _4915_/A3 _4499_/B _5060_/B _4689_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6307_ _7297_/Q _7296_/Q _6594_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold664 _4216_/Z _6754_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7287_ _7287_/D _7322_/RN _4144_/I1 _7287_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3519_ _4178_/S hold31/Z _3519_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold697 _6757_/Q hold697/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold686 _6916_/Q hold686/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6238_ hold94/I _6294_/A2 _6293_/A2 _7081_/Q _6240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_55__1403_ net579_205/I net579_221/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6169_ _6169_/A1 _6169_/A2 _6169_/A3 _6170_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _6848_/Q _4435_/A1 hold68/I _5557_/A2 _3948_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5540_ hold323/Z _6929_/Q _5540_/S _5540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5471_ _6925_/Q _4395_/C _5471_/B _5472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7210_ _7210_/D _7286_/RN _7210_/CLK _7210_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4422_ hold323/Z hold722/Z _4422_/S _4422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4353_ _4408_/A1 _6677_/A3 hold641/Z _5560_/A1 hold642/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7141_ _7141_/D _7243_/RN _7141_/CLK _7141_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_101_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7072_ _7072_/D _7322_/RN _7072_/CLK _7072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4284_ _4283_/Z hold678/Z _4286_/S _4284_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _5951_/B _6614_/B _7303_/Q _6065_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_420 net779_425/I _6816_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_431 net779_431/I _6801_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6925_ _6925_/D _7341_/RN _7331_/CLK _6925_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_82_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet779_442 net829_453/I _6785_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6_0__1403_ clkbuf_0__1403_/Z clkbuf_3_6_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6856_ _6856_/D _7325_/CLK _6856_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ hold331/Z hold2/Z _5807_/S _7163_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6787_ _6787_/D _7359_/RN _6787_/CLK _6787_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3999_ _7002_/Q hold18/I _4408_/A1 _5836_/A3 _4036_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_183_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ hold50/Z hold283/Z _5740_/S _5738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _5669_/A1 _4305_/C hold32/Z _5891_/A4 _5677_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_89_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7339_ _7339_/D _7341_/RN _4144_/I1 _7339_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold461 _7198_/Q hold461/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold472 _5879_/Z _7225_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold450 _7170_/Q hold450/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold483 _5888_/Z _7233_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold494 _6731_/Q hold494/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4971_ _4796_/Z _5327_/A2 _5327_/A3 _4971_/B2 _4972_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_149_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6710_ input75/Z _7012_/Q _4069_/C _6710_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_32_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _7019_/Q _4041_/A2 _4043_/B1 _6885_/Q _4040_/A2 _7035_/Q _3924_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6641_ _6898_/Q _6641_/A2 _6641_/B1 _6897_/Q _6643_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ _6730_/Q _3914_/B1 _4047_/B1 _7142_/Q _3853_/C _3854_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet729_383 net429_98/I _6861_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_361 net429_75/I _6911_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_372 net779_437/I _6900_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _6572_/A1 _6572_/A2 _6572_/A3 _6572_/A4 _6572_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xnet729_394 net779_425/I _6842_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3784_ _3784_/A1 _3784_/A2 _3784_/A3 _3784_/A4 _3785_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5523_ _5523_/A1 _5523_/A2 _5523_/A3 _5523_/A4 _5524_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_9_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5454_ _5454_/A1 _5454_/A2 _5455_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5385_ _5479_/A3 _5480_/A4 _5479_/A2 _5478_/A3 _5385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4405_ _5578_/B hold12/Z _4405_/A3 _5808_/A4 _4407_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_160_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7124_ _7124_/D _7286_/RN _7124_/CLK _7124_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4336_ hold38/Z hold329/Z _4337_/S _4336_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4267_ hold848/Z hold363/Z _4268_/S _4267_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7055_ _7055_/D _7243_/RN _7055_/CLK _7055_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6006_ _6807_/Q _6005_/Z _6006_/B1 _6343_/A4 _7298_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4198_ hold79/Z hold490/Z _4202_/S _4198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _6908_/D _7359_/RN _6908_/CLK _6908_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6839_ _6839_/D _7300_/RN _6839_/CLK _6839_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold280 _6947_/Q hold280/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold291 _6751_/Q hold291/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _5170_/A1 _5170_/A2 _5402_/A1 _5173_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4121_ _4119_/S _7279_/Q _4121_/B _4121_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4052_ _4051_/Z _3960_/S _6794_/Q _7356_/Q _4053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_92_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _5401_/A3 _4991_/B _4957_/B _4956_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3905_ _6850_/Q _6677_/A2 hold68/I _5557_/A2 _3945_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_177_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _5490_/B _5319_/A1 _5133_/B _5534_/A2 _4886_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6624_ _6624_/I0 _7327_/Q _6628_/S _7327_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3836_ _7132_/Q _4046_/B1 _4045_/A2 _7052_/Q input26/Z _4043_/A2 _3837_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6555_ _6555_/A1 _6555_/A2 _6555_/A3 _6555_/A4 _6556_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3767_ _7102_/Q _4006_/B1 _3919_/B1 _6748_/Q _3770_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5506_ _5506_/A1 _5506_/A2 _5319_/C _5507_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3698_ _7186_/Q _4014_/A2 _4006_/A2 _7080_/Q _3701_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6486_ hold63/I _6310_/Z _6335_/Z _7007_/Q _6494_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5437_ _5437_/A1 _5496_/A1 _5437_/A3 _5439_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xoutput330 _7327_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput341 _6863_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5368_ _5099_/C _5368_/A2 _5368_/A3 _4523_/C _5521_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_133_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4319_ _4318_/Z hold581/Z _4321_/S _4319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5299_ _4691_/C _5421_/C _5490_/C _5353_/A4 _5302_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7107_ _7107_/D input75/Z _7107_/CLK _7107_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7038_ _7038_/D _7315_/RN _7038_/CLK _7038_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0__1403_ clkbuf_4_9_0__1403_/I clkbuf_4_9_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_78_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4670_ _5099_/B _5099_/C _5460_/A3 _5172_/A1 _5442_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_175_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3621_ _3906_/A1 _3548_/B _5872_/A3 _3910_/A1 _4010_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_30_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6340_ _6340_/A1 _7294_/Q _7295_/Q _6610_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3552_ _3509_/Z _3521_/Z hold573/Z _3556_/B _4402_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6271_ _6778_/Q _6295_/A2 _6294_/A2 _6772_/Q _6273_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3483_ _3483_/A1 _3483_/A2 _4113_/A3 _3482_/B _7353_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5222_ _5222_/A1 _5499_/A1 _5499_/A2 _5263_/A2 _5222_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5153_ _5153_/A1 _5162_/A2 _5396_/A1 _5337_/A1 _5172_/A1 _5453_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4104_ _4104_/A1 _4104_/A2 _4104_/A3 _4116_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5084_ _5209_/A1 _5309_/B _5250_/B2 _5087_/B2 _5381_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4035_ _4035_/A1 _4035_/A2 _4035_/A3 _4035_/A4 _4035_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_53_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5986_ _6302_/A1 _6302_/A2 _7293_/Q _6807_/Q _5987_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4937_ _4963_/A2 _4963_/A3 _4957_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _5414_/A1 _5457_/A1 _4483_/B _4792_/B _4869_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_138_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3819_ _3819_/A1 _3809_/Z _3818_/Z _3819_/A4 _3819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6607_ _6607_/A1 _6607_/A2 _6607_/A3 _6612_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4799_ _3399_/I _5525_/A2 _5460_/A1 _4454_/Z _4802_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_165_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6538_ _5951_/B _7318_/Q _6614_/B _6539_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6469_ hold71/I _6324_/Z _6469_/B _6469_/C _6472_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput171 _4142_/ZN mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput182 _4140_/ZN mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput193 _3387_/ZN mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet479_108 net479_145/I _7179_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet479_119 net429_71/I _7168_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ hold79/Z hold281/Z _5844_/S _5840_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5771_ hold99/Z hold365/Z _5776_/S _5771_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4722_ _5295_/B2 _5322_/A2 _3399_/I _5220_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_147_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4653_ _5310_/B _4694_/B _5305_/B _4702_/B _5206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_174_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4584_ _4500_/B _5310_/B _4694_/B _5305_/B _5417_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold802 _6769_/Q hold802/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3604_ _3565_/B _3910_/A1 _3521_/Z _5872_/A4 _4008_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput73 pad_flash_io0_di input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput95 wb_adr_i[0] _3400_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold846 _6919_/Q hold846/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ _7298_/Q _6566_/A2 _6594_/A2 _6007_/B _6323_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold813 _6887_/Q hold813/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold824 _5778_/Z _7138_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput84 spimemio_flash_csb input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3535_ _3421_/B _6724_/Q _3536_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold835 _4268_/Z _6791_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold857 _4225_/Z _6760_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold868 _5670_/Z _7042_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold879 _6788_/Q hold879/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6254_ _6919_/Q _6265_/C _6299_/B _6299_/C _6275_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3466_ _6727_/Q _6726_/Q _6725_/Q _3960_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5205_ _5534_/A1 _5206_/B _5534_/B1 _5421_/B _5511_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3397_ _7292_/Q _6245_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_69_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _7015_/Q _6292_/A2 _6293_/B1 _7063_/Q _6193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5136_ _5438_/A1 _5135_/Z _5500_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _4515_/Z _5304_/A1 _5339_/A1 _5067_/B1 _5417_/A2 _5235_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_111_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ _4018_/A1 _4018_/A2 _4018_/A3 _4018_/A4 _4051_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_26_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5969_ _6231_/A1 _7290_/Q _6096_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15__1403_ clkbuf_4_10_0__1403_/Z net429_80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_178_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78__1403_ clkbuf_4_5_0__1403_/Z net779_425/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold109 _6842_/Q hold109/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _6941_/D input75/Z _6941_/CLK _6941_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6872_ _6872_/D _7286_/RN _6872_/CLK _6872_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5823_ hold59/Z hold170/Z _5826_/S _5823_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ hold79/Z hold178/Z _5758_/S _5754_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4705_ _5305_/C _4773_/B1 _4773_/C _4730_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_147_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5685_ hold38/Z hold209/Z hold19/Z _7056_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _4500_/B _5305_/B _4694_/B _4787_/B _5309_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold610 _4313_/Z _6820_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold621 _6987_/Q hold621/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_118_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7355_ _7355_/D _6709_/Z _4152_/I1 _7355_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4567_ _5460_/A1 _3399_/I _5133_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_162_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold632 _6918_/Q hold632/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6306_ _5951_/B _6614_/B _7313_/Q _6381_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold643 _4355_/Z _6852_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold654 _4349_/Z _6848_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold676 _4378_/Z _6871_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4498_ _4603_/A1 _4603_/A2 _4499_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7286_ _7286_/D _7286_/RN _4144_/I1 _7286_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3518_ _7365_/Q _6795_/Q _3520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold665 _6825_/Q hold665/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap373 _7243_/RN _7322_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold687 _4431_/Z _6916_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _7041_/Q _6295_/A2 _6290_/B1 _7049_/Q _6240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3449_ _6727_/Q _6725_/Q _6792_/Q _3492_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold698 _4220_/Z _6757_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _7118_/Q _6265_/C _6299_/B _6299_/C _6169_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_76_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _5406_/A1 _5277_/A2 _5130_/B1 _5534_/A2 _5526_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6099_ _7100_/Q _6294_/B1 _6293_/B1 _7060_/Q _6100_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_2__1403_ clkbuf_4_2_0__1403_/Z net429_72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5470_ _5470_/A1 _5509_/A3 _5470_/A3 _5470_/A4 _5471_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_145_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4421_ hold363/Z hold655/Z _4422_/S _4421_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7140_ _7140_/D _7243_/RN _7140_/CLK _7140_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4352_ hold741/Z hold323/Z _4352_/S _6850_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4283_ hold329/Z hold38/Z _4285_/S _4283_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7071_ _7071_/D _7322_/RN _7071_/CLK _7071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_140_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6022_ _6806_/Q _4062_/Z _6380_/C _6434_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_100_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_410 net779_410/I _6826_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_432 net779_435/I _6800_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6924_ _6924_/D _7341_/RN _6926_/CLK hold21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet779_421 net779_423/I _6815_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_443 net829_453/I _6784_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _6855_/D _7325_/CLK _6855_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5806_ hold415/Z hold38/Z _5807_/S _7162_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3998_ _6768_/Q _5891_/A4 hold185/I _5882_/A2 _4026_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6786_ _6786_/D _7359_/RN _6786_/CLK _6786_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5737_ hold59/Z hold276/Z _5740_/S _5737_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ hold2/Z _7041_/Q _5668_/S hold3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5599_ hold323/Z hold630/Z _5605_/S _5599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4619_ _4454_/Z _5462_/A2 _5421_/C _5534_/A2 _5195_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7338_ _7338_/D _7341_/RN _4144_/I1 _7338_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold451 _6998_/Q hold451/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold462 _5848_/Z _7198_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold440 _5835_/Z _7187_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7269_ _7269_/D _7315_/RN _7269_/CLK _7269_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold473 _6965_/Q hold473/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold484 _7062_/Q hold484/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold495 _4185_/Z _6731_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _5313_/A2 _5155_/B2 _4971_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ _7269_/Q _3921_/A2 _4037_/B1 _6872_/Q _3924_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _6640_/I0 _7332_/Q _6668_/S _7332_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3852_ _7206_/Q _4037_/A2 _4020_/B1 _7158_/Q _3854_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet729_362 net779_438/I _6910_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_384 _4150__3/I _6852_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6571_ _7358_/Q _6320_/Z _6325_/Z _6907_/Q _6572_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet729_373 net779_437/I _6899_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5522_ _5522_/A1 _5522_/A2 _5522_/A3 _5523_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3783_ _3783_/A1 _3783_/A2 _3783_/A3 _3784_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xnet729_395 net779_426/I _6841_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5453_ _5005_/Z _5529_/A2 _5529_/B1 _5335_/B _5453_/C _5454_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_145_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5384_ _5384_/A1 _5384_/A2 _5384_/B _5384_/C _5479_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4404_ hold813/Z hold323/Z _4404_/S _4404_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4335_ hold50/Z hold344/Z _4337_/S _4335_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7123_ _7123_/D _7243_/RN _7123_/CLK _7123_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _7054_/D _7243_/RN _7054_/CLK hold71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4266_ _5578_/B _5872_/A2 _3830_/B _4405_/A3 _4268_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6005_ _6343_/A4 _6007_/A2 _6005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4197_ hold99/Z hold492/Z _4202_/S _4197_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _6907_/D _7359_/RN _6907_/CLK _6907_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _6838_/D _7359_/RN _6838_/CLK _6838_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6769_ _6769_/D _7315_/RN _6769_/CLK _6769_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold270 _7120_/Q hold270/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold281 _7191_/Q hold281/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold292 _4211_/Z _6751_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4120_ _4119_/S input92/Z _4121_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4051_ _4051_/A1 _4051_/A2 _4051_/A3 _4050_/Z _4051_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_83_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _4789_/B _5030_/A2 _4953_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_91_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ _6910_/Q _5750_/A4 _5750_/A3 _4426_/A3 _3920_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4884_ _4454_/Z _5490_/B _5133_/B _5534_/A2 _4886_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6623_ _3859_/Z _7326_/Q _6628_/S _7326_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3835_ _7012_/Q _4038_/B1 _4041_/B1 input5/Z _3947_/B1 _7004_/Q _3837_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6554_ _7227_/Q _6317_/Z _6354_/Z hold42/I _6387_/Z _7065_/Q _6555_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3766_ _7216_/Q _4028_/A2 _3914_/B1 _6732_/Q _3770_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6485_ _6485_/A1 _6485_/A2 _6434_/S _6485_/B2 _7317_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5505_ hold67/I _4395_/C _5520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5436_ _5437_/A1 _5437_/A3 _5527_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3697_ _7128_/Q _3951_/B1 _3916_/B1 _7072_/Q _3701_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput331 _7328_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput320 _6855_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput342 _6864_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5367_ _5367_/A1 _5367_/A2 _5498_/C _5409_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_120_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4318_ hold91/Z hold38/Z _4320_/S _4318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7106_ _7106_/D _7315_/RN _7106_/CLK _7106_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5298_ _4698_/C _5417_/C _5344_/C _3399_/I _5300_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_113_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7037_ _7037_/D _7322_/RN _7037_/CLK _7037_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7300__378 _7300_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
X_4249_ hold363/Z hold594/Z _4250_/S _4249_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3620_ _3906_/A1 _3910_/A1 _3509_/Z _5872_/A3 _4010_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_30_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3551_ _3504_/Z _3523_/B _3554_/B _3548_/B _5564_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6270_ _6245_/B _6299_/B _6786_/Q _7292_/Q _6273_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3482_ _4113_/A3 _6792_/Q _3482_/B _3483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5221_ _5178_/Z _5345_/A1 _5346_/A2 _5221_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_102_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5152_ _5337_/A1 _5162_/A2 _5396_/A1 _5333_/B _5172_/A1 _5390_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_123_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4103_ _4103_/A1 _4103_/A2 _4103_/A3 _4103_/A4 _4104_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _5241_/A1 _5309_/B _5238_/B1 _5443_/B _5381_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4034_ _4034_/A1 _4034_/A2 _4034_/A3 _4034_/A4 _4035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5985_ _7290_/Q _7289_/Q _7292_/Q _7291_/Q _6142_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4936_ _5305_/C _5460_/A2 _5305_/B _4963_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_177_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _5417_/C _5350_/A2 _5475_/A1 _5416_/A2 _4869_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_21_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ _3818_/A1 _3818_/A2 _3818_/A3 _3817_/Z _3818_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6606_ _6606_/A1 _6606_/A2 _6606_/A3 _6606_/A4 _6607_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4798_ _5287_/A1 _5525_/A2 _4798_/B _4802_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_153_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6537_ _6537_/A1 _6537_/A2 _6992_/Q _6613_/A2 _6613_/C _6539_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_180_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3749_ input39/Z _4320_/S _3947_/B1 _7006_/Q _3752_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _6468_/A1 _6468_/A2 _6468_/A3 _6469_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5419_ _5308_/B _5533_/A3 _5419_/B _5419_/C _5514_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6399_ _7035_/Q _6312_/Z _6604_/A2 _7165_/Q _6400_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput194 _5877_/A2 mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput172 _3379_/ZN mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput183 _3369_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_38__1403_ clkbuf_4_14_0__1403_/Z net429_76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet479_109 net479_145/I _7178_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5770_ hold323/Z hold737/Z _5776_/S _5770_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _5457_/A1 _4843_/B1 _6898_/Q _5140_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4652_ _5380_/C _5534_/A1 _4591_/C _4499_/B _4656_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3603_ _5808_/A2 _3509_/Z _3504_/Z _5872_/A3 _4046_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4583_ _4773_/C _4693_/B _4787_/B _4702_/B _5353_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold803 _4235_/Z _6769_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7371_ _7371_/D _6723_/Z _3753_/A1 _7371_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput96 wb_adr_i[10] input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6322_ _7298_/Q _6594_/A2 _6594_/A4 _6007_/B _6322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xhold814 _4404_/Z _6887_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold836 _7389_/I hold836/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput85 spimemio_flash_io0_do input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold825 _6783_/Q hold825/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3534_ _6881_/Q hold115/Z _3542_/C _3868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xinput74 pad_flash_io1_di _3351_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold869 _7260_/Q hold869/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold847 _4436_/Z _6919_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold858 _7221_/Q hold858/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_107_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _6434_/S _6253_/A2 _6253_/B _7310_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3465_ _6727_/Q _6726_/Q _3469_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_171_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5204_ _5250_/A1 _5421_/B _5204_/B _5312_/C _5210_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _7289_/Q _6231_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_6184_ _6265_/C _7119_/Q _6245_/B _6245_/C _6194_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5135_ _5135_/A1 _5134_/Z _5135_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5066_ _4515_/Z _5304_/A1 _5473_/A1 _5296_/A3 _5066_/B2 _5068_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4017_ _7260_/Q _4017_/A2 _4017_/B1 input61/Z _4017_/C1 _6917_/Q _4018_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_84_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _6043_/A1 _7289_/Q _6266_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4919_ _5217_/B _4702_/B _5199_/A3 _5305_/B _5320_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_12_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5899_ hold2/Z hold55/Z _5899_/S hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_21__1403_ clkbuf_4_9_0__1403_/Z net429_64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _6940_/D input75/Z _6940_/CLK _6940_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_101__1403_ clkbuf_4_3_0__1403_/Z net829_452/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_84__1403_ clkbuf_4_5_0__1403_/Z net629_284/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _6871_/D _7286_/RN _6871_/CLK _6871_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5822_ hold79/Z hold267/Z _5826_/S _5822_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5753_ hold99/Z hold332/Z _5758_/S _5753_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4704_ _5305_/C _4698_/C _5462_/A2 _4773_/A2 _4702_/B _4839_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_175_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5684_ hold50/Z hold524/Z hold19/Z _7055_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4635_ _5443_/B _5460_/A1 _5214_/A4 _4454_/Z _4638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_8_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold600 _7277_/Q hold600/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4566_ _5296_/A3 _3399_/I _5475_/A1 _5162_/A2 _5063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_116_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold611 _6884_/Q hold611/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7354_ _7354_/D _6708_/Z _7364_/CLK _7354_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold633 _4434_/Z _6918_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap363 hold83/Z _5750_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold622 _7388_/I hold622/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6305_ _6305_/I0 _7312_/Q _6434_/S _7312_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3517_ _3421_/B hold182/Z hold183/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xmax_cap352 _5780_/A3 _5927_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold644 _6851_/Q hold644/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7285_ _7285_/D _7322_/RN _4144_/I1 _7285_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4497_ _4693_/B _5172_/A1 _4603_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_116_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold666 _6963_/Q _5576_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold655 _6909_/Q hold655/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap374 _7300_/RN _7243_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold677 _7051_/Q hold677/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold688 _6915_/Q hold688/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3353__1 _3353__1/I _6669_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3448_ _7365_/Q _3448_/I1 _3448_/S _7365_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6236_ _6236_/A1 _6236_/A2 _7293_/Q _6250_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold699 _6862_/Q hold699/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3379_ _7069_/Q _3379_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6167_ _6166_/Z _6167_/A2 _6167_/A3 _6170_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _5440_/A2 _5277_/A2 _5534_/B1 _5410_/B _5118_/C _5123_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_94_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _7076_/Q _6293_/A2 _6292_/A2 _7012_/Q _6100_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5049_ _5234_/A2 _5473_/A2 _5344_/B _5344_/C _5407_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_73_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet529_190 net579_213/I _7097_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4420_ _6677_/A3 _4426_/A3 _5750_/A3 hold83/Z _4422_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_132_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4351_ hold819/Z hold363/Z _4352_/S _6849_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4282_ _4281_/Z hold681/Z _4286_/S _4282_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7070_ _7070_/D _7322_/RN _7070_/CLK _7070_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6021_ _6613_/C _6807_/Q _6614_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_82_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_411 net779_411/I _6825_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_433 net779_435/I _6799_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6923_ _6923_/D _7341_/RN _6926_/CLK hold6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet779_444 net779_445/I _6783_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_422 net779_425/I _6814_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6854_ _6854_/D _7325_/CLK _6854_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6785_ _6785_/D _7359_/RN _6785_/CLK _6785_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3997_ _6784_/Q _5560_/A1 _5780_/A3 _5891_/A2 _4034_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5805_ hold177/Z hold50/Z _5807_/S _7161_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5736_ hold79/Z hold422/Z _5740_/S _5736_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5667_ hold38/Z hold441/Z _5668_/S _7040_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _4773_/C _4693_/B _4787_/B _4702_/B _5196_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5598_ hold363/Z hold708/Z _5605_/S _5598_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7337_ _7337_/D _7341_/RN _4144_/I1 _7337_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold452 _5620_/Z _6998_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold463 _7224_/Q hold463/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold441 _7040_/Q hold441/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4549_ _4641_/C _4787_/B _4499_/B _5095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_116_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold430 _5695_/Z _7065_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7268_ _7268_/D _7315_/RN _7268_/CLK _7268_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold474 _5582_/Z _6965_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold485 _5692_/Z _7062_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold496 _7038_/Q hold496/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6219_ _6219_/A1 _6219_/A2 _6219_/A3 _6219_/A4 _6219_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7199_ _7199_/D _7315_/RN _7199_/CLK _7199_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_38_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ input53/Z _4287_/A1 _4022_/B1 _6914_/Q _3920_/C _3924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ input58/Z _4303_/S _4285_/S input45/Z _4033_/A2 _7230_/Q _3854_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xnet729_352 net829_473/I _6920_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_374 net429_91/I _6887_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3782_ _7264_/Q _4017_/A2 _4015_/A2 _7046_/Q _3783_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet729_363 net729_367/I _6909_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6570_ _6884_/Q _6312_/Z _6337_/Z _6903_/Q _6572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _5534_/A1 _5534_/A2 _5075_/Z _5521_/B2 _5522_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet729_385 _4150__3/I _6851_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_396 net729_396/I _6840_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _5452_/A1 _5452_/A2 _5452_/A3 _5452_/A4 _5530_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_173_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4403_ hold885/Z hold363/Z _4404_/S _4403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5383_ _5442_/A2 _5383_/A2 _5484_/A2 _5383_/A4 _5386_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4334_ hold59/Z hold381/Z _4337_/S _4334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7122_ _7122_/D _7243_/RN _7122_/CLK _7122_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_141_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _7053_/D _7243_/RN _7053_/CLK _7053_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6004_ _6387_/A2 _6337_/A4 _6355_/A4 _6328_/A4 _6007_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4265_ hold323/Z hold827/Z _4265_/S _4265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4196_ hold323/Z hold795/Z _4202_/S _4196_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ _6906_/D _7359_/RN _6906_/CLK _6906_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6837_ _6837_/D _7359_/RN _6837_/CLK _6837_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6768_ _6768_/D _7315_/RN _6768_/CLK _6768_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5719_ hold59/Z hold235/Z _5722_/S _5719_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6699_ input75/Z _7012_/Q _4069_/C _6699_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_163_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold271 _5757_/Z _7120_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_163_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold260 _5637_/Z _7013_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold293 _7046_/Q hold293/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold282 _5840_/Z _7191_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4050_ _4035_/Z _4050_/A2 _4050_/A3 _4050_/A4 _4050_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_110_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _4789_/B _5030_/A2 _5401_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_91_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4883_ _4452_/Z _5490_/B _5216_/A2 _4773_/C _5195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3903_ _6920_/Q _4435_/A1 _5750_/A4 _5750_/A3 _3916_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6622_ _6622_/I0 _7325_/Q _6628_/S _7325_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3834_ _3834_/A1 _3834_/A2 _3834_/A3 _3834_/A4 _3834_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_177_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6553_ _7211_/Q _6316_/Z _6322_/Z _7121_/Q _6555_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3765_ _6998_/Q _3963_/A2 _3765_/B _3765_/C _3785_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5504_ _5504_/A1 _5503_/Z _5504_/B _5504_/C _5520_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6484_ _5951_/B _7316_/Q _4083_/B _6806_/Q _6485_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3696_ _3696_/A1 _3696_/A2 _3702_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5435_ _5435_/A1 _5435_/A2 _5435_/A3 _5437_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_145_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput310 _7323_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput332 _7329_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput321 _6856_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5366_ _4751_/B _5416_/A2 _5439_/A2 _5366_/B _5367_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_114_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4317_ _4316_/Z hold590/Z _4321_/S _4317_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5297_ _5183_/B _5297_/A2 _5515_/B1 _5421_/C _5302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_101_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7105_ _7105_/D _7322_/RN _7105_/CLK _7105_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4248_ _5550_/A1 _5863_/A4 _6677_/A1 _6677_/A3 _4250_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7036_ _7036_/D _7300_/RN _7036_/CLK _7036_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_142_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4179_ hold363/Z hold865/Z _4193_/S _4179_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3550_ _3521_/Z hold573/Z _5581_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_127_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5220_ _5220_/A1 _5344_/B _5220_/A3 _5338_/A2 _5346_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_127_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3481_ _3472_/B input58/Z _3483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5151_ _5333_/B _5162_/A2 _5396_/A1 _5391_/B _5172_/A1 _5529_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_96_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4102_ _4443_/A3 _4443_/A4 _4448_/A1 _4448_/A2 _4106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5082_ _5079_/Z _5246_/A1 _5444_/A1 _5082_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_97_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4033_ _7228_/Q _4033_/A2 _4033_/B1 _6772_/Q _4033_/C _4034_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5984_ _6245_/C _6245_/B _6302_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4935_ _3399_/I _4452_/Z _4454_/Z _4773_/C _4963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_52_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4866_ _5490_/B _4866_/A2 _5517_/A2 _5421_/A2 _5516_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4797_ _4961_/A2 _4961_/A3 _5171_/A2 _5326_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_6605_ _6777_/Q _6317_/Z _6354_/Z _6781_/Q _6387_/Z _6902_/Q _6606_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3817_ _3817_/A1 _3817_/A2 _3817_/A3 _3817_/A4 _3817_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_118_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6536_ _6613_/A2 _6530_/Z _6535_/Z _6537_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3748_ input48/Z _4285_/S _4041_/A2 _7022_/Q _3752_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ _7120_/Q _4010_/B1 _4042_/A2 _6766_/Q _3682_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6467_ _7134_/Q _6315_/Z _6316_/Z _7208_/Q _6468_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _5517_/A2 _5418_/A2 _5418_/B _5463_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6398_ _7141_/Q _6323_/Z _6334_/Z _7027_/Q _6352_/Z _7149_/Q _6400_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xoutput195 _3358_/ZN mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput173 _3378_/ZN mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput184 _3368_/ZN mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5349_ _5349_/I _6923_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _7019_/D _7243_/RN _7019_/CLK _7019_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_90_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4720_ _5216_/B _5216_/C _4843_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _4505_/Z _5061_/A3 _4499_/B _4591_/C _5482_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3602_ _3523_/B _3830_/C _3521_/Z _5808_/A4 _3919_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_162_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4582_ _4582_/A1 _4582_/A2 _5486_/A2 _4582_/A4 _4587_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7370_ _7370_/D _6722_/Z _3753_/A1 _7370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_44__1403_ clkbuf_4_15_0__1403_/Z net529_171/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput97 wb_adr_i[11] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold804 _6920_/Q hold804/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6321_ _7296_/Q _6594_/A2 _6540_/A4 _6355_/A4 _6321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xhold837 _5589_/Z _6970_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput86 spimemio_flash_io0_oeb input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3533_ _3542_/C _3532_/Z _3533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
Xhold826 _4256_/Z _6783_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput75 porb input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold815 _7019_/Q hold815/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold859 _5874_/Z _7221_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _6806_/Q _7309_/Q _6252_/B _6253_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3464_ _4114_/B2 _3464_/A2 _3464_/A3 _6794_/Q _3464_/B2 _7360_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xhold848 _6790_/Q hold848/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5203_ _5203_/A1 _5422_/A1 _5422_/A2 _5204_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6183_ _6183_/A1 _6183_/A2 _6183_/A3 _6182_/Z _6195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5134_ _5286_/A2 _5291_/C _5134_/A3 _5134_/A4 _5134_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_130_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3395_ _7290_/Q _6043_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_96_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5065_ _5482_/C _5065_/A2 _5087_/B2 _5371_/C _5373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4016_ _4016_/A1 _4016_/A2 _4016_/A3 _4016_/A4 _4051_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_25_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _6807_/Q _6006_/B1 _7289_/Q _7289_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4918_ _4918_/A1 _5508_/A4 _4918_/A3 _4924_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_178_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ hold38/Z hold141/Z _5899_/S _5898_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4849_ _4097_/B _4795_/B _5461_/A1 _5510_/A2 _5424_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_153_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _7040_/Q _6312_/Z _6355_/Z _7162_/Q _6520_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_250 net779_415/I _7037_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6870_ _6870_/D _6880_/CLK _6870_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_179_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5821_ hold99/Z hold367/Z _5826_/S _5821_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5752_ hold323/Z hold788/Z _5758_/S _5752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ _5294_/B _5462_/A2 _4698_/C _4500_/B _4730_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_148_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ hold59/Z hold71/Z hold19/Z _7054_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _4634_/A1 _5252_/A2 _4716_/B _4689_/A2 _5443_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4565_ _4500_/B _4693_/B _4787_/B _5305_/B _5296_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold601 _5938_/Z _7277_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_118_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold612 _4400_/Z _6884_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7353_ _7353_/D _6707_/Z _4152_/I1 _7353_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold645 _7253_/Q hold645/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3516_ _6881_/Q hold572/Z _3447_/B _3516_/B _3565_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xhold623 _4286_/Z _6804_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6304_ _6806_/Q _6304_/A2 _6304_/A3 _6304_/B _6305_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xhold634 _6904_/Q hold634/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7284_ _7284_/D _7315_/RN _7319_/CLK _7284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4496_ _5172_/A1 _4915_/A3 _5060_/B _4591_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_104_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold667 hold667/I hold667/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold678 _7387_/I hold678/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold656 _4421_/Z _6909_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap375 input75/Z _7300_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_104_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3447_ _7365_/Q _3421_/B _3447_/B _3448_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6235_ _6235_/A1 _6235_/A2 _6235_/A3 _6235_/A4 _6236_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold689 _4430_/Z _6915_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3378_ _7077_/Q _3378_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6166_ _6166_/A1 _6166_/A2 _6166_/A3 _6166_/A4 _6166_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _5117_/A1 _5360_/A1 _5360_/A2 _5118_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6097_ _7084_/Q _6289_/A2 _6292_/B1 _7068_/Q _7004_/Q _6295_/B1 _6100_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5048_ _4794_/Z _5182_/C _4483_/B _4716_/B _5346_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_85_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6999_ _6999_/D _7322_/RN _6999_/CLK _6999_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_139_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet529_191 net629_296/I _7096_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_180 net729_369/I _7107_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90__1403_ clkbuf_4_4_0__1403_/Z net829_493/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4350_ _5578_/B _5585_/A2 _5581_/A3 _5808_/A4 _4352_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_153_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4281_ hold344/Z hold50/Z _4285_/S _4281_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6020_ _4083_/B _6806_/Q _6380_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_79_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_434 net779_434/I _6798_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_412 net779_416/I _6824_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6922_ _6922_/D _7341_/RN _6926_/CLK hold31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet779_445 net779_445/I _6782_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_423 net779_423/I _6813_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6853_ _6853_/D _7325_/CLK _6853_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5804_ hold503/Z hold59/Z _5807_/S _7160_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3996_ _6788_/Q _5882_/A2 _5777_/A2 _4039_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6784_ _6784_/D _7359_/RN _6784_/CLK _6784_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5735_ hold99/Z hold583/Z _5740_/S _7100_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ hold50/Z hold410/Z _5668_/S _7039_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4617_ _4500_/B _5310_/B _4694_/B _5305_/B _5534_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5597_ _5936_/A1 _5812_/A1 _5597_/A3 _4305_/C _5605_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold420 _6771_/Q hold420/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold431 _7246_/Q hold431/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7336_ _7336_/D _7341_/RN _4144_/I1 _7336_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold442 _7184_/Q hold442/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold453 _7183_/Q hold453/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4548_ _5462_/A2 _5421_/C _5300_/A2 _5322_/A2 _5486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold486 _7044_/Q hold486/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4479_ _4711_/B _4483_/B _4795_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7267_ _7267_/D _7286_/RN _7267_/CLK _7267_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold464 _5878_/Z _7224_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold475 _7203_/Q hold475/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold497 _7280_/Q hold497/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6218_ _7000_/Q _6291_/C1 _6293_/B1 _7064_/Q _6219_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7198_ _7198_/D _7286_/RN _7198_/CLK _7198_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _7102_/Q _7292_/Q _7291_/Q _6266_/A2 _6156_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ _3850_/A1 _3850_/A2 _3850_/A3 _3850_/A4 _3850_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_189_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet729_353 net429_90/I _6919_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_375 net429_91/I _6886_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_364 net729_367/I _6908_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3781_ _7134_/Q _4046_/B1 _4045_/C2 input24/Z _3783_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5520_ _5520_/A1 _5520_/A2 _5520_/A3 _6926_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xnet729_397 net779_423/I _6839_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_386 net729_387/I _6850_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _5473_/A1 _5473_/A2 _5451_/B _5452_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5382_ _5382_/A1 _5382_/A2 _5382_/B1 _5382_/B2 _5382_/C _5383_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4402_ _4402_/A1 _5578_/B _4402_/A3 _4402_/A4 _4404_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_99_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4333_ hold79/Z hold158/Z _4337_/S _4333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7121_ _7121_/D _7286_/RN _7121_/CLK _7121_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4264_ hold363/Z hold879/Z _4265_/S _4264_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7052_ _7052_/D _7243_/RN _7052_/CLK _7052_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6003_ _4083_/B _7297_/Q _6339_/A1 _6003_/B _7297_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_140_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4195_ hold363/Z hold863/Z _4202_/S _4195_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6905_ _6905_/D _7359_/RN _6905_/CLK _6905_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6836_ _6836_/D _7359_/RN _6836_/CLK _6836_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6767_ _6767_/D _7286_/RN _6767_/CLK _6767_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5718_ hold79/Z hold455/Z _5722_/S _5718_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3979_ _6744_/Q _5891_/A4 _5550_/A1 _5566_/A1 _4026_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ input75/Z _7012_/Q _4069_/C _6698_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5649_ hold202/Z hold38/Z hold13/Z _7024_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold250 _7274_/Q hold250/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7319_ _7319_/D _7322_/RN _7319_/CLK _7319_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold261 _7135_/Q hold261/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold294 _5674_/Z _7046_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold272 _7016_/Q hold272/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold283 _7103_/Q hold283/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _4794_/Z _5171_/A2 _5331_/A3 _5342_/A2 _5475_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_36_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4882_ _4882_/A1 _5194_/C _4882_/A3 _4886_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_33_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3902_ _6753_/Q hold83/I _5557_/A2 _6677_/A2 _3943_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_178_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_14_0__1403_ clkbuf_3_7_0__1403_/Z clkbuf_4_14_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6621_ _4051_/Z _7324_/Q _6628_/S _7324_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3833_ _7028_/Q _4046_/A2 _4040_/B1 _6738_/Q _4040_/A2 _7036_/Q _3834_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_177_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3764_ _3764_/A1 _3764_/A2 _3765_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6552_ hold15/I _6308_/Z _6324_/Z _7057_/Q _6336_/Z _7105_/Q _6555_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5503_ _5503_/A1 _5503_/A2 _5503_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3695_ _7274_/Q _3921_/A2 _4019_/A2 _7250_/Q _3696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6483_ _6483_/A1 _6483_/A2 _6990_/Q _6613_/A2 _6613_/C _6485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5434_ _5434_/A1 _5434_/A2 _5435_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput300 _4062_/Z serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput311 _6873_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput322 _6874_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput333 _6875_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5365_ _5497_/A1 _5497_/A2 _5497_/B1 _5216_/C _5366_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7104_ _7104_/D _7322_/RN _7104_/CLK _7104_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4316_ hold127/Z hold50/Z _4320_/S _4316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5296_ _4691_/C _5416_/C _5296_/A3 _5296_/B1 _5417_/B _5297_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_114_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7035_ _7035_/D _7243_/RN _7035_/CLK _7035_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4247_ hold323/Z hold533/Z _4247_/S _4247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4178_ input58/Z hold362/Z _4178_/S _4178_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_142_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6819_ _6819_/D _7322_/RN _6819_/CLK _6819_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8__1403_ clkbuf_4_3_0__1403_/Z net779_445/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3480_ _3480_/A1 _3480_/A2 _7354_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5150_ _4698_/C _5344_/C _5326_/C _3399_/I _5397_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_170_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ _4101_/A1 _4101_/A2 _4448_/A3 _4448_/A4 _4103_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5081_ _5209_/A1 _5308_/B _5443_/B _5228_/A2 _5444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4032_ _7220_/Q hold7/I hold18/I _5882_/A2 _4033_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_84_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5983_ _7292_/Q _7291_/Q _6299_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_67__1403_ clkbuf_4_7_0__1403_/Z net579_217/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4934_ _4773_/C _4949_/A1 _4991_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4865_ _5417_/C _4694_/B _5310_/B _5294_/C _5517_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4796_ _5441_/A4 _4961_/A2 _4961_/A3 _4945_/A4 _4796_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6604_ _6783_/Q _6604_/A2 _6337_/Z _6904_/Q _6606_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3816_ input6/Z _4041_/B1 _4045_/A2 _7053_/Q _3817_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6535_ _6535_/A1 _6535_/A2 _6535_/A3 _6535_/A4 _6535_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3747_ _3746_/Z _6935_/Q _3961_/S _6935_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3678_ _7170_/Q _4047_/A2 _4038_/A2 _6992_/Q _3682_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6466_ _7248_/Q _6342_/Z _6355_/Z _7160_/Q _6468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5417_ _5417_/A1 _5417_/A2 _5417_/B _5417_/C _5418_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6397_ _7221_/Q _6317_/Z _6354_/Z _7213_/Q _6387_/Z _7059_/Q _6400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xoutput174 _3377_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput185 _5803_/A2 mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5348_ _5348_/A1 _5348_/A2 _5348_/A3 _4392_/Z hold6/I _5349_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xoutput196 _3357_/ZN mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ _5279_/A1 _5526_/A2 _5361_/A1 _5279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_102_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _7018_/D _7243_/RN _7018_/CLK _7018_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_29_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4650_ _5421_/C _5461_/A4 _5421_/B _5322_/A2 _4656_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3601_ _3548_/B _5872_/A3 _3910_/A1 _3504_/Z _4006_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_174_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4581_ _5102_/A1 _5475_/A1 _3399_/I _5162_/A2 _5413_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6320_ _7294_/Q _6594_/A3 _6387_/A1 _6387_/A2 _6320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput98 wb_adr_i[12] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput65 mgmt_gpio_in[36] _7399_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_156_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold805 _4437_/Z _6920_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput87 spimemio_flash_io1_do _7398_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3532_ _6881_/Q hold115/Z _3532_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold827 _6789_/Q hold827/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold816 _7173_/Q hold816/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput76 qspi_enabled _4119_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold838 _7390_/I hold838/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6251_ _5951_/B _6614_/B _7310_/Q _6253_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3463_ _7360_/Q _7356_/Q _3472_/B _3464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold849 _4267_/Z _6790_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5202_ _5534_/A1 _5421_/B _5534_/B1 _5309_/B _5422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ _6182_/A1 _6182_/A2 _6182_/A3 _6182_/A4 _6182_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5133_ _4454_/Z _5180_/B2 _5133_/B _5133_/C _5438_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_97_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3394_ _7293_/Q _6265_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_5064_ _5064_/A1 _5486_/A3 _5373_/A4 _5486_/A2 _5068_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _7042_/Q _4015_/A2 _4015_/B1 _6758_/Q _4015_/C1 _6886_/Q _4016_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_65_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _6805_/Q _6807_/Q _6006_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_12_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5897_ hold50/Z hold244/Z _5899_/S _5897_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4917_ _5461_/A4 _5213_/B _5218_/B _5322_/A2 _5508_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_12_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4848_ _4097_/B _4715_/B _4792_/B _5217_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4779_ _3399_/I _5277_/A2 _5460_/A1 _4454_/Z _4782_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_153_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6518_ _7128_/Q _6308_/Z _6322_/Z _7120_/Q _6520_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6449_ _7143_/Q _6323_/Z _6334_/Z hold90/I _6352_/Z _7151_/Q _6451_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_164_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50__1403_ clkbuf_4_15_0__1403_/Z net779_418/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet579_240 net579_240/I _7047_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_251 net779_426/I _7036_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ hold323/Z hold816/Z _5826_/S _7173_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ hold363/Z hold852/Z _5758_/S _5751_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4697_/Z _4518_/Z _4702_/B _4806_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xclkbuf_4_2_0__1403_ clkbuf_4_3_0__1403_/I clkbuf_4_2_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5682_ hold79/Z hold264/Z hold19/Z _7053_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4633_ _4633_/A1 _4633_/A2 _4633_/A3 _4638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold602 _7384_/I hold602/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_175_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7352_ _7352_/D _6706_/Z _4149_/B2 hold1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4564_ _4773_/C _5310_/B _4694_/B _4702_/B _5490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_128_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold613 _7383_/I hold613/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7283_ _7283_/D _7286_/RN _7283_/CLK _7283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold624 _7385_/I hold624/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6303_ _6806_/Q _7311_/Q _6304_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3515_ _6881_/Q hold17/Z _3554_/C _3523_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xmax_cap354 hold18/Z _5891_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xhold635 _4413_/Z _6904_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold646 _7245_/Q hold646/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap376 _3402_/I _4691_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_144_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4495_ _5310_/B _4694_/B _4915_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_116_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold668 hold668/I _6963_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold679 _4284_/Z _6803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap365 hold573/Z _3884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6234_ hold27/I _6290_/B1 _6291_/B1 _7155_/Q _6235_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold657 _6905_/Q hold657/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3446_ _3421_/B input58/Z _3447_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3377_ _7085_/Q _3377_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _7176_/Q _6291_/A2 _6292_/B1 _7192_/Q _6265_/C _6166_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _5417_/C _5359_/A1 _5416_/B _5324_/A4 _5274_/B _5360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_112_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6096_ _7036_/Q _6266_/A2 _6096_/B1 _7028_/Q _6299_/B _7020_/Q _6101_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_58_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5047_ _5047_/A1 _5047_/A2 _5051_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6998_ _6998_/D _7286_/RN _6998_/CLK _6998_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_26_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5949_ _6808_/Q _6806_/Q _6807_/Q _5952_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_13_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet529_170 net529_171/I _7117_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_181 net429_90/I _7106_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet529_192 net779_426/I _7095_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_153_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4280_ _4279_/Z hold624/Z _4286_/S _4280_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet779_402 net779_434/I _6834_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_435 net779_435/I _6797_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_413 net779_419/I _6823_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6921_ _6921_/D _7341_/RN _6926_/CLK hold17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet779_424 net779_425/I _6812_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6852_ _6852_/D _7359_/RN _6852_/CLK _6852_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_446 net429_75/I _6781_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5803_ _5807_/S _5803_/A2 _5803_/B hold757/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _6783_/D _7359_/RN _6783_/CLK _6783_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3995_ _6790_/Q _5560_/A1 _5836_/A3 _5827_/A3 _4029_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ hold323/Z hold717/Z _5740_/S _5734_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5665_ hold59/Z hold496/Z _5668_/S _7038_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _4500_/B _5305_/B _4694_/B _5310_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7335_ _7335_/D _7341_/RN _4144_/I1 _7335_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold410 _7039_/Q hold410/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5596_ hold2/Z hold413/Z _5596_/S _5596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold432 _5903_/Z _7246_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold443 _5832_/Z _7184_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold454 _5831_/Z _7183_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4547_ _5417_/C _5475_/A1 _3399_/I _5162_/A2 _5241_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold421 _4238_/Z _6771_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold487 _5672_/Z _7044_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7266_ _7266_/D _7286_/RN _7266_/CLK _7266_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ _4607_/A3 _4607_/A2 _5384_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold476 _6988_/Q hold476/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold465 _6741_/Q hold465/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7197_ _7197_/D _7315_/RN _7197_/CLK _7197_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_132_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold498 _5941_/Z _7280_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6217_ _7040_/Q _6295_/A2 _6292_/A2 _7016_/Q _6219_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3429_ _3421_/B hold81/Z _3531_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6148_ _6231_/A1 _6265_/B1 _7160_/Q _7290_/Q _6167_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6079_ _7149_/Q _6291_/B1 _6293_/B1 _7181_/Q _6080_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_354 net429_67/I _6918_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_365 net729_367/I _6907_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3780_ _5909_/A3 _5566_/A1 _4042_/A2 _6764_/Q _3783_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet729_398 net779_430/I _6838_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_376 net429_98/I _6885_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_387 net729_387/I _6849_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _5450_/A1 _5450_/A2 _5450_/B _5450_/C _5456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_145_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4401_ hold323/Z hold562/Z _4401_/S _4401_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5381_ _5381_/A1 _5381_/A2 _5381_/A3 _5381_/A4 _5484_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4332_ hold99/Z hold188/Z _4337_/S _4332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7120_ _7120_/D _7286_/RN _7120_/CLK _7120_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4263_ _5882_/A2 _5777_/A2 _6677_/A3 _4265_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_5_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7051_ _7051_/D _7243_/RN _7051_/CLK _7051_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6002_ _5999_/Z _7297_/Q _6003_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4194_ _5891_/A1 _5566_/A1 _5891_/A3 _5891_/A4 _4202_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_94_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _6904_/D input75/Z _6904_/CLK _6904_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6835_ _6835_/D _7359_/RN _6835_/CLK _6835_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6766_ _6766_/D _7286_/RN _6766_/CLK _6766_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _6728_/Q _5566_/A1 _6677_/A2 _4016_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ hold99/Z hold557/Z _5722_/S _7084_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6697_ _7359_/RN _7012_/Q _4069_/C _6697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7364_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5648_ hold530/Z hold50/Z hold13/Z _7023_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5579_ hold116/Z _5909_/A2 _6677_/A2 _4305_/C _5580_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold251 _5934_/Z _7274_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7318_ _7318_/D _7322_/RN _7322_/CLK _7318_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold262 _5774_/Z _7135_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold240 _5710_/Z _7078_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold273 _5640_/Z _7016_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7249_ _7249_/D _7286_/RN _7249_/CLK _7249_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold295 _7036_/Q hold295/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold284 _5738_/Z _7103_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_92_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _5473_/B _5326_/C _5325_/A2 _5395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_91_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4881_ _5417_/C _5416_/A2 _5475_/A2 _5359_/A1 _4882_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_33_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3901_ _4402_/A4 _5581_/A3 _5642_/A3 _4402_/A3 _3947_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_189_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6620_ _6895_/D _7341_/RN _6628_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_60_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ input22/Z _4045_/C2 _4019_/B1 _6947_/Q _3834_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6551_ _7137_/Q _6315_/Z _6342_/Z _7251_/Q _6551_/C _6555_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5502_ _5502_/A1 _5502_/A2 _5265_/Z _5504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3763_ _7192_/Q _3930_/A2 _3916_/B1 _7070_/Q _3764_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3694_ input59/Z _4287_/A1 _4038_/B1 _7016_/Q _3696_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6482_ _6482_/A1 _6482_/A2 _6481_/Z _6483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5433_ _5301_/B _5493_/A1 _5525_/A1 _5433_/B2 _5434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput301 _3736_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5364_ _5364_/A1 _5364_/A2 _5438_/A1 _5265_/Z _5367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_27__1403_ net429_73/I _4150__6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput334 _7330_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput323 _6857_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_107__1403_ clkbuf_4_1_0__1403_/Z net829_499/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput312 _6865_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4315_ _4314_/Z hold710/Z _4321_/S _6821_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7103_ _7103_/D _7322_/RN _7103_/CLK _7103_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5295_ _4691_/C _5353_/A4 _5462_/A2 _5295_/B2 _5296_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4246_ hold363/Z hold531/Z _4247_/S _4246_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7034_ _7034_/D _7243_/RN _7034_/CLK _7034_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_142_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ _5566_/A1 _6677_/A2 _5891_/A1 _4193_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_67_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _6818_/D _7322_/RN _6818_/CLK _6818_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6749_ _6749_/D _7243_/RN _6749_/CLK _6749_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_164_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ input97/Z input96/Z input99/Z input98/Z _4106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5080_ _5241_/A1 _5308_/B _5238_/B1 _5377_/B _5246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ input11/Z _4031_/A2 _4031_/B1 _6938_/Q _4031_/C _4034_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_77_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ _6805_/Q _6807_/Q _6245_/C _5982_/B1 _6291_/A2 _7292_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_18_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4933_ _4949_/A1 _4502_/B _4991_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_177_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ _5102_/A1 _5416_/A2 _4751_/B _4691_/C _4866_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4795_ _5414_/A1 _4795_/A2 _4795_/B _4795_/C _5171_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_119_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _6771_/Q _6323_/Z _6334_/Z _6883_/Q _6352_/Z _6775_/Q _6606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_32_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3815_ _7159_/Q _4020_/B1 _3947_/B1 _7005_/Q input23/Z _4045_/C2 _3817_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6534_ hold74/I _6335_/Z _6337_/Z _7072_/Q _6535_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _6934_/Q _3745_/Z _3960_/S _3746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6465_ _7184_/Q _6320_/Z _6325_/Z _7086_/Q _7038_/Q _6312_/Z _6468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5416_ _4751_/B _5416_/A2 _5416_/B _5416_/C _5418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3677_ _3673_/Z _3677_/A2 _3677_/A3 _3677_/A4 _3677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_161_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6396_ _6396_/A1 _6396_/A2 _6396_/A3 _6396_/A4 _6396_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xoutput175 _3376_/ZN mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput186 _5813_/A2 mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5347_ _6894_/Q _5320_/C _5347_/B1 _5430_/A2 _5347_/C _5348_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xoutput197 _3356_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5278_ _5421_/A2 _5525_/A2 _5278_/B _5278_/C _5361_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4229_ hold59/Z hold375/Z _4232_/S _4229_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7017_ _7017_/D _7322_/RN _7017_/CLK _7017_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_16_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_10__1403_ net479_128/I net729_359/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_79_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73__1403_ clkbuf_4_7_0__1403_/Z net679_333/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _5515_/A1 _5413_/A2 _5490_/C _5421_/C _4582_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3600_ _5808_/A2 _3509_/Z _3504_/Z _5808_/A3 _3951_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3531_ _3531_/A1 _3432_/B _4178_/S _3542_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput66 mgmt_gpio_in[37] _7400_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xinput88 spimemio_flash_io1_oeb input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold828 _4265_/Z _6789_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput77 ser_tx input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold806 _7237_/Q hold806/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold817 _6882_/Q hold817/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput99 wb_adr_i[13] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_171_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold839 _5590_/Z _6971_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6250_ _6250_/A1 _6250_/A2 _6806_/Q _6250_/C _6252_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3462_ _3421_/B _3472_/B _7360_/Q _3464_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_170_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _5413_/A2 _5497_/A1 _5309_/B _5421_/C _5422_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3393_ _7321_/Q _6590_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6181_ _7201_/Q _6293_/A2 _6289_/B1 hold76/I _6182_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5132_ _5132_/A1 _5494_/A1 _5501_/A1 _5137_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5063_ _5482_/C _5063_/A2 _5241_/B1 _5061_/Z _5373_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_84_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4014_ _7180_/Q _4014_/A2 _4014_/B1 _6782_/Q _4016_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _5965_/A1 _5963_/Z _5965_/A3 _5965_/B _7288_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_25_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5896_ hold59/Z hold379/Z _5899_/S _5896_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4916_ _5218_/B _5450_/A1 _4916_/B _4916_/C _4918_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4847_ _4711_/B _4929_/A3 _4929_/A2 _4483_/B _5218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_21_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4778_ _5287_/A1 _5277_/A2 _4778_/B _4782_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6517_ _7048_/Q _6609_/B1 _6341_/Z _7000_/Q _6520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3729_ _3729_/A1 _3729_/A2 _3729_/A3 _3729_/A4 _3743_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _7223_/Q _6317_/Z _6354_/Z _7215_/Q _6387_/Z _7061_/Q _6451_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_164_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6379_ _6379_/A1 _6613_/A2 _6365_/Z _6379_/A4 _6380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_241 _4150__46/I _7046_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet579_230 net629_266/I _7057_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _4305_/C _5750_/A2 _5750_/A3 _5750_/A4 _5758_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4701_ _4832_/A1 _4710_/A2 _5283_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5681_ hold99/Z hold608/Z hold19/Z _7052_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4632_ _5417_/C _5416_/C _5198_/A1 _4691_/C _4633_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_8_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold603 _4278_/Z _6800_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7351_ _7351_/D _6705_/Z _4149_/B2 hold37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4563_ _4693_/B _4787_/B _5306_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold614 _4276_/Z _6799_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4494_ _4693_/B _4787_/B _5461_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7282_ _7282_/D _7286_/RN _7282_/CLK _7282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold625 _4280_/Z _6801_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3514_ _6881_/Q hold572/Z _3447_/B _3554_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6302_ _6302_/A1 _6302_/A2 _6848_/Q _7293_/Q _6304_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xhold636 _6903_/Q hold636/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap377 _4762_/A4 _3399_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold647 _5902_/Z _7245_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3445_ hold571/Z _6795_/Q hold572/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6233_ _7235_/Q _6294_/A2 _6291_/C1 hold15/I _6235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold658 _6906_/Q hold658/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold669 _6752_/Q hold669/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3376_ _7093_/Q _3376_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6164_ _7216_/Q _6290_/A2 _6292_/A2 _6764_/Q _6293_/B1 _7184_/Q _6166_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _5193_/A1 _5268_/B _5134_/A4 _5274_/B _5473_/A2 _5360_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6095_ _6095_/A1 _6095_/A2 _6102_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5046_ _5098_/B1 _5344_/B _5177_/B1 _5473_/A2 _5046_/C _5047_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_111_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6997_ _6997_/D _7286_/RN _6997_/CLK _6997_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_25_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _6808_/Q _6806_/Q _5951_/B _5965_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5879_ hold471/Z hold50/Z _5881_/S _5879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet529_171 net529_171/I _7116_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet529_160 net629_284/I _7127_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_182 net529_184/I _7105_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet529_193 net429_87/I _7094_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150__50 net429_99/I _7237_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet779_403 net779_434/I _6833_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_414 net779_414/I _6822_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6920_ _6920_/D _7315_/RN _6920_/CLK _6920_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet779_425 net779_425/I _6811_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_436 net829_452/I _6791_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6851_ _6851_/D _7359_/RN _6851_/CLK _6851_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_447 net429_75/I _6780_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5802_ hold574/Z _5812_/A2 _4305_/C hold79/Z _5803_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6782_ _6782_/D _7359_/RN _6782_/CLK _6782_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3994_ _5564_/A1 _5566_/A1 _3993_/Z _4030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5733_ hold363/Z hold719/Z _5740_/S _5733_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5664_ hold79/Z hold406/Z _5668_/S _7037_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4615_ _4452_/Z _5421_/C _5320_/A1 _4773_/C _4620_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5595_ hold38/Z hold168/Z _5596_/S _5595_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7334_ _7334_/D _7341_/RN _4144_/I1 _7334_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4546_ _5214_/A4 _5460_/A1 _5322_/A2 _4751_/B _5417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_135_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold400 _7061_/Q hold400/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold411 _7077_/Q hold411/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold444 _7234_/Q hold444/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold433 _7226_/Q hold433/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold422 _7101_/Q hold422/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7265_ _7265_/D _7286_/RN _7265_/CLK _7265_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold477 _7222_/Q hold477/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4477_ _4792_/B _4523_/A2 _4523_/C _5099_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_145_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold455 _7085_/Q hold455/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold466 _4200_/Z _6741_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold499 _7278_/Q hold499/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7196_ _7196_/D _7315_/RN _7196_/CLK _7196_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6216_ _7112_/Q _6294_/A2 _6289_/B1 _7024_/Q _6219_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3428_ _7370_/Q _3428_/I1 _3448_/S _7370_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold488 _6928_/Q hold488/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3359_ _7223_/Q _5877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6147_ _6147_/A1 _6434_/S _6147_/B _7306_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6078_ _7221_/Q _6266_/A2 _6096_/B1 _7213_/Q _6299_/B _7205_/Q _6080_/B1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _5172_/A1 _5326_/C _5338_/A2 _4953_/Z _5032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_73_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet729_355 net429_64/I _6917_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_366 net729_367/I _6906_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_399 net429_72/I _6837_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_377 net729_387/I _6884_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_388 net729_389/I _6848_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4400_ hold363/Z hold611/Z _4401_/S _4400_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5380_ _5534_/A1 _5521_/B2 _5380_/B _5380_/C _5381_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4331_ hold323/Z hold626/Z _4337_/S _4331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4262_ hold323/Z hold619/Z _4262_/S _4262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7050_ _7050_/D _7243_/RN _7050_/CLK _7050_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6001_ _6001_/I _7296_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ hold2/Z hold210/Z _4193_/S _4193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _6903_/D input75/Z _6903_/CLK _6903_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6834_ _6834_/D _7286_/RN _6834_/CLK _6834_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6765_ _6765_/D _7286_/RN _6765_/CLK _6765_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3977_ _6940_/Q _5909_/A3 _5557_/A2 hold68/I _4021_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5716_ hold323/Z hold706/Z _5722_/S _5716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6696_ _7359_/RN _7012_/Q _4069_/C _6696_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_163_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ hold691/Z hold59/Z hold13/Z _7022_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5578_ hold667/Z _5578_/A2 _5578_/B hold668/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold252 _7282_/Q hold252/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4529_ _5490_/B _5460_/A1 _5214_/A4 _4454_/Z _5196_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_116_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7317_ _7317_/D _7322_/RN _7319_/CLK _7317_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold230 _5556_/Z _6950_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold241 _7110_/Q hold241/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold285 _6765_/Q hold285/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold274 _7249_/Q hold274/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7248_ _7248_/D _7315_/RN _7248_/CLK _7248_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold296 _5663_/Z _7036_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold263 _6957_/Q hold263/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7179_ hold26/Z _7300_/RN _7179_/CLK hold25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4880_ _5417_/C _5475_/A1 _5416_/A2 _5359_/A1 _5194_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3900_ _7261_/Q _5936_/A1 _5927_/A3 hold32/I _3934_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3831_ _7150_/Q _3981_/A2 _4042_/A2 _6762_/Q _7020_/Q _4041_/A2 _3834_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6550_ _6550_/A1 _6550_/A2 _6550_/A3 _6556_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3762_ _7184_/Q _4014_/A2 _4024_/A2 _7176_/Q _3764_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ _5501_/A1 _5501_/A2 _5502_/A2 _5528_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ _6613_/A2 _6481_/A2 _6481_/A3 _6481_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3693_ _3693_/A1 _3693_/A2 _3693_/A3 _3693_/A4 _3702_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5432_ _5432_/A1 _5432_/A2 _5432_/A3 _5496_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_160_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5363_ _5363_/A1 _5360_/Z _5432_/A2 _5495_/A1 _5364_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_126_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput335 _7331_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput324 _6858_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput302 _3670_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput313 _6866_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4314_ hold402/Z hold59/Z _4320_/S _4314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _7102_/D _7322_/RN _7102_/CLK _7102_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5294_ _5466_/A1 _5359_/A2 _5294_/B _5294_/C _5515_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_114_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ hold9/Z _7300_/RN _7033_/CLK _7033_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4245_ _5550_/A1 _5863_/A4 _5891_/A2 _6677_/A3 _4247_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4176_ hold309/Z hold101/Z _6881_/Q _4305_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_68_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6817_ _6817_/D _7322_/RN _6817_/CLK _6817_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6748_ _6748_/D _7300_/RN _6748_/CLK _6748_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_50_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6679_ hold323/Z hold753/Z _6679_/S _6679_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33__1403_ clkbuf_4_11_0__1403_/Z _4150__25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_113__1403_ net779_410/I net829_453/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_96__1403_ clkbuf_4_4_0__1403_/Z net429_87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_174_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _4030_/A1 _4030_/A2 _4031_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _5981_/A1 _6807_/Q _5982_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4932_ _4456_/Z _5199_/A3 _4932_/B _5336_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_80_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4863_ _5490_/B _5300_/B _5413_/B _4863_/B2 _4874_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6602_ _7359_/Q _6320_/Z _6325_/Z _6908_/Q _6885_/Q _6312_/Z _6606_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_60_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ _4961_/A2 _4961_/A3 _4794_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3814_ _7271_/Q _3921_/A2 _4287_/A1 input55/Z _3817_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _7194_/Q _6318_/Z _6334_/Z _7032_/Q _6535_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3745_ _3745_/A1 _3745_/A2 _3745_/A3 _3745_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
X_6464_ _6464_/A1 _6464_/A2 _6469_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5415_ _5369_/B _5300_/B _5300_/C _5415_/A4 _5518_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_133_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3676_ input32/Z _4043_/A2 _4041_/B1 input9/Z _3677_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6395_ _7197_/Q _6313_/Z _6331_/Z _7091_/Q _6335_/Z _7003_/Q _6396_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5346_ _5346_/A1 _5346_/A2 _5346_/A3 _5407_/B _5348_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xoutput176 _3375_/ZN mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput198 _3355_/ZN mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5277_ _5287_/A1 _5277_/A2 _5534_/B1 _5410_/B _5277_/C _5526_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xoutput187 _3365_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7016_ _7016_/D _7286_/RN _7016_/CLK _7016_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4228_ hold79/Z hold338/Z _4232_/S _4228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4159_ _4159_/A1 _7361_/Q _4159_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3530_ _6881_/Q hold10/Z _3530_/B hold11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput89 spimemio_flash_io2_do input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold807 _7148_/Q hold807/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput78 spi_csb input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold818 _4397_/Z _6882_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_170_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold829 _6761_/Q hold829/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3461_ _3461_/I _7361_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ _5534_/A1 _5309_/B _5200_/B _5200_/C _5203_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3392_ _7320_/Q _6565_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6180_ _7135_/Q _6295_/B1 _6291_/B1 _7153_/Q _6182_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5131_ _5440_/A2 _5216_/A2 _5493_/B _5501_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ _5241_/B1 _5369_/A1 _5061_/Z _5087_/B2 _5486_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _4013_/A1 _4013_/A2 _4011_/Z _4013_/A4 _4051_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _5964_/A1 _5964_/A2 _6808_/Q _5964_/B1 _7288_/Q _5965_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_80_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5895_ hold79/Z hold350/Z _5899_/S _5895_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4915_ _5324_/A4 _4702_/B _4915_/A3 _5305_/B _5450_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_61_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4846_ _4846_/A1 _4846_/A2 _5140_/B _5053_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _4777_/A1 _4777_/A2 _4777_/A3 _4777_/A4 _4778_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6516_ _7080_/Q _6338_/Z _6387_/Z _7064_/Q _6520_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3728_ _7193_/Q _3930_/A2 _4045_/C2 input25/Z _3729_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6447_ _6447_/A1 _6447_/A2 _6447_/A3 _6447_/A4 _6447_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3659_ _3659_/A1 _3643_/Z _3659_/A3 _3658_/Z _3659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_161_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _7066_/Q _6337_/Z _6347_/C _7236_/Q _6378_/C _6379_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5329_ _5329_/A1 _5327_/Z _5329_/B _5332_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_242 net629_271/I _7045_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_220 net629_298/I _7067_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_231 net729_389/I _7056_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_1__f__1085_ clkbuf_0__1085_/Z _6625_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ _5294_/B _4773_/B1 _4741_/C _4710_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_148_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ hold323/Z hold677/Z hold19/Z _7051_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ _5322_/A2 _5417_/C _5416_/C _5198_/A1 _4633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_30_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _5199_/A3 _5473_/A1 _4702_/B _5305_/B _5384_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7350_ _7350_/D _6704_/Z _4149_/B2 hold49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold626 _6832_/Q hold626/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4493_ _4603_/A1 _4787_/B _5060_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7281_ _7281_/D _7286_/RN _7281_/CLK _7281_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6301_ _7293_/Q _6301_/A2 _6301_/B _6304_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3513_ _6881_/Q hold17/Z _3516_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold615 _6953_/Q hold615/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold604 _6912_/Q hold604/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold648 _7244_/Q hold648/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold659 _6755_/Q hold659/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3444_ _3444_/A1 _3444_/A2 _7366_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xmax_cap345 _5669_/A1 _4408_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6232_ _7203_/Q _6293_/A2 _6293_/B1 _7187_/Q _6235_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold637 _4412_/Z _6903_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3375_ _7101_/Q _3375_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ _7200_/Q _6293_/A2 _6291_/B1 _7152_/Q _6166_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _5294_/C _5199_/A3 _5196_/B1 _5274_/B _5473_/A2 _5358_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6094_ _7092_/Q _6290_/A2 _6291_/C1 _6996_/Q _6095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5045_ _5417_/A2 _5344_/C _5344_/B _5177_/B1 _5324_/A4 _5458_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6996_ _6996_/D _7286_/RN _6996_/CLK _6996_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _4062_/Z _6806_/Q _5951_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_25_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5878_ hold463/Z hold59/Z _5881_/S _5878_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet529_172 net429_81/I _7115_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4829_ _5421_/A2 _5216_/B _4835_/A1 _4829_/A4 _5135_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet529_161 net429_71/I _7126_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_194 net779_415/I _7093_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_183 net629_297/I _7104_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150__40 _4150__40/I _7247_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__51 _4150__51/I _7236_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold1 hold1/I hold1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_79_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_404 net779_404/I _6832_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_415 net779_415/I _6821_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_426 net779_426/I _6810_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6850_ _6850_/D _7359_/RN _6850_/CLK _6850_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet779_448 net829_475/I _6779_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_437 net779_437/I _6790_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5801_ hold566/Z hold99/Z _5807_/S _7158_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ _6781_/D _7359_/RN _6781_/CLK _6781_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5732_ _5891_/A1 _5741_/A2 hold18/Z _5732_/A4 _5740_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3993_ _7362_/Q _7345_/Q _6955_/Q _3993_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_188_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5663_ hold99/Z hold295/Z _5668_/S _5663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4614_ _4452_/Z _5421_/C _5413_/A2 _4773_/C _5240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5594_ hold50/Z hold516/Z _5596_/S _5594_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7333_ _7333_/D _7341_/RN _4144_/I1 _7333_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4545_ _5295_/B2 _4691_/C _3399_/I _5162_/A2 _5517_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold401 _5691_/Z _7061_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold445 _5889_/Z _7234_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold434 _5880_/Z _7226_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold412 _5709_/Z _7077_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold423 _5736_/Z _7101_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _4485_/A4 _4447_/Z _4485_/A2 _4711_/B _4607_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold467 _7270_/Q hold467/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold478 _5875_/Z _7222_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7264_ _7264_/D _7286_/RN _7264_/CLK _7264_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold456 _5718_/Z _7085_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6215_ _7080_/Q _6293_/A2 _6294_/B1 _7104_/Q _6219_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold489 _5539_/Z _6928_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3427_ _3418_/Z hold82/I _3427_/B _3428_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7195_ hold45/Z _7243_/RN _7195_/CLK hold44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3358_ _7231_/Q _3358_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6146_ _6146_/A1 _6146_/A2 _6806_/Q _7305_/Q _6147_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ _6761_/Q _6299_/C _6265_/B1 _7165_/Q _6265_/C _6080_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_57_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5028_ _5028_/A1 _5028_/A2 _5028_/A3 _5032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6979_ _6979_/D _7286_/RN _6979_/CLK _6979_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet729_356 net729_357/I _6916_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_367 net729_367/I _6905_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet729_378 net429_99/I _6883_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_389 net729_389/I _6847_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4330_ hold363/Z hold711/Z _4337_/S _4330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ hold363/Z hold617/Z _4262_/S _4261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _5999_/Z _7296_/Q _6000_/B _6001_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ hold1/Z _7339_/Q _6881_/Q hold2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_67_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6902_ _6902_/D input75/Z _6902_/CLK _6902_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6833_ _6833_/D _7286_/RN _6833_/CLK _6833_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6764_ _6764_/D _7315_/RN _6764_/CLK _6764_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3976_ _6776_/Q hold185/I hold7/I _5882_/A2 _4012_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_11_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5715_ _4178_/Z hold908/Z _5722_/S _7082_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6695_ _7359_/RN _7012_/Q _4069_/C _6695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5646_ hold93/Z hold79/Z hold13/Z _7021_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _5750_/A3 _5777_/A2 _4178_/Z hold68/Z _5578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold220 _7134_/Q hold220/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold231 _7186_/Q hold231/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold253 _5943_/Z _7282_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4528_ _5417_/C _5162_/A2 _3399_/I _4698_/C _5534_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7316_ _7316_/D _7322_/RN _7319_/CLK _7316_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold242 _5746_/Z _7110_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4459_ _5214_/A4 _5295_/B2 _5322_/A2 _4693_/B _5030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7247_ _7247_/D _7315_/RN _7247_/CLK _7247_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold286 _4230_/Z _6765_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold275 _5906_/Z _7249_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold264 _7053_/Q hold264/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold297 _6828_/Q hold297/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7178_ hold47/Z _7300_/RN _7178_/CLK hold46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6129_ _7101_/Q _6294_/B1 _6291_/C1 _6997_/Q _6293_/B1 _7061_/Q _6132_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_56__1403_ net579_205/I net579_219/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3830_ _4405_/A3 _5872_/A3 _3830_/B _3830_/C _3853_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3761_ _3761_/A1 _3761_/A2 _3761_/A3 _3761_/A4 _3765_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5500_ _5500_/A1 _5440_/C _5500_/A3 _5502_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_173_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6480_ _7176_/Q _6310_/Z _6319_/Z _7256_/Q _7272_/Q _6610_/B1 _6481_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3692_ hold48/I _3771_/A2 _4024_/A2 hold46/I _3693_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5431_ _5431_/A1 _5431_/A2 _5431_/A3 _5432_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _5362_/A1 _4906_/C _5362_/A3 _5362_/A4 _5495_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput325 _6859_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput303 _4147_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput314 _6867_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4313_ _4312_/Z hold609/Z _4321_/S _4313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _7101_/D _7322_/RN _7101_/CLK _7101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput336 _6876_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5293_ _5293_/A1 _5293_/A2 _5440_/C _5348_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7032_ hold39/Z _7300_/RN _7032_/CLK _7032_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ hold323/Z hold832/Z _4244_/S _4244_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4175_ hold101/Z _4395_/A2 _4175_/B hold102/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_95_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6816_ _6816_/D _7300_/RN _6816_/CLK _7378_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6747_ _6747_/D input75/Z _6747_/CLK _6747_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3959_ _3915_/Z _3917_/Z _3959_/A3 _3959_/A4 _6622_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_149_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ hold363/Z hold841/Z _6679_/S _6678_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5629_ hold59/Z hold111/Z _5632_/S _5629_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_300 net629_301/I _6987_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _6302_/A1 _7291_/Q _6245_/C _5981_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4931_ _4456_/Z _5184_/A2 _4931_/B _5220_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_17_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4862_ _5228_/B _5460_/A1 _5214_/A4 _4454_/Z _5313_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_32_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6601_ _6601_/A1 _6601_/A2 _6601_/A3 _6607_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3813_ _7151_/Q _3981_/A2 _4024_/A2 _7175_/Q _3817_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4793_ _4793_/A1 _4793_/A2 _4711_/B _4961_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_165_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6532_ _7210_/Q _6316_/Z _6352_/Z hold52/I _6535_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3744_ _3720_/Z _3744_/A2 _3744_/A3 _3744_/A4 _3745_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3675_ _7258_/Q _3778_/A2 _4040_/A2 _7040_/Q _3677_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6463_ _7126_/Q _6308_/Z _6336_/Z _7102_/Q _6464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ _5414_/A1 _5414_/A2 _4483_/B _4792_/B _5415_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_127_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ _7229_/Q _6599_/A2 _6329_/Z _7011_/Q _6338_/Z _7075_/Q _6396_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xoutput177 _3374_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5345_ _5345_/A1 _5345_/A2 _5345_/A3 _5346_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_130_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput199 _4125_/ZN mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5276_ _5457_/A1 _5268_/B _5286_/A4 _5283_/A4 _5277_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_141_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput188 _3364_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4227_ hold99/Z hold508/Z _4232_/S _4227_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7015_ _7015_/D _7322_/RN _7015_/CLK _7015_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4158_ _4158_/A1 input73/Z _4158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _6355_/A4 _6343_/A4 _7299_/Q _7296_/Q _6340_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_55_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_167_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput68 mgmt_gpio_in[5] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold808 _7165_/Q hold808/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput79 spi_enabled _4128_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold819 _6849_/Q hold819/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3460_ _6796_/Q _3464_/A3 _7361_/Q _3461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3391_ _7319_/Q _6539_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5130_ _5406_/A1 _5287_/A2 _5130_/B1 _5206_/B _5494_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5061_ _4591_/C _4499_/B _5061_/A3 _5061_/A4 _5061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_96_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4012_ _7196_/Q _4012_/A2 _4012_/B1 _6786_/Q _4012_/C _4013_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5963_ _7285_/Q _7286_/Q _7287_/Q _7288_/Q _5963_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_80_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _5466_/A1 _5466_/A2 _5217_/B _5424_/A2 _5439_/A1 _4916_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_80_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ hold99/Z hold521/Z _5899_/S _5894_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4845_ _5497_/A2 _5322_/A2 _5295_/B2 _5133_/B _4846_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _3399_/I _5277_/A2 _5460_/A1 _5319_/A1 _4777_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6515_ _7088_/Q _6325_/Z _6326_/Z _7266_/Q _6521_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3727_ _7079_/Q _4006_/A2 _4010_/A2 _7087_/Q _3729_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _7199_/Q _6313_/Z _6331_/Z _7093_/Q _6335_/Z _7005_/Q _6447_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3658_ _3658_/A1 _3658_/A2 _3658_/A3 _3657_/Z _3658_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _6377_/A1 _6377_/A2 _6377_/A3 _6377_/A4 _6378_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_103_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3589_ _3884_/A1 _5808_/A2 _3521_/Z _5872_/A4 _3981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5328_ _5329_/A1 _5327_/Z _5398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ _5416_/B _5405_/A1 _5259_/B _5344_/C _5262_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_76_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_243 net579_243/I _7044_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_210 net779_415/I _7077_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_221 net579_221/I _7066_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_232 net629_286/I _7055_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_189_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4630_ _4630_/A1 _4630_/A2 _4630_/A3 _4630_/A4 _4633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_175_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4561_ _5322_/A2 _4751_/B _5162_/A2 _4762_/A4 _5473_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6300_ _7293_/Q _6297_/Z _6300_/B1 _6302_/A1 _6300_/C _6301_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xhold627 _4331_/Z _6832_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7280_ _7280_/D _7315_/RN _7280_/CLK _7280_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4492_ _3399_/I _5162_/A2 _4694_/B _4454_/Z _4603_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3512_ _3504_/Z _3509_/Z _5808_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold616 _5561_/Z _6953_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold605 _4425_/Z _6912_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold649 _5901_/Z _7244_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap368 _5490_/B _5421_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xmax_cap346 _5588_/A1 _5936_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xhold638 _7367_/Q hold638/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6231_ _6231_/A1 _6299_/C _7137_/Q _7290_/Q _6235_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3443_ _3448_/S _7365_/Q _3444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xmax_cap357 _5560_/A1 _5550_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_143_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _7208_/Q _6289_/A2 _6294_/B1 _7224_/Q _6166_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _5113_/A1 _5434_/A1 _5117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3374_ _7109_/Q _3374_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _7108_/Q _6294_/A2 _6290_/B1 _7044_/Q _6095_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _5406_/A1 _5450_/A2 _5401_/A2 _4974_/Z _5046_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _6995_/D _7243_/RN _6995_/CLK _6995_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5946_ _6808_/Q _4091_/B _5946_/B _7284_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _5881_/S _5877_/A2 _5877_/B hold576/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4828_ _5133_/C _5322_/A2 _5295_/B2 _5133_/B _4830_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_138_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet529_173 net429_81/I _7114_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_162 net629_301/I _7125_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4759_ _5491_/A1 _5491_/A2 _4759_/A3 _4759_/A4 _4760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet529_195 net579_221/I _7092_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_184 net529_184/I _7103_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _6613_/A2 _6429_/A2 _6429_/A3 _6428_/Z _6430_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_150_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150__41 _4150__46/I _7246_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__30 _4150__46/I _7257_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold2 hold2/I hold2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_54_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet779_405 net779_414/I _6831_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_416 net779_416/I _6820_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_427 net779_427/I _6809_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_438 net779_438/I _6789_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet779_449 net829_475/I _6778_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6780_ _6780_/D _7359_/RN _6780_/CLK _6780_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5800_ hold892/Z hold323/Z _5807_/S _7157_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3992_ _6909_/Q hold83/I _5557_/A2 _4426_/A3 _4036_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_95_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ hold2/Z hold121/Z _5731_/S _5731_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5662_ hold323/Z hold742/Z _5668_/S _7035_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ hold59/Z hold544/Z _5596_/S _5593_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4613_ _4613_/A1 _4613_/A2 _5074_/C _4620_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7332_ _7332_/D _7341_/RN _4144_/I1 _7332_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold402 _6982_/Q hold402/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4544_ _5322_/A2 _4751_/B _5475_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_117_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7263_ _7263_/D _7315_/RN _7263_/CLK _7263_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold413 _7396_/I hold413/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold435 _7069_/Q hold435/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold424 _6742_/Q hold424/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4475_ _4485_/A4 _4447_/Z _4485_/A2 _4711_/B _4523_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold468 _5930_/Z _7270_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold457 _7264_/Q hold457/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _7056_/Q _6291_/A2 _6295_/B1 hold74/I _6289_/A2 _7088_/Q _6220_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold446 _6749_/Q hold446/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold479 _7272_/Q hold479/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3426_ _3426_/A1 _6795_/Q _3426_/B hold81/I _3427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7194_ _7194_/D _7243_/RN _7194_/CLK _7194_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3357_ _7239_/Q _3357_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6145_ _6806_/Q _6145_/A2 _6146_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6076_ _6076_/I _6086_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _5238_/B1 _4796_/Z _5401_/A2 _5401_/A3 _5028_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6978_ _6978_/D _7286_/RN _6978_/CLK _6978_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ hold323/Z hold715/Z _5935_/S _5929_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2_0__1403_ clkbuf_0__1403_/Z clkbuf_4_5_0__1403_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_28_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16__1403_ clkbuf_4_10_0__1403_/Z _4150__40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_157_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet729_357 net729_357/I _6915_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_79__1403_ clkbuf_4_5_0__1403_/Z net779_423/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet729_379 net429_99/I _6882_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet729_368 net729_369/I _6904_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _5891_/A4 hold185/Z _5812_/A2 _6677_/A3 _4262_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4191_ hold38/Z hold306/Z _4193_/S _4191_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6901_ _6901_/D input75/Z _6901_/CLK _6901_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _6832_/D _7286_/RN _6832_/CLK _6832_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6763_ _6763_/D _7315_/RN _6763_/CLK _6763_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3975_ _6911_/Q _5560_/A1 _5732_/A4 _4423_/A2 _4005_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5714_ _5891_/A1 _5741_/A2 _5780_/A3 hold18/Z _5722_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_31_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6694_ _7359_/RN _7012_/Q _4069_/C _6694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ hold373/Z hold99/Z hold13/Z _7020_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5576_ _5585_/A2 _5576_/A2 _5576_/B hold667/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold210 _6735_/Q hold210/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold243 _7257_/Q hold243/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4527_ _4097_/B _4711_/B _4715_/B _5417_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold232 _5834_/Z _7186_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7315_ _7315_/D _7315_/RN _7319_/CLK _7315_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold221 _5773_/Z _7134_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7246_ _7246_/D _7286_/RN _7246_/CLK _7246_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4458_ _3399_/I _4694_/B _4787_/B _4454_/Z _4932_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold254 _7209_/Q hold254/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold265 _6944_/Q hold265/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold276 _7102_/Q hold276/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold287 _7017_/Q hold287/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ hold64/Z _7300_/RN _7177_/CLK hold63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold298 _7004_/Q hold298/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3409_ _6727_/Q _6726_/Q _6725_/Q _3409_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4389_ _6896_/Q _6897_/Q _6898_/Q _6666_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6128_ _6128_/A1 _6128_/A2 _6133_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ _6231_/A1 _6245_/C _7291_/Q _7290_/Q _6293_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3__1403_ clkbuf_4_3_0__1403_/Z net429_74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _6990_/Q _4038_/A2 _4020_/A2 _7240_/Q _3761_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _4395_/C _5430_/A2 _5430_/A3 _5430_/B _6924_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3691_ _7194_/Q _3930_/A2 _4020_/B1 _7162_/Q _3693_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5361_ _5361_/A1 _5361_/A2 _5361_/A3 _5361_/A4 _5432_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput326 _6860_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput304 _4146_/Z serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput315 _6868_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4312_ hold148/Z hold79/Z _4320_/S _4312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5292_ _5497_/A2 _5440_/A2 _5440_/B1 _5228_/B _5497_/C _5293_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7100_ _7100_/D _7322_/RN _7100_/CLK _7100_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_5_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput337 _6877_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _7031_/D _7300_/RN _7031_/CLK hold57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4243_ hold363/Z hold786/Z _4244_/S _4243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4174_ _7342_/Q _6881_/Q _4175_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _6815_/D _7300_/RN _6815_/CLK _6815_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6746_ _6746_/D input75/Z _6746_/CLK _6746_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3958_ _3958_/A1 _3958_/A2 _3958_/A3 _3958_/A4 _3959_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_129_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6677_ _6677_/A1 _6677_/A2 _6677_/A3 _6679_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3889_ _6900_/Q _5891_/A4 _5560_/A1 _4408_/A1 _3918_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ hold79/Z hold119/Z _5632_/S _5628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5559_ hold323/Z hold739/Z _5559_/S _5559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet629_301 net629_301/I _6986_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _7229_/D _7315_/RN _7229_/CLK _7229_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_105_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_183_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _5294_/B _4691_/C _4751_/B _3399_/I _4931_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_92_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _5439_/A1 _5344_/C _5359_/A2 _5350_/A2 _4863_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3812_ _7037_/Q _4040_/A2 _4037_/A2 _7207_/Q _3818_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6600_ _6789_/Q _6313_/Z _6331_/Z _6910_/Q _6335_/Z _6852_/Q _6601_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4792_ _4792_/A1 _4792_/A2 _4792_/B _4961_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_159_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6531_ _7104_/Q _6336_/Z _6342_/Z _7250_/Q _6535_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3743_ _3743_/A1 _3743_/A2 _3743_/A3 _3743_/A4 _3744_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xclkbuf_4_5_0__1403_ clkbuf_4_5_0__1403_/I clkbuf_4_5_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_146_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3674_ input69/Z _4303_/S _4285_/S input50/Z _4046_/A2 _7032_/Q _3677_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6462_ _7118_/Q _6594_/A2 _6594_/A3 _6594_/A4 _6464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5413_ _5228_/B _5413_/A2 _5413_/B _5413_/C _5414_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6393_ _7051_/Q _6324_/Z _6393_/B _6393_/C _6396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5344_ _5417_/A2 _5416_/B _5344_/B _5344_/C _5345_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput167 _4164_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5275_ _5360_/A1 _5273_/Z _5360_/A3 _5279_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput178 _6138_/A1 mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput189 _3363_/ZN mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4226_ hold323/Z hold829/Z _4232_/S _4226_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7014_ _7014_/D _7286_/RN _7014_/CLK _7014_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4157_ input85/Z input58/Z _7362_/Q _4157_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4088_ _6328_/A4 _7297_/Q _6566_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_83_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6729_ _6729_/D _7243_/RN _6729_/CLK _6729_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_165_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold809 _7139_/Q hold809/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput69 mgmt_gpio_in[6] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_124_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3390_ _7318_/Q _6512_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5060_ _4693_/B _5172_/A1 _5060_/B _5060_/C _5369_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_123_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4011_ _4011_/A1 _4011_/A2 _4011_/A3 _4011_/A4 _4011_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_84_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _5952_/B _6017_/A3 _5959_/B _5964_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_92_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4913_ _5461_/A4 _5206_/B _5218_/B _5322_/A2 _5507_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5893_ hold323/Z hold806/Z _5899_/S _7237_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4844_ _4844_/A1 _4844_/A2 _4846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _5268_/B _5305_/B _4839_/A3 _5286_/A4 _4775_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_147_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6514_ _7202_/Q _6313_/Z _6610_/A2 _7282_/Q _6521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3726_ _6991_/Q _4038_/A2 _4020_/B1 _7161_/Q _3729_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _7231_/Q _6599_/A2 _6329_/Z _7013_/Q _6338_/Z _7077_/Q _6447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3657_ _3654_/Z _3657_/A2 _3657_/A3 _3657_/A4 _3657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_173_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6376_ _7058_/Q _6376_/A2 _6387_/A1 _6540_/A4 _6377_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3588_ _5872_/A2 _3509_/Z _3504_/Z _5808_/A3 _4014_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5327_ _5384_/A2 _5327_/A2 _5327_/A3 _5327_/A4 _5327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_115_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _5099_/B _5099_/C _5344_/C _5405_/A1 _5481_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_102_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _5482_/C _5384_/A1 _5300_/B _5190_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4209_ hold446/Z hold50/Z _4211_/S _4209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_211 net629_297/I _7076_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_222 net629_272/I _7065_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_233 net629_266/I _7054_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_244 _4150__48/I _7043_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _5214_/A4 _5460_/A1 _5295_/B2 _4691_/C _5228_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_129_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold606 _6819_/Q hold606/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4491_ _4715_/B _5384_/B _4097_/B _5259_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_129_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold617 _6786_/Q hold617/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3511_ _3556_/B _3548_/B _5891_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xmax_cap369 _3400_/I _5162_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold628 _6881_/Q _4178_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_155_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3442_ _3421_/B _6792_/Q _7366_/Q _3444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold639 hold639/I hold639/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap358 hold185/Z _5560_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6230_ _6230_/A1 _6230_/A2 _6230_/A3 _6236_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_171_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3373_ _7117_/Q _6138_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6161_ _7134_/Q _6295_/B1 _6291_/C1 _7126_/Q _6167_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _5112_/A1 _5406_/A1 _5130_/B1 _5462_/A4 _5434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6092_ _6434_/S _6092_/A2 _6092_/B _7304_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _5038_/Z _5043_/A2 _5043_/A3 _5047_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0_wbbd_sck _7340_/Q clkbuf_0_wbbd_sck/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _6994_/D _7286_/RN _6994_/CLK _6994_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_81_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5945_ _5999_/I0 _6808_/Q _5945_/B _7284_/Q _5946_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5876_ hold574/Z _5882_/A2 hold310/Z hold79/Z hold575/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4827_ _5283_/A2 _5286_/A2 _5104_/B1 _5133_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_139_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet529_163 net629_301/I _7124_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet529_152 net679_333/I _7135_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _5441_/A4 _4835_/A1 _4758_/A3 _4758_/A4 _5104_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_147_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet529_174 net629_298/I _7113_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_196 net679_330/I _7091_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_185 net679_333/I _7102_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4689_ _5259_/B _4689_/A2 _4641_/C _5339_/A1 _4690_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3709_ _7249_/Q _4019_/A2 _4045_/A2 _7055_/Q _3711_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6428_ _6428_/A1 _6428_/A2 _6428_/A3 _6428_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_162_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6359_ _7204_/Q _6316_/Z _6609_/B1 _7042_/Q _6317_/Z _7220_/Q _6365_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_108_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150__42 net429_80/I _7245_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_39__1403_ clkbuf_4_14_0__1403_/Z net579_243/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4150__31 _4150__48/I _7256_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__20 net429_55/I _7267_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold3 hold3/I hold3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_119__1403_ clkbuf_4_2_0__1403_/Z net829_475/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet779_417 net779_419/I _6819_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_406 net779_431/I _6830_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_439 net829_455/I _6788_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_428 net779_430/I _6804_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ _6882_/Q _4408_/A1 _4426_/A3 _4048_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5730_ hold38/Z hold197/Z _5731_/S _5730_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7400_ _7400_/I _7400_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ hold363/Z hold790/Z _5668_/S _7034_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _4518_/Z _5417_/C _5475_/A1 _5359_/A1 _5074_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5592_ hold79/Z hold538/Z _5596_/S _5592_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4543_ _5295_/B2 _4691_/C _5319_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7331_ _7331_/D _7331_/CLK _7331_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7262_ _7262_/D _7315_/RN _7262_/CLK _7262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold436 _7118_/Q hold436/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold403 _5602_/Z _6982_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold414 _5596_/Z _6977_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold425 _4201_/Z _6742_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold458 _5923_/Z _7264_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4474_ _4523_/A2 _4792_/B _4607_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold469 _7281_/Q hold469/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6213_ _7072_/Q _6292_/B1 _6291_/B1 _7032_/Q _6220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold447 _4209_/Z _6749_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3425_ hold81/Z _6795_/Q _3425_/B hold82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7193_ _7193_/D _7243_/RN _7193_/CLK _7193_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3356_ _7247_/Q _3356_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6144_ _6302_/A1 _6302_/A2 _6989_/Q _7293_/Q _6145_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_58_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6075_ _7043_/Q _6290_/B1 _7293_/Q _6076_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xload_slew361 _5836_/A3 _5827_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xload_slew350 _5827_/A3 _5891_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_58_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _5482_/A2 _4796_/Z _5401_/A2 _5401_/A3 _5028_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0__1085_ _3785_/ZN clkbuf_0__1085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _6977_/D _7359_/RN _6977_/CLK _7396_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ hold363/Z hold747/Z _5935_/S _5928_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ hold59/Z hold356/Z _5862_/S _5859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_358 net729_359/I _6914_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet729_369 net729_369/I _6903_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4190_ hold37/Z _7338_/Q _6881_/Q hold38/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_113_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _6900_/D _7359_/RN _6900_/CLK _6900_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6831_ _6831_/D _7286_/RN _6831_/CLK _6831_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6762_ _6762_/D _7315_/RN _6762_/CLK _6762_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3974_ _6953_/Q _5560_/A1 _5732_/A4 _5566_/A1 _4007_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ hold2/Z hold438/Z _5713_/S _7081_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6693_ _7359_/RN _7012_/Q _4069_/C _6693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_176_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ hold815/Z hold323/Z hold13/Z _7019_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7314_ _7314_/D _7322_/RN _7319_/CLK _7314_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold200 _5748_/Z _7112_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold211 _4193_/Z _6735_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5575_ hold671/Z hold323/Z _5575_/S _6962_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold244 _7241_/Q hold244/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold233 _7210_/Q hold233/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4526_ _4483_/B _4792_/B _4929_/A3 _4929_/A2 _5490_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold222 _6961_/Q hold222/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7245_ _7245_/D _7315_/RN _7245_/CLK _7245_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4457_ _3399_/I _4751_/B _4691_/C _5460_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold255 _5860_/Z _7209_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold266 _5549_/Z _6944_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold277 _5737_/Z _7102_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold299 _5627_/Z _7004_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3408_ _7353_/Q _3472_/A2 _4063_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7176_ _7176_/D _7300_/RN _7176_/CLK _7176_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold288 _5641_/Z _7017_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6127_ _7077_/Q _6293_/A2 _6292_/A2 _7013_/Q _6128_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4388_ _6628_/I0 _6880_/Q _4388_/S _6880_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3339_ _7287_/Q _5959_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22__1403_ clkbuf_4_9_0__1403_/Z net429_83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6058_ _6058_/A1 _6058_/A2 _6058_/B1 _6058_/B2 _6063_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_102__1403_ clkbuf_4_1_0__1403_/Z net729_387/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _4796_/Z _4974_/Z _5024_/A4 _5336_/A3 _5010_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_73_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_85__1403_ net629_288/I net629_286/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3690_ hold53/I _4046_/B1 _4009_/B1 _7112_/Q _3693_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _5360_/A1 _5360_/A2 _5360_/A3 _5360_/A4 _5360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_114_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput305 _4163_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput316 _6869_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5291_ _5417_/A2 _5368_/A2 _5291_/B _5291_/C _5497_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_160_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _4310_/Z hold606/Z _4321_/S _4311_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput327 _7324_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput338 _6878_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7030_ hold60/Z _7300_/RN _7030_/CLK _7030_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4242_ _6677_/A1 _4426_/A3 _6677_/A3 _4244_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_141_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _7359_/RN _7012_/Q _4069_/C _4173_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_83_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _6814_/D _7300_/RN _6814_/CLK _7377_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3957_ _3957_/A1 _3957_/A2 _3957_/A3 _3957_/A4 _3958_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6745_ _6745_/D _7300_/RN _6745_/CLK _6745_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_137_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6676_ _5320_/C _6616_/Z _6676_/A3 _6676_/B _7341_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_149_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3888_ _5576_/A2 _5750_/A4 _3533_/Z _3986_/A3 _4042_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5627_ hold99/Z hold298/Z _5632_/S _5627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5558_ hold363/Z hold760/Z _5559_/S _5558_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4509_ _4603_/A1 _4603_/A2 _4641_/C _4591_/C _4688_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_117_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _7228_/D _7315_/RN _7228_/CLK _7228_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_120_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5489_ _5481_/Z _5489_/A2 _5504_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7159_ _7159_/D _7315_/RN _7159_/CLK _7159_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _5466_/A1 _5460_/A3 _5324_/A4 _5344_/C _5413_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_177_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3811_ _7239_/Q _4020_/A2 _4038_/B1 _7013_/Q _3818_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4791_ _4442_/Z _4444_/Z _4447_/Z _4790_/Z _4927_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_177_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _6530_/A1 _6530_/A2 _6530_/A3 _6530_/A4 _6530_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_32_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3742_ _3742_/A1 _3742_/A2 _3742_/A3 _3743_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6461_ _7264_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6472_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3673_ _3673_/A1 _3673_/A2 _3673_/A3 _3673_/A4 _3673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_173_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5412_ _5193_/C _5412_/A2 _5412_/A3 _5412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6392_ _6392_/A1 _6392_/A2 _6392_/A3 _6393_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5343_ _5343_/A1 _5343_/A2 _5405_/B _5343_/A4 _5345_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput168 _7373_/Z irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5274_ _5457_/A1 _5324_/A3 _5274_/B _5360_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput179 _3372_/ZN mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4225_ hold363/Z hold856/Z _4232_/S _4225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7013_ _7013_/D _7243_/RN _7013_/CLK _7013_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_68_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4156_ _4156_/I _4156_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4087_ _6007_/B _7298_/Q _6593_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_56_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4989_ _4989_/A1 _4989_/A2 _4989_/A3 _4996_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6728_ _6728_/D _7300_/RN _6728_/CLK _6728_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6659_ _6659_/A1 _6659_/A2 _6660_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _7082_/Q _4010_/A2 _4010_/B1 _7114_/Q _4011_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ _5961_/A1 _7288_/Q _5965_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4912_ _5066_/B2 _5344_/C _5313_/A1 _5182_/C _4912_/C _4916_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_52_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5892_ hold363/Z hold871/Z _5899_/S _7236_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4843_ _5344_/C _5359_/A2 _5291_/C _4843_/B1 _5339_/A1 _4844_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_61_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4774_ _5268_/B _5305_/B _4839_/A3 _5286_/A4 _5277_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_159_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6513_ hold46/I _6310_/Z _6347_/C _7242_/Q _6521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3725_ hold76/I _3771_/A2 _4009_/A2 _7063_/Q _3729_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6444_ _7053_/Q _6324_/Z _6444_/B _6444_/C _6447_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_161_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3656_ hold44/I _3930_/A2 _4047_/A2 hold27/I _4024_/A2 hold25/I _3657_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6375_ _6994_/Q _6376_/A2 _6594_/A4 _6540_/A4 _6377_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3587_ _3906_/A1 _5808_/A2 _3509_/Z _5872_/A3 _3771_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5326_ _5333_/A1 _5333_/A2 _5326_/B _5326_/C _5329_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_161_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5257_ _5257_/A1 _5480_/A4 _5262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4208_ hold396/Z hold59/Z _4211_/S _4208_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5188_ _5310_/A1 _5461_/A3 _4787_/B _4694_/B _5518_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4139_ _7012_/Q _7343_/Q _4069_/C _4140_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_223 net579_240/I _7064_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_212 net629_298/I _7075_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_234 net729_389/I _7053_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_189_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_245 _4150__51/I _7042_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3510_ _6881_/Q hold21/Z _3556_/C _3548_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_171_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold607 _4311_/Z _6819_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4490_ _4483_/B _4929_/A3 _4929_/A2 _5099_/B _5093_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold618 _4261_/Z _6786_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold629 _5937_/Z _7276_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3441_ _7367_/Q _3441_/I1 _3448_/S _7367_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3372_ _7125_/Q _3372_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6160_ _6160_/A1 _6160_/A2 _6160_/A3 _6160_/A4 _6170_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5111_ _5112_/A1 _5440_/A2 _5111_/B1 _5105_/C _5111_/C _5113_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6091_ _5951_/B _6614_/B _7304_/Q _6092_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _5461_/A1 _5515_/A1 _5510_/A2 _5450_/A2 _5043_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ _6993_/D _7322_/RN _6993_/CLK hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_19_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5944_ hold2/Z hold137/Z _5944_/S _5944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ hold477/Z hold99/Z _5881_/S _5875_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4826_ _5214_/A4 _5295_/B2 _5322_/A2 _5162_/A2 _5134_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xnet529_164 net429_71/I _7123_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_153 _4150__44/I _7134_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4757_ _5421_/A2 _5138_/B _4835_/A1 _5441_/A4 _4759_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet529_186 net579_221/I _7101_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_175 net629_296/I _7112_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet529_197 net429_87/I _7090_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _4688_/A1 _5384_/B _5098_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ input17/Z _4031_/A2 _3947_/B1 _7007_/Q _3711_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6427_ _7278_/Q _6610_/A2 _6347_/C _7238_/Q _6428_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3639_ _7275_/Q _3921_/A2 _4046_/A2 _7033_/Q _4047_/B1 _7147_/Q _3659_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_89_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6358_ _7098_/Q _6336_/Z _6352_/Z _7148_/Q _6370_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5309_ _5320_/A1 _5493_/A1 _5309_/B _5421_/C _5422_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _6908_/Q _6289_/A2 _6289_/B1 _6872_/Q _6297_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_153_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150__10 _4150__9/I _7277_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__43 net429_80/I _7244_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__32 net429_80/I _7255_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__21 _4150__22/I _7266_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold4 hold4/I hold4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_94_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_418 net779_418/I _6818_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_407 net779_430/I _6829_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet779_429 net779_430/I _6803_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3990_ _6964_/Q _3561_/B _5909_/A2 _6677_/A2 _4018_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5660_ _5891_/A1 _5678_/A2 _5891_/A3 _5732_/A4 _5668_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_176_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _4773_/C _4694_/B _4787_/B _4702_/B _5359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_31_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ hold99/Z hold546/Z _5596_/S _5591_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4542_ _5421_/C _5322_/A2 _5295_/B2 _5462_/A2 _5066_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_128_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7330_ _7330_/D _7331_/CLK _7330_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4473_ _4960_/A1 _4485_/A2 _4711_/B _5368_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7261_ _7261_/D _7315_/RN _7261_/CLK _7261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold426 _7199_/Q hold426/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold415 _7162_/Q hold415/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold404 _6746_/Q hold404/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold437 _5755_/Z _7118_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6212_ _7096_/Q _6290_/A2 _6290_/B1 _7048_/Q _6220_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3424_ _3426_/A1 _6795_/Q _3425_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold459 _6770_/Q hold459/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold448 _7001_/Q hold448/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _7192_/D _7243_/RN _7192_/CLK _7192_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3355_ _7255_/Q _3355_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ _7293_/Q _6143_/A2 _6143_/B _6143_/C _6146_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xload_slew351 _5827_/A3 _5882_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xload_slew362 hold641/Z _5836_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6074_ _6074_/A1 _6074_/A2 _6074_/A3 _6073_/Z _6074_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _5025_/A1 _5025_/A2 _5025_/B _5028_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _6976_/D _7359_/RN _6976_/CLK _7395_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5927_ _5936_/A1 hold18/Z _5927_/A3 _4305_/C _5935_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_70_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5858_ hold79/Z hold377/Z _5862_/S _5858_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4809_ _4809_/A1 _4809_/A2 _5431_/A1 _4809_/A4 _4815_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _6677_/A3 _5818_/A2 _5863_/A3 _5863_/A4 hold33/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_45__1403_ clkbuf_4_15_0__1403_/Z net779_404/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_175_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet729_359 net729_359/I _6913_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _6830_/D _7359_/RN _6830_/CLK _6830_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6761_ _6761_/D _7315_/RN _6761_/CLK _6761_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5712_ hold38/Z hold481/Z _5713_/S _7080_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3973_ _6919_/Q _4435_/A1 hold83/I _5557_/A2 _4005_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_189_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _7359_/RN _7012_/Q _4069_/C _6692_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5643_ hold780/Z hold363/Z hold13/Z _7018_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ hold222/Z hold38/Z _5575_/S _6961_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4525_ _4792_/B _4929_/A3 _4929_/A2 _4890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7313_ _7313_/D _7322_/RN _7319_/CLK _7313_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold201 _7152_/Q hold201/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold234 _5861_/Z _7210_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold223 _6838_/Q hold223/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold212 _6991_/Q hold212/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7244_ _7244_/D _7315_/RN _7244_/CLK _7244_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4456_ _3399_/I _4751_/B _4691_/C _4456_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold245 _5897_/Z _7241_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold278 _7265_/Q hold278/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold256 _7151_/Q hold256/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold267 _7175_/Q hold267/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold289 _7119_/Q hold289/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_98_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7175_ _7175_/D input75/Z _7175_/CLK _7175_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3407_ _7355_/Q _7354_/Q _3472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4387_ _6627_/I0 _6879_/Q _4388_/S _6879_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3338_ _7286_/Q _6017_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6126_ _7069_/Q _6292_/B1 _6291_/B1 hold90/I _6128_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6057_ _6057_/A1 _6057_/A2 _6057_/A3 _6057_/A4 _6058_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5008_ _5008_/A1 _5008_/A2 _5008_/A3 _5008_/A4 _5010_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_73_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6959_ _6959_/D _7300_/RN _6959_/CLK _6959_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold790 _7034_/Q hold790/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4152_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput306 _4158_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput317 _6870_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4310_ hold180/Z hold99/Z _4320_/S _4310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5290_ _5290_/A1 _5498_/C _5293_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput328 _7325_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_91__1403_ clkbuf_4_4_0__1403_/Z net429_95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput339 _6879_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ hold323/Z hold749/Z _4241_/S _4241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4172_ _4172_/A1 _6897_/Q _6890_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6813_ _6813_/D _7300_/RN _6813_/CLK _7376_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3956_ _7277_/Q _4027_/A2 _4027_/B1 _7253_/Q _3957_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6744_ _6744_/D _7300_/RN _6744_/CLK _6744_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _7341_/Q _6894_/Q _6675_/B _6676_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3887_ _5808_/A4 _5808_/A2 _3523_/B _3554_/B _4028_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5626_ hold323/Z hold683/Z _5632_/S _7003_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5557_ _5900_/A3 _5557_/A2 _5891_/A1 hold68/Z _5559_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_145_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ _5061_/A3 _4508_/A2 _4508_/A3 _4641_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_105_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ _5488_/A1 _5484_/Z _5523_/A3 _5489_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_160_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7227_ _7227_/D _7286_/RN _7227_/CLK _7227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4439_ _4483_/B _4792_/B _4929_/A3 _4929_/A2 _4795_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7158_ _7158_/D _7315_/RN _7158_/CLK _7158_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_59_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _7198_/Q _6293_/A2 _6292_/A2 _6762_/Q _6110_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7089_ hold89/Z _7322_/RN _7089_/CLK hold88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _4702_/B _5305_/B _4787_/B _5030_/A2 _4790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_33_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _6958_/Q _4045_/B1 _3855_/B1 _6943_/Q _6739_/Q _4040_/B1 _3818_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3741_ _7023_/Q _4041_/A2 _3778_/A2 _7257_/Q _3742_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3672_ input41/Z _4320_/S _4015_/A2 _7048_/Q _3673_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6460_ _6460_/A1 _6460_/A2 _6434_/S _6460_/B2 _7316_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5411_ _5417_/A2 _5457_/A1 _5417_/C _5533_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_115_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6391_ _7131_/Q _6315_/Z _6316_/Z _7205_/Q _6392_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5342_ _5440_/A2 _5342_/A2 _5450_/A2 _5401_/A2 _5405_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_127_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ _5435_/A1 _5271_/Z _5435_/A2 _5273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7012_ _7012_/D _7286_/RN _7012_/CLK _7012_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_88_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput169 _4165_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4224_ _4305_/C _5812_/A2 hold32/Z _5927_/A3 _4232_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_114_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4155_ _4158_/A1 input86/Z _4156_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _6387_/A2 _7294_/Q _6543_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4988_ _5238_/B1 _4796_/Z _5336_/A2 _5331_/A3 _4989_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6727_ _6727_/D _6682_/Z _7364_/CLK _6727_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3939_ _7237_/Q _4020_/A2 _3939_/B1 _6781_/Q input15/Z _4043_/A2 _3950_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6658_ _6896_/Q _6658_/A2 _6658_/B1 _6666_/B2 _6659_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ hold99/Z hold476/Z hold69/Z _6988_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6589_ _5951_/B _7320_/Q _4083_/B _6806_/Q _6590_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5960_ _5960_/A1 _5960_/A2 _7287_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_92_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4911_ _4691_/C _5461_/A4 _5510_/A2 _5184_/A2 _5182_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5891_ _5891_/A1 _5891_/A2 _5891_/A3 _5891_/A4 _5899_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4842_ _4842_/A1 _4842_/A2 _4842_/A3 _4842_/A4 _4844_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4773_ _4702_/B _4773_/A2 _4773_/B1 _5305_/C _4773_/C _5283_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_186_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _6512_/A1 _6512_/A2 _6434_/S _6512_/B2 _7318_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3724_ _7103_/Q _4006_/B1 _4008_/A2 _7095_/Q _4019_/B1 _6950_/Q _3744_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_173_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6443_ _6443_/A1 _6443_/A2 _6443_/A3 _6443_/A4 _6444_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_107_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _7137_/Q _4046_/B1 _4038_/A2 hold77/I _4020_/B1 _7163_/Q _3657_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6374_ _7002_/Q _6543_/A2 _6594_/A4 _6540_/A4 _6377_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3586_ _5909_/A2 hold68/Z _3868_/A1 _5808_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5325_ _5326_/C _5325_/A2 _4953_/Z _5396_/B1 _5476_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_114_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5256_ _5482_/B _5384_/B _5384_/C _5482_/A2 _5480_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_88_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ hold398/Z hold79/Z _4211_/S _4207_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5187_ _5304_/A1 _5234_/A2 _5416_/B _5268_/B _5310_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_84_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _6809_/Q input3/Z input1/Z _4138_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ _7360_/Q _7342_/Q _7012_/Q _4069_/C _4172_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_56_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet579_202 net579_219/I _7085_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_224 net629_272/I _7063_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_213 net579_213/I _7074_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_246 net779_426/I _7041_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_235 net629_286/I _7052_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_9__1403_ clkbuf_4_9_0__1403_/Z net429_91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold608 _7052_/Q hold608/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_183_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold619 _6787_/Q hold619/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3440_ _6795_/Q _3416_/Z _3440_/A3 _3440_/B _3441_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xmax_cap349 _5812_/A2 _6677_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3371_ _7133_/Q _3371_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _5417_/B _5268_/B _5134_/A4 _5473_/A2 _5272_/B _5435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6090_ _6090_/A1 _6090_/A2 _6806_/Q _7303_/Q _6092_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _5450_/A1 _5450_/A2 _5039_/Z _5525_/A1 _5043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6992_ hold70/Z _7286_/RN _6992_/CLK _6992_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5943_ hold38/Z hold252/Z _5944_/S _5943_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5874_ hold858/Z hold323/Z _5881_/S _5874_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _5460_/A1 _4751_/B _4691_/C _3399_/I _5216_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_33_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet529_154 net779_404/I _7133_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4756_ _4839_/A3 _4839_/A2 _4839_/A4 _5421_/A2 _5104_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet529_176 net629_301/I _7111_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_187 net579_207/I _7100_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_198 net579_217/I _7089_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_165 net829_457/I _7122_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ _5260_/C _5097_/B _4690_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3707_ input31/Z _4043_/A2 _4017_/B1 _7400_/I _3711_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ _7174_/Q _6310_/Z _6321_/Z _7020_/Q _6428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3638_ _3906_/A1 _5808_/A2 _3509_/Z _5872_/A3 _4047_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_161_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6357_ _7034_/Q _6312_/Z _6323_/Z _7140_/Q _6364_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3569_ _3504_/Z _3509_/Z _3884_/A1 _3554_/B _5909_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5308_ _5310_/A1 _5312_/A1 _5308_/B _5514_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6288_ _6284_/Z _6288_/A2 _6288_/A3 _6288_/A4 _6301_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _5395_/A1 _5380_/B _5239_/A3 _4796_/Z _5240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_124_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_68__1403_ clkbuf_4_7_0__1403_/Z net579_213/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150__33 net429_82/I _7254_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__22 _4150__22/I _7265_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__11 _4150__9/I _7276_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150__44 _4150__44/I _7243_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold5 hold5/I hold5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_0_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet779_408 net779_411/I _6828_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet779_419 net779_419/I _6817_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ _4500_/B _4693_/B _5310_/B _5305_/B _5410_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_175_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5590_ hold323/Z hold838/Z _5596_/S _5590_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4541_ _5417_/C _4691_/C _4751_/B _4518_/Z _5209_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7260_ _7260_/D _7315_/RN _7260_/CLK _7260_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4472_ _5305_/B _4960_/A1 _4452_/Z _5395_/A1 _4523_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_171_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold427 _5849_/Z _7199_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold416 _7273_/Q hold416/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold405 _4206_/Z _6746_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6211_ _7120_/Q _6265_/C _6299_/B _6299_/C _6221_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3423_ _3423_/I0 _7371_/Q _3423_/S _7371_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7191_ _7191_/D input75/Z _7191_/CLK _7191_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold449 _5623_/Z _7001_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold438 _7081_/Q hold438/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6142_ _6142_/A1 _6142_/A2 _6142_/B1 _6142_/B2 _6143_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3354_ _7314_/Q _6408_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6073_ _6073_/A1 _6073_/A2 _6073_/A3 _6073_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _4796_/Z _5401_/A2 _5401_/A3 _5024_/A4 _5025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6975_ _6975_/D _7359_/RN _6975_/CLK _7394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ hold2/Z hold162/Z _5926_/S _5926_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5857_ hold99/Z hold514/Z _5862_/S _5857_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _4691_/C _5287_/A1 _5284_/A2 _4809_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_166_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5788_ hold2/Z _7147_/Q hold23/Z hold24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4739_ _5214_/A4 _5295_/B2 _5322_/A2 _5162_/A2 _5406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _7044_/Q _6566_/A2 _6593_/A3 _6540_/A4 _6429_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7389_ _7389_/I _7389_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6760_ _6760_/D _7315_/RN _6760_/CLK _6760_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xclkbuf_leaf_51__1403_ clkbuf_4_15_0__1403_/Z net779_419/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ hold50/Z hold529/Z _5713_/S _7079_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3972_ _6770_/Q _5560_/A1 _5780_/A3 _6677_/A1 _4040_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6691_ _7359_/RN _7012_/Q _4069_/C _6691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_176_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5642_ hold102/I hold12/Z _5642_/A3 _5872_/A3 hold13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5573_ hold219/Z hold50/Z _5575_/S _6960_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4524_ _5441_/A4 _4607_/A3 _4607_/A2 _5441_/A3 _5304_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_129_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold202 _7024_/Q hold202/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7312_ _7312_/D _7322_/RN _7322_/CLK _7312_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold213 _7250_/Q hold213/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold224 _4337_/Z _6838_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold235 _7086_/Q hold235/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4455_ _4751_/B _4691_/C _4698_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_171_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold246 _7266_/Q hold246/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold257 _6943_/Q hold257/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold268 _5822_/Z _7175_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7243_ hold56/Z _7243_/RN _7243_/CLK hold55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3406_ _4787_/B _5310_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_12
Xhold279 _5924_/Z _7265_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7174_ _7174_/D _7300_/RN _7174_/CLK _7174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4386_ _3745_/Z _6878_/Q _4388_/S _6878_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3337_ _7285_/Q _5952_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_105_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6125_ _6125_/A1 _6268_/A1 _6125_/B _6125_/C _6142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6056_ _7204_/Q _6289_/A2 _6292_/B1 _7188_/Q _6057_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _5395_/A1 _5529_/B2 _5005_/Z _5138_/A2 _5008_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6958_ hold80/Z _7300_/RN _6958_/CLK _6958_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6889_ _6889_/D _7341_/RN _6926_/CLK _6895_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5909_ hold116/Z _5909_/A2 _5909_/A3 _4305_/C hold117/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_167_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold780 _7018_/Q hold780/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold791 _7212_/Q hold791/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput307 _4159_/ZN spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput329 _7326_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput318 _6853_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ hold363/Z hold882/Z _4241_/S _4240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4171_ _4172_/A1 _6894_/Q _6891_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6812_ _6812_/D _7300_/RN _6812_/CLK _7375_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3955_ input47/Z _4303_/S _4320_/S input72/Z _3957_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6743_ _6743_/D _7243_/RN _6743_/CLK _6743_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6674_ _6674_/A1 _6674_/A2 _6674_/A3 _6676_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_177_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ hold363/Z hold745/Z _5632_/S _7002_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3886_ _7205_/Q _5891_/A3 _5780_/A3 _5891_/A2 _3943_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5556_ hold50/Z _6950_/Q _5556_/S _5556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5487_ _5487_/A1 _5486_/Z _5487_/A3 _5487_/A4 _5523_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4507_ _5061_/A3 _4508_/A2 _4508_/A3 _5380_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7226_ _7226_/D _7315_/RN _7226_/CLK _7226_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4438_ _5320_/C _6894_/Q hold17/I _5054_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7157_ _7157_/D _7359_/RN _7157_/CLK _7157_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4369_ _4051_/Z _6863_/Q _4376_/S _6863_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_10_0__1403_ clkbuf_3_5_0__1403_/Z clkbuf_4_10_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6108_ _7150_/Q _6291_/B1 _6291_/C1 _7124_/Q _6110_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7088_ _7088_/D _7322_/RN _7088_/CLK _7088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6039_ _6043_/A1 _6245_/C _6245_/B _7289_/Q _6294_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_73_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_155_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3740_ hold86/I _3951_/B1 _3916_/B1 _7071_/Q _3742_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ input18/Z _4031_/A2 _4045_/B1 _3670_/Z _3673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _5517_/A1 _5421_/A2 _5410_/B _5421_/C _5412_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6390_ _7245_/Q _6342_/Z _6355_/Z _7157_/Q _6392_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5341_ _5525_/A1 _5039_/Z _5404_/B _5343_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ _5457_/A1 _5324_/A3 _5272_/B _5435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7011_ _7011_/D _7322_/RN _7011_/CLK _7011_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_141_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4223_ hold323/Z hold751/Z _4223_/S _4223_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4154_ _4154_/I _4154_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4085_ _6806_/Q _4092_/A2 _4091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _5482_/A2 _4796_/Z _5336_/A2 _5331_/A3 _4989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6726_ _6726_/D _6681_/Z _7364_/CLK _6726_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3938_ _7165_/Q _4047_/A2 _4020_/B1 _7157_/Q _3938_/C _3950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6657_ _6898_/Q _6657_/A2 _6657_/B1 _6897_/Q _6659_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3869_ _7083_/Q hold18/I _5780_/A3 _5741_/A2 _3917_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5608_ hold323/Z hold621/Z hold69/Z _6987_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6588_ _6847_/Q _6613_/A2 _6588_/B _6613_/C _6590_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_164_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5539_ hold363/Z hold488/Z _5540_/S _5539_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _7209_/D _7286_/RN _7209_/CLK _7209_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_108_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ hold2/Z hold125/Z _5890_/S _5890_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4910_ _4910_/A1 _4910_/A2 _4910_/A3 _4910_/A4 _4912_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_93_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _4691_/C _5323_/C _5216_/B _5216_/C _4842_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _3399_/I _5433_/B2 _5460_/A1 _4454_/Z _4777_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6511_ _5951_/B _7317_/Q _6614_/B _6512_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3723_ _5585_/A2 _3509_/Z _3504_/Z _4405_/A3 _4019_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_173_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _7133_/Q _6315_/Z _6316_/Z _7207_/Q _6443_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3654_ _3654_/A1 _3654_/A2 _3654_/A3 _3654_/A4 _3654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_174_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6373_ _7122_/Q _6308_/Z _6604_/A2 _7164_/Q _6373_/C _6379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3585_ _3533_/Z _3624_/A2 hold83/I hold11/Z _5812_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5324_ _5339_/A1 _5368_/A2 _5324_/A3 _5324_/A4 _5529_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_88_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _5255_/A1 _5484_/A1 _5442_/A2 _5255_/A4 _5257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_88_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4206_ hold404/Z hold99/Z _4211_/S _4206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5186_ _5482_/C _5413_/A2 _5497_/A1 _5105_/C _5306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_96_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4137_ _7361_/Q _4159_/A1 _4137_/B _4137_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4068_ _4148_/A1 _4068_/A2 input67/Z _6964_/Q _4115_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_83_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_225 _4150__15/I _7062_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_203 net579_219/I _7084_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_214 net579_217/I _7073_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_247 net629_291/I _7040_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_236 net629_266/I _7051_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6709_ input75/Z _7012_/Q _4069_/C _6709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_138_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28__1403_ net429_73/I net429_54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_108__1403_ clkbuf_4_1_0__1403_/Z net829_498/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_5_0__1403_ clkbuf_0__1403_/Z clkbuf_3_5_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_94_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold609 _7379_/I hold609/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3370_ _6763_/Q _3370_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _4788_/B _5450_/A2 _5401_/A2 _5040_/A4 _5177_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_112_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _6991_/D _7322_/RN _6991_/CLK _6991_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5942_ hold50/Z hold469/Z _5944_/S _5942_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5873_ hold901/Z hold363/Z _5881_/S _5873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4824_ _3399_/I _5493_/B _5460_/A1 _5180_/B2 _4830_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4755_ _5457_/A1 _5286_/A2 _4755_/A3 _4741_/C _5497_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xnet529_155 net829_493/I _7132_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet529_166 net629_271/I _7121_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3706_ _4405_/A3 _4402_/A4 _3986_/A3 _5872_/A4 _4017_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xnet529_188 net679_327/I _7099_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_177 net679_327/I _7110_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _4688_/A1 _5384_/B _5384_/C _5482_/A2 _5097_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet529_199 net579_217/I _7088_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6425_ _7254_/Q _6319_/Z _6328_/Z _6762_/Q _6610_/B1 _7270_/Q _6428_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_108_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3637_ input19/Z _4031_/A2 _4015_/A2 _7049_/Q _3637_/C _3661_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_115_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3568_ _4402_/A4 _3986_/A3 _3830_/B _5808_/A3 _4019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6356_ _7212_/Q _6354_/Z _6355_/Z _7156_/Q _6370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5307_ _5307_/A1 _5534_/C _5419_/B _5311_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6287_ _6789_/Q _6293_/A2 _6289_/A2 _6785_/Q _6288_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3499_ _7357_/Q _7342_/Q _3500_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5238_ _5517_/A1 _5301_/B _5238_/B1 _5445_/B1 _5238_/C _5375_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_88_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _5395_/A1 _5169_/A2 _5340_/A1 _5525_/A1 _5402_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150__34 net429_82/I _7253_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__12 net429_55/I _7275_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__23 net429_63/I _7264_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold6 hold6/I hold6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_58_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4150__45 net429_70/I _7242_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet779_409 net779_431/I _6827_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _5214_/A4 _5460_/A1 _5295_/B2 _5322_/A2 _5466_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_11_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ _5162_/A2 _5305_/B _4452_/Z _4456_/Z _4483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold417 _5933_/Z _7273_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold406 _7037_/Q hold406/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold428 _6990_/Q hold428/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6210_ _6210_/A1 _6210_/A2 _7293_/Q _6221_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3422_ _3422_/A1 _4060_/S _3421_/B _3426_/A1 _3423_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7190_ _7190_/D _7243_/RN _7190_/CLK _7190_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold439 _7187_/Q hold439/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6141_ _7293_/Q _6141_/A2 _6139_/Z _6294_/A2 _6140_/Z _6289_/B1 _6143_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_74__1403_ clkbuf_4_5_0__1403_/Z net629_266/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xload_slew364 _3556_/B _3906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xload_slew353 hold22/Z _5780_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6072_ _7003_/Q _6295_/B1 _6294_/B1 _7099_/Q _6073_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _5214_/A4 _5475_/A1 _5154_/A2 _5153_/A1 _5172_/A1 _5025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _6974_/D _7359_/RN _6974_/CLK _7393_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ hold38/Z hold246/Z _5926_/S _5925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ hold323/Z hold799/Z _5862_/S _7205_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4807_ _3399_/I _5284_/A2 _5460_/A1 _5319_/A1 _5431_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5787_ hold38/Z hold48/Z hold23/Z _7146_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4738_ _3399_/I _5112_/A1 _5460_/A1 _5319_/A1 _5354_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4669_ _4500_/B _4773_/C _5310_/B _4694_/B _5460_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_150_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6408_ _6408_/A1 _6408_/A2 _6434_/S _6408_/B2 _7314_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7388_ _7388_/I _7388_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6339_ _6339_/A1 _7299_/Q _7298_/Q _7297_/Q _6609_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _6778_/Q _5560_/A1 _5732_/A4 _6677_/A1 _4019_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_35_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5710_ hold59/Z hold239/Z _5713_/S _5710_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6690_ input75/Z _7012_/Q _4069_/C _6690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_86_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5641_ hold2/Z hold287/Z _5641_/S _5641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_8_0__1403_ clkbuf_4_9_0__1403_/I net479_128/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_117_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5572_ _6959_/Q hold99/Z _5575_/S _5572_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4523_ _4792_/B _4523_/A2 _5099_/C _4523_/C _5482_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7311_ _7311_/D _7322_/RN _7322_/CLK _7311_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold214 _5907_/Z _7250_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold203 _7088_/Q hold203/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold225 _7370_/Q hold225/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7242_ _7242_/D _7243_/RN _7242_/CLK _7242_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4454_ _4751_/B _4691_/C _4454_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xhold247 _5925_/Z _7266_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold236 _5719_/Z _7086_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold269 _6948_/Q hold269/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold258 _5548_/Z _6943_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3405_ _4694_/B _4693_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_20
XFILLER_131_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7173_ _7173_/D _7243_/RN _7173_/CLK _7173_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4385_ _4385_/I0 _6877_/Q _4388_/S _6877_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3336_ _6805_/Q _5999_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6124_ _7215_/Q _6290_/A2 _6291_/B1 _7151_/Q _6293_/B1 _7183_/Q _6125_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6055_ _7212_/Q _6290_/A2 _6291_/B1 _7148_/Q _6057_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _4788_/B _4796_/Z _5336_/A3 _5040_/A4 _5337_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _6957_/D _7243_/RN _6957_/CLK _6957_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ hold2/Z hold146/Z _5908_/S _5908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6888_ _6888_/D _7341_/RN _7341_/CLK _6888_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_139_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5839_ hold99/Z hold385/Z _5844_/S _5839_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold781 _6901_/Q hold781/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold770 _5565_/Z _6955_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold792 _5864_/Z _7212_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet829_490 net829_498/I _6737_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput308 _7399_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput319 _6854_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4170_ _4172_/A1 _6896_/Q _6893_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6811_ _6811_/D _7300_/RN _6811_/CLK _7374_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3954_ _5909_/A3 _5566_/A1 _4015_/A2 _7043_/Q _3957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6742_ _6742_/D _7300_/RN _6742_/CLK _6742_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6673_ _6896_/Q _6673_/A2 _6673_/A3 _6674_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3885_ _6939_/Q _5863_/A4 _5863_/A3 _5566_/A1 _3918_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5624_ _5678_/A2 _5891_/A1 _5827_/A1 _5891_/A3 _5632_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_164_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5555_ hold59/Z hold394/Z _5556_/S _6949_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4506_ _4508_/A2 _4508_/A3 _5061_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5486_ _5486_/A1 _5486_/A2 _5486_/A3 _5486_/A4 _5486_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_105_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7225_ _7225_/D _7286_/RN _7225_/CLK _7225_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4437_ hold323/Z hold804/Z _4437_/S _4437_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7156_ _7156_/D _7315_/RN _7156_/CLK _7156_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6107_ _7230_/Q _6294_/A2 _6290_/B1 _7166_/Q _6293_/B1 _7182_/Q _6110_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_86_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4368_ _6890_/Q _7341_/RN _4376_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_140_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7087_ _7087_/D _7322_/RN _7087_/CLK _7087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ hold61/Z hold50/Z _4303_/S _4299_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6038_ _7010_/Q _6292_/A2 _6289_/A2 _7082_/Q _6048_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ _7322_/Q _6961_/Q _6962_/Q _3670_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5340_ _5340_/A1 _5529_/A2 _5340_/B _5340_/C _5343_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5271_ _5355_/A1 _5492_/A4 _5351_/B _5492_/A1 _5271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_142_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7010_ _7010_/D _7286_/RN _7010_/CLK _7010_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_142_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ hold363/Z hold890/Z _4223_/S _4222_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4153_ _7361_/Q input88/Z _4154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4084_ _6805_/Q _6963_/Q _4091_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4986_ _4986_/A1 _4986_/A2 _4989_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6725_ _6725_/D _6680_/Z _4152_/I1 _6725_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3937_ _3937_/A1 _3937_/A2 _3938_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6656_ _6656_/I0 _7336_/Q _6668_/S _7336_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3868_ _3868_/A1 _4402_/A1 _5750_/A4 _3986_/A3 _4033_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_20_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ hold363/Z hold768/Z hold69/Z _6986_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3799_ _7167_/Q _4047_/A2 _4042_/A2 _6763_/Q _7133_/Q _4046_/B1 _3800_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6587_ _6581_/Z _6587_/A2 _6587_/A3 _6586_/Z _6588_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5538_ hold116/Z _5909_/A2 _5777_/A2 _6677_/A3 _5540_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_11_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7208_ _7208_/D _7315_/RN _7208_/CLK _7208_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_133_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _4392_/Z _5508_/A3 _5469_/A3 _5469_/A4 _5470_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7139_ _7139_/D _7359_/RN _7139_/CLK _7139_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4840_ _4454_/Z _5133_/B _5216_/C _5138_/B _4842_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4771_ _3399_/I _5433_/B2 _5460_/A1 _5180_/B2 _4777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_159_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6510_ _6510_/A1 _6510_/A2 _6991_/Q _6613_/A2 _6613_/C _6512_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_14_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3722_ _3504_/Z _3509_/Z _3523_/B _3521_/Z _4411_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _7247_/Q _6342_/Z _6355_/Z _7159_/Q _6443_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3653_ _7187_/Q _4014_/A2 _3963_/A2 _7001_/Q _3919_/B1 _6751_/Q _3654_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6372_ _6372_/A1 _6372_/A2 _6372_/A3 _6372_/A4 _6373_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5323_ _4456_/Z _5460_/A1 _5323_/B _5323_/C _5396_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_3584_ _3548_/B _5872_/A3 _5872_/A2 _3504_/Z _3914_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5254_ _5478_/A1 _4671_/B _5255_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5185_ _5250_/A1 _5353_/A3 _5462_/A4 _5534_/A1 _5190_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ hold764/Z hold323/Z _4211_/S _4205_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _7363_/Q input38/Z _4136_/B _7361_/Q _4137_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_110_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4067_ _7012_/Q _4069_/C _5597_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_25_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_215 net629_296/I _7072_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_204 net579_213/I _7083_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet579_226 net579_240/I _7061_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_248 net629_299/I _7039_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_237 net629_266/I _7050_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _3399_/I _5162_/A2 _4454_/Z _4796_/Z _5234_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6708_ _7359_/RN _7012_/Q _4069_/C _6708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6639_ _6639_/A1 _6639_/A2 _6640_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _6990_/D _7322_/RN _6990_/CLK _6990_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5941_ hold59/Z hold497/Z _5944_/S _5941_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_34__1403_ clkbuf_4_10_0__1403_/Z _4150__48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5872_ _5578_/B _5872_/A2 _5872_/A3 _5872_/A4 _5881_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_114__1403_ net779_410/I net779_451/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4823_ _4823_/A1 _4823_/A2 _4823_/A3 _4830_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_178_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_97__1403_ clkbuf_4_4_0__1403_/Z _4150__44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_187_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4754_ _4839_/A3 _4839_/A2 _4839_/A4 _5138_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xnet529_167 net579_243/I _7120_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_178 net779_419/I _7109_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_156 net429_95/I _7131_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3705_ _3704_/Z _6936_/Q _3961_/S _6936_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet529_189 net679_327/I _7098_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _5384_/B _5384_/C _5228_/B _5493_/A1 _5260_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _7190_/Q _6318_/Z _6608_/B1 _7108_/Q _6341_/Z _6996_/Q _6429_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3636_ _3636_/I _3637_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6355_ _7296_/Q _6543_/A2 _6594_/A3 _6355_/A4 _6355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3567_ _3504_/Z _3509_/Z _3521_/Z hold573/Z _5900_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5306_ _5306_/A1 _5306_/A2 _5306_/B _5306_/C _5419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6286_ _6777_/Q _6294_/B1 _6293_/B1 _7359_/Q _6288_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5237_ _5237_/A1 _5237_/A2 _5238_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3498_ _6725_/Q _3498_/A2 _3498_/B _7344_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _4796_/Z _5336_/A2 _5336_/A3 _5176_/A2 _5170_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _5382_/B2 _5182_/C _5099_/B _5099_/C _5100_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4119_ _6829_/Q input89/Z _4119_/S _4119_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4150__13 _4150__22/I _7274_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__24 net429_59/I _7263_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150__35 _4150__40/I _7252_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__46 _4150__46/I _7241_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold7 hold7/I hold7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_90_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ _4773_/C _5305_/C _4698_/C _4995_/A4 _4485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold407 _7093_/Q hold407/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold418 _6942_/Q hold418/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_99_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ _7371_/Q _3419_/Z _3421_/B _3422_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold429 _7065_/Q hold429/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6140_ hold93/I _7143_/Q _7293_/Q _6140_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3352_ _7322_/Q _6615_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6071_ _7011_/Q _6292_/A2 _6289_/A2 _7083_/Q _6073_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xload_slew343 _4423_/A2 _5741_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5022_ _4794_/Z _5171_/A2 _5401_/A2 _5401_/A3 _5154_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _6973_/D _7359_/RN _6973_/CLK _7392_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ hold50/Z hold278/Z _5926_/S _5924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _4178_/Z hold855/Z _5862_/S _7204_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4806_ _5283_/A2 _5268_/B _4806_/A3 _4730_/B _5284_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5786_ hold50/Z hold76/Z hold23/Z _7145_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4737_ _5460_/A1 _5322_/A2 _4751_/B _4762_/A4 _5405_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4668_ _4693_/B _4787_/B _4702_/B _5305_/B _5213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_108_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6407_ _5951_/B _7313_/Q _6614_/B _6408_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3619_ _3906_/A1 _5872_/A2 _3509_/Z _5808_/A3 _4012_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4599_ _5421_/C _5461_/A3 _5184_/A2 _5413_/A2 _5237_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7387_ _7387_/I _7387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6338_ _6593_/A3 _6387_/A1 _6343_/A4 _6007_/B _6338_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_103_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _6756_/Q _6295_/B1 _6291_/C1 _6752_/Q _6289_/B1 _6770_/Q _6273_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_28_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80__1403_ clkbuf_4_5_0__1403_/Z net729_396/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_100 net629_286/I _7187_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3970_ input93/Z _5891_/A4 _5759_/A3 _5566_/A1 _4007_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_44_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5640_ hold38/Z hold272/Z _5641_/S _5640_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5571_ _6958_/Q hold79/Z _5571_/S hold80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4522_ _5441_/A4 _4607_/A3 _4607_/A2 _5382_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7310_ _7310_/D _7322_/RN _7322_/CLK _7310_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4453_ _4702_/B _4694_/B _4787_/B _5305_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7241_ _7241_/D _7286_/RN _7241_/CLK _7241_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold215 _7258_/Q hold215/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold204 _5721_/Z _7088_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold226 hold226/I hold226/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3404_ _5305_/B _4773_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_20
Xhold248 _6766_/Q hold248/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet429_90 net429_90/I _7197_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold237 _7070_/Q hold237/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold259 _7013_/Q hold259/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7172_ _7172_/D input75/Z _7172_/CLK _7172_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4384_ _6624_/I0 _6876_/Q _4388_/S _6876_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3335_ _7012_/Q _4148_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6123_ _7207_/Q _6289_/A2 _6294_/B1 _7223_/Q _6125_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6054_ _7130_/Q _6295_/B1 _6290_/B1 _7164_/Q _6057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _4788_/B _4796_/Z _5336_/A3 _5040_/A4 _5005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6956_ _6956_/D _7359_/RN _6956_/CLK _7373_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ hold38/Z hold213/Z _5908_/S _5907_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6887_ _6887_/D _7315_/RN _6887_/CLK _6887_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ hold323/Z hold766/Z _5844_/S _5838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ hold363/Z hold821/Z _5776_/S _5769_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold760 _6951_/Q hold760/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold771 _6946_/Q hold771/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold782 _4409_/Z _6901_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold793 _7043_/Q hold793/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet829_480 net829_482/I _6747_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet829_491 net829_499/I _6736_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_183_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput309 _7400_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6810_ _6810_/D _7300_/RN _6810_/CLK _6810_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3953_ _7181_/Q _4014_/A2 _3953_/B1 _6902_/Q _4033_/A2 _7229_/Q _3957_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6741_ _6741_/D _7300_/RN _6741_/CLK _6741_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_16_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6672_ _6898_/Q _6672_/A2 _6673_/A2 _6674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3884_ _3884_/A1 _3830_/C _3521_/Z _5872_/A4 _4031_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_137_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5623_ hold2/Z hold448/Z _5623_/S _5623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5554_ hold79/Z hold269/Z _5556_/S _6948_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5485_ _5534_/A1 _5490_/C _5061_/Z _5521_/B2 _5486_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4505_ _4508_/A2 _4508_/A3 _4505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7224_ _7224_/D _7286_/RN _7224_/CLK _7224_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4436_ hold363/Z hold846/Z _4437_/S _4436_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7155_ hold34/Z _7300_/RN _7155_/CLK _7155_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4367_ hold323/Z hold699/Z _4367_/S _4367_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6106_ _6106_/A1 _6106_/A2 _6106_/A3 _6106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_86_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7086_ _7086_/D _7322_/RN _7086_/CLK _7086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_58_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ hold577/Z _4297_/Z _4304_/S _4298_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6037_ _6245_/C _6245_/B _7290_/Q _7289_/Q _6289_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_2217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6939_ _6939_/D _7359_/RN _6939_/CLK _6939_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_183_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold590 _6822_/Q hold590/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ _5268_/B _5270_/A2 _5286_/A4 _5270_/A4 _5492_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_142_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4221_ _5882_/A2 _6677_/A2 _6677_/A3 _4223_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_96_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ input83/Z _4152_/I1 _7361_/Q _4152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4083_ _4092_/A2 _6613_/C _4083_/B _6806_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4985_ _4796_/Z _5336_/A2 _5331_/A3 _5024_/A4 _4986_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_63_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6724_ _6724_/D _4173_/Z _3753_/A1 _6724_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3936_ _3924_/Z _3936_/A2 _3936_/A3 _3935_/Z _3958_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6655_ _6655_/A1 _6655_/A2 _6656_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3867_ _3868_/A1 hold68/I _4402_/A1 _4402_/A3 _4047_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_165_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6586_ _6613_/A2 _6586_/A2 _6586_/A3 _6586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5606_ _5750_/A3 _5750_/A2 _5891_/A1 hold68/Z hold69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3798_ _6747_/Q _3919_/B1 _3914_/B1 _6731_/Q _3798_/C _3820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_180_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _5537_/A1 _5537_/A2 _5537_/A3 _6927_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_160_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7207_ _7207_/D _7315_/RN _7207_/CLK _7207_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _5468_/A1 _5468_/A2 _5509_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5399_ _5399_/A1 _5452_/A2 _5476_/A2 _5400_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4419_ hold323/Z hold512/Z _4419_/S _4419_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7138_ _7138_/D _7359_/RN _7138_/CLK _7138_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7069_ _7069_/D _7322_/RN _7069_/CLK _7069_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _4770_/A1 _4770_/A2 _4770_/A3 _4770_/A4 _4777_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_1891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3721_ _6999_/Q _5678_/A2 _5827_/A1 _5759_/A3 _3744_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_158_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _7183_/Q _6320_/Z _6341_/Z _6997_/Q _6443_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3652_ input51/Z _4285_/S _4019_/A2 _7251_/Q _3654_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6371_ _7050_/Q _6324_/Z _6325_/Z _7082_/Q _6371_/C _6372_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3583_ _3533_/Z _5909_/A2 hold68/Z _5872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_61_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5322_ _5323_/C _5322_/A2 _5460_/A1 _4456_/Z _5333_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_115_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_57__1403_ net579_205/I net629_297/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5253_ _5253_/A1 _5253_/A2 _5253_/A3 _5442_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5184_ _5294_/C _5184_/A2 _5184_/A3 _5184_/B _5191_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_69_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4204_ hold844/Z hold363/Z _4211_/S _4204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _4135_/A1 _4135_/A2 _7363_/Q _4136_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4066_ _4148_/A1 hold535/Z input67/Z _4305_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xnet579_205 net579_205/I _7082_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_216 net579_217/I _7071_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet579_238 net429_76/I _7049_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_227 net579_240/I _7060_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_249 _4150__9/I _7038_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _5214_/A4 _5460_/A1 _4698_/C _5326_/C _5250_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_51_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4899_ _4691_/C _5490_/B _5309_/B _5353_/A4 _5431_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6707_ input75/Z _7012_/Q _4069_/C _6707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3919_ _6995_/Q _3963_/A2 _3919_/B1 _6745_/Q _3919_/C _3959_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6638_ _6896_/Q _6638_/A2 _6638_/B1 _6666_/B2 _6639_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _6770_/Q _6323_/Z _6334_/Z _6882_/Q _6352_/Z _6774_/Q _6572_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_180_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ hold79/Z hold548/Z _5944_/S _5940_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5871_ hold2/Z hold42/Z _5871_/S hold43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4822_ _5286_/A2 _5268_/B _5134_/A3 _5473_/A2 _4823_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_33_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4753_ _5216_/B _4829_/A4 _4753_/A3 _4835_/A1 _4759_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet529_168 net579_243/I _7119_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_179 net629_301/I _7108_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet529_157 net429_71/I _7130_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3704_ _6935_/Q _6627_/I0 _3960_/S _3704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4684_ _5214_/A4 _5295_/B2 _4691_/C _5162_/A2 _5359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _6423_/A1 _6423_/A2 _6423_/A3 _6423_/A4 _6430_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_134_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ _7267_/Q _4017_/A2 _4027_/B1 _7259_/Q input42/Z _4320_/S _3636_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_143_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6354_ _7297_/Q _7296_/Q _6376_/A2 _6594_/A3 _6354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3566_ _3523_/B _3554_/B _5808_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_170_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5305_ _5306_/A1 _5306_/A2 _5305_/B _5305_/C _5534_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6285_ _6773_/Q _6294_/A2 _6290_/B1 _6783_/Q _6291_/B1 _6775_/Q _6288_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3497_ _3496_/Z _3497_/A2 _7344_/Q _3498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5236_ _5395_/A1 _5445_/A2 _5441_/A3 _5236_/A4 _5237_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5167_ _5395_/A1 _5005_/Z _5169_/A2 _5525_/A1 _5167_/C _5170_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ _5099_/C _5368_/A2 _5098_/A3 _5098_/B1 _5259_/B _5262_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4118_ _6830_/Q input91/Z _4119_/S _4118_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _4044_/Z _4049_/A2 _4048_/Z _4049_/A4 _4050_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40__1403_ clkbuf_4_14_0__1403_/Z _4150__22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4150__25 _4150__25/I _7262_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__14 _4150__15/I _7273_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150__36 net429_76/I _7251_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__47 _4150__48/I _7240_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold8 hold8/I hold8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold408 _7202_/Q hold408/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _7371_/Q _7370_/Q hold81/I _3426_/B _4060_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xhold419 _5547_/Z _6942_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3351_ _3351_/I _4159_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xload_slew355 hold7/Z _5732_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6070_ _7035_/Q _6295_/A2 _6291_/C1 _6995_/Q _6292_/B1 _7067_/Q _6073_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew344 _4408_/A1 _5678_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5021_ _5326_/C _5030_/A2 _4789_/B _5338_/A2 _5389_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xload_slew366 _4305_/C _6677_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ _6972_/D _7359_/RN _6972_/CLK _7391_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5923_ hold59/Z hold457/Z _5926_/S _5923_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5854_ _4305_/C _5882_/A2 _5927_/A3 hold18/Z _5862_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _3399_/I _5280_/B _5460_/A1 _4454_/Z _4809_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5785_ hold59/Z hold176/Z hold23/Z _7144_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4736_ _5214_/A4 _5295_/B2 _3402_/I _5162_/A2 _5525_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4667_ _5095_/A2 _5384_/B _5384_/C _5228_/A2 _4671_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_134_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _6406_/A1 _6406_/A2 _6987_/Q _6613_/A2 _6613_/C _6408_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_7386_ _7386_/I _7386_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3618_ _3906_/A1 _3548_/B _5872_/A3 _5872_/A2 _4020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6337_ _7295_/Q _6387_/A1 _6540_/A4 _6337_/A4 _6337_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_4598_ _4598_/A1 _4598_/A2 _5071_/C _4601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3549_ _3509_/Z _3556_/B _5872_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_135_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6268_ _6268_/A1 _6268_/A2 _6268_/B1 _6268_/B2 _6268_/C _6274_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5219_ _5215_/Z _5219_/A2 _5320_/A1 _5320_/A2 _5320_/C _5224_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6199_ _6199_/I0 _7308_/Q _6434_/S _7308_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet429_101 net429_89/I _7186_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ hold263/Z hold59/Z _5575_/S _6957_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4521_ _4792_/B _4523_/A2 _4523_/C _4716_/B _5236_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4452_ _4702_/B _4694_/B _4787_/B _4452_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7240_ _7240_/D _7315_/RN _7240_/CLK _7240_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold216 _7071_/Q hold216/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold205 _7200_/Q hold205/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet429_80 net429_80/I _7207_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3403_ _4702_/B _4500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_12
XFILLER_171_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold249 _4231_/Z _6766_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet429_91 net429_91/I _7196_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold238 _7397_/I hold238/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold227 _3545_/B hold227/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ hold28/Z _7243_/RN _7171_/CLK hold27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4383_ _3859_/Z _6875_/Q _4388_/S _6875_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3334_ _6892_/Q _4109_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6122_ _6763_/Q _6299_/C _6265_/B1 _7167_/Q _6265_/C _6125_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6053_ _7228_/Q _6294_/A2 _6294_/B1 _7220_/Q _6057_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _5238_/B1 _5342_/A2 _4796_/Z _5336_/A3 _5008_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _6955_/D _7359_/RN _6955_/CLK _6955_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5906_ hold50/Z hold274/Z _5908_/S _5906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6886_ _6886_/D _7315_/RN _6886_/CLK _6886_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ hold363/Z hold874/Z _5844_/S _7188_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5768_ _5891_/A1 _6677_/A1 _5836_/A3 _5891_/A3 _5776_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4719_ _5291_/B _4835_/A1 _4483_/B _4716_/B _5497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_163_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5699_ hold99/Z hold556/Z hold84/Z _7068_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7369_ _7369_/D _6721_/Z _3753_/A1 hold81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold750 _4241_/Z _6773_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold761 _5558_/Z _6951_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold772 _6861_/Q hold772/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold794 _5671_/Z _7043_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold783 _6940_/Q hold783/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet829_481 net829_483/I _6746_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_470 net429_98/I _6757_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet829_492 net429_95/I _6735_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _6740_/D _7243_/RN _6740_/CLK _6740_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3952_ _3952_/A1 _3952_/A2 _3952_/A3 _3952_/A4 _3958_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_189_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6671_ _6897_/Q _6673_/A2 _6671_/A3 _6674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3883_ _6771_/Q _5560_/A1 _5780_/A3 _6677_/A1 _3925_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5622_ hold38/Z hold107/Z _5623_/S _5622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5553_ hold99/Z hold280/Z _5556_/S _6947_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4504_ _5162_/A2 _4452_/Z _4456_/Z _4773_/C _4508_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_129_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5484_ _5484_/A1 _5484_/A2 _5484_/A3 _5484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_172_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7223_ _7223_/D _7315_/RN _7223_/CLK _7223_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4435_ _4435_/A1 _5750_/A4 _5750_/A3 hold310/Z _4437_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_99_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7154_ _7154_/D _7300_/RN _7154_/CLK hold52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4366_ hold363/Z hold772/Z _4367_/S _4366_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _7174_/Q _6291_/A2 _6295_/B1 _7132_/Q _6292_/B1 _7190_/Q _6106_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7085_ _7085_/D _7322_/RN _7085_/CLK _7085_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ hold65/Z hold59/Z _4303_/S _4297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6036_ _6043_/A1 _6231_/A1 _7292_/Q _7291_/Q _6292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_74_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _6938_/D _7359_/RN _6938_/CLK _6938_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _6869_/D _7325_/CLK _6869_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold580 _4300_/Z _6814_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold591 _4317_/Z _6822_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ hold323/Z hold697/Z _4220_/S _4220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4151_ input84/Z input67/Z _7362_/Q _4151_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4082_ _5952_/B _4062_/Z _5964_/A2 _7286_/Q _4092_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4984_ _5405_/A1 _5473_/A2 _5024_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17__1403_ clkbuf_4_10_0__1403_/Z _4150__51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3935_ _3935_/A1 _3935_/A2 _3931_/Z _3934_/Z _3935_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6723_ _7359_/RN _7012_/Q _4069_/C _6723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_51_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6654_ _6896_/Q _6654_/A2 _6654_/B1 _6666_/B2 _6655_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5605_ hold2/Z hold35/Z _5605_/S hold36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3866_ _6908_/Q _5560_/A1 _5780_/A3 _5741_/A2 _3917_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6585_ _6786_/Q _6310_/Z _6321_/Z _6871_/Q _6610_/B1 _6917_/Q _6586_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3797_ _3797_/I _3798_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5536_ _5536_/A1 _5536_/A2 _5536_/B _5536_/C _5537_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5467_ _5509_/A1 _5467_/A2 _5467_/A3 _5506_/A2 _5470_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7206_ _7206_/D _7315_/RN _7206_/CLK _7206_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_172_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4418_ hold363/Z hold510/Z _4419_/S _4418_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5398_ _5398_/A1 _5398_/A2 _5476_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7137_ _7137_/D _7286_/RN _7137_/CLK _7137_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ hold323/Z hold653/Z _4349_/S _4349_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ _7068_/D _7322_/RN _7068_/CLK _7068_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _6019_/A1 _6019_/A2 _7302_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _3720_/A1 _3720_/A2 _3720_/A3 _3720_/A4 _3720_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_186_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3651_ input70/Z _4303_/S _4027_/A2 _7283_/Q _3654_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6370_ _6370_/A1 _6370_/A2 _6370_/A3 _6371_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3582_ _3624_/A2 hold83/I hold11/Z _3868_/A1 _5827_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_161_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5321_ _5468_/A1 _5469_/A3 _5430_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _5099_/B _5252_/A2 _5384_/A2 _5441_/A4 _5253_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5183_ _5510_/A2 _5183_/A2 _5183_/B _5184_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_4__1403_ clkbuf_4_2_0__1403_/Z _4150__3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4203_ _5578_/B _3830_/C _4405_/A3 _5808_/A4 _4211_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_84_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _6937_/Q _7012_/Q _4069_/C _4135_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4065_ input67/Z _6964_/Q _4069_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_83_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet579_206 net629_272/I _7081_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_239 net579_240/I _7048_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_217 net579_217/I _7070_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_228 net629_298/I _7059_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4967_ _5087_/B2 _4967_/A2 _5397_/A2 _5395_/A1 _4972_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6706_ _7286_/RN _7012_/Q _4069_/C _6706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4898_ _4898_/A1 _5200_/C _4898_/A3 _4898_/A4 _4901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3918_ _3918_/A1 _3918_/A2 _3919_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6637_ _6898_/Q _6637_/A2 _6637_/B1 _6897_/Q _6639_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3849_ _7124_/Q _3951_/B1 _4015_/A2 _7044_/Q _3850_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6568_ _6919_/Q _6594_/A2 _6594_/A3 _6594_/A4 _6579_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ _5519_/A1 _5536_/A1 _5536_/B _5520_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ hold86/I _6308_/Z _6336_/Z _7103_/Q _6503_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5870_ hold38/Z hold131/Z _5871_/S _5870_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ _5286_/A2 _5268_/B _5405_/A1 _5134_/A3 _4823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_2390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _5473_/A1 _5416_/B _4753_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xnet529_169 _4150__25/I _7118_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _5460_/A1 _5322_/A2 _4751_/B _3399_/I _5493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3703_ _3677_/Z _3703_/A2 _3703_/A3 _6627_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xnet529_158 net629_266/I _7129_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3634_ _4402_/A4 _3986_/A3 _5872_/A3 _3830_/B _4027_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6422_ _7222_/Q _6317_/Z _6354_/Z _7214_/Q _6387_/Z _7060_/Q _6423_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_108_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6353_ _7026_/Q _6566_/A2 _6376_/A2 _6540_/A4 _6377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3565_ _6881_/Q hold31/Z _3565_/B _3565_/C hold32/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_142_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _5304_/A1 _5466_/A1 _5359_/A2 _5268_/B _5312_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6284_ _6284_/A1 _6284_/A2 _6284_/A3 _6284_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3496_ _7345_/Q _6725_/Q _3496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5235_ _5235_/A1 _5235_/A2 _5235_/A3 _5242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5166_ _5337_/A1 _5333_/A1 _5166_/B _5167_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ _4117_/A1 _4117_/A2 _6894_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5097_ _5259_/B _5098_/B1 _5097_/B _5481_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ _4048_/A1 _4048_/A2 _4048_/A3 _4048_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_140_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5999_ _5999_/I0 _6339_/A1 _6807_/Q _5999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4150__15 _4150__15/I _7272_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput290 _6747_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4150__37 _4150__46/I _7250_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__48 _4150__48/I _7239_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__26 _4150__51/I _7261_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 hold9/I hold9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_74_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold409 _5852_/Z _7202_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3350_ _3350_/I _4101_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _5020_/A1 _5020_/A2 _5020_/A3 _5025_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xload_slew356 hold7/Z _5863_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew367 _4305_/C _5891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6971_ _6971_/D _7359_/RN _6971_/CLK _7390_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ hold79/Z hold340/Z _5926_/S _5922_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5853_ hold2/Z hold475/Z _5853_/S _7203_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4804_ _5287_/A1 _5280_/B _4804_/B _4809_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_167_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5784_ hold79/Z hold308/Z hold23/Z _7143_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _5322_/A2 _4751_/B _4762_/A4 _5396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _5172_/A1 _4689_/A2 _4641_/C _5304_/A1 _4673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_119_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4597_ _5417_/C _5294_/C _5417_/A2 _5199_/A3 _5071_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6405_ _6613_/A2 _6405_/A2 _6405_/A3 _6404_/Z _6406_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7385_ _7385_/I _7385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold910 _7156_/Q hold910/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3617_ _3906_/A1 _3548_/B _5872_/A3 _5585_/A2 _4038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6336_ _7297_/Q _7296_/Q _6543_/A2 _6540_/A4 _6336_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3548_ _6881_/Q hold6/Z _3548_/B _3548_/C hold7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_131_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6267_ _6780_/Q _6290_/A2 _6291_/B1 _6774_/Q _6293_/B1 _7358_/Q _6268_/C VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _6792_/Q _3482_/B _7354_/Q _3480_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5218_ _5413_/A2 _5493_/A1 _5218_/B _5228_/B _5219_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6198_ _6806_/Q _6198_/A2 _6198_/A3 _6198_/B _6199_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_28_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5149_ _5395_/A2 _4975_/Z _5149_/A3 _5176_/A2 _5525_/A1 _5157_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_97_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_13_0__1403_ clkbuf_3_6_0__1403_/Z net579_205/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_84_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4520_ _5214_/A4 _5460_/A1 _4751_/B _4691_/C _5439_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _4694_/B _4787_/B _5294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_117_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold217 _7087_/Q hold217/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold206 _5850_/Z _7200_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet429_81 net429_81/I _7206_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3402_ _3402_/I _5322_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_20
XFILLER_144_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7170_ _7170_/D _7315_/RN _7170_/CLK _7170_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_70 net429_70/I _7217_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold239 _7078_/Q hold239/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold228 hold228/I hold228/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6121_ _6121_/A1 _6268_/A1 _6121_/A3 _6265_/C _6142_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet429_92 net429_97/I _7195_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4382_ _6622_/I0 _6874_/Q _4388_/S _6874_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3333_ _6793_/Q _4095_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6052_ _6052_/A1 _6052_/A2 _6052_/A3 _6058_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _5482_/A2 _5342_/A2 _4796_/Z _5336_/A3 _5008_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6954_ _6954_/D _6954_/CLK _6954_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ hold59/Z hold501/Z _5908_/S _5905_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _6885_/D input75/Z _6885_/CLK _6885_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5836_ _6677_/A3 _5891_/A2 _5836_/A3 _5891_/A3 _5844_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_50_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5767_ hold2/Z hold15/Z _5767_/S hold16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4718_ _4829_/A4 _4718_/A2 _4718_/A3 _5291_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_108_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5698_ hold323/Z hold727/Z hold84/Z _7067_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4649_ _4649_/A1 _4649_/A2 _4649_/A3 _4656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold762 _6966_/Q hold762/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7368_ _7368_/D _6720_/Z _3753_/A1 _7368_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold751 _6759_/Q hold751/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold740 _5559_/Z _6952_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold773 _4366_/Z _6861_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7299_ _7299_/D _7322_/RN _7319_/CLK _7299_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_6319_ _6543_/A2 _6343_/A4 _7299_/Q _6594_/A4 _6319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_103_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold795 _6737_/Q hold795/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold784 _6954_/Q hold784/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet829_460 _4150__46/I _6767_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet829_471 net429_98/I _6756_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_493 net829_493/I _6734_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_482 net829_482/I _6745_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ input12/Z _4031_/A2 _3951_/B1 _7123_/Q _3951_/C _3952_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_50_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _6890_/Q _6670_/A2 _4393_/Z _7340_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_32_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3882_ _6952_/Q _5900_/A3 _5557_/A2 hold68/I _3937_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_177_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5621_ hold50/Z hold680/Z _5623_/S _6999_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5552_ hold323/Z hold771/Z _5556_/S _6946_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4503_ _4502_/C _5305_/B _4508_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_8_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5483_ _5483_/A1 _5483_/A2 _5484_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7222_ _7222_/D _7286_/RN _7222_/CLK _7222_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4434_ hold323/Z hold632/Z _4434_/S _4434_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7153_ _7153_/D _7243_/RN _7153_/CLK _7153_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4365_ _4408_/A1 _5777_/A2 _6677_/A3 _4367_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_140_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6104_ _7158_/Q _6295_/A2 _6294_/B1 _7222_/Q _6106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7084_ _7084_/D _7322_/RN _7084_/CLK _7084_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6035_ _6035_/A1 _6035_/A2 _6035_/A3 _6058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ hold588/Z _4295_/Z _4304_/S _4296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _6937_/D _6695_/Z _4152_/I1 _6937_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_6868_ _6868_/D _6880_/CLK _6868_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5819_ hold363/Z hold862/Z _5826_/S _7172_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _6799_/D _7286_/RN _6799_/CLK _7383_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold581 _6823_/Q hold581/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold570 hold570/I _7167_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold592 _7374_/I hold592/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f__1085_ clkbuf_0__1085_/Z _4385_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4081_ _5959_/B _7288_/Q _5964_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_110_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _5014_/A1 _5330_/B _4983_/B _4983_/C _4986_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3934_ _3934_/A1 _3934_/A2 _3934_/A3 _3934_/A4 _3934_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6722_ _7359_/RN _7012_/Q _4069_/C _6722_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_16_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6653_ _6898_/Q _6653_/A2 _6653_/B1 _6897_/Q _6655_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3865_ _4405_/A3 _4402_/A4 _4402_/A3 _3830_/B _3963_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_31_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5604_ hold38/Z hold91/Z _5605_/S hold92/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6584_ _6913_/Q _6610_/A2 _6328_/Z _7138_/Q _6347_/C _6768_/Q _6586_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3796_ _7231_/Q _4033_/A2 _4012_/A2 _7199_/Q _7183_/Q _4014_/A2 _3797_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5535_ _5535_/A1 _5535_/A2 _5412_/Z _5463_/Z _5536_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5466_ _5466_/A1 _5466_/A2 _5217_/B _5466_/B _5467_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7205_ _7205_/D _7315_/RN _7205_/CLK _7205_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_105_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4417_ _6677_/A3 _4423_/A2 _5780_/A3 _5560_/A1 _4419_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5397_ _5440_/A2 _5397_/A2 _5397_/B1 _4796_/Z _5397_/C _5398_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7136_ hold54/Z _7300_/RN _7136_/CLK hold53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4348_ hold363/Z hold704/Z _4349_/S _4348_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4279_ hold381/Z hold59/Z _4285_/S _4279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7067_ _7067_/D _7322_/RN _7067_/CLK _7067_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6018_ _6014_/Z _7302_/Q _6019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_1_0__1403_ clkbuf_4_1_0__1403_/I clkbuf_4_1_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_23__1403_ clkbuf_4_9_0__1403_/Z net829_473/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_103__1403_ clkbuf_4_1_0__1403_/Z net729_369/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_86__1403_ clkbuf_4_4_0__1403_/Z net429_93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3650_ hold15/I _3951_/B1 _3914_/B1 _6735_/Q _4012_/A2 _7203_/Q _3654_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_155_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3581_ _3906_/A1 _3830_/C _3509_/Z _5581_/A3 _4043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_127_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5320_ _5320_/A1 _5320_/A2 _5320_/B _5320_/C _5468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_114_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5251_ _5251_/A1 _5251_/A2 _5484_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4202_ hold2/Z hold360/Z _4202_/S _4202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5182_ _5182_/A1 _5296_/A3 _5417_/B _5416_/B _5182_/C _5183_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_95_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4133_ _5597_/A3 _6810_/Q _4135_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4064_ _7360_/Q _7342_/Q _4068_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xnet579_207 net579_207/I _7080_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_229 _4150__9/I _7058_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_218 net579_221/I _7069_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4966_ _5405_/A1 _5338_/A2 _5220_/A3 _5327_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6705_ _7286_/RN _7012_/Q _4069_/C _6705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_177_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4897_ _5417_/C _5199_/A3 _5306_/C _5416_/B _4898_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_20_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3917_ _3917_/A1 _3917_/A2 _3917_/A3 _3917_/A4 _3917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6636_ _6636_/A1 _6636_/A2 _4392_/Z _6668_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_177_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _7182_/Q _4014_/A2 _4012_/A2 _7198_/Q _3850_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3779_ _3779_/A1 _3779_/A2 _3784_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6567_ _6928_/Q _6593_/A2 _6593_/A3 _6594_/A4 _6575_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5518_ _5518_/A1 _5518_/A2 _5518_/A3 _5536_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _6494_/Z _6498_/A2 _6498_/A3 _6498_/A4 _6510_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _5449_/A1 _5262_/B _5472_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7119_ _7119_/D _7286_/RN _7119_/CLK _7119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/Z _3353__1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4820_ _5286_/A2 _5268_/B _5134_/A3 _5493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_2380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4751_ _5267_/A1 _5102_/B2 _4751_/B _5475_/B _4760_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_159_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet529_159 net579_240/I _7128_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4682_ _5460_/A1 _4751_/B _3399_/I _5353_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3702_ _3702_/A1 _3702_/A2 _3702_/A3 _3702_/A4 _3703_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_147_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6421_ _7036_/Q _6312_/Z _6604_/A2 _7166_/Q _6423_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3633_ _7227_/Q _3914_/A2 _4028_/A2 hold42/I _3661_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_146_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6352_ _7296_/Q _6376_/A2 _6594_/A3 _6355_/A4 _6352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3564_ _3556_/B _3548_/B _3830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5303_ _5482_/C _5320_/A1 _5493_/A1 _5105_/C _5306_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6283_ _6787_/Q _6291_/A2 _6295_/A2 _6779_/Q _6290_/A2 _6781_/Q _6284_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3495_ input58/Z _6727_/Q _6726_/Q _6792_/Q _3498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_170_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _5304_/A1 _5234_/A2 _5417_/B _5234_/B1 _4515_/Z _5235_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5165_ _5395_/A1 _5529_/B2 _5005_/Z _5525_/A1 _5165_/C _5166_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4116_ _6888_/Q _4116_/A2 _4106_/Z _4117_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5096_ _5096_/A1 _5478_/A1 _5096_/A3 _5100_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4047_ _7164_/Q _4047_/A2 _4047_/B1 _7140_/Q _4047_/C1 _6915_/Q _4048_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_25_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5998_ _7295_/Q _7294_/Q _7296_/Q _6339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4949_ _4949_/A1 _4502_/B _4963_/A2 _4963_/A3 _5473_/B _4967_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_166_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6619_ _6619_/I _7323_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput280 _6730_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150__16 net429_59/I _7271_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput291 _6748_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4150__49 net429_82/I _7238_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__27 _4150__51/I _7260_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__38 _4150__5/I _7249_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6970_ _6970_/D _7359_/RN _6970_/CLK _7389_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_65_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ hold99/Z hold553/Z _5926_/S _5921_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ hold38/Z hold408/Z _5853_/S _5852_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4803_ _4691_/C _5287_/A1 _5280_/B _5282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5783_ hold99/Z hold301/Z hold23/Z _7142_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4734_ _5214_/A4 _5295_/B2 _3402_/I _5138_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_159_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _4656_/Z _5253_/A3 _5091_/C _4673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7384_ _7384_/I _7384_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold900 _6994_/Q hold900/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4596_ _5417_/C _5294_/C _4694_/B _4787_/B _5301_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6404_ _6404_/A1 _6404_/A2 _6404_/A3 _6404_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3616_ _5557_/A2 hold68/Z _5585_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_150_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6335_ _7295_/Q _6594_/A4 _6540_/A4 _6337_/A4 _6335_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3547_ _5808_/A4 _4405_/A3 _4402_/A4 _3986_/A3 _4303_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_170_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _6776_/Q _6266_/A2 _6299_/B _6784_/Q _6268_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3478_ _3482_/B _3478_/A2 _3478_/B _7355_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5217_ _5234_/A2 _5359_/A2 _5217_/B _5344_/C _5320_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6197_ _6806_/Q _7307_/Q _6198_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5148_ _5326_/C _5325_/A2 _4953_/Z _5333_/A1 _5149_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_57_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5079_ _5079_/A1 _5522_/A1 _5378_/A1 _5378_/A2 _5079_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_57_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ _4442_/Z _4444_/Z _4447_/Z _4959_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_156_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold207 _7094_/Q hold207/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet429_82 net429_82/I _7205_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3401_ _4751_/B _5295_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_16
Xnet429_60 _4150__5/I _7227_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold218 _5720_/Z _7087_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold229 hold229/I _5556_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4381_ _4051_/Z _6873_/Q _4388_/S _6873_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet429_71 net429_71/I _7216_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6120_ _5951_/B _6614_/B _7306_/Q _6147_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xnet429_93 net429_93/I _7194_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3332_ _6792_/Q _3472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_112_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _7172_/Q _6291_/A2 _6295_/A2 _7156_/Q _6265_/C _6052_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _5002_/A1 _5002_/A2 _5008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6953_ _6953_/D _7243_/RN _6953_/CLK _6953_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_35_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ hold79/Z hold387/Z _5908_/S _5904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6884_ _6884_/D input75/Z _6884_/CLK _6884_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5835_ hold2/Z hold439/Z _5835_/S _5835_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5766_ hold38/Z hold371/Z _5767_/S _5766_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4717_ _4835_/A1 _4929_/A2 _4929_/A3 _4483_/B _5216_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_163_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5697_ hold363/Z hold889/Z hold84/Z _7066_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4648_ _4906_/A1 _3399_/I _5475_/A2 _5162_/A2 _5312_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_108_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold730 _7011_/Q hold730/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _5417_/C _5475_/A2 _3399_/I _5162_/A2 _5250_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_122_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7367_ _7367_/D _6719_/Z _3753_/A1 _7367_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold752 _4223_/Z _6759_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold763 _7149_/Q hold763/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold741 _6850_/Q hold741/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7298_ _7298_/D _7322_/RN _7319_/CLK _7298_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6318_ _7295_/Q _6594_/A3 _6387_/A1 _6337_/A4 _6318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold796 _4196_/Z _6737_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold774 _6756_/Q hold774/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold785 _5563_/Z _6954_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet829_461 _4150__22/I _6766_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet829_472 net829_473/I _6755_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6249_ _6302_/A1 _6302_/A2 hold77/I _7293_/Q _6250_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_130_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet829_483 net829_483/I _6744_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_494 net829_495/I _6733_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold90 hold90/I hold90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_63_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3950_ _3950_/A1 _3950_/A2 _3943_/Z _3950_/A4 _3958_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_189_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3881_ _5585_/A2 _3509_/Z _3504_/Z _5808_/A3 _4024_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_176_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5620_ hold59/Z hold451/Z _5623_/S _5620_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5551_ hold363/Z hold755/Z _5556_/S _6945_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _5162_/A2 _4702_/B _4502_/B _4502_/C _5061_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_117_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7221_ _7221_/D _7315_/RN _7221_/CLK _7221_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_129_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5482_ _5515_/A1 _5482_/A2 _5482_/B _5482_/C _5483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_6_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4433_ hold363/Z hold661/Z _4434_/S _4433_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4364_ _6628_/I0 _6860_/Q _4364_/S _6860_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7152_ _7152_/D _7243_/RN _7152_/CLK _7152_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_112_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6103_ _7214_/Q _6290_/A2 _6289_/A2 _7206_/Q _6106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7083_ _7083_/D _7322_/RN _7083_/CLK _7083_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4295_ hold109/Z hold79/Z _4303_/S _4295_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6034_ _7050_/Q _6291_/A2 _6295_/B1 _7002_/Q _7293_/Q _6035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6936_ _6936_/D _6694_/Z _7364_/CLK _6936_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_81_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _6867_/D _6880_/CLK _6867_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6798_ _6798_/D _7286_/RN _6798_/CLK _7382_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5818_ _6677_/A3 _5818_/A2 _5891_/A3 _5891_/A4 _5826_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_50_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5749_ hold2/Z hold94/Z _5749_/S hold95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold571 _7365_/Q hold571/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold560 _6911_/Q hold560/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold582 _4319_/Z _6823_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold593 _4294_/Z _6811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_46__1403_ clkbuf_4_15_0__1403_/Z net779_414/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _6017_/A3 _7285_/Q _5964_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _5395_/A1 _4975_/Z _5392_/A2 _5138_/A2 _4983_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3933_ _7245_/Q _4019_/A2 _4017_/B1 input62/Z _3963_/B1 _6852_/Q _3934_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6721_ _7359_/RN _7012_/Q _4069_/C _6721_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6652_ _6652_/I0 _7335_/Q _6668_/S _7335_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3864_ _6941_/Q _5909_/A3 _5557_/A2 hold68/I _3948_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5603_ hold50/Z hold127/Z _5605_/S _5603_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3795_ _3795_/A1 _3795_/A2 _3795_/A3 _3795_/A4 _3795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6583_ _6754_/Q _6319_/Z _6609_/B1 _6886_/Q _6587_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ _5534_/A1 _5534_/A2 _5534_/B1 _5410_/B _5534_/C _5535_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_172_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _5514_/A1 _5514_/A2 _5463_/Z _5514_/A3 _5467_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7204_ _7204_/D _7315_/RN _7204_/CLK _7204_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_105_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4416_ hold323/Z hold658/Z _4416_/S _6906_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5396_ _5396_/A1 _5330_/B _5396_/B1 _5475_/C _5396_/C _5452_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_132_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7135_ _7135_/D _7322_/RN _7135_/CLK _7135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4347_ _4435_/A1 hold68/Z _5557_/A2 _5891_/A1 _4349_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4278_ _4277_/Z hold602/Z _4286_/S _4278_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7066_ _7066_/D _7322_/RN _7066_/CLK _7066_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6017_ _7285_/Q _6017_/A2 _6017_/A3 _6808_/Q _6019_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/Z _4149_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6919_ _6919_/D _7315_/RN _6919_/CLK _6919_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold390 _5867_/Z _7215_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3580_ _5808_/A4 _4402_/A4 _3986_/A3 _5808_/A3 _4320_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_142_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5250_ _5250_/A1 _5421_/B _5250_/B1 _5250_/B2 _5251_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ hold38/Z hold424/Z _4202_/S _4201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5181_ _4691_/C _5461_/A4 _5319_/A1 _5133_/B _5182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ _6815_/Q input77/Z _4132_/S _4132_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4063_ _4063_/A1 _4063_/A2 _3409_/Z _3472_/B _6792_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet579_219 net579_219/I _7068_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet579_208 net629_264/I _7079_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4965_ _5142_/C _5155_/B2 _5326_/C _5329_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6704_ _7286_/RN _7012_/Q _4069_/C _6704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3916_ _7059_/Q _4009_/A2 _3916_/B1 _7067_/Q _3916_/C _3917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_149_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ _5417_/C _5199_/A3 _5457_/A1 _5306_/C _4898_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6635_ _6897_/Q _6635_/A2 _6635_/B1 _6898_/Q _6636_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_149_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3847_ _7060_/Q _4009_/A2 _4010_/A2 _7084_/Q _3847_/C _3850_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _6782_/Q _6566_/A2 _6593_/A3 _6594_/A3 _6572_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3778_ _7256_/Q _3778_/A2 _4045_/B1 _6957_/Q _3779_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5517_ _5517_/A1 _5517_/A2 _5517_/B _5518_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_92__1403_ clkbuf_4_4_0__1403_/Z net829_495/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6497_ _7055_/Q _6324_/Z _6331_/Z _7095_/Q _6498_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _5448_/A1 _5480_/A2 _5449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5379_ _5379_/A1 _5378_/Z _5383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7118_ _7118_/D _7286_/RN _7118_/CLK _7118_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7049_ _7049_/D _7286_/RN _7049_/CLK _7049_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _4829_/A4 _5406_/A1 _4750_/A3 _4835_/A1 _5491_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4681_ _4681_/A1 _5478_/A3 _4681_/A3 _5478_/A2 _4690_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3701_ _3701_/A1 _3701_/A2 _3701_/A3 _3701_/A4 _3702_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6420_ _7142_/Q _6323_/Z _6334_/Z _7028_/Q _6352_/Z _7150_/Q _6423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3632_ _5808_/A4 _4402_/A4 _5872_/A3 _4402_/A3 _4045_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6351_ _6351_/A1 _6351_/A2 _6351_/A3 _6613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_115_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5302_ _5302_/A1 _5412_/A2 _5302_/A3 _5302_/A4 _5307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3563_ _3505_/B _3503_/Z _3556_/C _3508_/Z hold641/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6282_ _7139_/Q _6292_/A2 _6291_/C1 _6753_/Q _6284_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3494_ _6726_/Q _3494_/A2 _3494_/B _7345_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5233_ _5241_/A1 _5353_/A3 _5241_/B1 _5371_/C _5233_/C _5446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5164_ _5164_/A1 _5164_/A2 _5164_/A3 _5163_/Z _5165_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_142_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ _6894_/Q _4115_/A2 _4117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _5093_/C _5095_/A2 _5323_/C _5096_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _7026_/Q _4046_/A2 _4046_/B1 _7130_/Q _4046_/C _4048_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_140_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5997_ _4083_/B _6387_/A2 _6337_/A4 _7296_/Q _6000_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4948_ _4991_/A1 _4991_/B _4991_/A2 _5325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_149_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ _4879_/A1 _4879_/A2 _4879_/A3 _4882_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _6618_/A1 _7323_/Q _6895_/D _6617_/B _6619_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ _7203_/Q _6313_/Z _6331_/Z _7097_/Q _6335_/Z hold29/I _6550_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_165_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput270 _6947_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput292 _6749_/Q pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput281 _6731_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4150__28 _4150__46/I _7259_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__17 _4150__25/I _7270_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__39 net429_61/I _7248_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xload_slew347 _5750_/A3 _5557_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5920_ hold323/Z hold800/Z _5926_/S _5920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ hold50/Z hold537/Z _5853_/S _7201_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4802_ _4802_/A1 _4802_/A2 _5361_/A3 _4804_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5782_ hold323/Z hold731/Z hold23/Z _7141_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4733_ _3399_/I _5112_/A1 _5460_/A1 _5180_/B2 _4764_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4664_ _5252_/A2 _4688_/A1 _5236_/A4 _5238_/B1 _5091_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6403_ _7277_/Q _6610_/A2 _6347_/C _7237_/Q _6404_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7383_ _7383_/I _7383_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold901 _7220_/Q hold901/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4595_ _4500_/B _4693_/B _5310_/B _5305_/B _5193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3615_ hold227/Z hold83/Z _3868_/A1 _3624_/A2 hold228/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6334_ _6566_/A2 _6387_/A2 _7294_/Q _6540_/A4 _6334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3546_ hold68/Z _3986_/A3 _3542_/C _3532_/Z _5588_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_135_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6265_ _7138_/Q _6299_/C _6265_/B1 _6782_/Q _6265_/C _6268_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_1_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ _5323_/B _5216_/A2 _5216_/B _5216_/C _5263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3477_ _3472_/B _3477_/A2 _7354_/Q _3478_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6196_ _6302_/A1 _6302_/A2 _6991_/Q _7293_/Q _6198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5147_ _5451_/B _5162_/A2 _5396_/A1 _5330_/B _5172_/A1 _5452_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_130_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _5209_/A1 _5534_/A2 _5377_/B _5228_/A2 _5378_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4029_ _4029_/A1 _4029_/A2 _4029_/A3 _4029_/A4 _4035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_44_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold208 _5728_/Z _7094_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3400_ _3400_/I _5460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_20
XFILLER_171_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet429_61 net429_61/I _7226_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_72 net429_72/I _7215_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold219 _6960_/Q hold219/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4380_ _6891_/Q _7341_/RN _4388_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet429_83 net429_83/I _7204_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_94 net429_97/I _7193_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3331_ _6794_/Q _4160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_124_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6050_ _7196_/Q _6293_/A2 _6292_/A2 _6760_/Q _6052_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _5342_/A2 _4796_/Z _5024_/A4 _5336_/A3 _5002_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _6952_/D _7300_/RN _6952_/CLK _6952_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5903_ hold99/Z hold431/Z _5908_/S _5903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6883_ _6883_/D input75/Z _6883_/CLK _6883_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5834_ hold38/Z hold231/Z _5835_/S _5834_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ hold50/Z hold86/Z _5767_/S hold87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4716_ _4758_/A3 _4758_/A4 _4716_/B _4829_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5696_ _5909_/A3 _5891_/A1 _5750_/A3 _5750_/A4 hold84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4647_ _5322_/A2 _5417_/C _5416_/C _4906_/A1 _4649_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_163_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7366_ _7366_/D _6718_/Z _3753_/A1 _7366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold720 _5733_/Z _7098_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4578_ _5482_/C _4577_/Z _5369_/B _4582_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _7297_/Q _7296_/Q _6543_/A2 _6594_/A3 _6317_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xhold753 _7359_/Q hold753/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold731 _7141_/Q hold731/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold764 _6745_/Q hold764/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold742 _7035_/Q hold742/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7297_ _7297_/D _7315_/RN _4144_/I1 _7297_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_131_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3529_ _4178_/S hold226/Z _3529_/B _3545_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_1_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold797 _6729_/Q hold797/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold775 _4219_/Z _6756_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold786 _6774_/Q hold786/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xnet829_462 net429_76/I _6765_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6248_ _6265_/C _6248_/A2 _6247_/Z _6289_/B1 _6248_/C _6250_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet829_473 net829_473/I _6754_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6179_ _6765_/Q _6292_/A2 _6293_/B1 _7185_/Q _6182_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet829_484 net829_496/I _6743_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_495 net829_495/I _6732_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold91 hold91/I hold91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold80 hold80/I hold80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_36_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_69__1403_ clkbuf_4_7_0__1403_/Z net679_327/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3880_ _6775_/Q _6677_/A1 _4426_/A3 _3940_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_188_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5550_ _5550_/A1 _5836_/A3 hold228/Z _6677_/A3 hold229/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4501_ _3399_/I _5162_/A2 _4452_/Z _4454_/Z _4502_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_129_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _5481_/A1 _5481_/A2 _5481_/A3 _5442_/Z _5481_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_8_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7220_ _7220_/D _7315_/RN _7220_/CLK _7220_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4432_ _5936_/A1 _4305_/C _5927_/A3 hold185/Z _4434_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4363_ _6627_/I0 _6859_/Q _4364_/S _6859_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7151_ _7151_/D input75/Z _7151_/CLK _7151_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6102_ _7052_/Q _6291_/A2 _6102_/B _6102_/C _6114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7082_ _7082_/D _7322_/RN _7082_/CLK _7082_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4294_ hold592/Z _4293_/Z _4304_/S _4294_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6033_ _6043_/A1 _7289_/Q _7292_/Q _7291_/Q _6295_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _6935_/D _6693_/Z _7364_/CLK _6935_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _6866_/D _6880_/CLK _6866_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6797_ _6797_/D _7286_/RN _6797_/CLK _7381_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5817_ hold27/Z hold2/Z _5817_/S hold28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5748_ hold38/Z hold199/Z _5749_/S _5748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ hold363/Z hold746/Z hold19/Z _7050_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold550 _6824_/Q hold550/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7349_ _7349_/D _6703_/Z _4149_/B2 hold58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold572 hold572/I hold572/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold561 _4424_/Z _6911_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold583 _7100_/Q hold583/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold594 _6778_/Q hold594/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_1_0__1403_ net479_128/I clkbuf_opt_1_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4981_ _4794_/Z _5171_/A2 _5336_/A2 _5331_/A3 _5451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_64_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3932_ input44/Z _4285_/S _3985_/B1 _6755_/Q _3934_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6720_ _7359_/RN _7012_/Q _4069_/C _6720_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6651_ _6651_/A1 _6651_/A2 _6652_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3863_ _6779_/Q _5560_/A1 _5732_/A4 _6677_/A1 _3945_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5602_ hold59/Z hold402/Z _5605_/S _5602_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6582_ _6790_/Q _6318_/Z _6608_/B1 _6915_/Q _6341_/Z _6849_/Q _6587_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_164_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5533_ _4787_/B _5310_/C _5533_/A3 _5535_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3794_ _6997_/Q _3963_/A2 _3951_/B1 _7125_/Q _3795_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _5421_/C _5464_/A2 _5533_/A3 _5309_/B _5464_/C _5514_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5395_ _5395_/A1 _5395_/A2 _4975_/Z _5440_/A2 _5396_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7203_ _7203_/D _7243_/RN _7203_/CLK _7203_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4415_ hold363/Z hold657/Z _4416_/S _6905_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4346_ hold2/Z hold4/Z _4346_/S hold5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7134_ _7134_/D _7243_/RN _7134_/CLK _7134_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4277_ hold158/Z hold79/Z _4285_/S _4277_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7065_ _7065_/D _7322_/RN _7065_/CLK _7065_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6016_ _6613_/C _4062_/Z _6014_/Z _6016_/B _7301_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_2007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_52__1403_ clkbuf_4_15_0__1403_/Z net629_301/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _6918_/D _7315_/RN _6918_/CLK _6918_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _6849_/D _7359_/RN _6849_/CLK _6849_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold380 _5896_/Z _7240_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold391 _7047_/Q hold391/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ hold50/Z hold465/Z _4202_/S _4200_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5180_ _5515_/A1 _5294_/B _5133_/B _5180_/B2 _5184_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4131_ _6817_/Q input67/Z _7364_/Q _4131_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4062_ _7301_/Q _6957_/Q _6962_/Q _4062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_49_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet579_209 net679_327/I _7078_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _5155_/B2 _4964_/A2 _4964_/A3 _4716_/B _5327_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_36_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6703_ _7286_/RN _7012_/Q _4069_/C _6703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3915_ _3915_/A1 _3915_/A2 _3915_/A3 _3915_/A4 _3915_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_149_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4895_ _5198_/A1 _4751_/B _5416_/A2 _4691_/C _5464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6634_ _6672_/A2 _6673_/A2 _6635_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3846_ _7100_/Q _4006_/B1 _4008_/A2 _7092_/Q _4010_/B1 _7116_/Q _3858_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6565_ _6565_/A1 _6565_/A2 _6434_/S _6565_/B2 _7320_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3777_ _7248_/Q _4019_/A2 _4017_/B1 _7399_/I _3779_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5516_ _5516_/A1 _5516_/A2 _5517_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6496_ _7087_/Q _6325_/Z _6329_/Z _7015_/Q _6498_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5447_ _5442_/Z _5488_/A1 _5523_/A2 _5448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_160_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _5378_/A1 _5378_/A2 _5378_/A3 _5378_/A4 _5378_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7117_ _7117_/D _7286_/RN _7117_/CLK _7117_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4329_ _5588_/A1 _5564_/A1 _5597_/A3 _6677_/A3 _4337_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_59_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7048_ _7048_/D _7315_/RN _7048_/CLK _7048_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _5909_/A3 _5566_/A1 _4008_/A2 _7096_/Q _3701_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_187_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4680_ _5384_/B _5384_/C _5228_/B _5497_/A1 _5478_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _4402_/A4 _5872_/A3 _4402_/A3 _3830_/B _3947_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_174_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6350_ _6349_/Z _6609_/B1 _6326_/Z _6351_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3562_ _4402_/A4 _5872_/A3 _5642_/A3 _4402_/A3 _4041_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5301_ _5461_/A4 _5497_/A1 _5493_/A1 _5301_/B _5412_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_52_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6281_ _6757_/Q _6295_/B1 _6292_/B1 _6791_/Q _6284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3493_ input58/Z _6727_/Q _6725_/Q _6792_/Q _3494_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5232_ _5417_/C _5234_/A2 _5417_/B _5234_/B1 _4515_/Z _5233_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5163_ _4796_/Z _5176_/A2 _5336_/A3 _5342_/A2 _5163_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_111_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4114_ _4114_/A1 _4160_/B _3421_/B _4114_/B2 _6794_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5094_ _5095_/A2 _5384_/B _5384_/C _5238_/B1 _5479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4045_ _7050_/Q _4045_/A2 _4045_/B1 _7284_/Q input20/Z _4045_/C2 _4049_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_64_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5996_ _6807_/Q _5996_/A2 _6006_/B1 _6387_/A2 _7295_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _4949_/A1 _4502_/B _4963_/A2 _4963_/A3 _5331_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_33_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4878_ _4452_/Z _5490_/B _5421_/A2 _4773_/C _4879_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6617_ _6895_/D _6888_/Q _6616_/Z _6617_/B _6618_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_137_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3829_ _7068_/Q _5750_/A4 _5909_/A3 _5750_/A3 _3847_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ _7235_/Q _6599_/A2 _6329_/Z _7017_/Q _6338_/Z _7081_/Q _6550_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _7280_/Q _6610_/A2 _6328_/Z _6764_/Q _6347_/C _7240_/Q _6481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_133_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput260 _6953_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput271 _6744_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput293 _6750_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput282 _6745_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150__29 _4150__46/I _7258_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4150__18 net429_59/I _7269_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xload_slew359 _5863_/A3 _5759_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xload_slew348 _6677_/A1 _5818_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_66_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_290 net429_57/I _6997_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5850_ hold59/Z hold205/Z _5853_/S _5850_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4801_ _3399_/I _5280_/B _5460_/A1 _5319_/A1 _5361_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ hold363/Z hold732/Z hold23/Z _7140_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4732_ _5268_/B _4787_/B _4832_/A1 _5270_/A2 _5272_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_4663_ _3399_/I _5162_/A2 _4688_/A1 _5180_/B2 _5382_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6402_ _7253_/Q _6319_/Z _6328_/Z _6761_/Q _6610_/B1 _7269_/Q _6404_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3614_ _3556_/B _3548_/B _5872_/A3 _5808_/A2 _4024_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7382_ _7382_/I _7382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold902 _5873_/Z _7220_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4594_ _4773_/C _4694_/B _4787_/B _4702_/B _5462_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_155_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6333_ _7298_/Q _6339_/A1 _7299_/Q _6355_/A4 _6608_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3545_ _6881_/Q _4060_/I0 _3545_/B _3986_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_170_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _6264_/I _6274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3476_ _4113_/A3 _7355_/Q _3477_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _5210_/Z _5424_/C _5507_/A2 _5468_/A2 _5215_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_85_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6195_ _7293_/Q _6195_/A2 _6195_/B _6198_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5146_ _5368_/A2 _5324_/A3 _5176_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ _5241_/A1 _5534_/A2 _5241_/B1 _5075_/Z _5378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4028_ _7212_/Q _4028_/A2 _4028_/B1 _7358_/Q _4029_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ _6245_/C _7291_/Q _7290_/Q _7289_/Q _6291_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_40_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_29__1403_ clkbuf_4_14_0__1403_/Z _4150__5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_109__1403_ net779_410/I net829_482/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_172_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet429_62 _4150__6/I _7225_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_73 net429_73/I _7214_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold209 _7056_/Q hold209/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3330_ _6795_/Q _3421_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
Xnet429_95 net429_95/I _7192_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_84 net429_86/I _7203_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _5014_/A1 _5391_/B _5000_/B _5000_/C _5002_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _6951_/D _7300_/RN _6951_/CLK _6951_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_35_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5902_ hold323/Z hold646/Z _5908_/S _5902_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6882_ _6882_/D input75/Z _6882_/CLK _6882_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5833_ hold50/Z hold143/Z _5835_/S _5833_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5764_ hold59/Z hold192/Z _5767_/S _5764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ _4792_/A1 _4730_/C _4715_/B _4758_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_163_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5695_ hold2/Z hold429/Z _5695_/S _5695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4646_ _4518_/Z _5417_/C _5475_/A1 _4906_/A1 _4649_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_30_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4577_ _5384_/A2 _5229_/A2 _4577_/A3 _5065_/A2 _4577_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
Xhold710 _7380_/I hold710/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7365_ _7365_/D _6717_/Z _3753_/A1 _7365_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold721 _7214_/Q hold721/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6316_ _7297_/Q _7296_/Q _6594_/A2 _6594_/A3 _6316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xhold754 _6679_/Z _7359_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold732 _7140_/Q hold732/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold743 _7123_/Q hold743/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7296_ _7296_/D _7315_/RN _4144_/I1 _7296_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_116_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ _6881_/Q hold10/Z _3529_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold765 _4205_/Z _6745_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold776 _6780_/Q hold776/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold787 _4243_/Z _6774_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet829_463 _4150__48/I _6764_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6247_ _7025_/Q _7147_/Q _7293_/Q _6247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold798 _4181_/Z _6729_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3459_ _7362_/Q _7345_/Q _3459_/S _7362_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet829_452 net829_452/I _6775_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet829_496 net829_496/I _6731_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_485 net829_499/I _6742_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_474 net829_475/I _6753_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6178_ _7161_/Q _6295_/A2 _6292_/B1 _7193_/Q _6182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5129_ _5440_/A2 _5287_/A2 _5534_/B1 _5421_/B _5129_/C _5132_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold92 hold92/I hold92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold70 hold70/I hold70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold81 hold81/I hold81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_63_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4500_ _5294_/B _5460_/A2 _4500_/B _4502_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_145_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5480_ _5262_/B _5480_/A2 _5479_/Z _5480_/A4 _5481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4431_ hold323/Z hold686/Z _4431_/S _4431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4362_ _3745_/Z _6858_/Q _4364_/S _6858_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7150_ _7150_/D _7300_/RN _7150_/CLK _7150_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_98_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6101_ _6121_/A3 _6101_/A2 _6101_/B _6102_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7081_ _7081_/D _7322_/RN _7081_/CLK _7081_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4293_ _6841_/Q hold99/Z _4303_/S _4293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6032_ _7106_/Q _6294_/A2 _6293_/A2 _7074_/Q _6035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _6934_/D _6692_/Z _3753_/A1 _6934_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_54_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _6865_/D _7325_/CLK _6865_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5816_ hold450/Z hold38/Z _5817_/S _7170_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6796_ _6796_/D _6687_/Z _7364_/CLK _6796_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5747_ hold50/Z hold96/Z _5749_/S hold97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5678_ _5891_/A1 _5678_/A2 _5891_/A3 _5891_/A4 hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_135_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4629_ _5462_/A2 _5421_/C _5319_/A1 _5308_/B _4630_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_12__1403_ clkbuf_opt_1_0__1403_/Z net779_431/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold551 _4321_/Z _6824_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7348_ _7348_/D _6702_/Z _4149_/B2 hold78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold540 _7378_/I hold540/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold562 _6885_/Q hold562/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_75__1403_ clkbuf_4_7_0__1403_/Z net729_389/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_173_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _7279_/D _7286_/RN _7279_/CLK _7279_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold573 _3565_/B hold573/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold595 _4249_/Z _6778_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold584 _6900_/Q hold584/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput160 wb_rstn_i _7341_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_63_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _5326_/C _5220_/A3 _5325_/A2 _5392_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_63_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3931_ _3931_/A1 _3931_/A2 _3931_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6650_ _6896_/Q _6650_/A2 _6650_/B1 _6666_/B2 _6651_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3862_ _7075_/Q _4006_/A2 _4010_/B1 _7115_/Q _3917_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5601_ hold79/Z hold148/Z _5605_/S _5601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6581_ _6572_/Z _6575_/Z _6579_/Z _6581_/A4 _6581_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_176_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3793_ input67/Z _4303_/S _4320_/S input38/Z _4017_/B1 input64/Z _3795_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5532_ hold10/I _4395_/C _5537_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ _5463_/A1 _5463_/A2 _5463_/A3 _5463_/A4 _5463_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_8_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5394_ _5394_/A1 _5332_/C _5399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _7202_/D _7286_/RN _7202_/CLK _7202_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4414_ _6677_/A3 _5777_/A2 _5557_/A2 hold83/Z _4416_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7133_ _7133_/D _7286_/RN _7133_/CLK _7133_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_125_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4345_ hold38/Z hold40/Z _4346_/S hold41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4276_ _4275_/Z hold613/Z _4286_/S _4276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7064_ _7064_/D _7315_/RN _7064_/CLK _7064_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6015_ _6014_/Z _7301_/Q _6016_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6917_ _6917_/D _7315_/RN _6917_/CLK _6917_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6848_ _6848_/D _7322_/RN _6848_/CLK _6848_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6779_ _6779_/D _7359_/RN _6779_/CLK _6779_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold381 _6835_/Q hold381/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold370 _4187_/Z _6732_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold392 _5675_/Z _7047_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ _6818_/Q _4149_/B2 _7363_/Q _4130_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4061_ _3423_/S _4060_/Z _4061_/B _6724_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4963_ _4991_/B _4963_/A2 _4963_/A3 _5183_/A2 _5155_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6702_ _7286_/RN _7012_/Q _4069_/C _6702_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3914_ _7221_/Q _3914_/A2 _3914_/B1 _6729_/Q _4033_/B1 _6773_/Q _3915_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_189_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ _6673_/A2 _6671_/A3 _6635_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4894_ _5308_/B _5322_/A2 _5490_/B _5353_/A4 _5282_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ _3845_/A1 _3845_/A2 _3845_/A3 _3845_/A4 _3845_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6564_ _5951_/B _7319_/Q _6614_/B _6565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3776_ _3776_/A1 _3776_/A2 _3776_/A3 _3776_/A4 _3784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5515_ _5515_/A1 _5517_/A2 _5515_/B1 _5490_/B _5516_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6495_ _7233_/Q _6599_/A2 _6608_/B1 hold96/I _6326_/Z _7265_/Q _6498_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5446_ _5446_/A1 _5446_/A2 _5372_/Z _5446_/A4 _5523_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_172_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5377_ _5515_/A1 _5482_/A2 _5377_/B _5378_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7116_ _7116_/D _7286_/RN _7116_/CLK _7116_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4328_ hold50/Z _6830_/Q _4328_/S _4328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7047_ _7047_/D _7315_/RN _7047_/CLK _7047_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4259_ hold323/Z hold352/Z _4259_/S _4259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1_0__1403_ clkbuf_0__1403_/Z clkbuf_4_3_0__1403_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3630_ _6767_/Q _5780_/A3 _5863_/A3 _6677_/A1 _3643_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3561_ _6881_/Q _4060_/I0 _3561_/B hold11/Z hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_155_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5300_ _5310_/A1 _5300_/A2 _5300_/B _5300_/C _5302_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6280_ _6434_/S _6280_/A2 _6280_/B _7311_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xnet679_350 net729_367/I _6929_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3492_ _3492_/A1 _7345_/Q _3494_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5231_ _5373_/A4 _5231_/A2 _5230_/Z _5235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _5333_/B _5162_/A2 _5396_/A1 _5161_/B _5172_/A1 _5164_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_130_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5093_ _5515_/A1 _5421_/A2 _5213_/B _5093_/C _5478_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_69_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4113_ _4114_/B2 _7355_/Q _4113_/A3 _7354_/Q _4114_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_111_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4044_ _4044_/A1 _4044_/A2 _4044_/A3 _4044_/A4 _4044_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_92_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5995_ _6543_/A2 _6376_/A2 _5996_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4946_ _5304_/A1 _5473_/A1 _5473_/B _5338_/A2 _5032_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4877_ _5462_/A4 _5322_/A2 _5490_/B _5353_/A4 _4879_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_165_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6616_ _6892_/Q _6895_/Q _6616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_137_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3828_ _7076_/Q hold22/I _5863_/A3 _4423_/A2 _3850_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6547_ _6547_/A1 _6547_/A2 _6547_/A3 _6547_/A4 _6556_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_152_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3759_ _7232_/Q _4033_/A2 _4010_/B1 _7118_/Q _3761_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6478_ _7022_/Q _6321_/Z _6609_/B1 _7046_/Q _6482_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5429_ hold21/I _4395_/C _5429_/B _5430_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput250 _4168_/Z pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput261 _6939_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput294 _6751_/Q pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput272 _6738_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput283 _6732_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4150__19 net429_59/I _7268_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet629_280 net629_281/I _7007_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_291 net629_291/I _6996_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _5268_/B _4787_/B _4832_/A1 _5283_/A4 _5280_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_2180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ _5891_/A1 _5818_/A2 _5780_/A3 _5891_/A3 hold23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4731_ _5268_/B _4787_/B _4832_/A1 _5270_/A2 _5112_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_175_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _4689_/A2 _4641_/C _5014_/A1 _3402_/I _5261_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6401_ _7189_/Q _6318_/Z _6608_/B1 _7107_/Q _6341_/Z _6995_/Q _6405_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3613_ _5808_/A4 _3830_/C _3523_/B _3554_/B _3914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7381_ _7381_/I _7381_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold903 _7381_/I hold903/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4593_ _4689_/A2 _5060_/C _5439_/A1 _5304_/A1 _4598_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_127_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6332_ _6343_/A4 _6339_/A1 _7299_/Q _7297_/Q _6604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3544_ _3624_/A2 hold11/Z _5909_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_116_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ _6886_/Q _6290_/B1 _7293_/Q _6264_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3475_ _6792_/Q _3482_/B _7355_/Q _3478_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5214_ _5319_/A1 _5228_/B _5218_/B _5214_/A4 _5468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_130_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6194_ _7290_/Q _7289_/Q _6194_/A3 _6193_/Z _7293_/Q _6195_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5145_ _4691_/C _5323_/C _5323_/B _5333_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_96_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _5209_/A1 _5410_/B _5087_/B2 _5075_/Z _5522_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4027_ _7276_/Q _4027_/A2 _4027_/B1 _7252_/Q _4027_/C _4029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ _5978_/I _7291_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _4794_/Z _4929_/A2 _4929_/A3 _4483_/B _5344_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_100_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet429_52 net429_89/I _7235_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_63 net429_63/I _7224_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet429_85 _4150__6/I _7202_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet429_74 net429_74/I _7213_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_96 net429_96/I _7191_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _6950_/D input75/Z _6950_/CLK _6950_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5901_ hold363/Z hold648/Z _5908_/S _5901_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6881_ _6881_/D _7341_/RN _7341_/CLK _6881_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_35_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ hold59/Z hold442/Z _5835_/S _5832_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ hold79/Z hold133/Z _5767_/S _5763_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4714_ _5305_/B _4793_/A1 _4945_/A4 _4730_/A2 _4758_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5694_ hold38/Z hold354/Z _5695_/S _5694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4645_ _4500_/B _4773_/C _4694_/B _4787_/B _4906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold711 _6831_/Q hold711/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_146_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4576_ _5102_/A1 _5475_/A2 _3399_/I _5162_/A2 _5229_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_7364_ _7364_/D _6716_/Z _7364_/CLK _7364_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold700 _4367_/Z _6862_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6315_ _7298_/Q _6543_/A2 _6594_/A4 _6007_/B _6315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _6881_/Q hold226/I _3530_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold722 _6910_/Q hold722/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold755 _6945_/Q hold755/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold744 _5761_/Z _7123_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold733 _6883_/Q hold733/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold788 _7115_/Q hold788/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _7295_/D _7315_/RN _7319_/CLK _7295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_115_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold766 _7189_/Q hold766/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold777 _4252_/Z _6780_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold799 _7205_/Q hold799/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6246_ _6246_/A1 _7289_/Q _7290_/Q _6248_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3458_ _3497_/A2 _6725_/Q _3459_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xnet829_453 net829_453/I _6774_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_464 net429_81/I _6763_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3389_ _7317_/Q _6485_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ hold63/I _6291_/A2 _6291_/C1 hold86/I _6294_/B1 _7225_/Q _6183_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xnet829_486 net829_499/I _6741_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_497 net429_95/I _6730_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_475 net829_475/I _6752_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5128_ _5128_/A1 _5431_/A2 _5128_/A3 _5362_/A4 _5129_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5059_ _5384_/A1 _5059_/A2 _5261_/A2 _5482_/C _5369_/C _5064_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xclkbuf_4_4_0__1403_ clkbuf_4_5_0__1403_/I clkbuf_4_4_0__1403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_38_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_35__1403_ clkbuf_4_10_0__1403_/Z net429_82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_115__1403_ net779_410/I net429_96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_98__1403_ clkbuf_4_4_0__1403_/Z net429_70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_186_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold82 hold82/I hold82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold60 hold60/I hold60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold71 hold71/I hold71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold93 hold93/I hold93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_63_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ hold363/Z hold688/Z _4431_/S _4430_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6100_ _6100_/A1 _6100_/A2 _6100_/A3 _6101_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4361_ _6625_/I0 _6857_/Q _4364_/S _6857_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7080_ _7080_/D _7322_/RN _7080_/CLK _7080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4292_ hold850/Z _4291_/Z _4304_/S _4292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6031_ _6043_/A1 _6231_/A1 _6245_/C _7291_/Q _6293_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _6933_/D _6691_/Z _7364_/CLK _6933_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_179_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _6864_/D _6880_/CLK _6864_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_179_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5815_ hold72/Z hold50/Z _5817_/S hold73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6795_ _6795_/D _6686_/Z _4152_/I1 _6795_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_50_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ hold59/Z hold241/Z _5749_/S _5746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5677_ hold2/Z hold150/Z _5677_/S _5677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4628_ _4773_/C _5310_/B _4694_/B _4702_/B _5198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold530 _7023_/Q hold530/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4559_ _5460_/A1 _5460_/A2 _5417_/C _5344_/C _5369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7347_ _7347_/D _6701_/Z _4149_/B2 hold98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold552 _7092_/Q hold552/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold541 _4304_/Z _6816_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold563 _4401_/Z _6885_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7278_ _7278_/D _7286_/RN _7278_/CLK _7278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold574 hold574/I hold574/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold596 _6779_/Q hold596/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold585 _4407_/Z _6900_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ hold42/I _6290_/A2 _6289_/A2 _7211_/Q hold25/I _6291_/A2 _6230_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_18_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput150 wb_dat_i[2] _6646_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput161 wb_sel_i[0] _6629_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3930_ _7189_/Q _3930_/A2 _4019_/B1 _6946_/Q _3931_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_81__1403_ clkbuf_4_5_0__1403_/Z net779_427/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3861_ _3860_/Z _6932_/Q _3961_/S _6932_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ hold99/Z hold180/Z _5605_/S _5600_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3792_ _7279_/Q _5936_/A1 hold7/I hold32/I _3795_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6580_ _6776_/Q _6317_/Z _6354_/Z _6780_/Q _6387_/Z _6901_/Q _6581_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _5503_/Z _5531_/A2 _5531_/B _5531_/C _5537_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5462_ _4751_/B _5462_/A2 _5490_/B _5462_/A4 _5463_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7201_ _7201_/D _7243_/RN _7201_/CLK _7201_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5393_ _5394_/A1 _5332_/C _5393_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4413_ hold323/Z hold634/Z _4413_/S _4413_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ hold50/Z hold61/Z _4346_/S hold62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7132_ _7132_/D _7243_/RN _7132_/CLK _7132_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ _7063_/D _7322_/RN _7063_/CLK _7063_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ hold188/Z hold99/Z _4285_/S _4275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6014_ _6014_/I0 _6014_/I1 _6808_/Q _6014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _6916_/D _7359_/RN _6916_/CLK _6916_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6847_ _6847_/D _7243_/RN _6847_/CLK _6847_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6778_ _6778_/D _7359_/RN _6778_/CLK _6778_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ hold50/Z _7095_/Q _5731_/S hold51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold371 _7128_/Q hold371/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold360 _6743_/Q hold360/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold382 _4334_/Z _6835_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold393 _6989_/Q hold393/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4060_ _4060_/I0 _3536_/B _4060_/S _4060_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _5338_/A2 _4787_/B _4694_/B _5324_/A4 _5397_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_51_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6701_ _7286_/RN _7012_/Q _4069_/C _6701_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4893_ _4915_/A3 _5417_/C _5306_/C _5134_/A4 _5200_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3913_ _7107_/Q _4009_/B1 _3913_/B1 _6912_/Q _3915_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6632_ _6894_/Q _6632_/A2 _6632_/B1 _6896_/Q _6636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_3844_ input13/Z _4031_/A2 _4009_/B1 _7108_/Q _3845_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _6556_/Z _6563_/A2 hold77/I _6613_/A2 _6613_/C _6565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3775_ _7078_/Q _4006_/A2 _4019_/B1 _6949_/Q _3776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5514_ _5514_/A1 _5514_/A2 _5514_/A3 _5514_/A4 _5519_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6494_ _6494_/A1 _6494_/A2 _6494_/A3 _6493_/Z _6494_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5445_ _5534_/A1 _5445_/A2 _5445_/B1 _5482_/A2 _5446_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7115_ _7115_/D _7315_/RN _7115_/CLK _7115_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5376_ _5376_/A1 _5376_/A2 _5523_/A1 _5379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_160_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ hold59/Z hold384/Z _4328_/S _6829_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _7046_/D _7315_/RN _7046_/CLK _7046_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4258_ hold363/Z _6784_/Q _4259_/S _4258_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4189_ hold50/Z hold327/Z _4193_/S _4189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold190 _7216_/Q hold190/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_93_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3560_ hold68/Z _3624_/A2 _3533_/Z _3545_/B _5669_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ _7346_/Q input58/Z _3491_/S _7346_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5230_ _5487_/A3 _5486_/A1 _5487_/A1 _5373_/A3 _5230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet679_340 net829_483/I _6947_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet679_351 net779_438/I _6928_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5161_ _5368_/A2 _5324_/A3 _5161_/B _5164_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _5092_/A1 _5442_/A1 _5096_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ _4112_/A1 _7345_/Q _7344_/Q _3421_/B _3409_/Z _6795_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_56_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ input4/Z _4043_/A2 _4043_/B1 _6884_/Q _4044_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5994_ _6337_/A4 _7295_/Q _6376_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4945_ _5441_/A4 _4794_/Z _5401_/A2 _4945_/A4 _5473_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_52_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _4876_/A1 _4876_/A2 _4876_/A3 _4879_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_177_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3827_ _7214_/Q hold7/I _5863_/A3 _5882_/A2 _3845_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6615_ _6615_/A1 _6615_/A2 _6434_/S _6615_/B2 _7322_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3758_ _7208_/Q _4037_/A2 _4010_/A2 _7086_/Q _3761_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6546_ _7187_/Q _6320_/Z _6325_/Z hold88/I _6547_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6477_ _7192_/Q _6318_/Z _6608_/B1 _7110_/Q _6341_/Z _6998_/Q _6482_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3689_ _6742_/Q _4040_/B1 _4010_/A2 _7088_/Q _3693_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5428_ _4392_/Z _5469_/A3 _5506_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput251 _4157_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput262 _6940_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput240 _7375_/Z mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5359_ _5359_/A1 _5359_/A2 _5268_/B _5405_/A1 _4775_/Z _5360_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_161_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput295 _6736_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput284 _6733_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput273 _6739_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _7029_/D _7300_/RN _7029_/CLK hold90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet629_270 net679_327/I _7017_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_281 net629_281/I _7006_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet629_292 net429_87/I _6995_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4730_ _4806_/A3 _4730_/A2 _4730_/B _4730_/C _5270_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_1491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _5295_/B2 _5322_/A2 _3399_/I _5162_/A2 _5339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_159_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7380_ _7380_/I _7380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3612_ _3523_/B _3554_/B _3556_/B _3548_/B _6677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6400_ _6396_/Z _6400_/A2 _6400_/A3 _6400_/A4 _6406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold904 _4272_/Z _6797_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_128_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4592_ _5384_/B _5099_/C _4689_/A2 _5060_/C _5445_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6331_ _7297_/Q _7296_/Q _6376_/A2 _6540_/A4 _6331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_116_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3543_ _5750_/A4 _3868_/A1 _4402_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_143_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _6258_/Z _6262_/A2 _6262_/A3 _6262_/A4 _6262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3474_ _3482_/B _4113_/A3 _3480_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5213_ _5517_/A1 _5413_/A2 _5213_/B _5218_/B _5507_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_103_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6193_ _6193_/A1 _6193_/A2 _6193_/A3 _6192_/Z _6193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5144_ _5387_/A1 _5450_/C _5450_/B _5144_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_130_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5075_ _5239_/A3 _4499_/B _4591_/C _5075_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_57_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4026_ _4026_/A1 _4026_/A2 _4027_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _5976_/Z _6807_/Q _7291_/Q _6006_/B1 _5978_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4928_ _4794_/Z _4929_/A2 _4929_/A3 _4483_/B _5450_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _5460_/A2 _4787_/B _4694_/B _5162_/A2 _5183_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_181_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6529_ _7226_/Q _6317_/Z _6323_/Z hold48/I _6530_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_58__1403_ net429_73/I net579_207/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet429_53 net429_54/I _7234_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_64 net429_64/I _7223_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet429_97 net429_97/I _7190_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_75 net429_75/I _7212_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_86 net429_86/I _7201_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5900_ hold116/Z _5909_/A2 _5900_/A3 _4305_/C _5908_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_47_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6880_ _6880_/D _6880_/CLK _6880_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_179_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ hold79/Z hold453/Z _5835_/S _5831_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5762_ hold99/Z hold320/Z _5767_/S _5762_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4713_ _4718_/A3 _4718_/A2 _4835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5693_ hold50/Z hold519/Z _5695_/S _5693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4644_ _4693_/B _5310_/B _4702_/B _5305_/B _5421_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold712 _4330_/Z _6831_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4575_ _5214_/A4 _5460_/A1 _5295_/B2 _3402_/I _5234_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7363_ _7363_/D _6715_/Z _4152_/I1 _7363_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold701 _6781_/Q hold701/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7294_ _7294_/D _7315_/RN _7319_/CLK _7294_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6314_ _6340_/A1 _7295_/Q _6337_/A4 _6610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3526_ hold225/Z _6795_/Q _7371_/Q hold226/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xhold723 _4422_/Z _6910_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold745 _7002_/Q hold745/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold734 _4398_/Z _6883_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold756 _7159_/Q _3367_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6245_ _6265_/C _7121_/Q _6245_/B _6245_/C _6246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xhold767 _5838_/Z _7189_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold778 _7090_/Q hold778/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold789 _5752_/Z _7115_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet829_454 _4150__3/I _6773_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3457_ _6727_/Q _6726_/Q _6792_/Q _3497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet829_465 net429_81/I _6762_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3388_ _7316_/Q _6460_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6176_ _7233_/Q _6294_/A2 _6289_/A2 _7209_/Q _6183_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet829_487 net829_499/I _6740_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_476 net829_482/I _6751_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5127_ _5406_/A1 _5284_/A2 _5130_/B1 _5421_/B _5362_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet829_498 net829_498/I _6729_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5058_ _5099_/C _5058_/A2 _5368_/A3 _4523_/C _5369_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_29_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4009_ _7058_/Q _4009_/A2 _4009_/B1 _7106_/Q _4009_/C _4011_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 hold50/I hold50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold83 hold83/I hold83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold61 hold61/I hold61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold72 hold72/I hold72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold94 hold94/I hold94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _6624_/I0 _6856_/Q _4364_/S _6856_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_41__1403_ clkbuf_4_14_0__1403_/Z net429_89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4291_ hold598/Z hold323/Z _4303_/S _4291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6030_ _6043_/A1 _6231_/A1 _6245_/C _6245_/B _6294_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6932_ _6932_/D _6690_/Z _7364_/CLK _6932_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_35_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _6863_/D _6880_/CLK _6863_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5814_ hold194/Z hold59/Z _5817_/S _5814_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ _6794_/D _6685_/Z _7364_/CLK _6794_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5745_ hold79/Z hold154/Z _5749_/S _5745_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5676_ hold38/Z hold348/Z _5677_/S _5676_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4627_ _4500_/B _4693_/B _4787_/B _5305_/B _5308_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_136_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold520 _5693_/Z _7063_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4558_ _4500_/B _4773_/C _4693_/B _5310_/B _5344_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7346_ _7346_/D _6700_/Z _4149_/B2 _7346_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold553 _7262_/Q hold553/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold542 _7060_/Q hold542/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold531 _6776_/Q hold531/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7277_ _7277_/D _7286_/RN _7277_/CLK _7277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold575 hold575/I _5877_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4489_ _5441_/A4 _5382_/A1 _5382_/A2 _5099_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_104_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3509_ _3556_/C _3508_/Z _3509_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
Xhold586 _6899_/Q hold586/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold564 _6938_/Q hold564/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold597 _4250_/Z _6779_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _7163_/Q _6295_/A2 _6294_/B1 _7227_/Q _6230_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ hold71/I _6291_/A2 _6292_/A2 _7014_/Q _6160_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput162 wb_sel_i[1] _6671_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput151 wb_dat_i[30] _6661_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput140 wb_dat_i[20] _6654_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ _6931_/Q _3859_/Z _3960_/S _3860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3791_ _7061_/Q _5750_/A4 _5900_/A3 _5750_/A3 _3819_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_82_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5530_ _5393_/Z _5530_/A2 _5530_/A3 _5530_/A4 _5531_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5461_ _5461_/A1 _5421_/C _5461_/A3 _5461_/A4 _5463_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4412_ hold363/Z hold636/Z _4413_/S _4412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7200_ _7200_/D _7243_/RN _7200_/CLK _7200_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5392_ _5395_/A1 _5392_/A2 _5529_/A1 _5525_/A1 _5392_/C _5394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_99_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4343_ hold59/Z hold65/Z _4346_/S hold66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7131_ _7131_/D _7243_/RN _7131_/CLK _7131_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4274_ _4273_/Z hold875/Z _4286_/S _4274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7062_ _7062_/D _7286_/RN _7062_/CLK _7062_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_140_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ _6805_/Q _6806_/Q _6807_/Q _6014_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6915_ _6915_/D _7359_/RN _6915_/CLK _6915_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6846_ hold5/Z _7300_/RN _6846_/CLK hold4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _6777_/D _7359_/RN _6777_/CLK _6777_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3989_ _6901_/Q _4408_/A1 _6677_/A2 _4030_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5728_ hold59/Z hold207/Z _5731_/S _5728_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ hold2/Z _7033_/Q hold8/Z hold9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold350 _7239_/Q hold350/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7329_ _7329_/D _7331_/CLK _7329_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold361 _4202_/Z _6743_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold383 _7255_/Q hold383/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold372 _5766_/Z _7128_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold394 _6949_/Q hold394/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_86_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _5441_/A4 _4961_/A2 _4961_/A3 _4927_/Z _5142_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_92_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _7286_/RN _7012_/Q _4069_/C _6700_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4892_ _4892_/A1 _4892_/A2 _5361_/A2 _4898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3912_ _7099_/Q _4006_/B1 _4008_/A2 _7091_/Q _3912_/C _3915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6631_ _6673_/A2 _6673_/A3 _6632_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3843_ _7190_/Q _3930_/A2 _3919_/B1 _6746_/Q _3845_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6562_ _6613_/A2 _6562_/A2 _6562_/A3 _6561_/Z _6563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3774_ _7062_/Q _4009_/A2 _4008_/A2 _7094_/Q _3776_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5513_ _5514_/A1 _5514_/A2 _5514_/A3 _5514_/A4 _5536_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6493_ _6493_/A1 _6493_/A2 _6493_/A3 _6493_/A4 _6493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_173_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5444_ _5444_/A1 _5246_/Z _5378_/Z _5444_/A4 _5488_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_172_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7114_ _7114_/D _7315_/RN _7114_/CLK _7114_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5375_ _5375_/A1 _5375_/A2 _5375_/A3 _5523_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4326_ hold79/Z hold297/Z _4328_/S _6828_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7045_ _7045_/D _7286_/RN _7045_/CLK _7045_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4257_ _5550_/A1 _5780_/A3 _5891_/A2 _6677_/A3 _4259_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_47_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4188_ hold49/Z _7337_/Q _6881_/Q hold50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_101_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6829_ _6829_/D _7359_/RN _6829_/CLK _6829_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold180 _6980_/Q hold180/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold191 _5868_/Z _7216_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3490_ hold98/I _7346_/Q _3491_/S _7347_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet679_341 net679_347/I _6946_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet679_330 net679_330/I _6957_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _5172_/A1 _5451_/B _5161_/B _5405_/A1 _5160_/C _5164_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5091_ _5382_/B1 _5382_/C _5091_/B1 _5259_/B _5091_/C _5442_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_96_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4111_ _6796_/Q _4110_/Z _6796_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ _6760_/Q _4042_/A2 _4042_/B1 _7138_/Q _4044_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5993_ _7295_/Q _7294_/Q _6594_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_92_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4944_ _5473_/A1 _5326_/C _5087_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_178_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _5417_/C _5294_/C _5199_/A3 _5416_/B _4876_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6614_ _5951_/B _7321_/Q _6614_/B _6615_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3826_ _7174_/Q _5891_/A4 _5891_/A3 _6677_/A1 _3834_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3757_ _7224_/Q _3914_/A2 _3981_/A2 _7152_/Q _3761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6545_ _7041_/Q _6312_/Z _6337_/Z _7073_/Q _6547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6476_ _6472_/Z _6476_/A2 _6476_/A3 _6476_/A4 _6483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3688_ _3688_/A1 _3688_/A2 _3688_/A3 _3688_/A4 _3702_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput230 _7394_/Z mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5427_ _5427_/A1 _5470_/A4 _5319_/C _5430_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput241 _7376_/Z mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput252 _4156_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5358_ _5358_/A1 _5360_/A2 _5360_/A3 _5358_/A4 _5526_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_160_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput285 _6734_/Q pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput274 _6740_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput263 _6941_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4309_ _4308_/Z hold872/Z _4321_/S _4309_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput296 _6737_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_48_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5289_ _5285_/Z _5364_/A1 _5494_/A2 _5265_/Z _5290_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7028_ _7028_/D _7300_/RN _7028_/CLK _7028_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_87_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18__1403_ clkbuf_4_10_0__1403_/Z net429_59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet629_271 net629_271/I _7016_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_260 net729_396/I _7027_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_293 net429_63/I _6994_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet629_282 net629_284/I _7005_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4660_ _5214_/A4 _5460_/A1 _4751_/B _3402_/I _5238_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_175_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ _3906_/A1 _3830_/C _3509_/Z _5808_/A3 _4045_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_162_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _7294_/Q _7297_/Q _6540_/A4 _6387_/A2 _6330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4591_ _4603_/A1 _4603_/A2 _5060_/C _4591_/C _5445_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_183_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3542_ _6881_/Q hold115/Z hold68/Z _3542_/C _3561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xhold905 _6809_/Q hold905/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_50_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ _6909_/Q _6290_/A2 _6292_/A2 _6861_/Q _6262_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3473_ _3468_/S _3470_/S _3473_/A3 _3473_/A4 _3482_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_170_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ _5421_/A2 _5406_/A1 _5218_/B _5213_/B _5424_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6192_ _6192_/A1 _6192_/A2 _6192_/A3 _6192_/A4 _6192_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5143_ _5324_/A3 _5473_/B _5344_/B _5338_/A2 _5450_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_124_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5074_ _5241_/B2 _5241_/B1 _5074_/B _5074_/C _5079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4025_ _4025_/A1 _4025_/A2 _4025_/A3 _4025_/A4 _4035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _7291_/Q _6299_/B _5976_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _4482_/Z _4483_/B _4927_/S _4927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ _5416_/C _5460_/A3 _5313_/A1 _4691_/C _5300_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_60_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3809_ _3809_/A1 _3809_/A2 _3809_/A3 _3809_/A4 _3809_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4789_ _4787_/B _5030_/A2 _4789_/B _5473_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_119_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ _7186_/Q _6320_/Z _6610_/B1 _7274_/Q _6530_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6459_ _5951_/B _7315_/Q _4083_/B _6806_/Q _6460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_125_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5__1403_ clkbuf_4_2_0__1403_/Z net729_367/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet429_54 net429_54/I _7233_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet429_76 net429_76/I _7211_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet429_65 _4150__5/I _7222_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet429_87 net429_87/I _7200_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet429_98 net429_98/I _7189_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ hold99/Z hold567/Z _5835_/S _5830_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ hold323/Z hold743/Z _5767_/S _5761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4712_ _4792_/B _5305_/B _4960_/A1 _4730_/A2 _4718_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_64__1403_ net629_288/I net629_264/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5692_ hold59/Z hold484/Z _5695_/S _5692_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4643_ _4643_/A1 _4643_/A2 _4643_/A3 _4649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4574_ _5322_/A2 _4751_/B _5162_/A2 _3399_/I _5413_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_128_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _7362_/D _6714_/Z _4152_/I1 _7362_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold702 _4253_/Z _6781_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6313_ _7297_/Q _6593_/A3 _6594_/A3 _6328_/A4 _6313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_7293_ _7293_/D _7322_/RN _7322_/CLK _7293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3525_ _3523_/B _3521_/Z _3906_/A1 _3548_/B _4435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold713 _7075_/Q hold713/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold724 _7026_/Q hold724/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold746 _7050_/Q hold746/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold735 _7091_/Q hold735/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold768 _6986_/Q hold768/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold757 hold757/I _7159_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6244_ _6240_/Z _6244_/A2 _6244_/A3 _6244_/A4 _6248_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold779 _5724_/Z _7090_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3456_ _4058_/A2 _6796_/Q _4095_/B _3456_/B _7363_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xnet829_466 _4150__25/I _6761_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_455 net829_455/I _6772_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ _7217_/Q _6290_/A2 _6290_/B1 hold72/I _6183_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet829_488 net829_499/I _6739_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet829_477 net829_482/I _6750_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3387_ _7005_/Q _3387_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5126_ _5440_/A2 _5284_/A2 _5534_/B1 _5309_/B _5128_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet829_499 net829_499/I _6728_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ _5228_/B _5421_/A2 _5183_/A2 _5510_/A2 _5058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4008_ _7090_/Q _4008_/A2 _4008_/B _4008_/C _4013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5959_ _5954_/B _5959_/A2 _5959_/B _5960_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold40 hold40/I hold40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold62 hold62/I hold62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold73 hold73/I hold73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold51 hold51/I hold51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_90_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold84 hold84/I hold84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_63_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold95 hold95/I hold95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_189_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4290_ hold905/Z _4289_/Z _4304_/S _4290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6931_ _6931_/D _6689_/Z _7364_/CLK _6931_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_54_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6862_ _6862_/D _7359_/RN _6862_/CLK _6862_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5813_ _5817_/S _5813_/A2 _5813_/B hold570/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6793_ _6793_/D _6684_/Z _7364_/CLK _6793_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5744_ hold99/Z hold313/Z _5749_/S _5744_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5675_ hold50/Z hold391/Z _5677_/S _5675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4626_ _5377_/B _5460_/A1 _5214_/A4 _4454_/Z _4630_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7345_ _7345_/D _6699_/Z _7364_/CLK _7345_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold510 _6907_/Q hold510/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold521 _7238_/Q hold521/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold554 _5921_/Z _7262_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4557_ _4702_/B _5305_/B _4694_/B _4787_/B _5228_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold543 _5690_/Z _7060_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold532 _4246_/Z _6776_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4488_ _4483_/B _4523_/A2 _4488_/B _4716_/B _5384_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xhold576 hold576/I _7223_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7276_ _7276_/D _7315_/RN _7276_/CLK _7276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_103_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3508_ _4178_/S hold21/Z _3508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold587 _4406_/Z _6899_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold565 _5542_/Z _6938_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_106_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3439_ _7366_/Q _7365_/Q _7367_/Q _3440_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6227_ _6767_/Q _6292_/A2 _6292_/B1 hold44/I _6230_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold598 _6840_/Q hold598/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6158_ _7086_/Q _6289_/A2 _6291_/C1 _6998_/Q _6293_/B1 _7062_/Q _6160_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _5109_/A1 _5354_/A1 _5111_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6089_ _6806_/Q _6089_/A2 _6090_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput130 wb_dat_i[11] _6649_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput152 wb_dat_i[31] _6665_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput141 wb_dat_i[21] _6658_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput163 wb_sel_i[2] _6673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3790_ _7085_/Q hold18/I hold22/I _4423_/A2 _3809_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ _5460_/A1 _5460_/A2 _5460_/A3 _5217_/B _5506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_75_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _5891_/A1 _4411_/A2 _5557_/A2 hold83/Z _4413_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5391_ _5473_/A1 _5473_/A2 _5391_/B _5392_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7130_ _7130_/D _7243_/RN _7130_/CLK _7130_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4342_ hold79/Z hold109/Z _4346_/S _4342_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4273_ hold626/Z hold323/Z _4285_/S _4273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7061_ _7061_/D _7315_/RN _7061_/CLK _7061_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _6017_/A2 _6012_/A2 _6014_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

