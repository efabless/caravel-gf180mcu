VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_defaults_block
  CLASS BLOCK ;
  FOREIGN gpio_defaults_block ;
  ORIGIN 0.430 0.430 ;
  SIZE 19.900 BY 16.540 ;
  PIN gpio_defaults[0]
    PORT
      LAYER Metal2 ;
        RECT 3.500 -0.420 3.780 1.235 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[4]
    PORT
      LAYER Metal2 ;
        RECT 10.220 -0.420 10.500 1.235 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[8]
    PORT
      LAYER Metal2 ;
        RECT 16.940 -0.420 17.220 1.235 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[7]
    PORT
      LAYER Metal2 ;
        RECT 15.260 -0.420 15.540 0.605 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[1]
    PORT
      LAYER Metal2 ;
        RECT 5.180 -0.420 5.460 0.485 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[5]
    PORT
      LAYER Metal2 ;
        RECT 11.900 -0.420 12.180 0.590 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[9]
    PORT
      LAYER Metal2 ;
        RECT 18.620 -0.420 18.900 6.285 ;
    END
  END gpio_defaults[9]
  PIN gpio_defaults[3]
    PORT
      LAYER Metal2 ;
        RECT 8.540 -0.420 8.820 2.200 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[2]
    PORT
      LAYER Metal2 ;
        RECT 6.860 -0.420 7.140 9.075 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[6]
    PORT
      LAYER Metal2 ;
        RECT 13.580 -0.420 13.860 9.075 ;
    END
  END gpio_defaults[6]
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 8.865 -0.265 11.895 15.960 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.330 -0.265 3.360 15.960 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0 0 19.900 16.540 ;
      LAYER Metal2 ;
        RECT 0 0 19.900 16.540 ;
      LAYER Metal3 ;
        RECT 0 0 19.900 16.540 ;
  END
END gpio_defaults_block
END LIBRARY

