magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< error_p >>
rect -160 509 -149 555
rect 54 509 65 555
<< nwell >>
rect -480 -786 480 786
<< mvpmos >>
rect -162 -524 -52 476
rect 52 -524 162 476
<< mvpdiff >>
rect -250 463 -162 476
rect -250 -511 -237 463
rect -191 -511 -162 463
rect -250 -524 -162 -511
rect -52 463 52 476
rect -52 -511 -23 463
rect 23 -511 52 463
rect -52 -524 52 -511
rect 162 463 250 476
rect 162 -511 191 463
rect 237 -511 250 463
rect 162 -524 250 -511
<< mvpdiffc >>
rect -237 -511 -191 463
rect -23 -511 23 463
rect 191 -511 237 463
<< mvnsubdiff >>
rect -394 628 394 700
rect -394 584 -322 628
rect -394 -584 -381 584
rect -335 -584 -322 584
rect 322 584 394 628
rect -394 -628 -322 -584
rect 322 -584 335 584
rect 381 -584 394 584
rect 322 -628 394 -584
rect -394 -641 394 -628
rect -394 -687 -278 -641
rect 278 -687 394 -641
rect -394 -700 394 -687
<< mvnsubdiffcont >>
rect -381 -584 -335 584
rect 335 -584 381 584
rect -278 -687 278 -641
<< polysilicon >>
rect -162 555 -52 568
rect -162 509 -149 555
rect -65 509 -52 555
rect -162 476 -52 509
rect 52 555 162 568
rect 52 509 65 555
rect 149 509 162 555
rect 52 476 162 509
rect -162 -568 -52 -524
rect 52 -568 162 -524
<< polycontact >>
rect -149 509 -65 555
rect 65 509 149 555
<< metal1 >>
rect -381 641 381 687
rect -381 584 -335 641
rect 335 584 381 641
rect -160 509 -149 555
rect -65 509 -54 555
rect 54 509 65 555
rect 149 509 160 555
rect -237 463 -191 474
rect -237 -522 -191 -511
rect -23 463 23 474
rect -23 -522 23 -511
rect 191 463 237 474
rect 191 -522 237 -511
rect -381 -641 -335 -584
rect 335 -641 381 -584
rect -381 -687 -278 -641
rect 278 -687 381 -641
<< properties >>
string FIXED_BBOX -348 -664 348 664
string gencell pmos_6p0
string library gf180mcu
string parameters w 5.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
