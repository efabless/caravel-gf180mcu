magic
tech gf180mcuC
magscale 1 10
timestamp 1669064184
<< metal1 >>
rect 6626 11230 6638 11282
rect 6690 11279 6702 11282
rect 7298 11279 7310 11282
rect 6690 11233 7310 11279
rect 6690 11230 6702 11233
rect 7298 11230 7310 11233
rect 7362 11230 7374 11282
rect 9090 11118 9102 11170
rect 9154 11167 9166 11170
rect 10546 11167 10558 11170
rect 9154 11121 10558 11167
rect 9154 11118 9166 11121
rect 10546 11118 10558 11121
rect 10610 11167 10622 11170
rect 11554 11167 11566 11170
rect 10610 11121 11566 11167
rect 10610 11118 10622 11121
rect 11554 11118 11566 11121
rect 11618 11118 11630 11170
rect 13346 11118 13358 11170
rect 13410 11167 13422 11170
rect 14466 11167 14478 11170
rect 13410 11121 14478 11167
rect 13410 11118 13422 11121
rect 14466 11118 14478 11121
rect 14530 11118 14542 11170
rect 224 11002 16848 11036
rect 224 10950 4210 11002
rect 4262 10950 4314 11002
rect 4366 10950 4418 11002
rect 4470 10950 8326 11002
rect 8378 10950 8430 11002
rect 8482 10950 8534 11002
rect 8586 10950 12442 11002
rect 12494 10950 12546 11002
rect 12598 10950 12650 11002
rect 12702 10950 16558 11002
rect 16610 10950 16662 11002
rect 16714 10950 16766 11002
rect 16818 10950 16848 11002
rect 224 10916 16848 10950
rect 11566 10834 11618 10846
rect 11566 10770 11618 10782
rect 12574 10834 12626 10846
rect 12574 10770 12626 10782
rect 2706 10558 2718 10610
rect 2770 10558 2782 10610
rect 7410 10558 7422 10610
rect 7474 10558 7486 10610
rect 10546 10558 10558 10610
rect 10610 10558 10622 10610
rect 13346 10558 13358 10610
rect 13410 10558 13422 10610
rect 3726 10498 3778 10510
rect 1026 10446 1038 10498
rect 1090 10446 1102 10498
rect 6626 10446 6638 10498
rect 6690 10446 6702 10498
rect 9090 10446 9102 10498
rect 9154 10446 9166 10498
rect 14242 10446 14254 10498
rect 14306 10446 14318 10498
rect 3726 10434 3778 10446
rect 224 10218 16688 10252
rect 224 10166 2152 10218
rect 2204 10166 2256 10218
rect 2308 10166 2360 10218
rect 2412 10166 6268 10218
rect 6320 10166 6372 10218
rect 6424 10166 6476 10218
rect 6528 10166 10384 10218
rect 10436 10166 10488 10218
rect 10540 10166 10592 10218
rect 10644 10166 14500 10218
rect 14552 10166 14604 10218
rect 14656 10166 14708 10218
rect 14760 10166 16688 10218
rect 224 10132 16688 10166
rect 16158 9938 16210 9950
rect 1922 9886 1934 9938
rect 1986 9886 1998 9938
rect 8194 9886 8206 9938
rect 8258 9886 8270 9938
rect 14130 9886 14142 9938
rect 14194 9886 14206 9938
rect 16158 9874 16210 9886
rect 12574 9826 12626 9838
rect 2930 9774 2942 9826
rect 2994 9774 3006 9826
rect 9202 9774 9214 9826
rect 9266 9774 9278 9826
rect 13346 9774 13358 9826
rect 13410 9774 13422 9826
rect 12574 9762 12626 9774
rect 10222 9714 10274 9726
rect 10222 9650 10274 9662
rect 4510 9602 4562 9614
rect 4510 9538 4562 9550
rect 6638 9602 6690 9614
rect 6638 9538 6690 9550
rect 224 9434 16848 9468
rect 224 9382 4210 9434
rect 4262 9382 4314 9434
rect 4366 9382 4418 9434
rect 4470 9382 8326 9434
rect 8378 9382 8430 9434
rect 8482 9382 8534 9434
rect 8586 9382 12442 9434
rect 12494 9382 12546 9434
rect 12598 9382 12650 9434
rect 12702 9382 16558 9434
rect 16610 9382 16662 9434
rect 16714 9382 16766 9434
rect 16818 9382 16848 9434
rect 224 9348 16848 9382
rect 4734 9266 4786 9278
rect 4734 9202 4786 9214
rect 15598 9042 15650 9054
rect 3378 8990 3390 9042
rect 3442 8990 3454 9042
rect 5282 8990 5294 9042
rect 5346 8990 5358 9042
rect 8754 8990 8766 9042
rect 8818 8990 8830 9042
rect 14578 8990 14590 9042
rect 14642 8990 14654 9042
rect 15598 8978 15650 8990
rect 2482 8878 2494 8930
rect 2546 8878 2558 8930
rect 7634 8878 7646 8930
rect 7698 8878 7710 8930
rect 10098 8878 10110 8930
rect 10162 8878 10174 8930
rect 13570 8878 13582 8930
rect 13634 8878 13646 8930
rect 224 8650 16688 8684
rect 224 8598 2152 8650
rect 2204 8598 2256 8650
rect 2308 8598 2360 8650
rect 2412 8598 6268 8650
rect 6320 8598 6372 8650
rect 6424 8598 6476 8650
rect 6528 8598 10384 8650
rect 10436 8598 10488 8650
rect 10540 8598 10592 8650
rect 10644 8598 14500 8650
rect 14552 8598 14604 8650
rect 14656 8598 14708 8650
rect 14760 8598 16688 8650
rect 224 8564 16688 8598
rect 3490 8430 3502 8482
rect 3554 8479 3566 8482
rect 4050 8479 4062 8482
rect 3554 8433 4062 8479
rect 3554 8430 3566 8433
rect 4050 8430 4062 8433
rect 4114 8430 4126 8482
rect 4510 8370 4562 8382
rect 1362 8318 1374 8370
rect 1426 8318 1438 8370
rect 8642 8318 8654 8370
rect 8706 8318 8718 8370
rect 15026 8318 15038 8370
rect 15090 8318 15102 8370
rect 4510 8306 4562 8318
rect 3726 8258 3778 8270
rect 10670 8258 10722 8270
rect 2706 8206 2718 8258
rect 2770 8206 2782 8258
rect 9650 8206 9662 8258
rect 9714 8206 9726 8258
rect 16146 8206 16158 8258
rect 16210 8206 16222 8258
rect 3726 8194 3778 8206
rect 10670 8194 10722 8206
rect 224 7866 16848 7900
rect 224 7814 4210 7866
rect 4262 7814 4314 7866
rect 4366 7814 4418 7866
rect 4470 7814 8326 7866
rect 8378 7814 8430 7866
rect 8482 7814 8534 7866
rect 8586 7814 12442 7866
rect 12494 7814 12546 7866
rect 12598 7814 12650 7866
rect 12702 7814 16558 7866
rect 16610 7814 16662 7866
rect 16714 7814 16766 7866
rect 16818 7814 16848 7866
rect 224 7780 16848 7814
rect 3826 7422 3838 7474
rect 3890 7422 3902 7474
rect 15474 7422 15486 7474
rect 15538 7422 15550 7474
rect 4734 7362 4786 7374
rect 2818 7310 2830 7362
rect 2882 7310 2894 7362
rect 4734 7298 4786 7310
rect 5182 7362 5234 7374
rect 5182 7298 5234 7310
rect 8542 7362 8594 7374
rect 14354 7310 14366 7362
rect 14418 7310 14430 7362
rect 8542 7298 8594 7310
rect 224 7082 16688 7116
rect 224 7030 2152 7082
rect 2204 7030 2256 7082
rect 2308 7030 2360 7082
rect 2412 7030 6268 7082
rect 6320 7030 6372 7082
rect 6424 7030 6476 7082
rect 6528 7030 10384 7082
rect 10436 7030 10488 7082
rect 10540 7030 10592 7082
rect 10644 7030 14500 7082
rect 14552 7030 14604 7082
rect 14656 7030 14708 7082
rect 14760 7030 16688 7082
rect 224 6996 16688 7030
rect 914 6750 926 6802
rect 978 6750 990 6802
rect 9538 6750 9550 6802
rect 9602 6750 9614 6802
rect 15922 6750 15934 6802
rect 15986 6750 15998 6802
rect 11566 6690 11618 6702
rect 2706 6638 2718 6690
rect 2770 6638 2782 6690
rect 5394 6638 5406 6690
rect 5458 6638 5470 6690
rect 10770 6638 10782 6690
rect 10834 6638 10846 6690
rect 14130 6638 14142 6690
rect 14194 6638 14206 6690
rect 11566 6626 11618 6638
rect 3726 6578 3778 6590
rect 3726 6514 3778 6526
rect 4846 6578 4898 6590
rect 13134 6578 13186 6590
rect 7186 6526 7198 6578
rect 7250 6526 7262 6578
rect 4846 6514 4898 6526
rect 13134 6514 13186 6526
rect 224 6298 16848 6332
rect 224 6246 4210 6298
rect 4262 6246 4314 6298
rect 4366 6246 4418 6298
rect 4470 6246 8326 6298
rect 8378 6246 8430 6298
rect 8482 6246 8534 6298
rect 8586 6246 12442 6298
rect 12494 6246 12546 6298
rect 12598 6246 12650 6298
rect 12702 6246 16558 6298
rect 16610 6246 16662 6298
rect 16714 6246 16766 6298
rect 16818 6246 16848 6298
rect 224 6212 16848 6246
rect 15262 6130 15314 6142
rect 15262 6066 15314 6078
rect 4722 5854 4734 5906
rect 4786 5854 4798 5906
rect 7298 5854 7310 5906
rect 7362 5854 7374 5906
rect 11106 5854 11118 5906
rect 11170 5854 11182 5906
rect 14242 5854 14254 5906
rect 14306 5854 14318 5906
rect 8542 5794 8594 5806
rect 15822 5794 15874 5806
rect 3266 5742 3278 5794
rect 3330 5742 3342 5794
rect 6626 5742 6638 5794
rect 6690 5742 6702 5794
rect 9874 5742 9886 5794
rect 9938 5742 9950 5794
rect 13010 5742 13022 5794
rect 13074 5742 13086 5794
rect 8542 5730 8594 5742
rect 15822 5730 15874 5742
rect 15474 5630 15486 5682
rect 15538 5679 15550 5682
rect 15810 5679 15822 5682
rect 15538 5633 15822 5679
rect 15538 5630 15550 5633
rect 15810 5630 15822 5633
rect 15874 5630 15886 5682
rect 224 5514 16688 5548
rect 224 5462 2152 5514
rect 2204 5462 2256 5514
rect 2308 5462 2360 5514
rect 2412 5462 6268 5514
rect 6320 5462 6372 5514
rect 6424 5462 6476 5514
rect 6528 5462 10384 5514
rect 10436 5462 10488 5514
rect 10540 5462 10592 5514
rect 10644 5462 14500 5514
rect 14552 5462 14604 5514
rect 14656 5462 14708 5514
rect 14760 5462 16688 5514
rect 224 5428 16688 5462
rect 12462 5234 12514 5246
rect 5730 5182 5742 5234
rect 5794 5182 5806 5234
rect 10210 5182 10222 5234
rect 10274 5182 10286 5234
rect 12462 5170 12514 5182
rect 12910 5234 12962 5246
rect 15026 5182 15038 5234
rect 15090 5182 15102 5234
rect 12910 5170 12962 5182
rect 3950 5122 4002 5134
rect 4610 5070 4622 5122
rect 4674 5070 4686 5122
rect 11218 5070 11230 5122
rect 11282 5070 11294 5122
rect 15698 5070 15710 5122
rect 15762 5070 15774 5122
rect 3950 5058 4002 5070
rect 224 4730 16848 4764
rect 224 4678 4210 4730
rect 4262 4678 4314 4730
rect 4366 4678 4418 4730
rect 4470 4678 8326 4730
rect 8378 4678 8430 4730
rect 8482 4678 8534 4730
rect 8586 4678 12442 4730
rect 12494 4678 12546 4730
rect 12598 4678 12650 4730
rect 12702 4678 16558 4730
rect 16610 4678 16662 4730
rect 16714 4678 16766 4730
rect 16818 4678 16848 4730
rect 224 4644 16848 4678
rect 15822 4562 15874 4574
rect 15822 4498 15874 4510
rect 7870 4338 7922 4350
rect 4274 4286 4286 4338
rect 4338 4286 4350 4338
rect 6850 4286 6862 4338
rect 6914 4286 6926 4338
rect 13906 4286 13918 4338
rect 13970 4286 13982 4338
rect 7870 4274 7922 4286
rect 14926 4226 14978 4238
rect 3154 4174 3166 4226
rect 3218 4174 3230 4226
rect 5842 4174 5854 4226
rect 5906 4174 5918 4226
rect 12114 4174 12126 4226
rect 12178 4174 12190 4226
rect 14926 4162 14978 4174
rect 224 3946 16688 3980
rect 224 3894 2152 3946
rect 2204 3894 2256 3946
rect 2308 3894 2360 3946
rect 2412 3894 6268 3946
rect 6320 3894 6372 3946
rect 6424 3894 6476 3946
rect 6528 3894 10384 3946
rect 10436 3894 10488 3946
rect 10540 3894 10592 3946
rect 10644 3894 14500 3946
rect 14552 3894 14604 3946
rect 14656 3894 14708 3946
rect 14760 3894 16688 3946
rect 224 3860 16688 3894
rect 11778 3726 11790 3778
rect 11842 3775 11854 3778
rect 12002 3775 12014 3778
rect 11842 3729 12014 3775
rect 11842 3726 11854 3729
rect 12002 3726 12014 3729
rect 12066 3726 12078 3778
rect 4510 3666 4562 3678
rect 11790 3666 11842 3678
rect 9426 3614 9438 3666
rect 9490 3614 9502 3666
rect 12786 3614 12798 3666
rect 12850 3614 12862 3666
rect 4510 3602 4562 3614
rect 11790 3602 11842 3614
rect 6526 3554 6578 3566
rect 15598 3554 15650 3566
rect 7074 3502 7086 3554
rect 7138 3502 7150 3554
rect 14578 3502 14590 3554
rect 14642 3502 14654 3554
rect 6526 3490 6578 3502
rect 15598 3490 15650 3502
rect 3950 3442 4002 3454
rect 3950 3378 4002 3390
rect 4958 3330 5010 3342
rect 4958 3266 5010 3278
rect 224 3162 16848 3196
rect 224 3110 4210 3162
rect 4262 3110 4314 3162
rect 4366 3110 4418 3162
rect 4470 3110 8326 3162
rect 8378 3110 8430 3162
rect 8482 3110 8534 3162
rect 8586 3110 12442 3162
rect 12494 3110 12546 3162
rect 12598 3110 12650 3162
rect 12702 3110 16558 3162
rect 16610 3110 16662 3162
rect 16714 3110 16766 3162
rect 16818 3110 16848 3162
rect 224 3076 16848 3110
rect 4274 2718 4286 2770
rect 4338 2718 4350 2770
rect 7522 2718 7534 2770
rect 7586 2718 7598 2770
rect 12002 2718 12014 2770
rect 12066 2718 12078 2770
rect 13122 2718 13134 2770
rect 13186 2718 13198 2770
rect 8542 2658 8594 2670
rect 3602 2606 3614 2658
rect 3666 2606 3678 2658
rect 5954 2606 5966 2658
rect 6018 2606 6030 2658
rect 10882 2606 10894 2658
rect 10946 2606 10958 2658
rect 14242 2606 14254 2658
rect 14306 2606 14318 2658
rect 8542 2594 8594 2606
rect 224 2378 16688 2412
rect 224 2326 2152 2378
rect 2204 2326 2256 2378
rect 2308 2326 2360 2378
rect 2412 2326 6268 2378
rect 6320 2326 6372 2378
rect 6424 2326 6476 2378
rect 6528 2326 10384 2378
rect 10436 2326 10488 2378
rect 10540 2326 10592 2378
rect 10644 2326 14500 2378
rect 14552 2326 14604 2378
rect 14656 2326 14708 2378
rect 14760 2326 16688 2378
rect 224 2292 16688 2326
rect 11790 2098 11842 2110
rect 2706 2046 2718 2098
rect 2770 2046 2782 2098
rect 5506 2046 5518 2098
rect 5570 2046 5582 2098
rect 13682 2046 13694 2098
rect 13746 2046 13758 2098
rect 11790 2034 11842 2046
rect 11342 1986 11394 1998
rect 3826 1934 3838 1986
rect 3890 1934 3902 1986
rect 6738 1934 6750 1986
rect 6802 1934 6814 1986
rect 12450 1934 12462 1986
rect 12514 1934 12526 1986
rect 11342 1922 11394 1934
rect 7646 1874 7698 1886
rect 7646 1810 7698 1822
rect 224 1594 16848 1628
rect 224 1542 4210 1594
rect 4262 1542 4314 1594
rect 4366 1542 4418 1594
rect 4470 1542 8326 1594
rect 8378 1542 8430 1594
rect 8482 1542 8534 1594
rect 8586 1542 12442 1594
rect 12494 1542 12546 1594
rect 12598 1542 12650 1594
rect 12702 1542 16558 1594
rect 16610 1542 16662 1594
rect 16714 1542 16766 1594
rect 16818 1542 16848 1594
rect 224 1508 16848 1542
<< via1 >>
rect 6638 11230 6690 11282
rect 7310 11230 7362 11282
rect 9102 11118 9154 11170
rect 10558 11118 10610 11170
rect 11566 11118 11618 11170
rect 13358 11118 13410 11170
rect 14478 11118 14530 11170
rect 4210 10950 4262 11002
rect 4314 10950 4366 11002
rect 4418 10950 4470 11002
rect 8326 10950 8378 11002
rect 8430 10950 8482 11002
rect 8534 10950 8586 11002
rect 12442 10950 12494 11002
rect 12546 10950 12598 11002
rect 12650 10950 12702 11002
rect 16558 10950 16610 11002
rect 16662 10950 16714 11002
rect 16766 10950 16818 11002
rect 11566 10782 11618 10834
rect 12574 10782 12626 10834
rect 2718 10558 2770 10610
rect 7422 10558 7474 10610
rect 10558 10558 10610 10610
rect 13358 10558 13410 10610
rect 1038 10446 1090 10498
rect 3726 10446 3778 10498
rect 6638 10446 6690 10498
rect 9102 10446 9154 10498
rect 14254 10446 14306 10498
rect 2152 10166 2204 10218
rect 2256 10166 2308 10218
rect 2360 10166 2412 10218
rect 6268 10166 6320 10218
rect 6372 10166 6424 10218
rect 6476 10166 6528 10218
rect 10384 10166 10436 10218
rect 10488 10166 10540 10218
rect 10592 10166 10644 10218
rect 14500 10166 14552 10218
rect 14604 10166 14656 10218
rect 14708 10166 14760 10218
rect 1934 9886 1986 9938
rect 8206 9886 8258 9938
rect 14142 9886 14194 9938
rect 16158 9886 16210 9938
rect 2942 9774 2994 9826
rect 9214 9774 9266 9826
rect 12574 9774 12626 9826
rect 13358 9774 13410 9826
rect 10222 9662 10274 9714
rect 4510 9550 4562 9602
rect 6638 9550 6690 9602
rect 4210 9382 4262 9434
rect 4314 9382 4366 9434
rect 4418 9382 4470 9434
rect 8326 9382 8378 9434
rect 8430 9382 8482 9434
rect 8534 9382 8586 9434
rect 12442 9382 12494 9434
rect 12546 9382 12598 9434
rect 12650 9382 12702 9434
rect 16558 9382 16610 9434
rect 16662 9382 16714 9434
rect 16766 9382 16818 9434
rect 4734 9214 4786 9266
rect 3390 8990 3442 9042
rect 5294 8990 5346 9042
rect 8766 8990 8818 9042
rect 14590 8990 14642 9042
rect 15598 8990 15650 9042
rect 2494 8878 2546 8930
rect 7646 8878 7698 8930
rect 10110 8878 10162 8930
rect 13582 8878 13634 8930
rect 2152 8598 2204 8650
rect 2256 8598 2308 8650
rect 2360 8598 2412 8650
rect 6268 8598 6320 8650
rect 6372 8598 6424 8650
rect 6476 8598 6528 8650
rect 10384 8598 10436 8650
rect 10488 8598 10540 8650
rect 10592 8598 10644 8650
rect 14500 8598 14552 8650
rect 14604 8598 14656 8650
rect 14708 8598 14760 8650
rect 3502 8430 3554 8482
rect 4062 8430 4114 8482
rect 1374 8318 1426 8370
rect 4510 8318 4562 8370
rect 8654 8318 8706 8370
rect 15038 8318 15090 8370
rect 2718 8206 2770 8258
rect 3726 8206 3778 8258
rect 9662 8206 9714 8258
rect 10670 8206 10722 8258
rect 16158 8206 16210 8258
rect 4210 7814 4262 7866
rect 4314 7814 4366 7866
rect 4418 7814 4470 7866
rect 8326 7814 8378 7866
rect 8430 7814 8482 7866
rect 8534 7814 8586 7866
rect 12442 7814 12494 7866
rect 12546 7814 12598 7866
rect 12650 7814 12702 7866
rect 16558 7814 16610 7866
rect 16662 7814 16714 7866
rect 16766 7814 16818 7866
rect 3838 7422 3890 7474
rect 15486 7422 15538 7474
rect 2830 7310 2882 7362
rect 4734 7310 4786 7362
rect 5182 7310 5234 7362
rect 8542 7310 8594 7362
rect 14366 7310 14418 7362
rect 2152 7030 2204 7082
rect 2256 7030 2308 7082
rect 2360 7030 2412 7082
rect 6268 7030 6320 7082
rect 6372 7030 6424 7082
rect 6476 7030 6528 7082
rect 10384 7030 10436 7082
rect 10488 7030 10540 7082
rect 10592 7030 10644 7082
rect 14500 7030 14552 7082
rect 14604 7030 14656 7082
rect 14708 7030 14760 7082
rect 926 6750 978 6802
rect 9550 6750 9602 6802
rect 15934 6750 15986 6802
rect 2718 6638 2770 6690
rect 5406 6638 5458 6690
rect 10782 6638 10834 6690
rect 11566 6638 11618 6690
rect 14142 6638 14194 6690
rect 3726 6526 3778 6578
rect 4846 6526 4898 6578
rect 7198 6526 7250 6578
rect 13134 6526 13186 6578
rect 4210 6246 4262 6298
rect 4314 6246 4366 6298
rect 4418 6246 4470 6298
rect 8326 6246 8378 6298
rect 8430 6246 8482 6298
rect 8534 6246 8586 6298
rect 12442 6246 12494 6298
rect 12546 6246 12598 6298
rect 12650 6246 12702 6298
rect 16558 6246 16610 6298
rect 16662 6246 16714 6298
rect 16766 6246 16818 6298
rect 15262 6078 15314 6130
rect 4734 5854 4786 5906
rect 7310 5854 7362 5906
rect 11118 5854 11170 5906
rect 14254 5854 14306 5906
rect 3278 5742 3330 5794
rect 6638 5742 6690 5794
rect 8542 5742 8594 5794
rect 9886 5742 9938 5794
rect 13022 5742 13074 5794
rect 15822 5742 15874 5794
rect 15486 5630 15538 5682
rect 15822 5630 15874 5682
rect 2152 5462 2204 5514
rect 2256 5462 2308 5514
rect 2360 5462 2412 5514
rect 6268 5462 6320 5514
rect 6372 5462 6424 5514
rect 6476 5462 6528 5514
rect 10384 5462 10436 5514
rect 10488 5462 10540 5514
rect 10592 5462 10644 5514
rect 14500 5462 14552 5514
rect 14604 5462 14656 5514
rect 14708 5462 14760 5514
rect 5742 5182 5794 5234
rect 10222 5182 10274 5234
rect 12462 5182 12514 5234
rect 12910 5182 12962 5234
rect 15038 5182 15090 5234
rect 3950 5070 4002 5122
rect 4622 5070 4674 5122
rect 11230 5070 11282 5122
rect 15710 5070 15762 5122
rect 4210 4678 4262 4730
rect 4314 4678 4366 4730
rect 4418 4678 4470 4730
rect 8326 4678 8378 4730
rect 8430 4678 8482 4730
rect 8534 4678 8586 4730
rect 12442 4678 12494 4730
rect 12546 4678 12598 4730
rect 12650 4678 12702 4730
rect 16558 4678 16610 4730
rect 16662 4678 16714 4730
rect 16766 4678 16818 4730
rect 15822 4510 15874 4562
rect 4286 4286 4338 4338
rect 6862 4286 6914 4338
rect 7870 4286 7922 4338
rect 13918 4286 13970 4338
rect 3166 4174 3218 4226
rect 5854 4174 5906 4226
rect 12126 4174 12178 4226
rect 14926 4174 14978 4226
rect 2152 3894 2204 3946
rect 2256 3894 2308 3946
rect 2360 3894 2412 3946
rect 6268 3894 6320 3946
rect 6372 3894 6424 3946
rect 6476 3894 6528 3946
rect 10384 3894 10436 3946
rect 10488 3894 10540 3946
rect 10592 3894 10644 3946
rect 14500 3894 14552 3946
rect 14604 3894 14656 3946
rect 14708 3894 14760 3946
rect 11790 3726 11842 3778
rect 12014 3726 12066 3778
rect 4510 3614 4562 3666
rect 9438 3614 9490 3666
rect 11790 3614 11842 3666
rect 12798 3614 12850 3666
rect 6526 3502 6578 3554
rect 7086 3502 7138 3554
rect 14590 3502 14642 3554
rect 15598 3502 15650 3554
rect 3950 3390 4002 3442
rect 4958 3278 5010 3330
rect 4210 3110 4262 3162
rect 4314 3110 4366 3162
rect 4418 3110 4470 3162
rect 8326 3110 8378 3162
rect 8430 3110 8482 3162
rect 8534 3110 8586 3162
rect 12442 3110 12494 3162
rect 12546 3110 12598 3162
rect 12650 3110 12702 3162
rect 16558 3110 16610 3162
rect 16662 3110 16714 3162
rect 16766 3110 16818 3162
rect 4286 2718 4338 2770
rect 7534 2718 7586 2770
rect 12014 2718 12066 2770
rect 13134 2718 13186 2770
rect 3614 2606 3666 2658
rect 5966 2606 6018 2658
rect 8542 2606 8594 2658
rect 10894 2606 10946 2658
rect 14254 2606 14306 2658
rect 2152 2326 2204 2378
rect 2256 2326 2308 2378
rect 2360 2326 2412 2378
rect 6268 2326 6320 2378
rect 6372 2326 6424 2378
rect 6476 2326 6528 2378
rect 10384 2326 10436 2378
rect 10488 2326 10540 2378
rect 10592 2326 10644 2378
rect 14500 2326 14552 2378
rect 14604 2326 14656 2378
rect 14708 2326 14760 2378
rect 2718 2046 2770 2098
rect 5518 2046 5570 2098
rect 11790 2046 11842 2098
rect 13694 2046 13746 2098
rect 3838 1934 3890 1986
rect 6750 1934 6802 1986
rect 11342 1934 11394 1986
rect 12462 1934 12514 1986
rect 7646 1822 7698 1874
rect 4210 1542 4262 1594
rect 4314 1542 4366 1594
rect 4418 1542 4470 1594
rect 8326 1542 8378 1594
rect 8430 1542 8482 1594
rect 8534 1542 8586 1594
rect 12442 1542 12494 1594
rect 12546 1542 12598 1594
rect 12650 1542 12702 1594
rect 16558 1542 16610 1594
rect 16662 1542 16714 1594
rect 16766 1542 16818 1594
<< metal2 >>
rect 560 12200 672 13000
rect 1008 12200 1120 13000
rect 1456 12200 1568 13000
rect 1904 12200 2016 13000
rect 2352 12200 2464 13000
rect 2800 12200 2912 13000
rect 3248 12200 3360 13000
rect 3696 12200 3808 13000
rect 4144 12200 4256 13000
rect 4592 12200 4704 13000
rect 5040 12200 5152 13000
rect 5488 12200 5600 13000
rect 5936 12200 6048 13000
rect 6384 12200 6496 13000
rect 6832 12200 6944 13000
rect 7280 12200 7392 13000
rect 7728 12200 7840 13000
rect 8176 12200 8288 13000
rect 8624 12200 8736 13000
rect 9072 12200 9184 13000
rect 9520 12200 9632 13000
rect 9968 12200 10080 13000
rect 10416 12200 10528 13000
rect 10864 12200 10976 13000
rect 11312 12200 11424 13000
rect 11760 12200 11872 13000
rect 12208 12200 12320 13000
rect 12656 12200 12768 13000
rect 13104 12200 13216 13000
rect 13552 12200 13664 13000
rect 14000 12200 14112 13000
rect 14448 12200 14560 13000
rect 14896 12200 15008 13000
rect 15344 12200 15456 13000
rect 15792 12200 15904 13000
rect 16240 12200 16352 13000
rect 588 8428 644 12200
rect 1036 10498 1092 12200
rect 1484 10724 1540 12200
rect 1036 10446 1038 10498
rect 1090 10446 1092 10498
rect 1036 10434 1092 10446
rect 1372 10668 1540 10724
rect 588 8372 980 8428
rect 924 6802 980 8372
rect 1372 8370 1428 10668
rect 1932 9938 1988 12200
rect 2380 10612 2436 12200
rect 2716 10612 2772 10622
rect 2380 10556 2548 10612
rect 2150 10220 2414 10230
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2150 10154 2414 10164
rect 1932 9886 1934 9938
rect 1986 9886 1988 9938
rect 1932 9874 1988 9886
rect 1372 8318 1374 8370
rect 1426 8318 1428 8370
rect 1372 8306 1428 8318
rect 1932 9492 1988 9502
rect 924 6750 926 6802
rect 978 6750 980 6802
rect 924 6738 980 6750
rect 1484 8260 1540 8270
rect 588 5124 644 5134
rect 588 800 644 5068
rect 1036 4340 1092 4350
rect 1036 800 1092 4284
rect 1484 800 1540 8204
rect 1932 800 1988 9436
rect 2492 8930 2548 10556
rect 2492 8878 2494 8930
rect 2546 8878 2548 8930
rect 2492 8866 2548 8878
rect 2604 10610 2772 10612
rect 2604 10558 2718 10610
rect 2770 10558 2772 10610
rect 2604 10556 2772 10558
rect 2604 10500 2660 10556
rect 2716 10546 2772 10556
rect 2150 8652 2414 8662
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2150 8586 2414 8596
rect 2150 7084 2414 7094
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2150 7018 2414 7028
rect 2492 5572 2548 5582
rect 2150 5516 2414 5526
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2150 5450 2414 5460
rect 2150 3948 2414 3958
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2150 3882 2414 3892
rect 2150 2380 2414 2390
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2150 2314 2414 2324
rect 2492 2212 2548 5516
rect 2604 4340 2660 10444
rect 2716 8260 2772 8270
rect 2716 8166 2772 8204
rect 2828 7362 2884 12200
rect 2940 9826 2996 9838
rect 2940 9774 2942 9826
rect 2994 9774 2996 9826
rect 2940 9492 2996 9774
rect 2940 9426 2996 9436
rect 2828 7310 2830 7362
rect 2882 7310 2884 7362
rect 2828 7298 2884 7310
rect 2716 6690 2772 6702
rect 2716 6638 2718 6690
rect 2770 6638 2772 6690
rect 2716 6580 2772 6638
rect 2716 5124 2772 6524
rect 2716 5058 2772 5068
rect 2828 6692 2884 6702
rect 2604 4274 2660 4284
rect 2380 2156 2548 2212
rect 2716 3332 2772 3342
rect 2380 800 2436 2156
rect 2716 2098 2772 3276
rect 2716 2046 2718 2098
rect 2770 2046 2772 2098
rect 2716 2034 2772 2046
rect 2828 800 2884 6636
rect 3164 6132 3220 6142
rect 3164 4226 3220 6076
rect 3276 5794 3332 12200
rect 3724 10724 3780 12200
rect 4172 11172 4228 12200
rect 3612 10668 3780 10724
rect 3948 11116 4228 11172
rect 3276 5742 3278 5794
rect 3330 5742 3332 5794
rect 3276 5730 3332 5742
rect 3388 9042 3444 9054
rect 3388 8990 3390 9042
rect 3442 8990 3444 9042
rect 3388 8484 3444 8990
rect 3500 8484 3556 8494
rect 3388 8482 3556 8484
rect 3388 8430 3502 8482
rect 3554 8430 3556 8482
rect 3388 8428 3556 8430
rect 3388 5572 3444 8428
rect 3500 8418 3556 8428
rect 3388 5506 3444 5516
rect 3164 4174 3166 4226
rect 3218 4174 3220 4226
rect 3164 4162 3220 4174
rect 3276 5348 3332 5358
rect 3276 800 3332 5292
rect 3612 2658 3668 10668
rect 3724 10500 3780 10510
rect 3724 10406 3780 10444
rect 3948 8372 4004 11116
rect 4208 11004 4472 11014
rect 4264 10948 4312 11004
rect 4368 10948 4416 11004
rect 4208 10938 4472 10948
rect 4508 9604 4564 9642
rect 4508 9538 4564 9548
rect 4208 9436 4472 9446
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4208 9370 4472 9380
rect 4060 8484 4116 8494
rect 4060 8482 4564 8484
rect 4060 8430 4062 8482
rect 4114 8430 4564 8482
rect 4060 8428 4564 8430
rect 4060 8418 4116 8428
rect 3948 8306 4004 8316
rect 4508 8370 4564 8428
rect 4508 8318 4510 8370
rect 4562 8318 4564 8370
rect 4508 8306 4564 8318
rect 3724 8260 3780 8270
rect 3724 8166 3780 8204
rect 4208 7868 4472 7878
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4208 7802 4472 7812
rect 3836 7474 3892 7486
rect 3836 7422 3838 7474
rect 3890 7422 3892 7474
rect 3836 6692 3892 7422
rect 3836 6626 3892 6636
rect 3724 6580 3780 6590
rect 3724 6486 3780 6524
rect 4208 6300 4472 6310
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4208 6234 4472 6244
rect 4620 6132 4676 12200
rect 4732 10724 4788 10734
rect 4732 9266 4788 10668
rect 4732 9214 4734 9266
rect 4786 9214 4788 9266
rect 4732 9044 4788 9214
rect 4732 8978 4788 8988
rect 4732 7362 4788 7374
rect 4732 7310 4734 7362
rect 4786 7310 4788 7362
rect 4732 6692 4788 7310
rect 4732 6626 4788 6636
rect 4844 6580 4900 6590
rect 4844 6486 4900 6524
rect 4620 6066 4676 6076
rect 4732 5908 4788 5918
rect 4732 5348 4788 5852
rect 4732 5282 4788 5292
rect 3948 5124 4004 5134
rect 4620 5124 4676 5134
rect 3948 5122 4676 5124
rect 3948 5070 3950 5122
rect 4002 5070 4622 5122
rect 4674 5070 4676 5122
rect 3948 5068 4676 5070
rect 3948 5058 4004 5068
rect 3948 3444 4004 3482
rect 3948 3378 4004 3388
rect 4060 3108 4116 5068
rect 4620 5058 4676 5068
rect 4208 4732 4472 4742
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4208 4666 4472 4676
rect 4284 4338 4340 4350
rect 4284 4286 4286 4338
rect 4338 4286 4340 4338
rect 4284 3668 4340 4286
rect 4508 3668 4564 3678
rect 4284 3666 4564 3668
rect 4284 3614 4510 3666
rect 4562 3614 4564 3666
rect 4284 3612 4564 3614
rect 4508 3388 4564 3612
rect 4844 3556 4900 3566
rect 4732 3444 4788 3454
rect 4508 3332 4676 3388
rect 3612 2606 3614 2658
rect 3666 2606 3668 2658
rect 3612 2594 3668 2606
rect 3948 3052 4116 3108
rect 4208 3164 4472 3174
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4208 3098 4472 3108
rect 3724 2548 3780 2558
rect 3724 800 3780 2492
rect 3836 1988 3892 1998
rect 3836 1894 3892 1932
rect 3948 1428 4004 3052
rect 4284 2770 4340 2782
rect 4284 2718 4286 2770
rect 4338 2718 4340 2770
rect 4284 2548 4340 2718
rect 4284 2482 4340 2492
rect 4208 1596 4472 1606
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4208 1530 4472 1540
rect 3948 1372 4228 1428
rect 4172 800 4228 1372
rect 4620 800 4676 3332
rect 4732 1988 4788 3388
rect 4844 2212 4900 3500
rect 4956 3330 5012 3342
rect 4956 3278 4958 3330
rect 5010 3278 5012 3330
rect 4956 2548 5012 3278
rect 5068 3332 5124 12200
rect 5292 9044 5348 9054
rect 5292 8950 5348 8988
rect 5180 7362 5236 7374
rect 5180 7310 5182 7362
rect 5234 7310 5236 7362
rect 5180 5908 5236 7310
rect 5404 6690 5460 6702
rect 5404 6638 5406 6690
rect 5458 6638 5460 6690
rect 5404 6580 5460 6638
rect 5404 6514 5460 6524
rect 5180 5842 5236 5852
rect 5068 3266 5124 3276
rect 4956 2482 5012 2492
rect 4844 2146 4900 2156
rect 5516 2098 5572 12200
rect 5964 10724 6020 12200
rect 5852 10668 6020 10724
rect 5740 8372 5796 8382
rect 5740 5234 5796 8316
rect 5740 5182 5742 5234
rect 5794 5182 5796 5234
rect 5740 5170 5796 5182
rect 5852 4226 5908 10668
rect 6412 10388 6468 12200
rect 6636 11282 6692 11294
rect 6636 11230 6638 11282
rect 6690 11230 6692 11282
rect 6636 10498 6692 11230
rect 6636 10446 6638 10498
rect 6690 10446 6692 10498
rect 6636 10434 6692 10446
rect 5852 4174 5854 4226
rect 5906 4174 5908 4226
rect 5852 4162 5908 4174
rect 5964 10332 6468 10388
rect 5964 2658 6020 10332
rect 6266 10220 6530 10230
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6266 10154 6530 10164
rect 6636 9604 6692 9614
rect 6636 9510 6692 9548
rect 6266 8652 6530 8662
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6860 8596 6916 12200
rect 7308 11282 7364 12200
rect 7308 11230 7310 11282
rect 7362 11230 7364 11282
rect 7308 11218 7364 11230
rect 6266 8586 6530 8596
rect 6748 8540 6916 8596
rect 7420 10610 7476 10622
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 9604 7476 10558
rect 6748 8372 6804 8540
rect 6636 8316 6804 8372
rect 6266 7084 6530 7094
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6266 7018 6530 7028
rect 6636 5794 6692 8316
rect 7196 6578 7252 6590
rect 7196 6526 7198 6578
rect 7250 6526 7252 6578
rect 7196 6468 7252 6526
rect 7196 6402 7252 6412
rect 6636 5742 6638 5794
rect 6690 5742 6692 5794
rect 6636 5730 6692 5742
rect 7308 5906 7364 5918
rect 7308 5854 7310 5906
rect 7362 5854 7364 5906
rect 7308 5796 7364 5854
rect 6266 5516 6530 5526
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6266 5450 6530 5460
rect 5964 2606 5966 2658
rect 6018 2606 6020 2658
rect 5964 2594 6020 2606
rect 6076 4340 6132 4350
rect 6076 2436 6132 4284
rect 6860 4340 6916 4350
rect 6860 4246 6916 4284
rect 6266 3948 6530 3958
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6266 3882 6530 3892
rect 6524 3556 6580 3566
rect 6524 3462 6580 3500
rect 7084 3556 7140 3566
rect 7084 3462 7140 3500
rect 7308 3388 7364 5740
rect 5516 2046 5518 2098
rect 5570 2046 5572 2098
rect 5516 2034 5572 2046
rect 5964 2380 6132 2436
rect 6860 3332 7364 3388
rect 6266 2380 6530 2390
rect 4732 1922 4788 1932
rect 5068 1988 5124 1998
rect 5068 800 5124 1932
rect 5516 1876 5572 1886
rect 5516 800 5572 1820
rect 5964 800 6020 2380
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6266 2314 6530 2324
rect 6412 2212 6468 2222
rect 6412 800 6468 2156
rect 6748 1986 6804 1998
rect 6748 1934 6750 1986
rect 6802 1934 6804 1986
rect 6748 1876 6804 1934
rect 6748 1810 6804 1820
rect 6860 800 6916 3332
rect 7420 2548 7476 9548
rect 7644 8932 7700 8942
rect 7644 8838 7700 8876
rect 7756 8372 7812 12200
rect 8204 9938 8260 12200
rect 8324 11004 8588 11014
rect 8380 10948 8428 11004
rect 8484 10948 8532 11004
rect 8324 10938 8588 10948
rect 8204 9886 8206 9938
rect 8258 9886 8260 9938
rect 8204 9874 8260 9886
rect 7756 8306 7812 8316
rect 8204 9716 8260 9726
rect 7756 6692 7812 6702
rect 7308 2492 7476 2548
rect 7532 2770 7588 2782
rect 7532 2718 7534 2770
rect 7586 2718 7588 2770
rect 7532 2660 7588 2718
rect 7308 800 7364 2492
rect 7532 2212 7588 2604
rect 7532 2146 7588 2156
rect 7644 1876 7700 1886
rect 7644 1782 7700 1820
rect 7756 800 7812 6636
rect 7868 4340 7924 4350
rect 7868 4246 7924 4284
rect 8204 800 8260 9660
rect 8324 9436 8588 9446
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8324 9370 8588 9380
rect 8652 9268 8708 12200
rect 9100 11170 9156 12200
rect 9100 11118 9102 11170
rect 9154 11118 9156 11170
rect 9100 11106 9156 11118
rect 9100 10498 9156 10510
rect 9100 10446 9102 10498
rect 9154 10446 9156 10498
rect 8652 9212 8932 9268
rect 8764 9042 8820 9054
rect 8764 8990 8766 9042
rect 8818 8990 8820 9042
rect 8652 8370 8708 8382
rect 8652 8318 8654 8370
rect 8706 8318 8708 8370
rect 8324 7868 8588 7878
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8324 7802 8588 7812
rect 8540 7362 8596 7374
rect 8540 7310 8542 7362
rect 8594 7310 8596 7362
rect 8540 6692 8596 7310
rect 8540 6626 8596 6636
rect 8324 6300 8588 6310
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8324 6234 8588 6244
rect 8540 5796 8596 5806
rect 8540 5702 8596 5740
rect 8324 4732 8588 4742
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8324 4666 8588 4676
rect 8324 3164 8588 3174
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8324 3098 8588 3108
rect 8540 2660 8596 2670
rect 8540 2566 8596 2604
rect 8324 1596 8588 1606
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8324 1530 8588 1540
rect 8652 800 8708 8318
rect 8764 6692 8820 8990
rect 8876 8260 8932 9212
rect 8876 8194 8932 8204
rect 8764 6626 8820 6636
rect 9100 800 9156 10446
rect 9212 9826 9268 9838
rect 9212 9774 9214 9826
rect 9266 9774 9268 9826
rect 9212 9716 9268 9774
rect 9212 9650 9268 9660
rect 9548 7252 9604 12200
rect 9660 8260 9716 8270
rect 9660 8166 9716 8204
rect 9548 7186 9604 7196
rect 9548 6802 9604 6814
rect 9548 6750 9550 6802
rect 9602 6750 9604 6802
rect 9436 3668 9492 3678
rect 9436 3574 9492 3612
rect 9548 800 9604 6750
rect 9996 5908 10052 12200
rect 10444 10388 10500 12200
rect 10556 11170 10612 11182
rect 10556 11118 10558 11170
rect 10610 11118 10612 11170
rect 10556 10610 10612 11118
rect 10556 10558 10558 10610
rect 10610 10558 10612 10610
rect 10556 10546 10612 10558
rect 10444 10322 10500 10332
rect 10382 10220 10646 10230
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10382 10154 10646 10164
rect 10220 9716 10276 9726
rect 10220 9622 10276 9660
rect 10108 8930 10164 8942
rect 10108 8878 10110 8930
rect 10162 8878 10164 8930
rect 10108 8372 10164 8878
rect 10382 8652 10646 8662
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10382 8586 10646 8596
rect 10108 8306 10164 8316
rect 10668 8260 10724 8270
rect 10668 8166 10724 8204
rect 10780 7252 10836 7262
rect 10382 7084 10646 7094
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10382 7018 10646 7028
rect 10780 6690 10836 7196
rect 10892 6804 10948 12200
rect 10892 6738 10948 6748
rect 11228 10388 11284 10398
rect 10780 6638 10782 6690
rect 10834 6638 10836 6690
rect 10780 6626 10836 6638
rect 9996 5842 10052 5852
rect 11116 5908 11172 5918
rect 11116 5814 11172 5852
rect 9884 5794 9940 5806
rect 9884 5742 9886 5794
rect 9938 5742 9940 5794
rect 9884 2884 9940 5742
rect 10382 5516 10646 5526
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10382 5450 10646 5460
rect 10220 5234 10276 5246
rect 10220 5182 10222 5234
rect 10274 5182 10276 5234
rect 9884 2828 10052 2884
rect 9996 800 10052 2828
rect 10220 2212 10276 5182
rect 11228 5236 11284 10332
rect 11340 7812 11396 12200
rect 11564 11170 11620 11182
rect 11564 11118 11566 11170
rect 11618 11118 11620 11170
rect 11564 10834 11620 11118
rect 11788 10948 11844 12200
rect 11788 10892 11956 10948
rect 11564 10782 11566 10834
rect 11618 10782 11620 10834
rect 11564 10770 11620 10782
rect 11788 10724 11844 10734
rect 11788 8932 11844 10668
rect 11788 8866 11844 8876
rect 11340 7756 11732 7812
rect 11564 7252 11620 7262
rect 11564 6690 11620 7196
rect 11564 6638 11566 6690
rect 11618 6638 11620 6690
rect 11564 6626 11620 6638
rect 11228 5122 11284 5180
rect 11228 5070 11230 5122
rect 11282 5070 11284 5122
rect 11228 5058 11284 5070
rect 10382 3948 10646 3958
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10382 3882 10646 3892
rect 11452 3444 11508 3454
rect 10892 2658 10948 2670
rect 10892 2606 10894 2658
rect 10946 2606 10948 2658
rect 10382 2380 10646 2390
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10382 2314 10646 2324
rect 10220 2156 10500 2212
rect 10444 800 10500 2156
rect 10892 800 10948 2606
rect 11340 1988 11396 1998
rect 11340 1894 11396 1932
rect 11452 1316 11508 3388
rect 11676 2772 11732 7756
rect 11900 7028 11956 10892
rect 11900 6962 11956 6972
rect 11788 6804 11844 6814
rect 11788 3778 11844 6748
rect 12124 4228 12180 4238
rect 11788 3726 11790 3778
rect 11842 3726 11844 3778
rect 11788 3666 11844 3726
rect 11788 3614 11790 3666
rect 11842 3614 11844 3666
rect 11788 3602 11844 3614
rect 11900 4226 12180 4228
rect 11900 4174 12126 4226
rect 12178 4174 12180 4226
rect 11900 4172 12180 4174
rect 11676 2100 11732 2716
rect 11788 2100 11844 2110
rect 11676 2098 11844 2100
rect 11676 2046 11790 2098
rect 11842 2046 11844 2098
rect 11676 2044 11844 2046
rect 11788 2034 11844 2044
rect 11900 1540 11956 4172
rect 12124 4162 12180 4172
rect 12012 3778 12068 3790
rect 12012 3726 12014 3778
rect 12066 3726 12068 3778
rect 12012 2770 12068 3726
rect 12012 2718 12014 2770
rect 12066 2718 12068 2770
rect 12012 2706 12068 2718
rect 12124 3668 12180 3678
rect 12124 2212 12180 3612
rect 12236 2996 12292 12200
rect 12684 11172 12740 12200
rect 12684 11116 12852 11172
rect 12440 11004 12704 11014
rect 12496 10948 12544 11004
rect 12600 10948 12648 11004
rect 12440 10938 12704 10948
rect 12572 10836 12628 10846
rect 12572 10742 12628 10780
rect 12572 9828 12628 9838
rect 12572 9734 12628 9772
rect 12440 9436 12704 9446
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12440 9370 12704 9380
rect 12440 7868 12704 7878
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12440 7802 12704 7812
rect 12440 6300 12704 6310
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12440 6234 12704 6244
rect 12460 5908 12516 5918
rect 12460 5234 12516 5852
rect 12460 5182 12462 5234
rect 12514 5182 12516 5234
rect 12460 5170 12516 5182
rect 12440 4732 12704 4742
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12440 4666 12704 4676
rect 12796 3892 12852 11116
rect 13132 8148 13188 12200
rect 13580 11284 13636 12200
rect 13580 11228 13748 11284
rect 13356 11170 13412 11182
rect 13356 11118 13358 11170
rect 13410 11118 13412 11170
rect 13356 10836 13412 11118
rect 13356 10610 13412 10780
rect 13356 10558 13358 10610
rect 13410 10558 13412 10610
rect 13356 10546 13412 10558
rect 13356 9828 13412 9838
rect 13356 9734 13412 9772
rect 13692 9044 13748 11228
rect 14028 9828 14084 12200
rect 14476 11170 14532 12200
rect 14476 11118 14478 11170
rect 14530 11118 14532 11170
rect 14476 11106 14532 11118
rect 14252 10498 14308 10510
rect 14252 10446 14254 10498
rect 14306 10446 14308 10498
rect 14028 9762 14084 9772
rect 14140 9938 14196 9950
rect 14140 9886 14142 9938
rect 14194 9886 14196 9938
rect 13692 8978 13748 8988
rect 13580 8930 13636 8942
rect 13580 8878 13582 8930
rect 13634 8878 13636 8930
rect 13132 8092 13300 8148
rect 13132 6580 13188 6590
rect 13132 6486 13188 6524
rect 13244 5908 13300 8092
rect 13244 5842 13300 5852
rect 13020 5794 13076 5806
rect 13020 5742 13022 5794
rect 13074 5742 13076 5794
rect 12908 5236 12964 5246
rect 12908 5142 12964 5180
rect 12796 3836 12964 3892
rect 12796 3666 12852 3678
rect 12796 3614 12798 3666
rect 12850 3614 12852 3666
rect 12440 3164 12704 3174
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12440 3098 12704 3108
rect 12236 2940 12516 2996
rect 12124 2146 12180 2156
rect 11340 1260 11508 1316
rect 11788 1484 11956 1540
rect 12236 2100 12292 2110
rect 11340 800 11396 1260
rect 11788 800 11844 1484
rect 12236 800 12292 2044
rect 12460 1988 12516 2940
rect 12460 1856 12516 1932
rect 12440 1596 12704 1606
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12440 1530 12704 1540
rect 12796 1428 12852 3614
rect 12908 3556 12964 3836
rect 12908 3490 12964 3500
rect 13020 2548 13076 5742
rect 13132 2772 13188 2782
rect 13132 2678 13188 2716
rect 13020 2492 13188 2548
rect 12684 1372 12852 1428
rect 12684 800 12740 1372
rect 13132 800 13188 2492
rect 13580 800 13636 8878
rect 13916 7028 13972 7038
rect 13916 4338 13972 6972
rect 14140 6916 14196 9886
rect 13916 4286 13918 4338
rect 13970 4286 13972 4338
rect 13916 4228 13972 4286
rect 13916 4162 13972 4172
rect 14028 6860 14196 6916
rect 13692 2100 13748 2110
rect 13692 2006 13748 2044
rect 14028 800 14084 6860
rect 14140 6690 14196 6702
rect 14140 6638 14142 6690
rect 14194 6638 14196 6690
rect 14140 6580 14196 6638
rect 14140 6514 14196 6524
rect 14252 6244 14308 10446
rect 14498 10220 14762 10230
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14498 10154 14762 10164
rect 14924 9940 14980 12200
rect 14924 9874 14980 9884
rect 14588 9044 14644 9054
rect 14588 8950 14644 8988
rect 14498 8652 14762 8662
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14498 8586 14762 8596
rect 15372 8428 15428 12200
rect 15596 9044 15652 9054
rect 15596 8950 15652 8988
rect 15820 8428 15876 12200
rect 16156 9940 16212 9950
rect 15036 8372 15092 8382
rect 15372 8372 15540 8428
rect 15820 8372 15988 8428
rect 15036 8370 15204 8372
rect 15036 8318 15038 8370
rect 15090 8318 15204 8370
rect 15036 8316 15204 8318
rect 15036 8306 15092 8316
rect 14140 6188 14308 6244
rect 14364 7362 14420 7374
rect 14364 7310 14366 7362
rect 14418 7310 14420 7362
rect 14140 4900 14196 6188
rect 14252 5908 14308 5918
rect 14252 5814 14308 5852
rect 14364 5124 14420 7310
rect 14498 7084 14762 7094
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14498 7018 14762 7028
rect 14498 5516 14762 5526
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14498 5450 14762 5460
rect 14364 5058 14420 5068
rect 15036 5234 15092 5246
rect 15036 5182 15038 5234
rect 15090 5182 15092 5234
rect 14140 4844 14420 4900
rect 14252 3444 14308 3454
rect 14252 2658 14308 3388
rect 14252 2606 14254 2658
rect 14306 2606 14308 2658
rect 14252 2594 14308 2606
rect 14364 2212 14420 4844
rect 14924 4228 14980 4238
rect 14924 4134 14980 4172
rect 15036 4116 15092 5182
rect 15036 4050 15092 4060
rect 14498 3948 14762 3958
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 15148 3892 15204 8316
rect 15484 7474 15540 8372
rect 15484 7422 15486 7474
rect 15538 7422 15540 7474
rect 15260 6132 15316 6142
rect 15260 6038 15316 6076
rect 15484 5682 15540 7422
rect 15932 7028 15988 8372
rect 16156 8258 16212 9884
rect 16156 8206 16158 8258
rect 16210 8206 16212 8258
rect 16156 8194 16212 8206
rect 15484 5630 15486 5682
rect 15538 5630 15540 5682
rect 15484 5618 15540 5630
rect 15708 6972 15988 7028
rect 14498 3882 14762 3892
rect 14924 3836 15204 3892
rect 15372 5124 15428 5134
rect 14588 3556 14644 3566
rect 14588 3462 14644 3500
rect 14498 2380 14762 2390
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14498 2314 14762 2324
rect 14364 2156 14532 2212
rect 14476 800 14532 2156
rect 14924 800 14980 3836
rect 15372 800 15428 5068
rect 15708 5122 15764 6972
rect 15932 6802 15988 6814
rect 15932 6750 15934 6802
rect 15986 6750 15988 6802
rect 15820 5794 15876 5806
rect 15820 5742 15822 5794
rect 15874 5742 15876 5794
rect 15820 5682 15876 5742
rect 15820 5630 15822 5682
rect 15874 5630 15876 5682
rect 15820 5618 15876 5630
rect 15708 5070 15710 5122
rect 15762 5070 15764 5122
rect 15708 4564 15764 5070
rect 15820 4564 15876 4574
rect 15708 4562 15876 4564
rect 15708 4510 15822 4562
rect 15874 4510 15876 4562
rect 15708 4508 15876 4510
rect 15820 4498 15876 4508
rect 15820 4116 15876 4126
rect 15596 3556 15652 3566
rect 15596 3462 15652 3500
rect 15820 800 15876 4060
rect 15932 3444 15988 6750
rect 16044 6580 16100 6590
rect 16268 6580 16324 12200
rect 16556 11004 16820 11014
rect 16612 10948 16660 11004
rect 16716 10948 16764 11004
rect 16556 10938 16820 10948
rect 16556 9436 16820 9446
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16556 9370 16820 9380
rect 16556 7868 16820 7878
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16556 7802 16820 7812
rect 16100 6524 16324 6580
rect 16044 6514 16100 6524
rect 16556 6300 16820 6310
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16556 6234 16820 6244
rect 16556 4732 16820 4742
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16556 4666 16820 4676
rect 15932 3388 16324 3444
rect 16268 800 16324 3388
rect 16556 3164 16820 3174
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16556 3098 16820 3108
rect 16556 1596 16820 1606
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16556 1530 16820 1540
rect 560 0 672 800
rect 1008 0 1120 800
rect 1456 0 1568 800
rect 1904 0 2016 800
rect 2352 0 2464 800
rect 2800 0 2912 800
rect 3248 0 3360 800
rect 3696 0 3808 800
rect 4144 0 4256 800
rect 4592 0 4704 800
rect 5040 0 5152 800
rect 5488 0 5600 800
rect 5936 0 6048 800
rect 6384 0 6496 800
rect 6832 0 6944 800
rect 7280 0 7392 800
rect 7728 0 7840 800
rect 8176 0 8288 800
rect 8624 0 8736 800
rect 9072 0 9184 800
rect 9520 0 9632 800
rect 9968 0 10080 800
rect 10416 0 10528 800
rect 10864 0 10976 800
rect 11312 0 11424 800
rect 11760 0 11872 800
rect 12208 0 12320 800
rect 12656 0 12768 800
rect 13104 0 13216 800
rect 13552 0 13664 800
rect 14000 0 14112 800
rect 14448 0 14560 800
rect 14896 0 15008 800
rect 15344 0 15456 800
rect 15792 0 15904 800
rect 16240 0 16352 800
<< via2 >>
rect 2150 10218 2206 10220
rect 2150 10166 2152 10218
rect 2152 10166 2204 10218
rect 2204 10166 2206 10218
rect 2150 10164 2206 10166
rect 2254 10218 2310 10220
rect 2254 10166 2256 10218
rect 2256 10166 2308 10218
rect 2308 10166 2310 10218
rect 2254 10164 2310 10166
rect 2358 10218 2414 10220
rect 2358 10166 2360 10218
rect 2360 10166 2412 10218
rect 2412 10166 2414 10218
rect 2358 10164 2414 10166
rect 1932 9436 1988 9492
rect 1484 8204 1540 8260
rect 588 5068 644 5124
rect 1036 4284 1092 4340
rect 2604 10444 2660 10500
rect 2150 8650 2206 8652
rect 2150 8598 2152 8650
rect 2152 8598 2204 8650
rect 2204 8598 2206 8650
rect 2150 8596 2206 8598
rect 2254 8650 2310 8652
rect 2254 8598 2256 8650
rect 2256 8598 2308 8650
rect 2308 8598 2310 8650
rect 2254 8596 2310 8598
rect 2358 8650 2414 8652
rect 2358 8598 2360 8650
rect 2360 8598 2412 8650
rect 2412 8598 2414 8650
rect 2358 8596 2414 8598
rect 2150 7082 2206 7084
rect 2150 7030 2152 7082
rect 2152 7030 2204 7082
rect 2204 7030 2206 7082
rect 2150 7028 2206 7030
rect 2254 7082 2310 7084
rect 2254 7030 2256 7082
rect 2256 7030 2308 7082
rect 2308 7030 2310 7082
rect 2254 7028 2310 7030
rect 2358 7082 2414 7084
rect 2358 7030 2360 7082
rect 2360 7030 2412 7082
rect 2412 7030 2414 7082
rect 2358 7028 2414 7030
rect 2150 5514 2206 5516
rect 2150 5462 2152 5514
rect 2152 5462 2204 5514
rect 2204 5462 2206 5514
rect 2150 5460 2206 5462
rect 2254 5514 2310 5516
rect 2254 5462 2256 5514
rect 2256 5462 2308 5514
rect 2308 5462 2310 5514
rect 2254 5460 2310 5462
rect 2358 5514 2414 5516
rect 2358 5462 2360 5514
rect 2360 5462 2412 5514
rect 2412 5462 2414 5514
rect 2358 5460 2414 5462
rect 2492 5516 2548 5572
rect 2150 3946 2206 3948
rect 2150 3894 2152 3946
rect 2152 3894 2204 3946
rect 2204 3894 2206 3946
rect 2150 3892 2206 3894
rect 2254 3946 2310 3948
rect 2254 3894 2256 3946
rect 2256 3894 2308 3946
rect 2308 3894 2310 3946
rect 2254 3892 2310 3894
rect 2358 3946 2414 3948
rect 2358 3894 2360 3946
rect 2360 3894 2412 3946
rect 2412 3894 2414 3946
rect 2358 3892 2414 3894
rect 2150 2378 2206 2380
rect 2150 2326 2152 2378
rect 2152 2326 2204 2378
rect 2204 2326 2206 2378
rect 2150 2324 2206 2326
rect 2254 2378 2310 2380
rect 2254 2326 2256 2378
rect 2256 2326 2308 2378
rect 2308 2326 2310 2378
rect 2254 2324 2310 2326
rect 2358 2378 2414 2380
rect 2358 2326 2360 2378
rect 2360 2326 2412 2378
rect 2412 2326 2414 2378
rect 2358 2324 2414 2326
rect 2716 8258 2772 8260
rect 2716 8206 2718 8258
rect 2718 8206 2770 8258
rect 2770 8206 2772 8258
rect 2716 8204 2772 8206
rect 2940 9436 2996 9492
rect 2716 6524 2772 6580
rect 2716 5068 2772 5124
rect 2828 6636 2884 6692
rect 2604 4284 2660 4340
rect 2716 3276 2772 3332
rect 3164 6076 3220 6132
rect 3388 5516 3444 5572
rect 3276 5292 3332 5348
rect 3724 10498 3780 10500
rect 3724 10446 3726 10498
rect 3726 10446 3778 10498
rect 3778 10446 3780 10498
rect 3724 10444 3780 10446
rect 4208 11002 4264 11004
rect 4208 10950 4210 11002
rect 4210 10950 4262 11002
rect 4262 10950 4264 11002
rect 4208 10948 4264 10950
rect 4312 11002 4368 11004
rect 4312 10950 4314 11002
rect 4314 10950 4366 11002
rect 4366 10950 4368 11002
rect 4312 10948 4368 10950
rect 4416 11002 4472 11004
rect 4416 10950 4418 11002
rect 4418 10950 4470 11002
rect 4470 10950 4472 11002
rect 4416 10948 4472 10950
rect 4508 9602 4564 9604
rect 4508 9550 4510 9602
rect 4510 9550 4562 9602
rect 4562 9550 4564 9602
rect 4508 9548 4564 9550
rect 4208 9434 4264 9436
rect 4208 9382 4210 9434
rect 4210 9382 4262 9434
rect 4262 9382 4264 9434
rect 4208 9380 4264 9382
rect 4312 9434 4368 9436
rect 4312 9382 4314 9434
rect 4314 9382 4366 9434
rect 4366 9382 4368 9434
rect 4312 9380 4368 9382
rect 4416 9434 4472 9436
rect 4416 9382 4418 9434
rect 4418 9382 4470 9434
rect 4470 9382 4472 9434
rect 4416 9380 4472 9382
rect 3948 8316 4004 8372
rect 3724 8258 3780 8260
rect 3724 8206 3726 8258
rect 3726 8206 3778 8258
rect 3778 8206 3780 8258
rect 3724 8204 3780 8206
rect 4208 7866 4264 7868
rect 4208 7814 4210 7866
rect 4210 7814 4262 7866
rect 4262 7814 4264 7866
rect 4208 7812 4264 7814
rect 4312 7866 4368 7868
rect 4312 7814 4314 7866
rect 4314 7814 4366 7866
rect 4366 7814 4368 7866
rect 4312 7812 4368 7814
rect 4416 7866 4472 7868
rect 4416 7814 4418 7866
rect 4418 7814 4470 7866
rect 4470 7814 4472 7866
rect 4416 7812 4472 7814
rect 3836 6636 3892 6692
rect 3724 6578 3780 6580
rect 3724 6526 3726 6578
rect 3726 6526 3778 6578
rect 3778 6526 3780 6578
rect 3724 6524 3780 6526
rect 4208 6298 4264 6300
rect 4208 6246 4210 6298
rect 4210 6246 4262 6298
rect 4262 6246 4264 6298
rect 4208 6244 4264 6246
rect 4312 6298 4368 6300
rect 4312 6246 4314 6298
rect 4314 6246 4366 6298
rect 4366 6246 4368 6298
rect 4312 6244 4368 6246
rect 4416 6298 4472 6300
rect 4416 6246 4418 6298
rect 4418 6246 4470 6298
rect 4470 6246 4472 6298
rect 4416 6244 4472 6246
rect 4732 10668 4788 10724
rect 4732 8988 4788 9044
rect 4732 6636 4788 6692
rect 4844 6578 4900 6580
rect 4844 6526 4846 6578
rect 4846 6526 4898 6578
rect 4898 6526 4900 6578
rect 4844 6524 4900 6526
rect 4620 6076 4676 6132
rect 4732 5906 4788 5908
rect 4732 5854 4734 5906
rect 4734 5854 4786 5906
rect 4786 5854 4788 5906
rect 4732 5852 4788 5854
rect 4732 5292 4788 5348
rect 3948 3442 4004 3444
rect 3948 3390 3950 3442
rect 3950 3390 4002 3442
rect 4002 3390 4004 3442
rect 3948 3388 4004 3390
rect 4208 4730 4264 4732
rect 4208 4678 4210 4730
rect 4210 4678 4262 4730
rect 4262 4678 4264 4730
rect 4208 4676 4264 4678
rect 4312 4730 4368 4732
rect 4312 4678 4314 4730
rect 4314 4678 4366 4730
rect 4366 4678 4368 4730
rect 4312 4676 4368 4678
rect 4416 4730 4472 4732
rect 4416 4678 4418 4730
rect 4418 4678 4470 4730
rect 4470 4678 4472 4730
rect 4416 4676 4472 4678
rect 4844 3500 4900 3556
rect 4732 3388 4788 3444
rect 4208 3162 4264 3164
rect 4208 3110 4210 3162
rect 4210 3110 4262 3162
rect 4262 3110 4264 3162
rect 4208 3108 4264 3110
rect 4312 3162 4368 3164
rect 4312 3110 4314 3162
rect 4314 3110 4366 3162
rect 4366 3110 4368 3162
rect 4312 3108 4368 3110
rect 4416 3162 4472 3164
rect 4416 3110 4418 3162
rect 4418 3110 4470 3162
rect 4470 3110 4472 3162
rect 4416 3108 4472 3110
rect 3724 2492 3780 2548
rect 3836 1986 3892 1988
rect 3836 1934 3838 1986
rect 3838 1934 3890 1986
rect 3890 1934 3892 1986
rect 3836 1932 3892 1934
rect 4284 2492 4340 2548
rect 4208 1594 4264 1596
rect 4208 1542 4210 1594
rect 4210 1542 4262 1594
rect 4262 1542 4264 1594
rect 4208 1540 4264 1542
rect 4312 1594 4368 1596
rect 4312 1542 4314 1594
rect 4314 1542 4366 1594
rect 4366 1542 4368 1594
rect 4312 1540 4368 1542
rect 4416 1594 4472 1596
rect 4416 1542 4418 1594
rect 4418 1542 4470 1594
rect 4470 1542 4472 1594
rect 4416 1540 4472 1542
rect 5292 9042 5348 9044
rect 5292 8990 5294 9042
rect 5294 8990 5346 9042
rect 5346 8990 5348 9042
rect 5292 8988 5348 8990
rect 5404 6524 5460 6580
rect 5180 5852 5236 5908
rect 5068 3276 5124 3332
rect 4956 2492 5012 2548
rect 4844 2156 4900 2212
rect 5740 8316 5796 8372
rect 6266 10218 6322 10220
rect 6266 10166 6268 10218
rect 6268 10166 6320 10218
rect 6320 10166 6322 10218
rect 6266 10164 6322 10166
rect 6370 10218 6426 10220
rect 6370 10166 6372 10218
rect 6372 10166 6424 10218
rect 6424 10166 6426 10218
rect 6370 10164 6426 10166
rect 6474 10218 6530 10220
rect 6474 10166 6476 10218
rect 6476 10166 6528 10218
rect 6528 10166 6530 10218
rect 6474 10164 6530 10166
rect 6636 9602 6692 9604
rect 6636 9550 6638 9602
rect 6638 9550 6690 9602
rect 6690 9550 6692 9602
rect 6636 9548 6692 9550
rect 6266 8650 6322 8652
rect 6266 8598 6268 8650
rect 6268 8598 6320 8650
rect 6320 8598 6322 8650
rect 6266 8596 6322 8598
rect 6370 8650 6426 8652
rect 6370 8598 6372 8650
rect 6372 8598 6424 8650
rect 6424 8598 6426 8650
rect 6370 8596 6426 8598
rect 6474 8650 6530 8652
rect 6474 8598 6476 8650
rect 6476 8598 6528 8650
rect 6528 8598 6530 8650
rect 6474 8596 6530 8598
rect 7420 9548 7476 9604
rect 6266 7082 6322 7084
rect 6266 7030 6268 7082
rect 6268 7030 6320 7082
rect 6320 7030 6322 7082
rect 6266 7028 6322 7030
rect 6370 7082 6426 7084
rect 6370 7030 6372 7082
rect 6372 7030 6424 7082
rect 6424 7030 6426 7082
rect 6370 7028 6426 7030
rect 6474 7082 6530 7084
rect 6474 7030 6476 7082
rect 6476 7030 6528 7082
rect 6528 7030 6530 7082
rect 6474 7028 6530 7030
rect 7196 6412 7252 6468
rect 7308 5740 7364 5796
rect 6266 5514 6322 5516
rect 6266 5462 6268 5514
rect 6268 5462 6320 5514
rect 6320 5462 6322 5514
rect 6266 5460 6322 5462
rect 6370 5514 6426 5516
rect 6370 5462 6372 5514
rect 6372 5462 6424 5514
rect 6424 5462 6426 5514
rect 6370 5460 6426 5462
rect 6474 5514 6530 5516
rect 6474 5462 6476 5514
rect 6476 5462 6528 5514
rect 6528 5462 6530 5514
rect 6474 5460 6530 5462
rect 6076 4284 6132 4340
rect 6860 4338 6916 4340
rect 6860 4286 6862 4338
rect 6862 4286 6914 4338
rect 6914 4286 6916 4338
rect 6860 4284 6916 4286
rect 6266 3946 6322 3948
rect 6266 3894 6268 3946
rect 6268 3894 6320 3946
rect 6320 3894 6322 3946
rect 6266 3892 6322 3894
rect 6370 3946 6426 3948
rect 6370 3894 6372 3946
rect 6372 3894 6424 3946
rect 6424 3894 6426 3946
rect 6370 3892 6426 3894
rect 6474 3946 6530 3948
rect 6474 3894 6476 3946
rect 6476 3894 6528 3946
rect 6528 3894 6530 3946
rect 6474 3892 6530 3894
rect 6524 3554 6580 3556
rect 6524 3502 6526 3554
rect 6526 3502 6578 3554
rect 6578 3502 6580 3554
rect 6524 3500 6580 3502
rect 7084 3554 7140 3556
rect 7084 3502 7086 3554
rect 7086 3502 7138 3554
rect 7138 3502 7140 3554
rect 7084 3500 7140 3502
rect 4732 1932 4788 1988
rect 5068 1932 5124 1988
rect 5516 1820 5572 1876
rect 6266 2378 6322 2380
rect 6266 2326 6268 2378
rect 6268 2326 6320 2378
rect 6320 2326 6322 2378
rect 6266 2324 6322 2326
rect 6370 2378 6426 2380
rect 6370 2326 6372 2378
rect 6372 2326 6424 2378
rect 6424 2326 6426 2378
rect 6370 2324 6426 2326
rect 6474 2378 6530 2380
rect 6474 2326 6476 2378
rect 6476 2326 6528 2378
rect 6528 2326 6530 2378
rect 6474 2324 6530 2326
rect 6412 2156 6468 2212
rect 6748 1820 6804 1876
rect 7644 8930 7700 8932
rect 7644 8878 7646 8930
rect 7646 8878 7698 8930
rect 7698 8878 7700 8930
rect 7644 8876 7700 8878
rect 8324 11002 8380 11004
rect 8324 10950 8326 11002
rect 8326 10950 8378 11002
rect 8378 10950 8380 11002
rect 8324 10948 8380 10950
rect 8428 11002 8484 11004
rect 8428 10950 8430 11002
rect 8430 10950 8482 11002
rect 8482 10950 8484 11002
rect 8428 10948 8484 10950
rect 8532 11002 8588 11004
rect 8532 10950 8534 11002
rect 8534 10950 8586 11002
rect 8586 10950 8588 11002
rect 8532 10948 8588 10950
rect 7756 8316 7812 8372
rect 8204 9660 8260 9716
rect 7756 6636 7812 6692
rect 7532 2604 7588 2660
rect 7532 2156 7588 2212
rect 7644 1874 7700 1876
rect 7644 1822 7646 1874
rect 7646 1822 7698 1874
rect 7698 1822 7700 1874
rect 7644 1820 7700 1822
rect 7868 4338 7924 4340
rect 7868 4286 7870 4338
rect 7870 4286 7922 4338
rect 7922 4286 7924 4338
rect 7868 4284 7924 4286
rect 8324 9434 8380 9436
rect 8324 9382 8326 9434
rect 8326 9382 8378 9434
rect 8378 9382 8380 9434
rect 8324 9380 8380 9382
rect 8428 9434 8484 9436
rect 8428 9382 8430 9434
rect 8430 9382 8482 9434
rect 8482 9382 8484 9434
rect 8428 9380 8484 9382
rect 8532 9434 8588 9436
rect 8532 9382 8534 9434
rect 8534 9382 8586 9434
rect 8586 9382 8588 9434
rect 8532 9380 8588 9382
rect 8324 7866 8380 7868
rect 8324 7814 8326 7866
rect 8326 7814 8378 7866
rect 8378 7814 8380 7866
rect 8324 7812 8380 7814
rect 8428 7866 8484 7868
rect 8428 7814 8430 7866
rect 8430 7814 8482 7866
rect 8482 7814 8484 7866
rect 8428 7812 8484 7814
rect 8532 7866 8588 7868
rect 8532 7814 8534 7866
rect 8534 7814 8586 7866
rect 8586 7814 8588 7866
rect 8532 7812 8588 7814
rect 8540 6636 8596 6692
rect 8324 6298 8380 6300
rect 8324 6246 8326 6298
rect 8326 6246 8378 6298
rect 8378 6246 8380 6298
rect 8324 6244 8380 6246
rect 8428 6298 8484 6300
rect 8428 6246 8430 6298
rect 8430 6246 8482 6298
rect 8482 6246 8484 6298
rect 8428 6244 8484 6246
rect 8532 6298 8588 6300
rect 8532 6246 8534 6298
rect 8534 6246 8586 6298
rect 8586 6246 8588 6298
rect 8532 6244 8588 6246
rect 8540 5794 8596 5796
rect 8540 5742 8542 5794
rect 8542 5742 8594 5794
rect 8594 5742 8596 5794
rect 8540 5740 8596 5742
rect 8324 4730 8380 4732
rect 8324 4678 8326 4730
rect 8326 4678 8378 4730
rect 8378 4678 8380 4730
rect 8324 4676 8380 4678
rect 8428 4730 8484 4732
rect 8428 4678 8430 4730
rect 8430 4678 8482 4730
rect 8482 4678 8484 4730
rect 8428 4676 8484 4678
rect 8532 4730 8588 4732
rect 8532 4678 8534 4730
rect 8534 4678 8586 4730
rect 8586 4678 8588 4730
rect 8532 4676 8588 4678
rect 8324 3162 8380 3164
rect 8324 3110 8326 3162
rect 8326 3110 8378 3162
rect 8378 3110 8380 3162
rect 8324 3108 8380 3110
rect 8428 3162 8484 3164
rect 8428 3110 8430 3162
rect 8430 3110 8482 3162
rect 8482 3110 8484 3162
rect 8428 3108 8484 3110
rect 8532 3162 8588 3164
rect 8532 3110 8534 3162
rect 8534 3110 8586 3162
rect 8586 3110 8588 3162
rect 8532 3108 8588 3110
rect 8540 2658 8596 2660
rect 8540 2606 8542 2658
rect 8542 2606 8594 2658
rect 8594 2606 8596 2658
rect 8540 2604 8596 2606
rect 8324 1594 8380 1596
rect 8324 1542 8326 1594
rect 8326 1542 8378 1594
rect 8378 1542 8380 1594
rect 8324 1540 8380 1542
rect 8428 1594 8484 1596
rect 8428 1542 8430 1594
rect 8430 1542 8482 1594
rect 8482 1542 8484 1594
rect 8428 1540 8484 1542
rect 8532 1594 8588 1596
rect 8532 1542 8534 1594
rect 8534 1542 8586 1594
rect 8586 1542 8588 1594
rect 8532 1540 8588 1542
rect 8876 8204 8932 8260
rect 8764 6636 8820 6692
rect 9212 9660 9268 9716
rect 9660 8258 9716 8260
rect 9660 8206 9662 8258
rect 9662 8206 9714 8258
rect 9714 8206 9716 8258
rect 9660 8204 9716 8206
rect 9548 7196 9604 7252
rect 9436 3666 9492 3668
rect 9436 3614 9438 3666
rect 9438 3614 9490 3666
rect 9490 3614 9492 3666
rect 9436 3612 9492 3614
rect 10444 10332 10500 10388
rect 10382 10218 10438 10220
rect 10382 10166 10384 10218
rect 10384 10166 10436 10218
rect 10436 10166 10438 10218
rect 10382 10164 10438 10166
rect 10486 10218 10542 10220
rect 10486 10166 10488 10218
rect 10488 10166 10540 10218
rect 10540 10166 10542 10218
rect 10486 10164 10542 10166
rect 10590 10218 10646 10220
rect 10590 10166 10592 10218
rect 10592 10166 10644 10218
rect 10644 10166 10646 10218
rect 10590 10164 10646 10166
rect 10220 9714 10276 9716
rect 10220 9662 10222 9714
rect 10222 9662 10274 9714
rect 10274 9662 10276 9714
rect 10220 9660 10276 9662
rect 10382 8650 10438 8652
rect 10382 8598 10384 8650
rect 10384 8598 10436 8650
rect 10436 8598 10438 8650
rect 10382 8596 10438 8598
rect 10486 8650 10542 8652
rect 10486 8598 10488 8650
rect 10488 8598 10540 8650
rect 10540 8598 10542 8650
rect 10486 8596 10542 8598
rect 10590 8650 10646 8652
rect 10590 8598 10592 8650
rect 10592 8598 10644 8650
rect 10644 8598 10646 8650
rect 10590 8596 10646 8598
rect 10108 8316 10164 8372
rect 10668 8258 10724 8260
rect 10668 8206 10670 8258
rect 10670 8206 10722 8258
rect 10722 8206 10724 8258
rect 10668 8204 10724 8206
rect 10780 7196 10836 7252
rect 10382 7082 10438 7084
rect 10382 7030 10384 7082
rect 10384 7030 10436 7082
rect 10436 7030 10438 7082
rect 10382 7028 10438 7030
rect 10486 7082 10542 7084
rect 10486 7030 10488 7082
rect 10488 7030 10540 7082
rect 10540 7030 10542 7082
rect 10486 7028 10542 7030
rect 10590 7082 10646 7084
rect 10590 7030 10592 7082
rect 10592 7030 10644 7082
rect 10644 7030 10646 7082
rect 10590 7028 10646 7030
rect 10892 6748 10948 6804
rect 11228 10332 11284 10388
rect 9996 5852 10052 5908
rect 11116 5906 11172 5908
rect 11116 5854 11118 5906
rect 11118 5854 11170 5906
rect 11170 5854 11172 5906
rect 11116 5852 11172 5854
rect 10382 5514 10438 5516
rect 10382 5462 10384 5514
rect 10384 5462 10436 5514
rect 10436 5462 10438 5514
rect 10382 5460 10438 5462
rect 10486 5514 10542 5516
rect 10486 5462 10488 5514
rect 10488 5462 10540 5514
rect 10540 5462 10542 5514
rect 10486 5460 10542 5462
rect 10590 5514 10646 5516
rect 10590 5462 10592 5514
rect 10592 5462 10644 5514
rect 10644 5462 10646 5514
rect 10590 5460 10646 5462
rect 11788 10668 11844 10724
rect 11788 8876 11844 8932
rect 11564 7196 11620 7252
rect 11228 5180 11284 5236
rect 10382 3946 10438 3948
rect 10382 3894 10384 3946
rect 10384 3894 10436 3946
rect 10436 3894 10438 3946
rect 10382 3892 10438 3894
rect 10486 3946 10542 3948
rect 10486 3894 10488 3946
rect 10488 3894 10540 3946
rect 10540 3894 10542 3946
rect 10486 3892 10542 3894
rect 10590 3946 10646 3948
rect 10590 3894 10592 3946
rect 10592 3894 10644 3946
rect 10644 3894 10646 3946
rect 10590 3892 10646 3894
rect 11452 3388 11508 3444
rect 10382 2378 10438 2380
rect 10382 2326 10384 2378
rect 10384 2326 10436 2378
rect 10436 2326 10438 2378
rect 10382 2324 10438 2326
rect 10486 2378 10542 2380
rect 10486 2326 10488 2378
rect 10488 2326 10540 2378
rect 10540 2326 10542 2378
rect 10486 2324 10542 2326
rect 10590 2378 10646 2380
rect 10590 2326 10592 2378
rect 10592 2326 10644 2378
rect 10644 2326 10646 2378
rect 10590 2324 10646 2326
rect 11340 1986 11396 1988
rect 11340 1934 11342 1986
rect 11342 1934 11394 1986
rect 11394 1934 11396 1986
rect 11340 1932 11396 1934
rect 11900 6972 11956 7028
rect 11788 6748 11844 6804
rect 11676 2716 11732 2772
rect 12124 3612 12180 3668
rect 12440 11002 12496 11004
rect 12440 10950 12442 11002
rect 12442 10950 12494 11002
rect 12494 10950 12496 11002
rect 12440 10948 12496 10950
rect 12544 11002 12600 11004
rect 12544 10950 12546 11002
rect 12546 10950 12598 11002
rect 12598 10950 12600 11002
rect 12544 10948 12600 10950
rect 12648 11002 12704 11004
rect 12648 10950 12650 11002
rect 12650 10950 12702 11002
rect 12702 10950 12704 11002
rect 12648 10948 12704 10950
rect 12572 10834 12628 10836
rect 12572 10782 12574 10834
rect 12574 10782 12626 10834
rect 12626 10782 12628 10834
rect 12572 10780 12628 10782
rect 12572 9826 12628 9828
rect 12572 9774 12574 9826
rect 12574 9774 12626 9826
rect 12626 9774 12628 9826
rect 12572 9772 12628 9774
rect 12440 9434 12496 9436
rect 12440 9382 12442 9434
rect 12442 9382 12494 9434
rect 12494 9382 12496 9434
rect 12440 9380 12496 9382
rect 12544 9434 12600 9436
rect 12544 9382 12546 9434
rect 12546 9382 12598 9434
rect 12598 9382 12600 9434
rect 12544 9380 12600 9382
rect 12648 9434 12704 9436
rect 12648 9382 12650 9434
rect 12650 9382 12702 9434
rect 12702 9382 12704 9434
rect 12648 9380 12704 9382
rect 12440 7866 12496 7868
rect 12440 7814 12442 7866
rect 12442 7814 12494 7866
rect 12494 7814 12496 7866
rect 12440 7812 12496 7814
rect 12544 7866 12600 7868
rect 12544 7814 12546 7866
rect 12546 7814 12598 7866
rect 12598 7814 12600 7866
rect 12544 7812 12600 7814
rect 12648 7866 12704 7868
rect 12648 7814 12650 7866
rect 12650 7814 12702 7866
rect 12702 7814 12704 7866
rect 12648 7812 12704 7814
rect 12440 6298 12496 6300
rect 12440 6246 12442 6298
rect 12442 6246 12494 6298
rect 12494 6246 12496 6298
rect 12440 6244 12496 6246
rect 12544 6298 12600 6300
rect 12544 6246 12546 6298
rect 12546 6246 12598 6298
rect 12598 6246 12600 6298
rect 12544 6244 12600 6246
rect 12648 6298 12704 6300
rect 12648 6246 12650 6298
rect 12650 6246 12702 6298
rect 12702 6246 12704 6298
rect 12648 6244 12704 6246
rect 12460 5852 12516 5908
rect 12440 4730 12496 4732
rect 12440 4678 12442 4730
rect 12442 4678 12494 4730
rect 12494 4678 12496 4730
rect 12440 4676 12496 4678
rect 12544 4730 12600 4732
rect 12544 4678 12546 4730
rect 12546 4678 12598 4730
rect 12598 4678 12600 4730
rect 12544 4676 12600 4678
rect 12648 4730 12704 4732
rect 12648 4678 12650 4730
rect 12650 4678 12702 4730
rect 12702 4678 12704 4730
rect 12648 4676 12704 4678
rect 13356 10780 13412 10836
rect 13356 9826 13412 9828
rect 13356 9774 13358 9826
rect 13358 9774 13410 9826
rect 13410 9774 13412 9826
rect 13356 9772 13412 9774
rect 14028 9772 14084 9828
rect 13692 8988 13748 9044
rect 13132 6578 13188 6580
rect 13132 6526 13134 6578
rect 13134 6526 13186 6578
rect 13186 6526 13188 6578
rect 13132 6524 13188 6526
rect 13244 5852 13300 5908
rect 12908 5234 12964 5236
rect 12908 5182 12910 5234
rect 12910 5182 12962 5234
rect 12962 5182 12964 5234
rect 12908 5180 12964 5182
rect 12440 3162 12496 3164
rect 12440 3110 12442 3162
rect 12442 3110 12494 3162
rect 12494 3110 12496 3162
rect 12440 3108 12496 3110
rect 12544 3162 12600 3164
rect 12544 3110 12546 3162
rect 12546 3110 12598 3162
rect 12598 3110 12600 3162
rect 12544 3108 12600 3110
rect 12648 3162 12704 3164
rect 12648 3110 12650 3162
rect 12650 3110 12702 3162
rect 12702 3110 12704 3162
rect 12648 3108 12704 3110
rect 12124 2156 12180 2212
rect 12236 2044 12292 2100
rect 12460 1986 12516 1988
rect 12460 1934 12462 1986
rect 12462 1934 12514 1986
rect 12514 1934 12516 1986
rect 12460 1932 12516 1934
rect 12440 1594 12496 1596
rect 12440 1542 12442 1594
rect 12442 1542 12494 1594
rect 12494 1542 12496 1594
rect 12440 1540 12496 1542
rect 12544 1594 12600 1596
rect 12544 1542 12546 1594
rect 12546 1542 12598 1594
rect 12598 1542 12600 1594
rect 12544 1540 12600 1542
rect 12648 1594 12704 1596
rect 12648 1542 12650 1594
rect 12650 1542 12702 1594
rect 12702 1542 12704 1594
rect 12648 1540 12704 1542
rect 12908 3500 12964 3556
rect 13132 2770 13188 2772
rect 13132 2718 13134 2770
rect 13134 2718 13186 2770
rect 13186 2718 13188 2770
rect 13132 2716 13188 2718
rect 13916 6972 13972 7028
rect 13916 4172 13972 4228
rect 13692 2098 13748 2100
rect 13692 2046 13694 2098
rect 13694 2046 13746 2098
rect 13746 2046 13748 2098
rect 13692 2044 13748 2046
rect 14140 6524 14196 6580
rect 14498 10218 14554 10220
rect 14498 10166 14500 10218
rect 14500 10166 14552 10218
rect 14552 10166 14554 10218
rect 14498 10164 14554 10166
rect 14602 10218 14658 10220
rect 14602 10166 14604 10218
rect 14604 10166 14656 10218
rect 14656 10166 14658 10218
rect 14602 10164 14658 10166
rect 14706 10218 14762 10220
rect 14706 10166 14708 10218
rect 14708 10166 14760 10218
rect 14760 10166 14762 10218
rect 14706 10164 14762 10166
rect 14924 9884 14980 9940
rect 14588 9042 14644 9044
rect 14588 8990 14590 9042
rect 14590 8990 14642 9042
rect 14642 8990 14644 9042
rect 14588 8988 14644 8990
rect 14498 8650 14554 8652
rect 14498 8598 14500 8650
rect 14500 8598 14552 8650
rect 14552 8598 14554 8650
rect 14498 8596 14554 8598
rect 14602 8650 14658 8652
rect 14602 8598 14604 8650
rect 14604 8598 14656 8650
rect 14656 8598 14658 8650
rect 14602 8596 14658 8598
rect 14706 8650 14762 8652
rect 14706 8598 14708 8650
rect 14708 8598 14760 8650
rect 14760 8598 14762 8650
rect 14706 8596 14762 8598
rect 15596 9042 15652 9044
rect 15596 8990 15598 9042
rect 15598 8990 15650 9042
rect 15650 8990 15652 9042
rect 15596 8988 15652 8990
rect 16156 9938 16212 9940
rect 16156 9886 16158 9938
rect 16158 9886 16210 9938
rect 16210 9886 16212 9938
rect 16156 9884 16212 9886
rect 14252 5906 14308 5908
rect 14252 5854 14254 5906
rect 14254 5854 14306 5906
rect 14306 5854 14308 5906
rect 14252 5852 14308 5854
rect 14498 7082 14554 7084
rect 14498 7030 14500 7082
rect 14500 7030 14552 7082
rect 14552 7030 14554 7082
rect 14498 7028 14554 7030
rect 14602 7082 14658 7084
rect 14602 7030 14604 7082
rect 14604 7030 14656 7082
rect 14656 7030 14658 7082
rect 14602 7028 14658 7030
rect 14706 7082 14762 7084
rect 14706 7030 14708 7082
rect 14708 7030 14760 7082
rect 14760 7030 14762 7082
rect 14706 7028 14762 7030
rect 14498 5514 14554 5516
rect 14498 5462 14500 5514
rect 14500 5462 14552 5514
rect 14552 5462 14554 5514
rect 14498 5460 14554 5462
rect 14602 5514 14658 5516
rect 14602 5462 14604 5514
rect 14604 5462 14656 5514
rect 14656 5462 14658 5514
rect 14602 5460 14658 5462
rect 14706 5514 14762 5516
rect 14706 5462 14708 5514
rect 14708 5462 14760 5514
rect 14760 5462 14762 5514
rect 14706 5460 14762 5462
rect 14364 5068 14420 5124
rect 14252 3388 14308 3444
rect 14924 4226 14980 4228
rect 14924 4174 14926 4226
rect 14926 4174 14978 4226
rect 14978 4174 14980 4226
rect 14924 4172 14980 4174
rect 15036 4060 15092 4116
rect 14498 3946 14554 3948
rect 14498 3894 14500 3946
rect 14500 3894 14552 3946
rect 14552 3894 14554 3946
rect 14498 3892 14554 3894
rect 14602 3946 14658 3948
rect 14602 3894 14604 3946
rect 14604 3894 14656 3946
rect 14656 3894 14658 3946
rect 14602 3892 14658 3894
rect 14706 3946 14762 3948
rect 14706 3894 14708 3946
rect 14708 3894 14760 3946
rect 14760 3894 14762 3946
rect 14706 3892 14762 3894
rect 15260 6130 15316 6132
rect 15260 6078 15262 6130
rect 15262 6078 15314 6130
rect 15314 6078 15316 6130
rect 15260 6076 15316 6078
rect 15372 5068 15428 5124
rect 14588 3554 14644 3556
rect 14588 3502 14590 3554
rect 14590 3502 14642 3554
rect 14642 3502 14644 3554
rect 14588 3500 14644 3502
rect 14498 2378 14554 2380
rect 14498 2326 14500 2378
rect 14500 2326 14552 2378
rect 14552 2326 14554 2378
rect 14498 2324 14554 2326
rect 14602 2378 14658 2380
rect 14602 2326 14604 2378
rect 14604 2326 14656 2378
rect 14656 2326 14658 2378
rect 14602 2324 14658 2326
rect 14706 2378 14762 2380
rect 14706 2326 14708 2378
rect 14708 2326 14760 2378
rect 14760 2326 14762 2378
rect 14706 2324 14762 2326
rect 15820 4060 15876 4116
rect 15596 3554 15652 3556
rect 15596 3502 15598 3554
rect 15598 3502 15650 3554
rect 15650 3502 15652 3554
rect 15596 3500 15652 3502
rect 16556 11002 16612 11004
rect 16556 10950 16558 11002
rect 16558 10950 16610 11002
rect 16610 10950 16612 11002
rect 16556 10948 16612 10950
rect 16660 11002 16716 11004
rect 16660 10950 16662 11002
rect 16662 10950 16714 11002
rect 16714 10950 16716 11002
rect 16660 10948 16716 10950
rect 16764 11002 16820 11004
rect 16764 10950 16766 11002
rect 16766 10950 16818 11002
rect 16818 10950 16820 11002
rect 16764 10948 16820 10950
rect 16556 9434 16612 9436
rect 16556 9382 16558 9434
rect 16558 9382 16610 9434
rect 16610 9382 16612 9434
rect 16556 9380 16612 9382
rect 16660 9434 16716 9436
rect 16660 9382 16662 9434
rect 16662 9382 16714 9434
rect 16714 9382 16716 9434
rect 16660 9380 16716 9382
rect 16764 9434 16820 9436
rect 16764 9382 16766 9434
rect 16766 9382 16818 9434
rect 16818 9382 16820 9434
rect 16764 9380 16820 9382
rect 16556 7866 16612 7868
rect 16556 7814 16558 7866
rect 16558 7814 16610 7866
rect 16610 7814 16612 7866
rect 16556 7812 16612 7814
rect 16660 7866 16716 7868
rect 16660 7814 16662 7866
rect 16662 7814 16714 7866
rect 16714 7814 16716 7866
rect 16660 7812 16716 7814
rect 16764 7866 16820 7868
rect 16764 7814 16766 7866
rect 16766 7814 16818 7866
rect 16818 7814 16820 7866
rect 16764 7812 16820 7814
rect 16044 6524 16100 6580
rect 16556 6298 16612 6300
rect 16556 6246 16558 6298
rect 16558 6246 16610 6298
rect 16610 6246 16612 6298
rect 16556 6244 16612 6246
rect 16660 6298 16716 6300
rect 16660 6246 16662 6298
rect 16662 6246 16714 6298
rect 16714 6246 16716 6298
rect 16660 6244 16716 6246
rect 16764 6298 16820 6300
rect 16764 6246 16766 6298
rect 16766 6246 16818 6298
rect 16818 6246 16820 6298
rect 16764 6244 16820 6246
rect 16556 4730 16612 4732
rect 16556 4678 16558 4730
rect 16558 4678 16610 4730
rect 16610 4678 16612 4730
rect 16556 4676 16612 4678
rect 16660 4730 16716 4732
rect 16660 4678 16662 4730
rect 16662 4678 16714 4730
rect 16714 4678 16716 4730
rect 16660 4676 16716 4678
rect 16764 4730 16820 4732
rect 16764 4678 16766 4730
rect 16766 4678 16818 4730
rect 16818 4678 16820 4730
rect 16764 4676 16820 4678
rect 16556 3162 16612 3164
rect 16556 3110 16558 3162
rect 16558 3110 16610 3162
rect 16610 3110 16612 3162
rect 16556 3108 16612 3110
rect 16660 3162 16716 3164
rect 16660 3110 16662 3162
rect 16662 3110 16714 3162
rect 16714 3110 16716 3162
rect 16660 3108 16716 3110
rect 16764 3162 16820 3164
rect 16764 3110 16766 3162
rect 16766 3110 16818 3162
rect 16818 3110 16820 3162
rect 16764 3108 16820 3110
rect 16556 1594 16612 1596
rect 16556 1542 16558 1594
rect 16558 1542 16610 1594
rect 16610 1542 16612 1594
rect 16556 1540 16612 1542
rect 16660 1594 16716 1596
rect 16660 1542 16662 1594
rect 16662 1542 16714 1594
rect 16714 1542 16716 1594
rect 16660 1540 16716 1542
rect 16764 1594 16820 1596
rect 16764 1542 16766 1594
rect 16766 1542 16818 1594
rect 16818 1542 16820 1594
rect 16764 1540 16820 1542
<< metal3 >>
rect 4198 10948 4208 11004
rect 4264 10948 4312 11004
rect 4368 10948 4416 11004
rect 4472 10948 4482 11004
rect 8314 10948 8324 11004
rect 8380 10948 8428 11004
rect 8484 10948 8532 11004
rect 8588 10948 8598 11004
rect 12430 10948 12440 11004
rect 12496 10948 12544 11004
rect 12600 10948 12648 11004
rect 12704 10948 12714 11004
rect 16546 10948 16556 11004
rect 16612 10948 16660 11004
rect 16716 10948 16764 11004
rect 16820 10948 16830 11004
rect 12562 10780 12572 10836
rect 12628 10780 13356 10836
rect 13412 10780 13422 10836
rect 0 10724 800 10752
rect 16200 10724 17000 10752
rect 0 10668 4732 10724
rect 4788 10668 4798 10724
rect 11778 10668 11788 10724
rect 11844 10668 17000 10724
rect 0 10640 800 10668
rect 16200 10640 17000 10668
rect 2594 10444 2604 10500
rect 2660 10444 3724 10500
rect 3780 10444 3790 10500
rect 10434 10332 10444 10388
rect 10500 10332 11228 10388
rect 11284 10332 11294 10388
rect 2140 10164 2150 10220
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2414 10164 2424 10220
rect 6256 10164 6266 10220
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6530 10164 6540 10220
rect 10372 10164 10382 10220
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10646 10164 10656 10220
rect 14488 10164 14498 10220
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14762 10164 14772 10220
rect 14914 9884 14924 9940
rect 14980 9884 16156 9940
rect 16212 9884 16222 9940
rect 12562 9772 12572 9828
rect 12628 9772 13356 9828
rect 13412 9772 14028 9828
rect 14084 9772 14094 9828
rect 8194 9660 8204 9716
rect 8260 9660 9212 9716
rect 9268 9660 10220 9716
rect 10276 9660 10286 9716
rect 2940 9548 4508 9604
rect 4564 9548 4574 9604
rect 6626 9548 6636 9604
rect 6692 9548 7420 9604
rect 7476 9548 7486 9604
rect 2940 9492 2996 9548
rect 1922 9436 1932 9492
rect 1988 9436 2940 9492
rect 2996 9436 3006 9492
rect 4198 9380 4208 9436
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4472 9380 4482 9436
rect 8314 9380 8324 9436
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8588 9380 8598 9436
rect 12430 9380 12440 9436
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12704 9380 12714 9436
rect 16546 9380 16556 9436
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16820 9380 16830 9436
rect 4722 8988 4732 9044
rect 4788 8988 5292 9044
rect 5348 8988 5358 9044
rect 13682 8988 13692 9044
rect 13748 8988 14588 9044
rect 14644 8988 15596 9044
rect 15652 8988 15662 9044
rect 7634 8876 7644 8932
rect 7700 8876 11788 8932
rect 11844 8876 11854 8932
rect 2140 8596 2150 8652
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2414 8596 2424 8652
rect 6256 8596 6266 8652
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6530 8596 6540 8652
rect 10372 8596 10382 8652
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10646 8596 10656 8652
rect 14488 8596 14498 8652
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14762 8596 14772 8652
rect 3938 8316 3948 8372
rect 4004 8316 5740 8372
rect 5796 8316 5806 8372
rect 7746 8316 7756 8372
rect 7812 8316 10108 8372
rect 10164 8316 10174 8372
rect 1474 8204 1484 8260
rect 1540 8204 2716 8260
rect 2772 8204 3724 8260
rect 3780 8204 3790 8260
rect 8866 8204 8876 8260
rect 8932 8204 9660 8260
rect 9716 8204 10668 8260
rect 10724 8204 10734 8260
rect 4198 7812 4208 7868
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4472 7812 4482 7868
rect 8314 7812 8324 7868
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8588 7812 8598 7868
rect 12430 7812 12440 7868
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12704 7812 12714 7868
rect 16546 7812 16556 7868
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16820 7812 16830 7868
rect 9538 7196 9548 7252
rect 9604 7196 10780 7252
rect 10836 7196 11564 7252
rect 11620 7196 11630 7252
rect 2140 7028 2150 7084
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2414 7028 2424 7084
rect 6256 7028 6266 7084
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6530 7028 6540 7084
rect 10372 7028 10382 7084
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10646 7028 10656 7084
rect 14488 7028 14498 7084
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14762 7028 14772 7084
rect 11890 6972 11900 7028
rect 11956 6972 13916 7028
rect 13972 6972 13982 7028
rect 10882 6748 10892 6804
rect 10948 6748 11788 6804
rect 11844 6748 11854 6804
rect 2818 6636 2828 6692
rect 2884 6636 3836 6692
rect 3892 6636 4732 6692
rect 4788 6636 4798 6692
rect 7746 6636 7756 6692
rect 7812 6636 8540 6692
rect 8596 6636 8764 6692
rect 8820 6636 8830 6692
rect 2706 6524 2716 6580
rect 2772 6524 3724 6580
rect 3780 6524 3790 6580
rect 4834 6524 4844 6580
rect 4900 6524 5404 6580
rect 5460 6524 5470 6580
rect 13122 6524 13132 6580
rect 13188 6524 14140 6580
rect 14196 6524 16044 6580
rect 16100 6524 16110 6580
rect 0 6468 800 6496
rect 4844 6468 4900 6524
rect 16200 6468 17000 6496
rect 0 6412 4900 6468
rect 7186 6412 7196 6468
rect 7252 6412 17000 6468
rect 0 6384 800 6412
rect 16200 6384 17000 6412
rect 4198 6244 4208 6300
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4472 6244 4482 6300
rect 8314 6244 8324 6300
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8588 6244 8598 6300
rect 12430 6244 12440 6300
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12704 6244 12714 6300
rect 16546 6244 16556 6300
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16820 6244 16830 6300
rect 3154 6076 3164 6132
rect 3220 6076 4620 6132
rect 4676 6076 4686 6132
rect 15092 6076 15260 6132
rect 15316 6076 15326 6132
rect 15092 5908 15148 6076
rect 4722 5852 4732 5908
rect 4788 5852 5180 5908
rect 5236 5852 5246 5908
rect 9986 5852 9996 5908
rect 10052 5852 11116 5908
rect 11172 5852 12460 5908
rect 12516 5852 12526 5908
rect 13234 5852 13244 5908
rect 13300 5852 14252 5908
rect 14308 5852 15148 5908
rect 7298 5740 7308 5796
rect 7364 5740 8540 5796
rect 8596 5740 8606 5796
rect 2482 5516 2492 5572
rect 2548 5516 3388 5572
rect 3444 5516 3454 5572
rect 2140 5460 2150 5516
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2414 5460 2424 5516
rect 6256 5460 6266 5516
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6530 5460 6540 5516
rect 10372 5460 10382 5516
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10646 5460 10656 5516
rect 14488 5460 14498 5516
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14762 5460 14772 5516
rect 3266 5292 3276 5348
rect 3332 5292 4732 5348
rect 4788 5292 4798 5348
rect 11218 5180 11228 5236
rect 11284 5180 12908 5236
rect 12964 5180 12974 5236
rect 578 5068 588 5124
rect 644 5068 2716 5124
rect 2772 5068 2782 5124
rect 14354 5068 14364 5124
rect 14420 5068 15372 5124
rect 15428 5068 15438 5124
rect 4198 4676 4208 4732
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4472 4676 4482 4732
rect 8314 4676 8324 4732
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8588 4676 8598 4732
rect 12430 4676 12440 4732
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12704 4676 12714 4732
rect 16546 4676 16556 4732
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16820 4676 16830 4732
rect 1026 4284 1036 4340
rect 1092 4284 2604 4340
rect 2660 4284 2670 4340
rect 6066 4284 6076 4340
rect 6132 4284 6860 4340
rect 6916 4284 7868 4340
rect 7924 4284 7934 4340
rect 13906 4172 13916 4228
rect 13972 4172 14924 4228
rect 14980 4172 14990 4228
rect 15026 4060 15036 4116
rect 15092 4060 15820 4116
rect 15876 4060 15886 4116
rect 2140 3892 2150 3948
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2414 3892 2424 3948
rect 6256 3892 6266 3948
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6530 3892 6540 3948
rect 10372 3892 10382 3948
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10646 3892 10656 3948
rect 14488 3892 14498 3948
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14762 3892 14772 3948
rect 9426 3612 9436 3668
rect 9492 3612 12124 3668
rect 12180 3612 12190 3668
rect 4834 3500 4844 3556
rect 4900 3500 6524 3556
rect 6580 3500 7084 3556
rect 7140 3500 7150 3556
rect 12898 3500 12908 3556
rect 12964 3500 14588 3556
rect 14644 3500 15596 3556
rect 15652 3500 15662 3556
rect 3938 3388 3948 3444
rect 4004 3388 4732 3444
rect 4788 3388 4798 3444
rect 11442 3388 11452 3444
rect 11508 3388 14252 3444
rect 14308 3388 14318 3444
rect 2706 3276 2716 3332
rect 2772 3276 5068 3332
rect 5124 3276 5134 3332
rect 4198 3108 4208 3164
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4472 3108 4482 3164
rect 8314 3108 8324 3164
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8588 3108 8598 3164
rect 12430 3108 12440 3164
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12704 3108 12714 3164
rect 16546 3108 16556 3164
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16820 3108 16830 3164
rect 11666 2716 11676 2772
rect 11732 2716 13132 2772
rect 13188 2716 13198 2772
rect 7522 2604 7532 2660
rect 7588 2604 8540 2660
rect 8596 2604 8606 2660
rect 3714 2492 3724 2548
rect 3780 2492 4284 2548
rect 4340 2492 4956 2548
rect 5012 2492 5022 2548
rect 2140 2324 2150 2380
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2414 2324 2424 2380
rect 6256 2324 6266 2380
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6530 2324 6540 2380
rect 10372 2324 10382 2380
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10646 2324 10656 2380
rect 14488 2324 14498 2380
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14762 2324 14772 2380
rect 0 2212 800 2240
rect 16200 2212 17000 2240
rect 0 2156 4844 2212
rect 4900 2156 4910 2212
rect 6402 2156 6412 2212
rect 6468 2156 7532 2212
rect 7588 2156 7598 2212
rect 12114 2156 12124 2212
rect 12180 2156 17000 2212
rect 0 2128 800 2156
rect 16200 2128 17000 2156
rect 12226 2044 12236 2100
rect 12292 2044 13692 2100
rect 13748 2044 13758 2100
rect 3826 1932 3836 1988
rect 3892 1932 4732 1988
rect 4788 1932 5068 1988
rect 5124 1932 5134 1988
rect 11330 1932 11340 1988
rect 11396 1932 12460 1988
rect 12516 1932 12526 1988
rect 5506 1820 5516 1876
rect 5572 1820 6748 1876
rect 6804 1820 7644 1876
rect 7700 1820 7710 1876
rect 4198 1540 4208 1596
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4472 1540 4482 1596
rect 8314 1540 8324 1596
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8588 1540 8598 1596
rect 12430 1540 12440 1596
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12704 1540 12714 1596
rect 16546 1540 16556 1596
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16820 1540 16830 1596
<< via3 >>
rect 4208 10948 4264 11004
rect 4312 10948 4368 11004
rect 4416 10948 4472 11004
rect 8324 10948 8380 11004
rect 8428 10948 8484 11004
rect 8532 10948 8588 11004
rect 12440 10948 12496 11004
rect 12544 10948 12600 11004
rect 12648 10948 12704 11004
rect 16556 10948 16612 11004
rect 16660 10948 16716 11004
rect 16764 10948 16820 11004
rect 2150 10164 2206 10220
rect 2254 10164 2310 10220
rect 2358 10164 2414 10220
rect 6266 10164 6322 10220
rect 6370 10164 6426 10220
rect 6474 10164 6530 10220
rect 10382 10164 10438 10220
rect 10486 10164 10542 10220
rect 10590 10164 10646 10220
rect 14498 10164 14554 10220
rect 14602 10164 14658 10220
rect 14706 10164 14762 10220
rect 4208 9380 4264 9436
rect 4312 9380 4368 9436
rect 4416 9380 4472 9436
rect 8324 9380 8380 9436
rect 8428 9380 8484 9436
rect 8532 9380 8588 9436
rect 12440 9380 12496 9436
rect 12544 9380 12600 9436
rect 12648 9380 12704 9436
rect 16556 9380 16612 9436
rect 16660 9380 16716 9436
rect 16764 9380 16820 9436
rect 2150 8596 2206 8652
rect 2254 8596 2310 8652
rect 2358 8596 2414 8652
rect 6266 8596 6322 8652
rect 6370 8596 6426 8652
rect 6474 8596 6530 8652
rect 10382 8596 10438 8652
rect 10486 8596 10542 8652
rect 10590 8596 10646 8652
rect 14498 8596 14554 8652
rect 14602 8596 14658 8652
rect 14706 8596 14762 8652
rect 4208 7812 4264 7868
rect 4312 7812 4368 7868
rect 4416 7812 4472 7868
rect 8324 7812 8380 7868
rect 8428 7812 8484 7868
rect 8532 7812 8588 7868
rect 12440 7812 12496 7868
rect 12544 7812 12600 7868
rect 12648 7812 12704 7868
rect 16556 7812 16612 7868
rect 16660 7812 16716 7868
rect 16764 7812 16820 7868
rect 2150 7028 2206 7084
rect 2254 7028 2310 7084
rect 2358 7028 2414 7084
rect 6266 7028 6322 7084
rect 6370 7028 6426 7084
rect 6474 7028 6530 7084
rect 10382 7028 10438 7084
rect 10486 7028 10542 7084
rect 10590 7028 10646 7084
rect 14498 7028 14554 7084
rect 14602 7028 14658 7084
rect 14706 7028 14762 7084
rect 4208 6244 4264 6300
rect 4312 6244 4368 6300
rect 4416 6244 4472 6300
rect 8324 6244 8380 6300
rect 8428 6244 8484 6300
rect 8532 6244 8588 6300
rect 12440 6244 12496 6300
rect 12544 6244 12600 6300
rect 12648 6244 12704 6300
rect 16556 6244 16612 6300
rect 16660 6244 16716 6300
rect 16764 6244 16820 6300
rect 2150 5460 2206 5516
rect 2254 5460 2310 5516
rect 2358 5460 2414 5516
rect 6266 5460 6322 5516
rect 6370 5460 6426 5516
rect 6474 5460 6530 5516
rect 10382 5460 10438 5516
rect 10486 5460 10542 5516
rect 10590 5460 10646 5516
rect 14498 5460 14554 5516
rect 14602 5460 14658 5516
rect 14706 5460 14762 5516
rect 4208 4676 4264 4732
rect 4312 4676 4368 4732
rect 4416 4676 4472 4732
rect 8324 4676 8380 4732
rect 8428 4676 8484 4732
rect 8532 4676 8588 4732
rect 12440 4676 12496 4732
rect 12544 4676 12600 4732
rect 12648 4676 12704 4732
rect 16556 4676 16612 4732
rect 16660 4676 16716 4732
rect 16764 4676 16820 4732
rect 2150 3892 2206 3948
rect 2254 3892 2310 3948
rect 2358 3892 2414 3948
rect 6266 3892 6322 3948
rect 6370 3892 6426 3948
rect 6474 3892 6530 3948
rect 10382 3892 10438 3948
rect 10486 3892 10542 3948
rect 10590 3892 10646 3948
rect 14498 3892 14554 3948
rect 14602 3892 14658 3948
rect 14706 3892 14762 3948
rect 4208 3108 4264 3164
rect 4312 3108 4368 3164
rect 4416 3108 4472 3164
rect 8324 3108 8380 3164
rect 8428 3108 8484 3164
rect 8532 3108 8588 3164
rect 12440 3108 12496 3164
rect 12544 3108 12600 3164
rect 12648 3108 12704 3164
rect 16556 3108 16612 3164
rect 16660 3108 16716 3164
rect 16764 3108 16820 3164
rect 2150 2324 2206 2380
rect 2254 2324 2310 2380
rect 2358 2324 2414 2380
rect 6266 2324 6322 2380
rect 6370 2324 6426 2380
rect 6474 2324 6530 2380
rect 10382 2324 10438 2380
rect 10486 2324 10542 2380
rect 10590 2324 10646 2380
rect 14498 2324 14554 2380
rect 14602 2324 14658 2380
rect 14706 2324 14762 2380
rect 4208 1540 4264 1596
rect 4312 1540 4368 1596
rect 4416 1540 4472 1596
rect 8324 1540 8380 1596
rect 8428 1540 8484 1596
rect 8532 1540 8588 1596
rect 12440 1540 12496 1596
rect 12544 1540 12600 1596
rect 12648 1540 12704 1596
rect 16556 1540 16612 1596
rect 16660 1540 16716 1596
rect 16764 1540 16820 1596
<< metal4 >>
rect 2122 10220 2442 11036
rect 2122 10164 2150 10220
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2414 10164 2442 10220
rect 2122 8652 2442 10164
rect 2122 8596 2150 8652
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2414 8596 2442 8652
rect 2122 7084 2442 8596
rect 2122 7028 2150 7084
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2414 7028 2442 7084
rect 2122 5516 2442 7028
rect 2122 5460 2150 5516
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2414 5460 2442 5516
rect 2122 3948 2442 5460
rect 2122 3892 2150 3948
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2414 3892 2442 3948
rect 2122 2380 2442 3892
rect 2122 2324 2150 2380
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2414 2324 2442 2380
rect 2122 1508 2442 2324
rect 4180 11004 4500 11036
rect 4180 10948 4208 11004
rect 4264 10948 4312 11004
rect 4368 10948 4416 11004
rect 4472 10948 4500 11004
rect 4180 9436 4500 10948
rect 4180 9380 4208 9436
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4472 9380 4500 9436
rect 4180 7868 4500 9380
rect 4180 7812 4208 7868
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4472 7812 4500 7868
rect 4180 6300 4500 7812
rect 4180 6244 4208 6300
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4472 6244 4500 6300
rect 4180 4732 4500 6244
rect 4180 4676 4208 4732
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4472 4676 4500 4732
rect 4180 3164 4500 4676
rect 4180 3108 4208 3164
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4472 3108 4500 3164
rect 4180 1596 4500 3108
rect 4180 1540 4208 1596
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4472 1540 4500 1596
rect 4180 1508 4500 1540
rect 6238 10220 6558 11036
rect 6238 10164 6266 10220
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6530 10164 6558 10220
rect 6238 8652 6558 10164
rect 6238 8596 6266 8652
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6530 8596 6558 8652
rect 6238 7084 6558 8596
rect 6238 7028 6266 7084
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6530 7028 6558 7084
rect 6238 5516 6558 7028
rect 6238 5460 6266 5516
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6530 5460 6558 5516
rect 6238 3948 6558 5460
rect 6238 3892 6266 3948
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6530 3892 6558 3948
rect 6238 2380 6558 3892
rect 6238 2324 6266 2380
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6530 2324 6558 2380
rect 6238 1508 6558 2324
rect 8296 11004 8616 11036
rect 8296 10948 8324 11004
rect 8380 10948 8428 11004
rect 8484 10948 8532 11004
rect 8588 10948 8616 11004
rect 8296 9436 8616 10948
rect 8296 9380 8324 9436
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8588 9380 8616 9436
rect 8296 7868 8616 9380
rect 8296 7812 8324 7868
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8588 7812 8616 7868
rect 8296 6300 8616 7812
rect 8296 6244 8324 6300
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8588 6244 8616 6300
rect 8296 4732 8616 6244
rect 8296 4676 8324 4732
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8588 4676 8616 4732
rect 8296 3164 8616 4676
rect 8296 3108 8324 3164
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8588 3108 8616 3164
rect 8296 1596 8616 3108
rect 8296 1540 8324 1596
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8588 1540 8616 1596
rect 8296 1508 8616 1540
rect 10354 10220 10674 11036
rect 10354 10164 10382 10220
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10646 10164 10674 10220
rect 10354 8652 10674 10164
rect 10354 8596 10382 8652
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10646 8596 10674 8652
rect 10354 7084 10674 8596
rect 10354 7028 10382 7084
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10646 7028 10674 7084
rect 10354 5516 10674 7028
rect 10354 5460 10382 5516
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10646 5460 10674 5516
rect 10354 3948 10674 5460
rect 10354 3892 10382 3948
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10646 3892 10674 3948
rect 10354 2380 10674 3892
rect 10354 2324 10382 2380
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10646 2324 10674 2380
rect 10354 1508 10674 2324
rect 12412 11004 12732 11036
rect 12412 10948 12440 11004
rect 12496 10948 12544 11004
rect 12600 10948 12648 11004
rect 12704 10948 12732 11004
rect 12412 9436 12732 10948
rect 12412 9380 12440 9436
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12704 9380 12732 9436
rect 12412 7868 12732 9380
rect 12412 7812 12440 7868
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12704 7812 12732 7868
rect 12412 6300 12732 7812
rect 12412 6244 12440 6300
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12704 6244 12732 6300
rect 12412 4732 12732 6244
rect 12412 4676 12440 4732
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12704 4676 12732 4732
rect 12412 3164 12732 4676
rect 12412 3108 12440 3164
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12704 3108 12732 3164
rect 12412 1596 12732 3108
rect 12412 1540 12440 1596
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12704 1540 12732 1596
rect 12412 1508 12732 1540
rect 14470 10220 14790 11036
rect 14470 10164 14498 10220
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14762 10164 14790 10220
rect 14470 8652 14790 10164
rect 14470 8596 14498 8652
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14762 8596 14790 8652
rect 14470 7084 14790 8596
rect 14470 7028 14498 7084
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14762 7028 14790 7084
rect 14470 5516 14790 7028
rect 14470 5460 14498 5516
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14762 5460 14790 5516
rect 14470 3948 14790 5460
rect 14470 3892 14498 3948
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14762 3892 14790 3948
rect 14470 2380 14790 3892
rect 14470 2324 14498 2380
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14762 2324 14790 2380
rect 14470 1508 14790 2324
rect 16528 11004 16848 11036
rect 16528 10948 16556 11004
rect 16612 10948 16660 11004
rect 16716 10948 16764 11004
rect 16820 10948 16848 11004
rect 16528 9436 16848 10948
rect 16528 9380 16556 9436
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16820 9380 16848 9436
rect 16528 7868 16848 9380
rect 16528 7812 16556 7868
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16820 7812 16848 7868
rect 16528 6300 16848 7812
rect 16528 6244 16556 6300
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16820 6244 16848 6300
rect 16528 4732 16848 6244
rect 16528 4676 16556 4732
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16820 4676 16848 4732
rect 16528 3164 16848 4676
rect 16528 3108 16556 3164
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16820 3108 16848 3164
rect 16528 1596 16848 3108
rect 16528 1540 16556 1596
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16820 1540 16848 1596
rect 16528 1508 16848 1540
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[0\]_I OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 10640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[1\]_I
timestamp 1666464484
transform 1 0 11536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[2\]_I
timestamp 1666464484
transform 1 0 11536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[3\]_I
timestamp 1666464484
transform 1 0 12432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[4\]_I
timestamp 1666464484
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[5\]_I
timestamp 1666464484
transform 1 0 11760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[6\]_I
timestamp 1666464484
transform -1 0 11872 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[7\]_I
timestamp 1666464484
transform 1 0 14896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[8\]_I
timestamp 1666464484
transform -1 0 11424 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[9\]_I
timestamp 1666464484
transform 1 0 15568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[10\]_I
timestamp 1666464484
transform 1 0 15232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[11\]_I
timestamp 1666464484
transform 1 0 15568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[12\]_I
timestamp 1666464484
transform -1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[13\]_I
timestamp 1666464484
transform -1 0 12656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[14\]_I
timestamp 1666464484
transform 1 0 16128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[15\]_I
timestamp 1666464484
transform 1 0 15792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[16\]_I
timestamp 1666464484
transform 1 0 15792 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[17\]_I
timestamp 1666464484
transform -1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[18\]_I
timestamp 1666464484
transform 1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[19\]_I
timestamp 1666464484
transform 1 0 4816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[20\]_I
timestamp 1666464484
transform 1 0 4704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[21\]_I
timestamp 1666464484
transform 1 0 3696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[22\]_I
timestamp 1666464484
transform 1 0 3696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[23\]_I
timestamp 1666464484
transform 1 0 3696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[24\]_I
timestamp 1666464484
transform 1 0 4480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[25\]_I
timestamp 1666464484
transform 1 0 4480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[26\]_I
timestamp 1666464484
transform 1 0 4704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[27\]_I
timestamp 1666464484
transform 1 0 5152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[28\]_I
timestamp 1666464484
transform 1 0 4928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[29\]_I
timestamp 1666464484
transform -1 0 4032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[30\]_I
timestamp 1666464484
transform 1 0 4480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[31\]_I
timestamp 1666464484
transform -1 0 4032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[32\]_I
timestamp 1666464484
transform 1 0 7616 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[33\]_I
timestamp 1666464484
transform 1 0 7840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[34\]_I
timestamp 1666464484
transform 1 0 8512 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[35\]_I
timestamp 1666464484
transform 1 0 8512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[36\]_I
timestamp 1666464484
transform 1 0 6608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[37\]_I
timestamp 1666464484
transform 1 0 8512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[38\]_I
timestamp 1666464484
transform 1 0 10192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 10416 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[1\]
timestamp 1666464484
transform -1 0 11312 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[2\]
timestamp 1666464484
transform -1 0 11312 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[3\]
timestamp 1666464484
transform -1 0 11872 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[4\]
timestamp 1666464484
transform -1 0 11984 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[5\]
timestamp 1666464484
transform -1 0 12768 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[6\]
timestamp 1666464484
transform 1 0 12992 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[7\]
timestamp 1666464484
transform -1 0 14672 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[8\]
timestamp 1666464484
transform 1 0 12320 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[9\]
timestamp 1666464484
transform -1 0 15344 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[10\]
timestamp 1666464484
transform -1 0 15008 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[11\]
timestamp 1666464484
transform -1 0 15344 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[12\]
timestamp 1666464484
transform 1 0 12880 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[13\]
timestamp 1666464484
transform 1 0 12880 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[14\]
timestamp 1666464484
transform -1 0 16352 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[15\]
timestamp 1666464484
transform -1 0 16016 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[16\]
timestamp 1666464484
transform -1 0 16352 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[17\]
timestamp 1666464484
transform 1 0 13440 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[18\]
timestamp 1666464484
transform 1 0 6944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[19\]
timestamp 1666464484
transform 1 0 5264 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[20\]
timestamp 1666464484
transform 1 0 5152 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[21\]
timestamp 1666464484
transform -1 0 3472 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[22\]
timestamp 1666464484
transform -1 0 3472 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[23\]
timestamp 1666464484
transform -1 0 3472 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[24\]
timestamp 1666464484
transform -1 0 3696 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[25\]
timestamp 1666464484
transform -1 0 4144 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[26\]
timestamp 1666464484
transform -1 0 4480 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[27\]
timestamp 1666464484
transform -1 0 4928 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[28\]
timestamp 1666464484
transform -1 0 4928 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[29\]
timestamp 1666464484
transform 1 0 4480 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[30\]
timestamp 1666464484
transform -1 0 4480 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[31\]
timestamp 1666464484
transform -1 0 4032 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[32\]
timestamp 1666464484
transform -1 0 7392 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[33\]
timestamp 1666464484
transform -1 0 7616 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[34\]
timestamp 1666464484
transform -1 0 8064 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[35\]
timestamp 1666464484
transform -1 0 8064 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[36\]
timestamp 1666464484
transform -1 0 7952 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[37\]
timestamp 1666464484
transform 1 0 8512 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[38\]
timestamp 1666464484
transform -1 0 9968 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 448 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 896 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4032 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1666464484
transform 1 0 4368 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64
timestamp 1666464484
transform 1 0 7392 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1666464484
transform 1 0 7840 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 8288 0 1 1568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 10080 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96
timestamp 1666464484
transform 1 0 10976 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100
timestamp 1666464484
transform 1 0 11424 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1666464484
transform 1 0 11872 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1666464484
transform 1 0 12208 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134
timestamp 1666464484
transform 1 0 15232 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 15680 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1666464484
transform 1 0 16128 0 1 1568
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1666464484
transform 1 0 16352 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2
timestamp 1666464484
transform 1 0 448 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_10
timestamp 1666464484
transform 1 0 1344 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_14
timestamp 1666464484
transform 1 0 1792 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1666464484
transform 1 0 4928 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1666464484
transform 1 0 8064 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1666464484
transform 1 0 8400 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_76
timestamp 1666464484
transform 1 0 8736 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_84
timestamp 1666464484
transform 1 0 9632 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_112
timestamp 1666464484
transform 1 0 12768 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_140
timestamp 1666464484
transform 1 0 15904 0 -1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1666464484
transform 1 0 16352 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_2
timestamp 1666464484
transform 1 0 448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_18
timestamp 1666464484
transform 1 0 2240 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_26
timestamp 1666464484
transform 1 0 3136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_30
timestamp 1666464484
transform 1 0 3584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 4032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1666464484
transform 1 0 4368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_40
timestamp 1666464484
transform 1 0 4704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_44
timestamp 1666464484
transform 1 0 5152 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_52
timestamp 1666464484
transform 1 0 6048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_58
timestamp 1666464484
transform 1 0 6720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_86
timestamp 1666464484
transform 1 0 9856 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_102
timestamp 1666464484
transform 1 0 11648 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 11984 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1666464484
transform 1 0 12320 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_135
timestamp 1666464484
transform 1 0 15344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_139
timestamp 1666464484
transform 1 0 15792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_143
timestamp 1666464484
transform 1 0 16240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_2
timestamp 1666464484
transform 1 0 448 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_10
timestamp 1666464484
transform 1 0 1344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_38
timestamp 1666464484
transform 1 0 4480 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_66
timestamp 1666464484
transform 1 0 7616 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 8064 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_73
timestamp 1666464484
transform 1 0 8400 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_89
timestamp 1666464484
transform 1 0 10192 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_97
timestamp 1666464484
transform 1 0 11088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_101
timestamp 1666464484
transform 1 0 11536 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_129
timestamp 1666464484
transform 1 0 14672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_133
timestamp 1666464484
transform 1 0 15120 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_137
timestamp 1666464484
transform 1 0 15568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1666464484
transform 1 0 16016 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1666464484
transform 1 0 16352 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_2
timestamp 1666464484
transform 1 0 448 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_18
timestamp 1666464484
transform 1 0 2240 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_26
timestamp 1666464484
transform 1 0 3136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_30
timestamp 1666464484
transform 1 0 3584 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 4032 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1666464484
transform 1 0 4368 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_64
timestamp 1666464484
transform 1 0 7392 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_72
timestamp 1666464484
transform 1 0 8288 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_76
timestamp 1666464484
transform 1 0 8736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_78
timestamp 1666464484
transform 1 0 8960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 11984 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1666464484
transform 1 0 12320 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_111
timestamp 1666464484
transform 1 0 12656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_115
timestamp 1666464484
transform 1 0 13104 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_117
timestamp 1666464484
transform 1 0 13328 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_144
timestamp 1666464484
transform 1 0 16352 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_2
timestamp 1666464484
transform 1 0 448 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_10
timestamp 1666464484
transform 1 0 1344 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_14
timestamp 1666464484
transform 1 0 1792 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_42
timestamp 1666464484
transform 1 0 4928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 8064 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1666464484
transform 1 0 8400 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_76
timestamp 1666464484
transform 1 0 8736 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_104
timestamp 1666464484
transform 1 0 11872 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_132
timestamp 1666464484
transform 1 0 15008 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_136
timestamp 1666464484
transform 1 0 15456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_138
timestamp 1666464484
transform 1 0 15680 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 16016 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1666464484
transform 1 0 16352 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1666464484
transform 1 0 448 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3472 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_33
timestamp 1666464484
transform 1 0 3920 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_37
timestamp 1666464484
transform 1 0 4368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_43
timestamp 1666464484
transform 1 0 5040 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_71
timestamp 1666464484
transform 1 0 8176 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_99
timestamp 1666464484
transform 1 0 11312 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_103
timestamp 1666464484
transform 1 0 11760 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 11984 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_108
timestamp 1666464484
transform 1 0 12320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_112
timestamp 1666464484
transform 1 0 12768 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_116
timestamp 1666464484
transform 1 0 13216 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_144
timestamp 1666464484
transform 1 0 16352 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_2
timestamp 1666464484
transform 1 0 448 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_10
timestamp 1666464484
transform 1 0 1344 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_38
timestamp 1666464484
transform 1 0 4480 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_42
timestamp 1666464484
transform 1 0 4928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_46
timestamp 1666464484
transform 1 0 5376 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_62
timestamp 1666464484
transform 1 0 7168 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1666464484
transform 1 0 8064 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1666464484
transform 1 0 8400 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_76 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 8736 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_108
timestamp 1666464484
transform 1 0 12320 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_112
timestamp 1666464484
transform 1 0 12768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_114
timestamp 1666464484
transform 1 0 12992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1666464484
transform 1 0 16016 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1666464484
transform 1 0 16352 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1666464484
transform 1 0 448 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_29
timestamp 1666464484
transform 1 0 3472 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_33
timestamp 1666464484
transform 1 0 3920 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1666464484
transform 1 0 4368 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_40
timestamp 1666464484
transform 1 0 4704 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_56
timestamp 1666464484
transform 1 0 6496 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_64
timestamp 1666464484
transform 1 0 7392 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_91
timestamp 1666464484
transform 1 0 10416 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_95
timestamp 1666464484
transform 1 0 10864 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1666464484
transform 1 0 11760 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 11984 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_108
timestamp 1666464484
transform 1 0 12320 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_116
timestamp 1666464484
transform 1 0 13216 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_144
timestamp 1666464484
transform 1 0 16352 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_2
timestamp 1666464484
transform 1 0 448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_6
timestamp 1666464484
transform 1 0 896 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_8
timestamp 1666464484
transform 1 0 1120 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_35
timestamp 1666464484
transform 1 0 4144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_39
timestamp 1666464484
transform 1 0 4592 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_42
timestamp 1666464484
transform 1 0 4928 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 8064 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_73
timestamp 1666464484
transform 1 0 8400 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_100
timestamp 1666464484
transform 1 0 11424 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_108
timestamp 1666464484
transform 1 0 12320 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_135
timestamp 1666464484
transform 1 0 15344 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_139
timestamp 1666464484
transform 1 0 15792 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 16016 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1666464484
transform 1 0 16352 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_2
timestamp 1666464484
transform 1 0 448 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_4
timestamp 1666464484
transform 1 0 672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_31
timestamp 1666464484
transform 1 0 3696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1666464484
transform 1 0 4368 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_40
timestamp 1666464484
transform 1 0 4704 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_56
timestamp 1666464484
transform 1 0 6496 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_59
timestamp 1666464484
transform 1 0 6832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_87
timestamp 1666464484
transform 1 0 9968 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_91
timestamp 1666464484
transform 1 0 10416 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_99
timestamp 1666464484
transform 1 0 11312 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_103
timestamp 1666464484
transform 1 0 11760 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 11984 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_108
timestamp 1666464484
transform 1 0 12320 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_111
timestamp 1666464484
transform 1 0 12656 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_139
timestamp 1666464484
transform 1 0 15792 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_141
timestamp 1666464484
transform 1 0 16016 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_144
timestamp 1666464484
transform 1 0 16352 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1666464484
transform 1 0 448 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_29
timestamp 1666464484
transform 1 0 3472 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_33
timestamp 1666464484
transform 1 0 3920 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_37
timestamp 1666464484
transform 1 0 4368 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_41
timestamp 1666464484
transform 1 0 4816 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1666464484
transform 1 0 7952 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_72
timestamp 1666464484
transform 1 0 8288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_99
timestamp 1666464484
transform 1 0 11312 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_103
timestamp 1666464484
transform 1 0 11760 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_107
timestamp 1666464484
transform 1 0 12208 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_111
timestamp 1666464484
transform 1 0 12656 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1666464484
transform 1 0 15792 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_142
timestamp 1666464484
transform 1 0 16128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1666464484
transform 1 0 16352 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 224 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 16688 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 224 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 16688 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 16688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 16688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 16688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 16688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 16688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 16688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 4144 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1666464484
transform 1 0 8064 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1666464484
transform 1 0 11984 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1666464484
transform 1 0 15904 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1666464484
transform 1 0 8176 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1666464484
transform 1 0 16128 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1666464484
transform 1 0 4144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1666464484
transform 1 0 12096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1666464484
transform 1 0 8176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1666464484
transform 1 0 16128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1666464484
transform 1 0 4144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1666464484
transform 1 0 12096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1666464484
transform 1 0 8176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1666464484
transform 1 0 16128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1666464484
transform 1 0 4144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1666464484
transform 1 0 12096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1666464484
transform 1 0 8176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1666464484
transform 1 0 16128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1666464484
transform 1 0 4144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1666464484
transform 1 0 12096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1666464484
transform 1 0 8176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1666464484
transform 1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1666464484
transform 1 0 4144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1666464484
transform 1 0 12096 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1666464484
transform 1 0 4144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1666464484
transform 1 0 8064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1666464484
transform 1 0 11984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1666464484
transform 1 0 15904 0 -1 10976
box -86 -86 310 870
<< labels >>
flabel metal4 s 2122 1508 2442 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 6238 1508 6558 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 10354 1508 10674 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 14470 1508 14790 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 4180 1508 4500 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 8296 1508 8616 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 12412 1508 12732 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 16528 1508 16848 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal2 s 560 0 672 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[0]
port 2 nsew signal input
flabel metal2 s 5040 0 5152 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[10]
port 3 nsew signal input
flabel metal2 s 5488 0 5600 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[11]
port 4 nsew signal input
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[12]
port 5 nsew signal input
flabel metal2 s 6384 0 6496 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[13]
port 6 nsew signal input
flabel metal2 s 6832 0 6944 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[14]
port 7 nsew signal input
flabel metal2 s 7280 0 7392 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[15]
port 8 nsew signal input
flabel metal2 s 7728 0 7840 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[16]
port 9 nsew signal input
flabel metal2 s 8176 0 8288 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[17]
port 10 nsew signal input
flabel metal2 s 1008 0 1120 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[1]
port 11 nsew signal input
flabel metal2 s 1456 0 1568 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[2]
port 12 nsew signal input
flabel metal2 s 1904 0 2016 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[3]
port 13 nsew signal input
flabel metal2 s 2352 0 2464 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[4]
port 14 nsew signal input
flabel metal2 s 2800 0 2912 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[5]
port 15 nsew signal input
flabel metal2 s 3248 0 3360 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[6]
port 16 nsew signal input
flabel metal2 s 3696 0 3808 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[7]
port 17 nsew signal input
flabel metal2 s 4144 0 4256 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[8]
port 18 nsew signal input
flabel metal2 s 4592 0 4704 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[9]
port 19 nsew signal input
flabel metal2 s 560 12200 672 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[0]
port 20 nsew signal tristate
flabel metal2 s 5040 12200 5152 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[10]
port 21 nsew signal tristate
flabel metal2 s 5488 12200 5600 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[11]
port 22 nsew signal tristate
flabel metal2 s 5936 12200 6048 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[12]
port 23 nsew signal tristate
flabel metal2 s 6384 12200 6496 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[13]
port 24 nsew signal tristate
flabel metal2 s 6832 12200 6944 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[14]
port 25 nsew signal tristate
flabel metal2 s 7280 12200 7392 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[15]
port 26 nsew signal tristate
flabel metal2 s 7728 12200 7840 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[16]
port 27 nsew signal tristate
flabel metal2 s 8176 12200 8288 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[17]
port 28 nsew signal tristate
flabel metal2 s 1008 12200 1120 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[1]
port 29 nsew signal tristate
flabel metal2 s 1456 12200 1568 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[2]
port 30 nsew signal tristate
flabel metal2 s 1904 12200 2016 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[3]
port 31 nsew signal tristate
flabel metal2 s 2352 12200 2464 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[4]
port 32 nsew signal tristate
flabel metal2 s 2800 12200 2912 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[5]
port 33 nsew signal tristate
flabel metal2 s 3248 12200 3360 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[6]
port 34 nsew signal tristate
flabel metal2 s 3696 12200 3808 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[7]
port 35 nsew signal tristate
flabel metal2 s 4144 12200 4256 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[8]
port 36 nsew signal tristate
flabel metal2 s 4592 12200 4704 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[9]
port 37 nsew signal tristate
flabel metal3 s 0 2128 800 2240 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[0]
port 38 nsew signal input
flabel metal3 s 0 6384 800 6496 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[1]
port 39 nsew signal input
flabel metal3 s 0 10640 800 10752 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[2]
port 40 nsew signal input
flabel metal3 s 16200 2128 17000 2240 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[0]
port 41 nsew signal tristate
flabel metal3 s 16200 6384 17000 6496 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[1]
port 42 nsew signal tristate
flabel metal3 s 16200 10640 17000 10752 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[2]
port 43 nsew signal tristate
flabel metal2 s 8624 12200 8736 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[0]
port 44 nsew signal input
flabel metal2 s 13104 12200 13216 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[10]
port 45 nsew signal input
flabel metal2 s 13552 12200 13664 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[11]
port 46 nsew signal input
flabel metal2 s 14000 12200 14112 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[12]
port 47 nsew signal input
flabel metal2 s 14448 12200 14560 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[13]
port 48 nsew signal input
flabel metal2 s 14896 12200 15008 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[14]
port 49 nsew signal input
flabel metal2 s 15344 12200 15456 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[15]
port 50 nsew signal input
flabel metal2 s 15792 12200 15904 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[16]
port 51 nsew signal input
flabel metal2 s 16240 12200 16352 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[17]
port 52 nsew signal input
flabel metal2 s 9072 12200 9184 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[1]
port 53 nsew signal input
flabel metal2 s 9520 12200 9632 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[2]
port 54 nsew signal input
flabel metal2 s 9968 12200 10080 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[3]
port 55 nsew signal input
flabel metal2 s 10416 12200 10528 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[4]
port 56 nsew signal input
flabel metal2 s 10864 12200 10976 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[5]
port 57 nsew signal input
flabel metal2 s 11312 12200 11424 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[6]
port 58 nsew signal input
flabel metal2 s 11760 12200 11872 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[7]
port 59 nsew signal input
flabel metal2 s 12208 12200 12320 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[8]
port 60 nsew signal input
flabel metal2 s 12656 12200 12768 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[9]
port 61 nsew signal input
flabel metal2 s 8624 0 8736 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[0]
port 62 nsew signal tristate
flabel metal2 s 13104 0 13216 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[10]
port 63 nsew signal tristate
flabel metal2 s 13552 0 13664 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[11]
port 64 nsew signal tristate
flabel metal2 s 14000 0 14112 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[12]
port 65 nsew signal tristate
flabel metal2 s 14448 0 14560 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[13]
port 66 nsew signal tristate
flabel metal2 s 14896 0 15008 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[14]
port 67 nsew signal tristate
flabel metal2 s 15344 0 15456 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[15]
port 68 nsew signal tristate
flabel metal2 s 15792 0 15904 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[16]
port 69 nsew signal tristate
flabel metal2 s 16240 0 16352 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[17]
port 70 nsew signal tristate
flabel metal2 s 9072 0 9184 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[1]
port 71 nsew signal tristate
flabel metal2 s 9520 0 9632 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[2]
port 72 nsew signal tristate
flabel metal2 s 9968 0 10080 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[3]
port 73 nsew signal tristate
flabel metal2 s 10416 0 10528 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[4]
port 74 nsew signal tristate
flabel metal2 s 10864 0 10976 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[5]
port 75 nsew signal tristate
flabel metal2 s 11312 0 11424 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[6]
port 76 nsew signal tristate
flabel metal2 s 11760 0 11872 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[7]
port 77 nsew signal tristate
flabel metal2 s 12208 0 12320 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[8]
port 78 nsew signal tristate
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[9]
port 79 nsew signal tristate
rlabel metal1 8456 10192 8456 10192 0 VDD
rlabel via1 8536 10976 8536 10976 0 VSS
rlabel metal2 2744 5880 2744 5880 0 mgmt_gpio_in[0]
rlabel metal3 4480 1960 4480 1960 0 mgmt_gpio_in[10]
rlabel metal2 6776 1904 6776 1904 0 mgmt_gpio_in[11]
rlabel metal2 6048 2408 6048 2408 0 mgmt_gpio_in[12]
rlabel metal2 7560 2464 7560 2464 0 mgmt_gpio_in[13]
rlabel metal2 6888 2058 6888 2058 0 mgmt_gpio_in[14]
rlabel metal2 7336 1638 7336 1638 0 mgmt_gpio_in[15]
rlabel metal2 8568 7000 8568 7000 0 mgmt_gpio_in[16]
rlabel metal2 9240 9744 9240 9744 0 mgmt_gpio_in[17]
rlabel metal2 1064 2534 1064 2534 0 mgmt_gpio_in[1]
rlabel metal3 2128 8232 2128 8232 0 mgmt_gpio_in[2]
rlabel metal2 2968 9632 2968 9632 0 mgmt_gpio_in[3]
rlabel metal2 2520 3864 2520 3864 0 mgmt_gpio_in[4]
rlabel metal2 2856 3710 2856 3710 0 mgmt_gpio_in[5]
rlabel metal2 3304 3038 3304 3038 0 mgmt_gpio_in[6]
rlabel metal2 4312 2632 4312 2632 0 mgmt_gpio_in[7]
rlabel metal2 4032 3080 4032 3080 0 mgmt_gpio_in[8]
rlabel metal2 4648 2058 4648 2058 0 mgmt_gpio_in[9]
rlabel metal2 952 7588 952 7588 0 mgmt_gpio_in_buf[0]
rlabel metal3 3920 3304 3920 3304 0 mgmt_gpio_in_buf[10]
rlabel metal2 5544 7154 5544 7154 0 mgmt_gpio_in_buf[11]
rlabel metal2 5880 7448 5880 7448 0 mgmt_gpio_in_buf[12]
rlabel metal2 6216 10360 6216 10360 0 mgmt_gpio_in_buf[13]
rlabel metal2 6664 7056 6664 7056 0 mgmt_gpio_in_buf[14]
rlabel metal2 6664 10864 6664 10864 0 mgmt_gpio_in_buf[15]
rlabel metal2 10136 8624 10136 8624 0 mgmt_gpio_in_buf[16]
rlabel metal2 8232 11074 8232 11074 0 mgmt_gpio_in_buf[17]
rlabel metal2 1064 11354 1064 11354 0 mgmt_gpio_in_buf[1]
rlabel metal2 1456 10696 1456 10696 0 mgmt_gpio_in_buf[2]
rlabel metal2 1960 11074 1960 11074 0 mgmt_gpio_in_buf[3]
rlabel metal2 2520 9744 2520 9744 0 mgmt_gpio_in_buf[4]
rlabel metal2 2856 9786 2856 9786 0 mgmt_gpio_in_buf[5]
rlabel metal2 3304 9002 3304 9002 0 mgmt_gpio_in_buf[6]
rlabel metal2 3696 10696 3696 10696 0 mgmt_gpio_in_buf[7]
rlabel metal2 5768 6776 5768 6776 0 mgmt_gpio_in_buf[8]
rlabel metal2 3192 5152 3192 5152 0 mgmt_gpio_in_buf[9]
rlabel metal3 2814 2184 2814 2184 0 mgmt_gpio_oeb[0]
rlabel metal3 5152 6552 5152 6552 0 mgmt_gpio_oeb[1]
rlabel metal2 4760 9968 4760 9968 0 mgmt_gpio_oeb[2]
rlabel metal3 14210 2184 14210 2184 0 mgmt_gpio_oeb_buf[0]
rlabel metal2 7224 6496 7224 6496 0 mgmt_gpio_oeb_buf[1]
rlabel metal2 11816 9800 11816 9800 0 mgmt_gpio_oeb_buf[2]
rlabel metal3 9296 8232 9296 8232 0 mgmt_gpio_out[0]
rlabel metal3 15204 6104 15204 6104 0 mgmt_gpio_out[10]
rlabel metal3 14168 9016 14168 9016 0 mgmt_gpio_out[11]
rlabel metal3 13720 9800 13720 9800 0 mgmt_gpio_out[12]
rlabel metal2 13384 10864 13384 10864 0 mgmt_gpio_out[13]
rlabel metal2 16184 9072 16184 9072 0 mgmt_gpio_out[14]
rlabel metal2 15512 6552 15512 6552 0 mgmt_gpio_out[15]
rlabel metal2 15736 6048 15736 6048 0 mgmt_gpio_out[16]
rlabel metal2 16184 6552 16184 6552 0 mgmt_gpio_out[17]
rlabel metal2 10584 10864 10584 10864 0 mgmt_gpio_out[1]
rlabel metal2 10808 6944 10808 6944 0 mgmt_gpio_out[2]
rlabel metal3 10584 5880 10584 5880 0 mgmt_gpio_out[3]
rlabel metal2 11256 7728 11256 7728 0 mgmt_gpio_out[4]
rlabel metal2 11816 5208 11816 5208 0 mgmt_gpio_out[5]
rlabel metal2 11760 2072 11760 2072 0 mgmt_gpio_out[6]
rlabel metal2 13944 5656 13944 5656 0 mgmt_gpio_out[7]
rlabel metal2 12488 2464 12488 2464 0 mgmt_gpio_out[8]
rlabel metal3 13776 3528 13776 3528 0 mgmt_gpio_out[9]
rlabel metal2 8680 4550 8680 4550 0 mgmt_gpio_out_buf[0]
rlabel metal2 13160 1638 13160 1638 0 mgmt_gpio_out_buf[10]
rlabel metal2 13608 4830 13608 4830 0 mgmt_gpio_out_buf[11]
rlabel metal2 14112 6888 14112 6888 0 mgmt_gpio_out_buf[12]
rlabel metal2 14504 1470 14504 1470 0 mgmt_gpio_out_buf[13]
rlabel metal2 14952 2310 14952 2310 0 mgmt_gpio_out_buf[14]
rlabel metal2 15400 2926 15400 2926 0 mgmt_gpio_out_buf[15]
rlabel metal2 15848 2422 15848 2422 0 mgmt_gpio_out_buf[16]
rlabel metal2 16296 2086 16296 2086 0 mgmt_gpio_out_buf[17]
rlabel metal2 9128 5614 9128 5614 0 mgmt_gpio_out_buf[1]
rlabel metal2 9576 3766 9576 3766 0 mgmt_gpio_out_buf[2]
rlabel metal2 10024 1806 10024 1806 0 mgmt_gpio_out_buf[3]
rlabel metal2 10472 1470 10472 1470 0 mgmt_gpio_out_buf[4]
rlabel metal2 10920 1694 10920 1694 0 mgmt_gpio_out_buf[5]
rlabel metal2 11368 1022 11368 1022 0 mgmt_gpio_out_buf[6]
rlabel metal2 11816 1134 11816 1134 0 mgmt_gpio_out_buf[7]
rlabel metal2 12264 1414 12264 1414 0 mgmt_gpio_out_buf[8]
rlabel metal2 12712 1078 12712 1078 0 mgmt_gpio_out_buf[9]
<< properties >>
string FIXED_BBOX 0 0 17000 13000
<< end >>
