* NGSPICE file created from caravel.ext - technology: gf180mcuC

* Black-box entry subcircuit for gpio_control_block abstract view
.subckt gpio_control_block VDD VSS gpio_defaults[0] gpio_defaults[1] gpio_defaults[2]
+ gpio_defaults[3] gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_drive_sel[0]
+ pad_gpio_drive_sel[1] pad_gpio_in pad_gpio_inen pad_gpio_out pad_gpio_outen pad_gpio_pulldown_sel
+ pad_gpio_pullup_sel pad_gpio_schmitt_sel pad_gpio_slew_sel resetn resetn_out serial_clock
+ serial_clock_out serial_data_in serial_data_out serial_load serial_load_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero
.ends

* Black-box entry subcircuit for gpio_defaults_block abstract view
.subckt gpio_defaults_block gpio_defaults[0] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3]
+ gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8]
+ gpio_defaults[9] VDD VSS
.ends

* Black-box entry subcircuit for digital_pll abstract view
.subckt digital_pll VDD VSS clockp[0] clockp[1] dco div[0] div[1] div[2] div[3] div[4]
+ enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__fill10 abstract view
.subckt gf180mcu_fd_io__fill10 DVDD DVSS VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__in_s abstract view
.subckt gf180mcu_fd_io__in_s DVDD DVSS PAD PD PU VDD VSS Y
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__dvss abstract view
.subckt gf180mcu_fd_io__dvss DVDD DVSS VDD
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__dvdd abstract view
.subckt gf180mcu_fd_io__dvdd DVDD DVSS VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__fill5 abstract view
.subckt gf180mcu_fd_io__fill5 DVDD DVSS VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__bi_t abstract view
.subckt gf180mcu_fd_io__bi_t A CS DVDD DVSS IE OE PAD PD PDRV0 PDRV1 PU SL VDD VSS Y
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__in_c abstract view
.subckt gf180mcu_fd_io__in_c DVDD DVSS PAD PD PU VDD VSS Y
.ends

* Black-box entry subcircuit for gf180mcu_fd_io__cor abstract view
.subckt gf180mcu_fd_io__cor DVDD DVSS VDD VSS
.ends

.subckt chip_io clock clock_core flash_clk flash_clk_core flash_clk_oe_core flash_csb
+ flash_csb_core flash_csb_oe_core flash_io0 flash_io0_di_core flash_io0_do_core flash_io0_ie_core
+ flash_io0_oe_core flash_io1 flash_io1_di_core flash_io1_do_core flash_io1_ie_core
+ flash_io1_oe_core gpio gpio_drive_select_core[0] gpio_drive_select_core[1] gpio_in_core
+ gpio_inen_core gpio_out_core gpio_outen_core gpio_pd_select gpio_pu_select gpio_schmitt_select
+ gpio_slew_select mprj_io[0] mprj_io[10] mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14]
+ mprj_io[15] mprj_io[16] mprj_io[17] mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20]
+ mprj_io[21] mprj_io[22] mprj_io[23] mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27]
+ mprj_io[28] mprj_io[29] mprj_io[2] mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33]
+ mprj_io[34] mprj_io[35] mprj_io[36] mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5]
+ mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9] mprj_io_drive_sel[0] mprj_io_drive_sel[10]
+ mprj_io_drive_sel[11] mprj_io_drive_sel[12] mprj_io_drive_sel[13] mprj_io_drive_sel[14]
+ mprj_io_drive_sel[15] mprj_io_drive_sel[16] mprj_io_drive_sel[17] mprj_io_drive_sel[18]
+ mprj_io_drive_sel[19] mprj_io_drive_sel[1] mprj_io_drive_sel[20] mprj_io_drive_sel[21]
+ mprj_io_drive_sel[22] mprj_io_drive_sel[23] mprj_io_drive_sel[24] mprj_io_drive_sel[25]
+ mprj_io_drive_sel[26] mprj_io_drive_sel[27] mprj_io_drive_sel[28] mprj_io_drive_sel[29]
+ mprj_io_drive_sel[2] mprj_io_drive_sel[30] mprj_io_drive_sel[31] mprj_io_drive_sel[32]
+ mprj_io_drive_sel[33] mprj_io_drive_sel[34] mprj_io_drive_sel[35] mprj_io_drive_sel[36]
+ mprj_io_drive_sel[37] mprj_io_drive_sel[38] mprj_io_drive_sel[39] mprj_io_drive_sel[3]
+ mprj_io_drive_sel[40] mprj_io_drive_sel[41] mprj_io_drive_sel[42] mprj_io_drive_sel[43]
+ mprj_io_drive_sel[44] mprj_io_drive_sel[45] mprj_io_drive_sel[46] mprj_io_drive_sel[47]
+ mprj_io_drive_sel[48] mprj_io_drive_sel[49] mprj_io_drive_sel[4] mprj_io_drive_sel[51]
+ mprj_io_drive_sel[525] mprj_io_drive_sel[52] mprj_io_drive_sel[53] mprj_io_drive_sel[54]
+ mprj_io_drive_sel[55] mprj_io_drive_sel[56] mprj_io_drive_sel[57] mprj_io_drive_sel[58]
+ mprj_io_drive_sel[59] mprj_io_drive_sel[5] mprj_io_drive_sel[61] mprj_io_drive_sel[62]
+ mprj_io_drive_sel[63] mprj_io_drive_sel[64] mprj_io_drive_sel[65] mprj_io_drive_sel[66]
+ mprj_io_drive_sel[67] mprj_io_drive_sel[68] mprj_io_drive_sel[69] mprj_io_drive_sel[6]
+ mprj_io_drive_sel[70] mprj_io_drive_sel[71] mprj_io_drive_sel[72] mprj_io_drive_sel[73]
+ mprj_io_drive_sel[74] mprj_io_drive_sel[75] mprj_io_drive_sel[7] mprj_io_drive_sel[8]
+ mprj_io_drive_sel[9] mprj_io_in[0] mprj_io_in[10] mprj_io_in[11] mprj_io_in[12]
+ mprj_io_in[13] mprj_io_in[14] mprj_io_in[15] mprj_io_in[16] mprj_io_in[17] mprj_io_in[18]
+ mprj_io_in[19] mprj_io_in[1] mprj_io_in[20] mprj_io_in[21] mprj_io_in[22] mprj_io_in[23]
+ mprj_io_in[24] mprj_io_in[25] mprj_io_in[26] mprj_io_in[27] mprj_io_in[28] mprj_io_in[29]
+ mprj_io_in[2] mprj_io_in[30] mprj_io_in[31] mprj_io_in[32] mprj_io_in[33] mprj_io_in[34]
+ mprj_io_in[35] mprj_io_in[36] mprj_io_in[37] mprj_io_in[3] mprj_io_in[4] mprj_io_in[5]
+ mprj_io_in[6] mprj_io_in[7] mprj_io_in[8] mprj_io_in[9] mprj_io_inen[0] mprj_io_inen[10]
+ mprj_io_inen[11] mprj_io_inen[12] mprj_io_inen[13] mprj_io_inen[14] mprj_io_inen[15]
+ mprj_io_inen[16] mprj_io_inen[17] mprj_io_inen[18] mprj_io_inen[19] mprj_io_inen[1]
+ mprj_io_inen[20] mprj_io_inen[21] mprj_io_inen[22] mprj_io_inen[23] mprj_io_inen[24]
+ mprj_io_inen[25] mprj_io_inen[26] mprj_io_inen[27] mprj_io_inen[28] mprj_io_inen[29]
+ mprj_io_inen[2] mprj_io_inen[30] mprj_io_inen[31] mprj_io_inen[32] mprj_io_inen[33]
+ mprj_io_inen[34] mprj_io_inen[35] mprj_io_inen[36] mprj_io_inen[37] mprj_io_inen[3]
+ mprj_io_inen[4] mprj_io_inen[5] mprj_io_inen[6] mprj_io_inen[7] mprj_io_inen[8]
+ mprj_io_inen[9] mprj_io_out[0] mprj_io_out[10] mprj_io_out[11] mprj_io_out[12] mprj_io_out[13]
+ mprj_io_out[14] mprj_io_out[15] mprj_io_out[16] mprj_io_out[17] mprj_io_out[18]
+ mprj_io_out[19] mprj_io_out[1] mprj_io_out[20] mprj_io_out[21] mprj_io_out[22] mprj_io_out[23]
+ mprj_io_out[24] mprj_io_out[25] mprj_io_out[26] mprj_io_out[27] mprj_io_out[28]
+ mprj_io_out[29] mprj_io_out[2] mprj_io_out[30] mprj_io_out[31] mprj_io_out[32] mprj_io_out[33]
+ mprj_io_out[34] mprj_io_out[35] mprj_io_out[36] mprj_io_out[37] mprj_io_out[3] mprj_io_out[4]
+ mprj_io_out[5] mprj_io_out[6] mprj_io_out[7] mprj_io_out[8] mprj_io_out[9] mprj_io_outen[0]
+ mprj_io_outen[10] mprj_io_outen[11] mprj_io_outen[12] mprj_io_outen[13] mprj_io_outen[14]
+ mprj_io_outen[15] mprj_io_outen[16] mprj_io_outen[17] mprj_io_outen[18] mprj_io_outen[19]
+ mprj_io_outen[1] mprj_io_outen[20] mprj_io_outen[21] mprj_io_outen[22] mprj_io_outen[23]
+ mprj_io_outen[24] mprj_io_outen[25] mprj_io_outen[26] mprj_io_outen[27] mprj_io_outen[28]
+ mprj_io_outen[29] mprj_io_outen[2] mprj_io_outen[30] mprj_io_outen[31] mprj_io_outen[32]
+ mprj_io_outen[33] mprj_io_outen[34] mprj_io_outen[35] mprj_io_outen[36] mprj_io_outen[37]
+ mprj_io_outen[3] mprj_io_outen[4] mprj_io_outen[5] mprj_io_outen[6] mprj_io_outen[7]
+ mprj_io_outen[8] mprj_io_outen[9] mprj_io_pd_select[0] mprj_io_pd_select[10] mprj_io_pd_select[11]
+ mprj_io_pd_select[12] mprj_io_pd_select[13] mprj_io_pd_select[14] mprj_io_pd_select[15]
+ mprj_io_pd_select[16] mprj_io_pd_select[17] mprj_io_pd_select[18] mprj_io_pd_select[19]
+ mprj_io_pd_select[1] mprj_io_pd_select[20] mprj_io_pd_select[21] mprj_io_pd_select[22]
+ mprj_io_pd_select[23] mprj_io_pd_select[24] mprj_io_pd_select[25] mprj_io_pd_select[26]
+ mprj_io_pd_select[27] mprj_io_pd_select[28] mprj_io_pd_select[29] mprj_io_pd_select[2]
+ mprj_io_pd_select[30] mprj_io_pd_select[31] mprj_io_pd_select[32] mprj_io_pd_select[33]
+ mprj_io_pd_select[34] mprj_io_pd_select[35] mprj_io_pd_select[36] mprj_io_pd_select[37]
+ mprj_io_pd_select[3] mprj_io_pd_select[4] mprj_io_pd_select[5] mprj_io_pd_select[6]
+ mprj_io_pd_select[7] mprj_io_pd_select[8] mprj_io_pd_select[9] mprj_io_pu_select[0]
+ mprj_io_pu_select[10] mprj_io_pu_select[11] mprj_io_pu_select[12] mprj_io_pu_select[13]
+ mprj_io_pu_select[14] mprj_io_pu_select[15] mprj_io_pu_select[16] mprj_io_pu_select[17]
+ mprj_io_pu_select[18] mprj_io_pu_select[19] mprj_io_pu_select[1] mprj_io_pu_select[20]
+ mprj_io_pu_select[21] mprj_io_pu_select[22] mprj_io_pu_select[23] mprj_io_pu_select[24]
+ mprj_io_pu_select[25] mprj_io_pu_select[26] mprj_io_pu_select[27] mprj_io_pu_select[28]
+ mprj_io_pu_select[29] mprj_io_pu_select[2] mprj_io_pu_select[30] mprj_io_pu_select[31]
+ mprj_io_pu_select[32] mprj_io_pu_select[33] mprj_io_pu_select[34] mprj_io_pu_select[35]
+ mprj_io_pu_select[36] mprj_io_pu_select[37] mprj_io_pu_select[3] mprj_io_pu_select[4]
+ mprj_io_pu_select[5] mprj_io_pu_select[6] mprj_io_pu_select[7] mprj_io_pu_select[8]
+ mprj_io_pu_select[9] mprj_io_schmitt_select[0] mprj_io_schmitt_select[10] mprj_io_schmitt_select[11]
+ mprj_io_schmitt_select[12] mprj_io_schmitt_select[13] mprj_io_schmitt_select[14]
+ mprj_io_schmitt_select[15] mprj_io_schmitt_select[16] mprj_io_schmitt_select[17]
+ mprj_io_schmitt_select[18] mprj_io_schmitt_select[19] mprj_io_schmitt_select[1]
+ mprj_io_schmitt_select[20] mprj_io_schmitt_select[21] mprj_io_schmitt_select[22]
+ mprj_io_schmitt_select[23] mprj_io_schmitt_select[24] mprj_io_schmitt_select[25]
+ mprj_io_schmitt_select[26] mprj_io_schmitt_select[27] mprj_io_schmitt_select[28]
+ mprj_io_schmitt_select[29] mprj_io_schmitt_select[2] mprj_io_schmitt_select[30]
+ mprj_io_schmitt_select[31] mprj_io_schmitt_select[32] mprj_io_schmitt_select[33]
+ mprj_io_schmitt_select[34] mprj_io_schmitt_select[35] mprj_io_schmitt_select[36]
+ mprj_io_schmitt_select[37] mprj_io_schmitt_select[3] mprj_io_schmitt_select[4] mprj_io_schmitt_select[5]
+ mprj_io_schmitt_select[6] mprj_io_schmitt_select[7] mprj_io_schmitt_select[8] mprj_io_schmitt_select[9]
+ mprj_io_slew_select[0] mprj_io_slew_select[10] mprj_io_slew_select[11] mprj_io_slew_select[12]
+ mprj_io_slew_select[13] mprj_io_slew_select[14] mprj_io_slew_select[15] mprj_io_slew_select[16]
+ mprj_io_slew_select[17] mprj_io_slew_select[18] mprj_io_slew_select[19] mprj_io_slew_select[1]
+ mprj_io_slew_select[20] mprj_io_slew_select[21] mprj_io_slew_select[22] mprj_io_slew_select[23]
+ mprj_io_slew_select[24] mprj_io_slew_select[25] mprj_io_slew_select[26] mprj_io_slew_select[27]
+ mprj_io_slew_select[28] mprj_io_slew_select[29] mprj_io_slew_select[2] mprj_io_slew_select[30]
+ mprj_io_slew_select[31] mprj_io_slew_select[32] mprj_io_slew_select[33] mprj_io_slew_select[34]
+ mprj_io_slew_select[35] mprj_io_slew_select[36] mprj_io_slew_select[37] mprj_io_slew_select[3]
+ mprj_io_slew_select[4] mprj_io_slew_select[5] mprj_io_slew_select[6] mprj_io_slew_select[7]
+ mprj_io_slew_select[8] mprj_io_slew_select[9] resetb resetb_core vdd vss gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__cor_3/VDD
Xgf180mcu_fd_io__fill10_513 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_524 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_535 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_546 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_557 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_568 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_579 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_502 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_94 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_83 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_72 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_61 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_50 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_398 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_387 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_376 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_365 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_354 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_343 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_332 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_321 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_310 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_140 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_151 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_162 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_173 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_184 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_195 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_909 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_706 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_717 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_728 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_739 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_514 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_525 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_536 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_547 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_558 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_569 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_503 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_95 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_84 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_73 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_62 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_51 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_40 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_399 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_388 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_377 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_366 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_355 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_344 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_333 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_322 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_311 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_300 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_130 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_141 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_152 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_163 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_174 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_185 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_196 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_707 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_718 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_729 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_515 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_526 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_537 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_504 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_548 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_559 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_96 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_85 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_74 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_63 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_52 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_41 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_30 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_389 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_378 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_367 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_356 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_345 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_334 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_323 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_312 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_301 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_890 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_120 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_131 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_142 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_153 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_164 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_175 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_186 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_197 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_708 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_719 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_516 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_527 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_538 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_549 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_505 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_97 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_86 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_75 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_64 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_53 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_42 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_31 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_20 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_379 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_368 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_357 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_346 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_335 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_324 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_313 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_302 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_880 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_891 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_110 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_121 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_132 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_143 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_154 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_165 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_176 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_187 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_198 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_709 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_517 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_528 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_539 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_506 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_87 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_65 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_76 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_54 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_43 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_32 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_21 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_10 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_98 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_303 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_369 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_358 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_347 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_336 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_325 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_314 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_870 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_881 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_892 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__in_s_0 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS resetb gf180mcu_fd_io__in_s_0/PD gf180mcu_fd_io__in_s_0/PU
+ gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS resetb_core gf180mcu_fd_io__in_s
Xgf180mcu_fd_io__fill10_100 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_111 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_122 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_133 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_144 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_155 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_166 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_177 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_188 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_199 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvss_0 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_518 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_529 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_507 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_44 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_33 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_22 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_11 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_66 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_77 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_55 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_88 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_99 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_359 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_348 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_337 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_326 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_315 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_304 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_860 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_882 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_893 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_871 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_101 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_112 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_123 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_134 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_145 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_156 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_167 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_178 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_690 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_189 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvss_1 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_519 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_508 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_67 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_45 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_56 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_34 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_23 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_12 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_78 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_89 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_349 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_338 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_327 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_316 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_305 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_850 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_861 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_872 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_883 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_894 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_102 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_113 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_124 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_135 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_146 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_157 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_168 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_179 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_680 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_691 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvss_2 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_509 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_68 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_46 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_57 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_35 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_24 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_13 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_79 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_339 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_328 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_317 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_306 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_840 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_851 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_862 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_873 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_884 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_895 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_0 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_103 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_114 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_125 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_136 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_147 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_158 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_169 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_670 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_681 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_692 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill5_0 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill5
Xgf180mcu_fd_io__dvss_3 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_69 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_58 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_47 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_36 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_25 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_14 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_329 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_318 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_307 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_830 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_841 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_852 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_863 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_874 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_885 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_896 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_1 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_104 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_115 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_126 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_137 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_148 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_159 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_660 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_671 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_682 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_693 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill5_1 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill5
Xgf180mcu_fd_io__fill10_490 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvss_4 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_59 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_48 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_37 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_26 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_15 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_319 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_308 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_820 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_831 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_842 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_853 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_864 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_875 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_2 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_897 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_886 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_105 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_116 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_127 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_138 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_149 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_650 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_661 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_672 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_683 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_694 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill5_2 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill5
Xgf180mcu_fd_io__fill10_491 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_480 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_0 flash_csb_core gf180mcu_fd_io__bi_t_0/CS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__bi_t_0/IE
+ flash_csb_oe_core flash_csb gf180mcu_fd_io__bi_t_0/PD gf180mcu_fd_io__bi_t_0/PDRV0 gf180mcu_fd_io__bi_t_0/PDRV1
+ gf180mcu_fd_io__bi_t_0/PU gf180mcu_fd_io__bi_t_0/SL gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__bi_t_0/Y gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__dvss_5 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_49 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_38 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_27 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_16 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_309 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_810 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_821 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_832 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_843 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_854 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_865 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_876 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_887 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_898 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_3 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_106 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_117 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_128 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_139 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_640 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_651 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_662 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_673 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_684 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_695 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_492 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_481 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_470 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_1 flash_clk_core gf180mcu_fd_io__bi_t_1/CS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__bi_t_1/IE
+ flash_clk_oe_core flash_clk gf180mcu_fd_io__bi_t_1/PD gf180mcu_fd_io__bi_t_1/PDRV0 gf180mcu_fd_io__bi_t_1/PDRV1
+ gf180mcu_fd_io__bi_t_1/PU gf180mcu_fd_io__bi_t_1/SL gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__bi_t_1/Y gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__dvss_6 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_39 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_28 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_17 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_811 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_822 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_833 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_844 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_855 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_866 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_877 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_888 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_899 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_800 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_4 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_630 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_107 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_118 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_129 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_641 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_652 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_663 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_674 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_685 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_696 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_493 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_482 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_471 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_460 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_2 flash_io0_do_core gf180mcu_fd_io__bi_t_2/CS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS flash_io0_ie_core
+ flash_io0_oe_core flash_io0 gf180mcu_fd_io__bi_t_2/PD gf180mcu_fd_io__bi_t_2/PDRV0 gf180mcu_fd_io__bi_t_2/PDRV1
+ gf180mcu_fd_io__bi_t_2/PU gf180mcu_fd_io__bi_t_2/SL gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS flash_io0_di_core
+ gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_290 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_29 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_18 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_801 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_812 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_823 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_834 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_845 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_867 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_878 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_889 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_856 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_5 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_108 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_119 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_620 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_631 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_642 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_653 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_664 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_675 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_686 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_697 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_494 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_483 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_472 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_461 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_450 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_3 flash_io1_do_core gf180mcu_fd_io__bi_t_3/CS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS flash_io1_ie_core
+ flash_io1_oe_core flash_io1 gf180mcu_fd_io__bi_t_3/PD gf180mcu_fd_io__bi_t_3/PDRV0 gf180mcu_fd_io__bi_t_3/PDRV1
+ gf180mcu_fd_io__bi_t_3/PU gf180mcu_fd_io__bi_t_3/SL gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS flash_io1_di_core
+ gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__dvss_8 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_280 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_291 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_19 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_802 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_813 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_824 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_835 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_846 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_857 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_868 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_879 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_109 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_610 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_621 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_632 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_643 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_654 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_665 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_676 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_687 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_698 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_495 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_484 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_473 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_462 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_451 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_440 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_4 gpio_out_core gpio_schmitt_select gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gpio_inen_core
+ gpio_outen_core gpio gpio_pd_select gpio_drive_select_core[0] gpio_drive_select_core[1]
+ gpio_pu_select gpio_slew_select gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gpio_in_core gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__dvss_9 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__dvss
Xgf180mcu_fd_io__fill10_292 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_270 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_281 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1040 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_803 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_814 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_825 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_836 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_858 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_869 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_847 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_7 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_600 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_611 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_622 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_633 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_644 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_655 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_666 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_677 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_688 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_699 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_496 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_485 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_474 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_463 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_452 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_441 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_430 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_5 mprj_io_out[0] mprj_io_schmitt_select[0] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[0] mprj_io_outen[0] mprj_io[0] mprj_io_pd_select[0] mprj_io_drive_sel[0]
+ mprj_io_drive_sel[1] mprj_io_pu_select[0] mprj_io_slew_select[0] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[0] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_260 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_271 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_282 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_293 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1041 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1030 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_8 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_804 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_815 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_826 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_837 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_848 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_859 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_601 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_612 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_623 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_634 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_645 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_656 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_667 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_678 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_689 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_497 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_486 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_475 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_464 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_453 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_442 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_431 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_420 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_6 mprj_io_out[1] mprj_io_schmitt_select[1] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[1] mprj_io_outen[1] mprj_io[1] mprj_io_pd_select[1] mprj_io_drive_sel[2]
+ mprj_io_drive_sel[3] mprj_io_pu_select[1] mprj_io_slew_select[1] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[1] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_294 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1042 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_250 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1031 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1020 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_261 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_272 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_283 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_805 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_816 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_838 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_849 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_827 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__dvdd_9 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__dvdd
Xgf180mcu_fd_io__fill10_602 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_613 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_624 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_635 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_646 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_657 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_668 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_679 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_498 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_487 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_476 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_465 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_454 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_443 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_432 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_421 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_410 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_7 mprj_io_out[2] mprj_io_schmitt_select[2] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[2] mprj_io_outen[2] mprj_io[2] mprj_io_pd_select[2] mprj_io_drive_sel[5]
+ mprj_io_drive_sel[4] mprj_io_pu_select[2] mprj_io_slew_select[2] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[2] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_295 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_240 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_251 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1010 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_262 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_273 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_284 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_0 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1043 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1032 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1021 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_806 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_817 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_828 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_839 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_603 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_614 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_625 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_636 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_647 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_658 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_669 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_499 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_488 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_477 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_466 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_455 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_444 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_433 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_422 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_411 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_400 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_8 mprj_io_out[3] mprj_io_schmitt_select[3] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[3] mprj_io_outen[3] mprj_io[3] mprj_io_pd_select[3] mprj_io_drive_sel[7]
+ mprj_io_drive_sel[6] mprj_io_pu_select[3] mprj_io_slew_select[3] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[3] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_296 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_230 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_241 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_252 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_263 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_274 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_285 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1044 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1033 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1022 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1011 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1000 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_807 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_829 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_818 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_604 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_615 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_626 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_637 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_648 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_659 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_412 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_401 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_489 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_478 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_467 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_456 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_445 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_434 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_423 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_9 mprj_io_out[4] mprj_io_schmitt_select[4] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[4] mprj_io_outen[4] mprj_io[4] mprj_io_pd_select[4] mprj_io_drive_sel[9]
+ mprj_io_drive_sel[8] mprj_io_pu_select[4] mprj_io_slew_select[4] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[4] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_990 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_297 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_220 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_231 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_242 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_253 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_264 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_275 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_286 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_2 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1045 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1034 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1001 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_808 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_819 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_605 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_616 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_627 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_638 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_649 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_479 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_468 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_457 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_446 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_435 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_424 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_413 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_402 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_980 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_991 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_210 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_221 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_232 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_243 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_254 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_265 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_276 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_287 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_298 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_3 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1046 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1035 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1024 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1013 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1002 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_809 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_606 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_617 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_628 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_639 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_469 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_458 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_447 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_436 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_425 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_414 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_403 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_970 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_981 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_992 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_40 mprj_io_out[33] mprj_io_schmitt_select[33] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[33] mprj_io_outen[33] mprj_io[33] mprj_io_pd_select[33] mprj_io_drive_sel[66]
+ mprj_io_drive_sel[67] mprj_io_pu_select[33] mprj_io_slew_select[33] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[33] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_299 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1047 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_200 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_211 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_222 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_233 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_244 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_255 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1036 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1025 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1014 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_266 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_277 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1003 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_288 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_4 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_607 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_618 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_629 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_459 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_448 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_437 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_426 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_415 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_404 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_960 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_971 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_982 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_993 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_30 mprj_io_out[28] mprj_io_schmitt_select[28] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[28] mprj_io_outen[28] mprj_io[28] mprj_io_pd_select[28] mprj_io_drive_sel[56]
+ mprj_io_drive_sel[57] mprj_io_pu_select[28] mprj_io_slew_select[28] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[28] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_41 mprj_io_out[34] mprj_io_schmitt_select[34] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[34] mprj_io_outen[34] mprj_io[34] mprj_io_pd_select[34] mprj_io_drive_sel[68]
+ mprj_io_drive_sel[69] mprj_io_pu_select[34] mprj_io_slew_select[34] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[34] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_289 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_201 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_212 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_223 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_234 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_245 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_256 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1026 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1015 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_267 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_278 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1004 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_790 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_5 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_608 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_619 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_449 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_438 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_427 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_416 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_405 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_950 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_961 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_972 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_983 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_994 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_20 mprj_io_out[13] mprj_io_schmitt_select[13] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[13] mprj_io_outen[13] mprj_io[12] mprj_io_pd_select[13] mprj_io_drive_sel[26]
+ mprj_io_drive_sel[27] mprj_io_pu_select[13] mprj_io_slew_select[13] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[13] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_31 mprj_io_out[29] mprj_io_schmitt_select[29] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[29] mprj_io_outen[29] mprj_io[29] mprj_io_pd_select[29] mprj_io_drive_sel[58]
+ mprj_io_drive_sel[59] mprj_io_pu_select[29] mprj_io_slew_select[29] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[29] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_42 mprj_io_out[36] mprj_io_schmitt_select[36] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[36] mprj_io_outen[36] mprj_io[36] mprj_io_pd_select[36] mprj_io_drive_sel[72]
+ mprj_io_drive_sel[73] mprj_io_pu_select[36] mprj_io_slew_select[36] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[36] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_202 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_213 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_224 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_235 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_246 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_257 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_268 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_279 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_780 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_791 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_6 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1038 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1027 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1016 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1005 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_609 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_428 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_417 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_406 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_439 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_940 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_951 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_962 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_973 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_21 mprj_io_out[20] mprj_io_schmitt_select[20] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[20] mprj_io_outen[20] mprj_io[20] mprj_io_pd_select[20] mprj_io_drive_sel[40]
+ mprj_io_drive_sel[41] mprj_io_pu_select[20] mprj_io_slew_select[20] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[20] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_32 mprj_io_out[30] mprj_io_schmitt_select[30] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[30] mprj_io_outen[30] mprj_io[30] mprj_io_pd_select[30] mprj_io_drive_sel[63]
+ mprj_io_drive_sel[61] mprj_io_pu_select[30] mprj_io_slew_select[30] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[30] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_10 mprj_io_out[5] mprj_io_schmitt_select[5] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[5] mprj_io_outen[5] mprj_io[5] mprj_io_pd_select[5] mprj_io_drive_sel[11]
+ mprj_io_drive_sel[10] mprj_io_pu_select[5] mprj_io_slew_select[5] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[5] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_995 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_203 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_214 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_225 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_236 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_247 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_258 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_269 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_770 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_781 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_792 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_7 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1039 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1028 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1017 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1006 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_429 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_418 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_407 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_22 mprj_io_out[12] mprj_io_schmitt_select[12] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[12] mprj_io_outen[12] mprj_io[13] mprj_io_pd_select[12] mprj_io_drive_sel[25]
+ mprj_io_drive_sel[24] mprj_io_pu_select[12] mprj_io_slew_select[12] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[12] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_33 mprj_io_out[25] mprj_io_schmitt_select[25] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[25] mprj_io_outen[25] mprj_io[25] mprj_io_pd_select[25] mprj_io_drive_sel[525]
+ mprj_io_drive_sel[51] mprj_io_pu_select[25] mprj_io_slew_select[25] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[25] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_930 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_941 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_952 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_963 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_11 mprj_io_out[6] mprj_io_schmitt_select[6] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[6] mprj_io_outen[6] mprj_io[6] mprj_io_pd_select[6] mprj_io_drive_sel[13]
+ mprj_io_drive_sel[12] mprj_io_pu_select[6] mprj_io_slew_select[6] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[6] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_974 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_985 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_996 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_204 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_215 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_226 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_237 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_259 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_248 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_760 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_771 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_782 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_793 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_8 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1029 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1018 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1007 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_590 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_419 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_408 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_920 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_931 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_942 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_953 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_964 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_975 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_997 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_986 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_12 mprj_io_out[18] mprj_io_schmitt_select[18] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[18] mprj_io_outen[18] mprj_io[18] mprj_io_pd_select[18] mprj_io_drive_sel[36]
+ mprj_io_drive_sel[37] mprj_io_pu_select[18] mprj_io_slew_select[18] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[18] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_23 mprj_io_out[21] mprj_io_schmitt_select[21] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[21] mprj_io_outen[21] mprj_io[21] mprj_io_pd_select[21] mprj_io_drive_sel[42]
+ mprj_io_drive_sel[43] mprj_io_pu_select[21] mprj_io_slew_select[21] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[21] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_34 mprj_io_out[26] mprj_io_schmitt_select[26] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[26] mprj_io_outen[26] mprj_io[26] mprj_io_pd_select[26] mprj_io_drive_sel[52]
+ mprj_io_drive_sel[53] mprj_io_pu_select[26] mprj_io_slew_select[26] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[26] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_750 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_205 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_216 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_227 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_238 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_249 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1019 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1008 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_772 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_783 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_794 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_9 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_761 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_580 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_591 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_409 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_910 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_921 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_932 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_943 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_965 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_976 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_987 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_13 mprj_io_out[22] mprj_io_schmitt_select[22] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[22] mprj_io_outen[22] mprj_io[22] mprj_io_pd_select[22] mprj_io_drive_sel[44]
+ mprj_io_drive_sel[45] mprj_io_pu_select[22] mprj_io_slew_select[22] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[22] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_24 mprj_io_out[14] mprj_io_schmitt_select[14] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[14] mprj_io_outen[14] mprj_io[14] mprj_io_pd_select[14] mprj_io_drive_sel[28]
+ mprj_io_drive_sel[29] mprj_io_pu_select[14] mprj_io_slew_select[14] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[14] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_35 mprj_io_out[27] mprj_io_schmitt_select[27] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[27] mprj_io_outen[27] mprj_io[27] mprj_io_pd_select[27] mprj_io_drive_sel[54]
+ mprj_io_drive_sel[55] mprj_io_pu_select[27] mprj_io_slew_select[27] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[27] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_206 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_217 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_228 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_239 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_1009 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_740 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_751 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_762 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_784 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_795 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_773 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_570 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_581 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_592 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_900 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_911 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_922 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_933 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_944 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_955 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_966 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_977 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_999 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_988 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_25 mprj_io_out[15] mprj_io_schmitt_select[15] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[15] mprj_io_outen[15] mprj_io[15] mprj_io_pd_select[15] mprj_io_drive_sel[30]
+ mprj_io_drive_sel[31] mprj_io_pu_select[15] mprj_io_slew_select[15] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[15] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_14 mprj_io_out[19] mprj_io_schmitt_select[19] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[19] mprj_io_outen[19] mprj_io[19] mprj_io_pd_select[19] mprj_io_drive_sel[38]
+ mprj_io_drive_sel[39] mprj_io_pu_select[19] mprj_io_slew_select[19] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[19] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_36 mprj_io_out[31] mprj_io_schmitt_select[31] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[31] mprj_io_outen[31] mprj_io[31] mprj_io_pd_select[31] mprj_io_drive_sel[62]
+ mprj_io_drive_sel[63] mprj_io_pu_select[31] mprj_io_slew_select[31] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[31] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_207 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_218 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_229 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_730 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_741 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_752 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_763 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_774 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_796 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_785 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_560 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_571 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_582 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_593 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_390 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_912 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_923 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_934 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_945 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_956 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_967 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_978 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_901 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_989 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_26 mprj_io_out[16] mprj_io_schmitt_select[16] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[16] mprj_io_outen[16] mprj_io[16] mprj_io_pd_select[16] mprj_io_drive_sel[32]
+ mprj_io_drive_sel[33] mprj_io_pu_select[16] mprj_io_slew_select[16] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[16] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_15 mprj_io_out[7] mprj_io_schmitt_select[7] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[7] mprj_io_outen[7] mprj_io[7] mprj_io_pd_select[7] mprj_io_drive_sel[15]
+ mprj_io_drive_sel[14] mprj_io_pu_select[7] mprj_io_slew_select[7] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[7] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_37 mprj_io_out[37] mprj_io_schmitt_select[37] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[37] mprj_io_outen[37] mprj_io[37] mprj_io_pd_select[37] mprj_io_drive_sel[74]
+ mprj_io_drive_sel[75] mprj_io_pu_select[37] mprj_io_slew_select[37] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[37] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_208 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_219 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_720 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_731 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_742 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_753 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_764 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_775 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_786 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_797 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_550 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_561 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_572 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_583 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_594 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_391 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_380 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_27 mprj_io_out[17] mprj_io_schmitt_select[17] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[17] mprj_io_outen[17] mprj_io[17] mprj_io_pd_select[17] mprj_io_drive_sel[34]
+ mprj_io_drive_sel[35] mprj_io_pu_select[17] mprj_io_slew_select[17] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[17] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_16 mprj_io_out[8] mprj_io_schmitt_select[8] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[8] mprj_io_outen[8] mprj_io[8] mprj_io_pd_select[8] mprj_io_drive_sel[17]
+ mprj_io_drive_sel[16] mprj_io_pu_select[8] mprj_io_slew_select[8] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[8] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_902 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_913 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_924 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_935 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_946 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_957 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_968 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_979 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_38 mprj_io_out[35] mprj_io_schmitt_select[35] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[35] mprj_io_outen[35] mprj_io[35] mprj_io_pd_select[35] mprj_io_drive_sel[70]
+ mprj_io_drive_sel[71] mprj_io_pu_select[35] mprj_io_slew_select[35] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[35] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__in_c_0 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS clock gf180mcu_fd_io__in_c_0/PD gf180mcu_fd_io__in_c_0/PU
+ gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS clock_core gf180mcu_fd_io__in_c
Xgf180mcu_fd_io__fill10_209 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_710 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_721 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_732 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_743 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_754 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_765 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_776 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_787 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_798 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_540 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_551 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_562 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_573 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_584 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_595 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_392 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_381 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_370 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__cor_0 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor
Xgf180mcu_fd_io__fill10_903 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_914 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_936 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_947 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_958 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_925 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_28 mprj_io_out[23] mprj_io_schmitt_select[23] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[23] mprj_io_outen[23] mprj_io[23] mprj_io_pd_select[23] mprj_io_drive_sel[46]
+ mprj_io_drive_sel[47] mprj_io_pu_select[23] mprj_io_slew_select[23] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[23] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_17 mprj_io_out[9] mprj_io_schmitt_select[9] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[9] mprj_io_outen[9] mprj_io[9] mprj_io_pd_select[9] mprj_io_drive_sel[19]
+ mprj_io_drive_sel[18] mprj_io_pu_select[9] mprj_io_slew_select[9] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[9] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_39 mprj_io_out[32] mprj_io_schmitt_select[32] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[32] mprj_io_outen[32] mprj_io[32] mprj_io_pd_select[32] mprj_io_drive_sel[64]
+ mprj_io_drive_sel[65] mprj_io_pu_select[32] mprj_io_slew_select[32] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[32] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_700 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_711 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_722 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_733 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_744 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_755 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_766 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_777 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_788 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_799 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_530 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_541 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_552 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_563 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_574 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_585 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_596 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_393 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_382 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_371 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_360 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__cor_1 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor
Xgf180mcu_fd_io__fill10_190 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_904 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_915 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_926 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_937 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_948 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_959 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_29 mprj_io_out[24] mprj_io_schmitt_select[24] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[24] mprj_io_outen[24] mprj_io[24] mprj_io_pd_select[24] mprj_io_drive_sel[48]
+ mprj_io_drive_sel[49] mprj_io_pu_select[24] mprj_io_slew_select[24] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[24] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__bi_t_18 mprj_io_out[10] mprj_io_schmitt_select[10] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[10] mprj_io_outen[10] mprj_io[10] mprj_io_pd_select[10] mprj_io_drive_sel[21]
+ mprj_io_drive_sel[20] mprj_io_pu_select[10] mprj_io_slew_select[10] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[10] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_701 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_712 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_723 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_734 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_745 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_756 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_767 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_778 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_789 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_520 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_531 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_553 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_542 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_564 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_575 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_586 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_597 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_90 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__cor_2 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor
Xgf180mcu_fd_io__fill10_394 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_383 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_372 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_361 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_350 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_180 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_191 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_905 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_927 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_938 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_949 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_916 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__bi_t_19 mprj_io_out[11] mprj_io_schmitt_select[11] gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ mprj_io_inen[11] mprj_io_outen[11] mprj_io[11] mprj_io_pd_select[11] mprj_io_drive_sel[23]
+ mprj_io_drive_sel[22] mprj_io_pu_select[11] mprj_io_slew_select[11] gf180mcu_fd_io__cor_3/VDD
+ gf180mcu_fd_io__cor_3/VSS mprj_io_in[11] gf180mcu_fd_io__bi_t
Xgf180mcu_fd_io__fill10_702 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_713 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_724 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_735 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_746 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_757 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_768 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_779 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_521 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_510 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_532 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_543 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_554 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_565 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_576 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_587 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_598 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_80 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_91 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__cor_3 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor
Xgf180mcu_fd_io__fill10_395 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_384 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_373 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_362 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_351 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_340 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_170 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_181 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_192 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_906 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_917 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_928 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_703 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_714 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_725 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_736 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_747 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_758 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_769 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_522 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_533 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_544 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_555 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_566 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_577 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_588 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_599 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_511 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_500 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_81 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_70 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_92 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_396 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_385 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_374 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_363 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_352 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_341 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_330 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_160 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_171 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_182 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_193 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_907 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_918 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_929 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_704 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_715 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_726 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_737 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_748 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_759 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_523 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_534 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_545 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_556 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_567 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_578 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_589 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_512 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_501 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_82 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_71 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_60 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_93 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_397 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_386 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_375 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_364 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_353 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_342 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_331 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_320 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_150 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_161 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_172 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_183 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_194 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_908 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_919 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_705 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_716 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_727 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_738 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
Xgf180mcu_fd_io__fill10_749 gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS gf180mcu_fd_io__cor_3/VDD gf180mcu_fd_io__cor_3/VSS
+ gf180mcu_fd_io__fill10
.ends

* Black-box entry subcircuit for mgmt_core_wrapper abstract view
.subckt mgmt_core_wrapper VDD VSS core_clk core_rstn debug_in debug_mode debug_oeb
+ debug_out flash_clk flash_csb flash_io0_di flash_io0_do flash_io0_oeb flash_io1_di
+ flash_io1_do flash_io1_oeb flash_io2_di flash_io2_do flash_io2_oeb flash_io3_di
+ flash_io3_do flash_io3_oeb gpio_in_pad gpio_inenb_pad gpio_mode0_pad gpio_mode1_pad
+ gpio_out_pad gpio_outenb_pad hk_ack_i hk_cyc_o hk_dat_i[0] hk_dat_i[10] hk_dat_i[11]
+ hk_dat_i[12] hk_dat_i[13] hk_dat_i[14] hk_dat_i[15] hk_dat_i[16] hk_dat_i[17] hk_dat_i[18]
+ hk_dat_i[19] hk_dat_i[1] hk_dat_i[20] hk_dat_i[21] hk_dat_i[22] hk_dat_i[23] hk_dat_i[24]
+ hk_dat_i[25] hk_dat_i[26] hk_dat_i[27] hk_dat_i[28] hk_dat_i[29] hk_dat_i[2] hk_dat_i[30]
+ hk_dat_i[31] hk_dat_i[3] hk_dat_i[4] hk_dat_i[5] hk_dat_i[6] hk_dat_i[7] hk_dat_i[8]
+ hk_dat_i[9] hk_stb_o irq[0] irq[1] irq[2] irq[3] irq[4] irq[5] la_iena[0] la_iena[10]
+ la_iena[11] la_iena[12] la_iena[13] la_iena[14] la_iena[15] la_iena[16] la_iena[17]
+ la_iena[18] la_iena[19] la_iena[1] la_iena[20] la_iena[21] la_iena[22] la_iena[23]
+ la_iena[24] la_iena[25] la_iena[26] la_iena[27] la_iena[28] la_iena[29] la_iena[2]
+ la_iena[30] la_iena[31] la_iena[32] la_iena[33] la_iena[34] la_iena[35] la_iena[36]
+ la_iena[37] la_iena[38] la_iena[39] la_iena[3] la_iena[40] la_iena[41] la_iena[42]
+ la_iena[43] la_iena[44] la_iena[45] la_iena[46] la_iena[47] la_iena[48] la_iena[49]
+ la_iena[4] la_iena[50] la_iena[51] la_iena[52] la_iena[53] la_iena[54] la_iena[55]
+ la_iena[56] la_iena[57] la_iena[58] la_iena[59] la_iena[5] la_iena[60] la_iena[61]
+ la_iena[62] la_iena[63] la_iena[6] la_iena[7] la_iena[8] la_iena[9] la_input[0]
+ la_input[10] la_input[11] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16]
+ la_input[17] la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22]
+ la_input[23] la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29]
+ la_input[2] la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35]
+ la_input[36] la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41]
+ la_input[42] la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48]
+ la_input[49] la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54]
+ la_input[55] la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60]
+ la_input[61] la_input[62] la_input[63] la_input[6] la_input[7] la_input[8] la_input[9]
+ la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15]
+ la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21]
+ la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28]
+ la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40]
+ la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5]
+ la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8]
+ la_oenb[9] la_output[0] la_output[10] la_output[11] la_output[12] la_output[13]
+ la_output[14] la_output[15] la_output[16] la_output[17] la_output[18] la_output[19]
+ la_output[1] la_output[20] la_output[21] la_output[22] la_output[23] la_output[24]
+ la_output[25] la_output[26] la_output[27] la_output[28] la_output[29] la_output[2]
+ la_output[30] la_output[31] la_output[32] la_output[33] la_output[34] la_output[35]
+ la_output[36] la_output[37] la_output[38] la_output[39] la_output[3] la_output[40]
+ la_output[41] la_output[42] la_output[43] la_output[44] la_output[45] la_output[46]
+ la_output[47] la_output[48] la_output[49] la_output[4] la_output[50] la_output[51]
+ la_output[52] la_output[53] la_output[54] la_output[55] la_output[56] la_output[57]
+ la_output[58] la_output[59] la_output[5] la_output[60] la_output[61] la_output[62]
+ la_output[63] la_output[6] la_output[7] la_output[8] la_output[9] mprj_ack_i mprj_adr_o[0]
+ mprj_adr_o[10] mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15]
+ mprj_adr_o[16] mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20]
+ mprj_adr_o[21] mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26]
+ mprj_adr_o[27] mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31]
+ mprj_adr_o[3] mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8]
+ mprj_adr_o[9] mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12]
+ mprj_dat_i[13] mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18]
+ mprj_dat_i[19] mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23]
+ mprj_dat_i[24] mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29]
+ mprj_dat_i[2] mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5]
+ mprj_dat_i[6] mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10]
+ mprj_dat_o[11] mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16]
+ mprj_dat_o[17] mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21]
+ mprj_dat_o[22] mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27]
+ mprj_dat_o[28] mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3]
+ mprj_dat_o[4] mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9]
+ mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2] mprj_sel_o[3] mprj_stb_o mprj_wb_iena
+ mprj_we_o qspi_enabled ser_rx ser_tx spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb trap uart_enabled user_irq_ena[0] user_irq_ena[1] user_irq_ena[2]
.ends

* Black-box entry subcircuit for simple_por abstract view
.subckt simple_por vdd vss porb por
.ends

* Black-box entry subcircuit for caravel_clocking abstract view
.subckt caravel_clocking VDD VSS core_clk ext_clk ext_clk_sel ext_reset pll_clk pll_clk90
+ resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
.ends

* Black-box entry subcircuit for spare_logic_block abstract view
.subckt spare_logic_block VDD VSS spare_xfq[0] spare_xfq[1] spare_xi[0] spare_xi[1]
+ spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0] spare_xna[1]
+ spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12] spare_xz[13]
+ spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19] spare_xz[1]
+ spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25] spare_xz[26]
+ spare_xz[27] spare_xz[28] spare_xz[29] spare_xz[2] spare_xz[30] spare_xz[3] spare_xz[4]
+ spare_xz[5] spare_xz[6] spare_xz[7] spare_xz[8] spare_xz[9]
.ends

* Black-box entry subcircuit for user_id_programming abstract view
.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VDD VSS
.ends

* Black-box entry subcircuit for mgmt_protect abstract view
.subckt mgmt_protect VDD VSS caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0]
+ la_data_in_core[10] la_data_in_core[11] la_data_in_core[12] la_data_in_core[13]
+ la_data_in_core[14] la_data_in_core[15] la_data_in_core[16] la_data_in_core[17]
+ la_data_in_core[18] la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21]
+ la_data_in_core[22] la_data_in_core[23] la_data_in_core[24] la_data_in_core[25]
+ la_data_in_core[26] la_data_in_core[27] la_data_in_core[28] la_data_in_core[29]
+ la_data_in_core[2] la_data_in_core[30] la_data_in_core[31] la_data_in_core[32] la_data_in_core[33]
+ la_data_in_core[34] la_data_in_core[35] la_data_in_core[36] la_data_in_core[37]
+ la_data_in_core[38] la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41]
+ la_data_in_core[42] la_data_in_core[43] la_data_in_core[44] la_data_in_core[45]
+ la_data_in_core[46] la_data_in_core[47] la_data_in_core[48] la_data_in_core[49]
+ la_data_in_core[4] la_data_in_core[50] la_data_in_core[51] la_data_in_core[52] la_data_in_core[53]
+ la_data_in_core[54] la_data_in_core[55] la_data_in_core[56] la_data_in_core[57]
+ la_data_in_core[58] la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61]
+ la_data_in_core[62] la_data_in_core[63] la_data_in_core[6] la_data_in_core[7] la_data_in_core[8]
+ la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[10] la_data_in_mprj[11] la_data_in_mprj[12]
+ la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15] la_data_in_mprj[16]
+ la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19] la_data_in_mprj[1] la_data_in_mprj[20]
+ la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23] la_data_in_mprj[24]
+ la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27] la_data_in_mprj[28]
+ la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31] la_data_in_mprj[32]
+ la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35] la_data_in_mprj[36]
+ la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39] la_data_in_mprj[3] la_data_in_mprj[40]
+ la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43] la_data_in_mprj[44]
+ la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47] la_data_in_mprj[48]
+ la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51] la_data_in_mprj[52]
+ la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55] la_data_in_mprj[56]
+ la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59] la_data_in_mprj[5] la_data_in_mprj[60]
+ la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63] la_data_in_mprj[6] la_data_in_mprj[7]
+ la_data_in_mprj[8] la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[10] la_data_out_core[11]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[6] la_data_out_core[7] la_data_out_core[8]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[10] la_data_out_mprj[11]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[6] la_data_out_mprj[7] la_data_out_mprj[8]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[10] la_iena_mprj[11] la_iena_mprj[12]
+ la_iena_mprj[13] la_iena_mprj[14] la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17]
+ la_iena_mprj[18] la_iena_mprj[19] la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21]
+ la_iena_mprj[22] la_iena_mprj[23] la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26]
+ la_iena_mprj[27] la_iena_mprj[28] la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30]
+ la_iena_mprj[31] la_iena_mprj[32] la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35]
+ la_iena_mprj[36] la_iena_mprj[37] la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3]
+ la_iena_mprj[40] la_iena_mprj[41] la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44]
+ la_iena_mprj[45] la_iena_mprj[46] la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49]
+ la_iena_mprj[4] la_iena_mprj[50] la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53]
+ la_iena_mprj[54] la_iena_mprj[55] la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58]
+ la_iena_mprj[59] la_iena_mprj[5] la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62]
+ la_iena_mprj[63] la_iena_mprj[6] la_iena_mprj[7] la_iena_mprj[8] la_iena_mprj[9]
+ la_oenb_core[0] la_oenb_core[10] la_oenb_core[11] la_oenb_core[12] la_oenb_core[13]
+ la_oenb_core[14] la_oenb_core[15] la_oenb_core[16] la_oenb_core[17] la_oenb_core[18]
+ la_oenb_core[19] la_oenb_core[1] la_oenb_core[20] la_oenb_core[21] la_oenb_core[22]
+ la_oenb_core[23] la_oenb_core[24] la_oenb_core[25] la_oenb_core[26] la_oenb_core[27]
+ la_oenb_core[28] la_oenb_core[29] la_oenb_core[2] la_oenb_core[30] la_oenb_core[31]
+ la_oenb_core[32] la_oenb_core[33] la_oenb_core[34] la_oenb_core[35] la_oenb_core[36]
+ la_oenb_core[37] la_oenb_core[38] la_oenb_core[39] la_oenb_core[3] la_oenb_core[40]
+ la_oenb_core[41] la_oenb_core[42] la_oenb_core[43] la_oenb_core[44] la_oenb_core[45]
+ la_oenb_core[46] la_oenb_core[47] la_oenb_core[48] la_oenb_core[49] la_oenb_core[4]
+ la_oenb_core[50] la_oenb_core[51] la_oenb_core[52] la_oenb_core[53] la_oenb_core[54]
+ la_oenb_core[55] la_oenb_core[56] la_oenb_core[57] la_oenb_core[58] la_oenb_core[59]
+ la_oenb_core[5] la_oenb_core[60] la_oenb_core[61] la_oenb_core[62] la_oenb_core[63]
+ la_oenb_core[6] la_oenb_core[7] la_oenb_core[8] la_oenb_core[9] la_oenb_mprj[0]
+ la_oenb_mprj[10] la_oenb_mprj[11] la_oenb_mprj[12] la_oenb_mprj[13] la_oenb_mprj[14]
+ la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18] la_oenb_mprj[19]
+ la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22] la_oenb_mprj[23]
+ la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27] la_oenb_mprj[28]
+ la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31] la_oenb_mprj[32]
+ la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36] la_oenb_mprj[37]
+ la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40] la_oenb_mprj[41]
+ la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45] la_oenb_mprj[46]
+ la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4] la_oenb_mprj[50]
+ la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54] la_oenb_mprj[55]
+ la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59] la_oenb_mprj[5]
+ la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63] la_oenb_mprj[6]
+ la_oenb_mprj[7] la_oenb_mprj[8] la_oenb_mprj[9] mprj_ack_i_core mprj_ack_i_user
+ mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12] mprj_adr_o_core[13]
+ mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16] mprj_adr_o_core[17]
+ mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21]
+ mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24] mprj_adr_o_core[25]
+ mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28] mprj_adr_o_core[29]
+ mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3] mprj_adr_o_core[4]
+ mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8] mprj_adr_o_core[9]
+ mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12] mprj_adr_o_user[13]
+ mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16] mprj_adr_o_user[17]
+ mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21]
+ mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24] mprj_adr_o_user[25]
+ mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28] mprj_adr_o_user[29]
+ mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3] mprj_adr_o_user[4]
+ mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8] mprj_adr_o_user[9]
+ mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0] mprj_dat_i_core[10] mprj_dat_i_core[11]
+ mprj_dat_i_core[12] mprj_dat_i_core[13] mprj_dat_i_core[14] mprj_dat_i_core[15]
+ mprj_dat_i_core[16] mprj_dat_i_core[17] mprj_dat_i_core[18] mprj_dat_i_core[19]
+ mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21] mprj_dat_i_core[22] mprj_dat_i_core[23]
+ mprj_dat_i_core[24] mprj_dat_i_core[25] mprj_dat_i_core[26] mprj_dat_i_core[27]
+ mprj_dat_i_core[28] mprj_dat_i_core[29] mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31]
+ mprj_dat_i_core[3] mprj_dat_i_core[4] mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7]
+ mprj_dat_i_core[8] mprj_dat_i_core[9] mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11]
+ mprj_dat_i_user[12] mprj_dat_i_user[13] mprj_dat_i_user[14] mprj_dat_i_user[15]
+ mprj_dat_i_user[16] mprj_dat_i_user[17] mprj_dat_i_user[18] mprj_dat_i_user[19]
+ mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21] mprj_dat_i_user[22] mprj_dat_i_user[23]
+ mprj_dat_i_user[24] mprj_dat_i_user[25] mprj_dat_i_user[26] mprj_dat_i_user[27]
+ mprj_dat_i_user[28] mprj_dat_i_user[29] mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31]
+ mprj_dat_i_user[3] mprj_dat_i_user[4] mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7]
+ mprj_dat_i_user[8] mprj_dat_i_user[9] mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11]
+ mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14] mprj_dat_o_core[15]
+ mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18] mprj_dat_o_core[19]
+ mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22] mprj_dat_o_core[23]
+ mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26] mprj_dat_o_core[27]
+ mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31]
+ mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7]
+ mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11]
+ mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14] mprj_dat_o_user[15]
+ mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18] mprj_dat_o_user[19]
+ mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22] mprj_dat_o_user[23]
+ mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26] mprj_dat_o_user[27]
+ mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31]
+ mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7]
+ mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user_clock user_clock2 user_irq[0] user_irq[1] user_irq[2] user_irq_core[0] user_irq_core[1]
+ user_irq_core[2] user_irq_ena[0] user_irq_ena[1] user_irq_ena[2] user_reset
.ends

* Black-box entry subcircuit for gpio_defaults_block_009 abstract view
.subckt gpio_defaults_block_009 gpio_defaults[0] gpio_defaults[1] gpio_defaults[2]
+ gpio_defaults[3] gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[9] VDD VSS
.ends

* Black-box entry subcircuit for gpio_defaults_block_007 abstract view
.subckt gpio_defaults_block_007 gpio_defaults[0] gpio_defaults[1] gpio_defaults[2]
+ gpio_defaults[3] gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[9] VDD VSS
.ends

* Black-box entry subcircuit for user_project_wrapper abstract view
.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for housekeeping abstract view
.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
.ends

.subckt caravel clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb vdd vss
Xgpio_control_in_2\[0\] soc/VDD soc/VSS gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[1]
+ gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3] gpio_defaults_block_6/gpio_defaults[4]
+ gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6] gpio_defaults_block_6/gpio_defaults[7]
+ gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9] housekeeping/mgmt_gpio_in[19]
+ gpio_control_in_2\[0\]/zero housekeeping/mgmt_gpio_out[19] gpio_control_in_2\[0\]/one
+ padframe/mprj_io_drive_sel[38] padframe/mprj_io_drive_sel[39] padframe/mprj_io_in[19]
+ padframe/mprj_io_inen[19] padframe/mprj_io_out[19] padframe/mprj_io_outen[19] padframe/mprj_io_pd_select[19]
+ padframe/mprj_io_pu_select[19] padframe/mprj_io_schmitt_select[19] padframe/mprj_io_slew_select[19]
+ gpio_control_in_2\[0\]/resetn gpio_control_in_2\[0\]/resetn_out gpio_control_in_2\[0\]/serial_clock
+ gpio_control_in_2\[0\]/serial_clock_out gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[0\]/serial_data_out
+ gpio_control_in_2\[0\]/serial_load gpio_control_in_2\[0\]/serial_load_out mprj/io_in[19]
+ mprj/io_oeb[19] mprj/io_out[19] gpio_control_in_2\[0\]/zero gpio_control_block
Xgpio_defaults_block_11 gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[1]
+ gpio_defaults_block_11/gpio_defaults[2] gpio_defaults_block_11/gpio_defaults[3]
+ gpio_defaults_block_11/gpio_defaults[4] gpio_defaults_block_11/gpio_defaults[5]
+ gpio_defaults_block_11/gpio_defaults[6] gpio_defaults_block_11/gpio_defaults[7]
+ gpio_defaults_block_11/gpio_defaults[8] gpio_defaults_block_11/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_22 gpio_defaults_block_22/gpio_defaults[0] gpio_defaults_block_22/gpio_defaults[1]
+ gpio_defaults_block_22/gpio_defaults[2] gpio_defaults_block_22/gpio_defaults[3]
+ gpio_defaults_block_22/gpio_defaults[4] gpio_defaults_block_22/gpio_defaults[5]
+ gpio_defaults_block_22/gpio_defaults[6] gpio_defaults_block_22/gpio_defaults[7]
+ gpio_defaults_block_22/gpio_defaults[8] gpio_defaults_block_22/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1\[6\] soc/VDD soc/VSS gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[1]
+ gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3] gpio_defaults_block_1/gpio_defaults[4]
+ gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6] gpio_defaults_block_1/gpio_defaults[7]
+ gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9] housekeeping/mgmt_gpio_in[14]
+ gpio_control_in_1\[6\]/zero housekeeping/mgmt_gpio_out[14] gpio_control_in_1\[6\]/one
+ padframe/mprj_io_drive_sel[28] padframe/mprj_io_drive_sel[29] padframe/mprj_io_in[14]
+ padframe/mprj_io_inen[14] padframe/mprj_io_out[14] padframe/mprj_io_outen[14] padframe/mprj_io_pd_select[14]
+ padframe/mprj_io_pu_select[14] padframe/mprj_io_schmitt_select[14] padframe/mprj_io_slew_select[14]
+ gpio_control_in_1\[6\]/resetn gpio_control_in_1\[7\]/resetn gpio_control_in_1\[6\]/serial_clock
+ gpio_control_in_1\[7\]/serial_clock gpio_control_in_1\[6\]/serial_data_in gpio_control_in_1\[7\]/serial_data_in
+ gpio_control_in_1\[6\]/serial_load gpio_control_in_1\[7\]/serial_load mprj/io_in[14]
+ mprj/io_oeb[14] mprj/io_out[14] gpio_control_in_1\[6\]/zero gpio_control_block
Xgpio_defaults_block_12 gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[1]
+ gpio_defaults_block_12/gpio_defaults[2] gpio_defaults_block_12/gpio_defaults[3]
+ gpio_defaults_block_12/gpio_defaults[4] gpio_defaults_block_12/gpio_defaults[5]
+ gpio_defaults_block_12/gpio_defaults[6] gpio_defaults_block_12/gpio_defaults[7]
+ gpio_defaults_block_12/gpio_defaults[8] gpio_defaults_block_12/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_23 gpio_defaults_block_23/gpio_defaults[0] gpio_defaults_block_23/gpio_defaults[1]
+ gpio_defaults_block_23/gpio_defaults[2] gpio_defaults_block_23/gpio_defaults[3]
+ gpio_defaults_block_23/gpio_defaults[4] gpio_defaults_block_23/gpio_defaults[5]
+ gpio_defaults_block_23/gpio_defaults[6] gpio_defaults_block_23/gpio_defaults[7]
+ gpio_defaults_block_23/gpio_defaults[8] gpio_defaults_block_23/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xpll soc/VDD soc/VSS pll/clockp[0] pll/clockp[1] pll/dco pll/div[0] pll/div[1] pll/div[2]
+ pll/div[3] pll/div[4] pll/enable pll/ext_trim[0] pll/ext_trim[10] pll/ext_trim[11]
+ pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14] pll/ext_trim[15] pll/ext_trim[16]
+ pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19] pll/ext_trim[1] pll/ext_trim[20]
+ pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23] pll/ext_trim[24] pll/ext_trim[25]
+ pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4] pll/ext_trim[5] pll/ext_trim[6]
+ pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9] pll/osc pll/resetb digital_pll
Xpadframe clock pll/osc flash_clk padframe/flash_clk_core padframe/flash_clk_oe_core
+ flash_csb padframe/flash_csb_core padframe/flash_csb_oe_core flash_io0 padframe/flash_io0_di_core
+ padframe/flash_io0_do_core padframe/flash_io0_ie_core padframe/flash_io0_oe_core
+ flash_io1 padframe/flash_io1_di_core padframe/flash_io1_do_core padframe/flash_io1_ie_core
+ padframe/flash_io1_oe_core gpio soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_in_pad
+ soc/gpio_inenb_pad soc/gpio_out_pad soc/gpio_outenb_pad padframe/gpio_pd_select
+ padframe/gpio_pu_select padframe/gpio_schmitt_select padframe/gpio_slew_select mprj_io[0]
+ mprj_io[10] mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16]
+ mprj_io[17] mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22]
+ mprj_io[23] mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29]
+ mprj_io[2] mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35]
+ mprj_io[36] mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8]
+ mprj_io[9] padframe/mprj_io_drive_sel[0] padframe/mprj_io_drive_sel[10] padframe/mprj_io_drive_sel[11]
+ padframe/mprj_io_drive_sel[12] padframe/mprj_io_drive_sel[13] padframe/mprj_io_drive_sel[14]
+ padframe/mprj_io_drive_sel[15] padframe/mprj_io_drive_sel[16] padframe/mprj_io_drive_sel[17]
+ padframe/mprj_io_drive_sel[18] padframe/mprj_io_drive_sel[19] padframe/mprj_io_drive_sel[1]
+ padframe/mprj_io_drive_sel[20] padframe/mprj_io_drive_sel[21] padframe/mprj_io_drive_sel[22]
+ padframe/mprj_io_drive_sel[23] padframe/mprj_io_drive_sel[24] padframe/mprj_io_drive_sel[25]
+ padframe/mprj_io_drive_sel[26] padframe/mprj_io_drive_sel[27] padframe/mprj_io_drive_sel[28]
+ padframe/mprj_io_drive_sel[29] padframe/mprj_io_drive_sel[2] padframe/mprj_io_drive_sel[30]
+ padframe/mprj_io_drive_sel[31] padframe/mprj_io_drive_sel[32] padframe/mprj_io_drive_sel[33]
+ padframe/mprj_io_drive_sel[34] padframe/mprj_io_drive_sel[35] padframe/mprj_io_drive_sel[36]
+ padframe/mprj_io_drive_sel[37] padframe/mprj_io_drive_sel[38] padframe/mprj_io_drive_sel[39]
+ padframe/mprj_io_drive_sel[3] padframe/mprj_io_drive_sel[40] padframe/mprj_io_drive_sel[41]
+ padframe/mprj_io_drive_sel[42] padframe/mprj_io_drive_sel[43] padframe/mprj_io_drive_sel[44]
+ padframe/mprj_io_drive_sel[45] padframe/mprj_io_drive_sel[46] padframe/mprj_io_drive_sel[47]
+ padframe/mprj_io_drive_sel[48] padframe/mprj_io_drive_sel[49] padframe/mprj_io_drive_sel[4]
+ padframe/mprj_io_drive_sel[51] padframe/mprj_io_drive_sel[525] padframe/mprj_io_drive_sel[52]
+ padframe/mprj_io_drive_sel[53] padframe/mprj_io_drive_sel[54] padframe/mprj_io_drive_sel[55]
+ padframe/mprj_io_drive_sel[56] padframe/mprj_io_drive_sel[57] padframe/mprj_io_drive_sel[58]
+ padframe/mprj_io_drive_sel[59] padframe/mprj_io_drive_sel[5] padframe/mprj_io_drive_sel[61]
+ padframe/mprj_io_drive_sel[62] padframe/mprj_io_drive_sel[63] padframe/mprj_io_drive_sel[64]
+ padframe/mprj_io_drive_sel[65] padframe/mprj_io_drive_sel[66] padframe/mprj_io_drive_sel[67]
+ padframe/mprj_io_drive_sel[68] padframe/mprj_io_drive_sel[69] padframe/mprj_io_drive_sel[6]
+ padframe/mprj_io_drive_sel[70] padframe/mprj_io_drive_sel[71] padframe/mprj_io_drive_sel[72]
+ padframe/mprj_io_drive_sel[73] padframe/mprj_io_drive_sel[74] padframe/mprj_io_drive_sel[75]
+ padframe/mprj_io_drive_sel[7] padframe/mprj_io_drive_sel[8] padframe/mprj_io_drive_sel[9]
+ padframe/mprj_io_in[0] padframe/mprj_io_in[10] padframe/mprj_io_in[11] padframe/mprj_io_in[12]
+ padframe/mprj_io_in[13] padframe/mprj_io_in[14] padframe/mprj_io_in[15] padframe/mprj_io_in[16]
+ padframe/mprj_io_in[17] padframe/mprj_io_in[18] padframe/mprj_io_in[19] padframe/mprj_io_in[1]
+ padframe/mprj_io_in[20] padframe/mprj_io_in[21] padframe/mprj_io_in[22] padframe/mprj_io_in[23]
+ padframe/mprj_io_in[24] padframe/mprj_io_in[25] padframe/mprj_io_in[26] padframe/mprj_io_in[27]
+ padframe/mprj_io_in[28] padframe/mprj_io_in[29] padframe/mprj_io_in[2] padframe/mprj_io_in[30]
+ padframe/mprj_io_in[31] padframe/mprj_io_in[32] padframe/mprj_io_in[33] padframe/mprj_io_in[34]
+ padframe/mprj_io_in[35] padframe/mprj_io_in[36] padframe/mprj_io_in[37] padframe/mprj_io_in[3]
+ padframe/mprj_io_in[4] padframe/mprj_io_in[5] padframe/mprj_io_in[6] padframe/mprj_io_in[7]
+ padframe/mprj_io_in[8] padframe/mprj_io_in[9] padframe/mprj_io_inen[0] padframe/mprj_io_inen[10]
+ padframe/mprj_io_inen[11] padframe/mprj_io_inen[12] padframe/mprj_io_inen[13] padframe/mprj_io_inen[14]
+ padframe/mprj_io_inen[15] padframe/mprj_io_inen[16] padframe/mprj_io_inen[17] padframe/mprj_io_inen[18]
+ padframe/mprj_io_inen[19] padframe/mprj_io_inen[1] padframe/mprj_io_inen[20] padframe/mprj_io_inen[21]
+ padframe/mprj_io_inen[22] padframe/mprj_io_inen[23] padframe/mprj_io_inen[24] padframe/mprj_io_inen[25]
+ padframe/mprj_io_inen[26] padframe/mprj_io_inen[27] padframe/mprj_io_inen[28] padframe/mprj_io_inen[29]
+ padframe/mprj_io_inen[2] padframe/mprj_io_inen[30] padframe/mprj_io_inen[31] padframe/mprj_io_inen[32]
+ padframe/mprj_io_inen[33] padframe/mprj_io_inen[34] padframe/mprj_io_inen[35] padframe/mprj_io_inen[36]
+ padframe/mprj_io_inen[37] padframe/mprj_io_inen[3] padframe/mprj_io_inen[4] padframe/mprj_io_inen[5]
+ padframe/mprj_io_inen[6] padframe/mprj_io_inen[7] padframe/mprj_io_inen[8] padframe/mprj_io_inen[9]
+ padframe/mprj_io_out[0] padframe/mprj_io_out[10] padframe/mprj_io_out[11] padframe/mprj_io_out[12]
+ padframe/mprj_io_out[13] padframe/mprj_io_out[14] padframe/mprj_io_out[15] padframe/mprj_io_out[16]
+ padframe/mprj_io_out[17] padframe/mprj_io_out[18] padframe/mprj_io_out[19] padframe/mprj_io_out[1]
+ padframe/mprj_io_out[20] padframe/mprj_io_out[21] padframe/mprj_io_out[22] padframe/mprj_io_out[23]
+ padframe/mprj_io_out[24] padframe/mprj_io_out[25] padframe/mprj_io_out[26] padframe/mprj_io_out[27]
+ padframe/mprj_io_out[28] padframe/mprj_io_out[29] padframe/mprj_io_out[2] padframe/mprj_io_out[30]
+ padframe/mprj_io_out[31] padframe/mprj_io_out[32] padframe/mprj_io_out[33] padframe/mprj_io_out[34]
+ padframe/mprj_io_out[35] padframe/mprj_io_out[36] padframe/mprj_io_out[37] padframe/mprj_io_out[3]
+ padframe/mprj_io_out[4] padframe/mprj_io_out[5] padframe/mprj_io_out[6] padframe/mprj_io_out[7]
+ padframe/mprj_io_out[8] padframe/mprj_io_out[9] padframe/mprj_io_outen[0] padframe/mprj_io_outen[10]
+ padframe/mprj_io_outen[11] padframe/mprj_io_outen[12] padframe/mprj_io_outen[13]
+ padframe/mprj_io_outen[14] padframe/mprj_io_outen[15] padframe/mprj_io_outen[16]
+ padframe/mprj_io_outen[17] padframe/mprj_io_outen[18] padframe/mprj_io_outen[19]
+ padframe/mprj_io_outen[1] padframe/mprj_io_outen[20] padframe/mprj_io_outen[21]
+ padframe/mprj_io_outen[22] padframe/mprj_io_outen[23] padframe/mprj_io_outen[24]
+ padframe/mprj_io_outen[25] padframe/mprj_io_outen[26] padframe/mprj_io_outen[27]
+ padframe/mprj_io_outen[28] padframe/mprj_io_outen[29] padframe/mprj_io_outen[2]
+ padframe/mprj_io_outen[30] padframe/mprj_io_outen[31] padframe/mprj_io_outen[32]
+ padframe/mprj_io_outen[33] padframe/mprj_io_outen[34] padframe/mprj_io_outen[35]
+ padframe/mprj_io_outen[36] padframe/mprj_io_outen[37] padframe/mprj_io_outen[3]
+ padframe/mprj_io_outen[4] padframe/mprj_io_outen[5] padframe/mprj_io_outen[6] padframe/mprj_io_outen[7]
+ padframe/mprj_io_outen[8] padframe/mprj_io_outen[9] padframe/mprj_io_pd_select[0]
+ padframe/mprj_io_pd_select[10] padframe/mprj_io_pd_select[11] padframe/mprj_io_pd_select[12]
+ padframe/mprj_io_pd_select[13] padframe/mprj_io_pd_select[14] padframe/mprj_io_pd_select[15]
+ padframe/mprj_io_pd_select[16] padframe/mprj_io_pd_select[17] padframe/mprj_io_pd_select[18]
+ padframe/mprj_io_pd_select[19] padframe/mprj_io_pd_select[1] padframe/mprj_io_pd_select[20]
+ padframe/mprj_io_pd_select[21] padframe/mprj_io_pd_select[22] padframe/mprj_io_pd_select[23]
+ padframe/mprj_io_pd_select[24] padframe/mprj_io_pd_select[25] padframe/mprj_io_pd_select[26]
+ padframe/mprj_io_pd_select[27] padframe/mprj_io_pd_select[28] padframe/mprj_io_pd_select[29]
+ padframe/mprj_io_pd_select[2] padframe/mprj_io_pd_select[30] padframe/mprj_io_pd_select[31]
+ padframe/mprj_io_pd_select[32] padframe/mprj_io_pd_select[33] padframe/mprj_io_pd_select[34]
+ padframe/mprj_io_pd_select[35] padframe/mprj_io_pd_select[36] padframe/mprj_io_pd_select[37]
+ padframe/mprj_io_pd_select[3] padframe/mprj_io_pd_select[4] padframe/mprj_io_pd_select[5]
+ padframe/mprj_io_pd_select[6] padframe/mprj_io_pd_select[7] padframe/mprj_io_pd_select[8]
+ padframe/mprj_io_pd_select[9] padframe/mprj_io_pu_select[0] padframe/mprj_io_pu_select[10]
+ padframe/mprj_io_pu_select[11] padframe/mprj_io_pu_select[12] padframe/mprj_io_pu_select[13]
+ padframe/mprj_io_pu_select[14] padframe/mprj_io_pu_select[15] padframe/mprj_io_pu_select[16]
+ padframe/mprj_io_pu_select[17] padframe/mprj_io_pu_select[18] padframe/mprj_io_pu_select[19]
+ padframe/mprj_io_pu_select[1] padframe/mprj_io_pu_select[20] padframe/mprj_io_pu_select[21]
+ padframe/mprj_io_pu_select[22] padframe/mprj_io_pu_select[23] padframe/mprj_io_pu_select[24]
+ padframe/mprj_io_pu_select[25] padframe/mprj_io_pu_select[26] padframe/mprj_io_pu_select[27]
+ padframe/mprj_io_pu_select[28] padframe/mprj_io_pu_select[29] padframe/mprj_io_pu_select[2]
+ padframe/mprj_io_pu_select[30] padframe/mprj_io_pu_select[31] padframe/mprj_io_pu_select[32]
+ padframe/mprj_io_pu_select[33] padframe/mprj_io_pu_select[34] padframe/mprj_io_pu_select[35]
+ padframe/mprj_io_pu_select[36] padframe/mprj_io_pu_select[37] padframe/mprj_io_pu_select[3]
+ padframe/mprj_io_pu_select[4] padframe/mprj_io_pu_select[5] padframe/mprj_io_pu_select[6]
+ padframe/mprj_io_pu_select[7] padframe/mprj_io_pu_select[8] padframe/mprj_io_pu_select[9]
+ padframe/mprj_io_schmitt_select[0] padframe/mprj_io_schmitt_select[10] padframe/mprj_io_schmitt_select[11]
+ padframe/mprj_io_schmitt_select[12] padframe/mprj_io_schmitt_select[13] padframe/mprj_io_schmitt_select[14]
+ padframe/mprj_io_schmitt_select[15] padframe/mprj_io_schmitt_select[16] padframe/mprj_io_schmitt_select[17]
+ padframe/mprj_io_schmitt_select[18] padframe/mprj_io_schmitt_select[19] padframe/mprj_io_schmitt_select[1]
+ padframe/mprj_io_schmitt_select[20] padframe/mprj_io_schmitt_select[21] padframe/mprj_io_schmitt_select[22]
+ padframe/mprj_io_schmitt_select[23] padframe/mprj_io_schmitt_select[24] padframe/mprj_io_schmitt_select[25]
+ padframe/mprj_io_schmitt_select[26] padframe/mprj_io_schmitt_select[27] padframe/mprj_io_schmitt_select[28]
+ padframe/mprj_io_schmitt_select[29] padframe/mprj_io_schmitt_select[2] padframe/mprj_io_schmitt_select[30]
+ padframe/mprj_io_schmitt_select[31] padframe/mprj_io_schmitt_select[32] padframe/mprj_io_schmitt_select[33]
+ padframe/mprj_io_schmitt_select[34] padframe/mprj_io_schmitt_select[35] padframe/mprj_io_schmitt_select[36]
+ padframe/mprj_io_schmitt_select[37] padframe/mprj_io_schmitt_select[3] padframe/mprj_io_schmitt_select[4]
+ padframe/mprj_io_schmitt_select[5] padframe/mprj_io_schmitt_select[6] padframe/mprj_io_schmitt_select[7]
+ padframe/mprj_io_schmitt_select[8] padframe/mprj_io_schmitt_select[9] padframe/mprj_io_slew_select[0]
+ padframe/mprj_io_slew_select[10] padframe/mprj_io_slew_select[11] padframe/mprj_io_slew_select[12]
+ padframe/mprj_io_slew_select[13] padframe/mprj_io_slew_select[14] padframe/mprj_io_slew_select[15]
+ padframe/mprj_io_slew_select[16] padframe/mprj_io_slew_select[17] padframe/mprj_io_slew_select[18]
+ padframe/mprj_io_slew_select[19] padframe/mprj_io_slew_select[1] padframe/mprj_io_slew_select[20]
+ padframe/mprj_io_slew_select[21] padframe/mprj_io_slew_select[22] padframe/mprj_io_slew_select[23]
+ padframe/mprj_io_slew_select[24] padframe/mprj_io_slew_select[25] padframe/mprj_io_slew_select[26]
+ padframe/mprj_io_slew_select[27] padframe/mprj_io_slew_select[28] padframe/mprj_io_slew_select[29]
+ padframe/mprj_io_slew_select[2] padframe/mprj_io_slew_select[30] padframe/mprj_io_slew_select[31]
+ padframe/mprj_io_slew_select[32] padframe/mprj_io_slew_select[33] padframe/mprj_io_slew_select[34]
+ padframe/mprj_io_slew_select[35] padframe/mprj_io_slew_select[36] padframe/mprj_io_slew_select[37]
+ padframe/mprj_io_slew_select[3] padframe/mprj_io_slew_select[4] padframe/mprj_io_slew_select[5]
+ padframe/mprj_io_slew_select[6] padframe/mprj_io_slew_select[7] padframe/mprj_io_slew_select[8]
+ padframe/mprj_io_slew_select[9] resetb pll/resetb vdd vss soc/VSS soc/VDD chip_io
Xgpio_defaults_block_13 gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[1]
+ gpio_defaults_block_13/gpio_defaults[2] gpio_defaults_block_13/gpio_defaults[3]
+ gpio_defaults_block_13/gpio_defaults[4] gpio_defaults_block_13/gpio_defaults[5]
+ gpio_defaults_block_13/gpio_defaults[6] gpio_defaults_block_13/gpio_defaults[7]
+ gpio_defaults_block_13/gpio_defaults[8] gpio_defaults_block_13/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_24 gpio_defaults_block_24/gpio_defaults[0] gpio_defaults_block_24/gpio_defaults[1]
+ gpio_defaults_block_24/gpio_defaults[2] gpio_defaults_block_24/gpio_defaults[3]
+ gpio_defaults_block_24/gpio_defaults[4] gpio_defaults_block_24/gpio_defaults[5]
+ gpio_defaults_block_24/gpio_defaults[6] gpio_defaults_block_24/gpio_defaults[7]
+ gpio_defaults_block_24/gpio_defaults[8] gpio_defaults_block_24/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[14\] soc/VDD soc/VSS gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[1]
+ gpio_defaults_block_27/gpio_defaults[2] gpio_defaults_block_27/gpio_defaults[3]
+ gpio_defaults_block_27/gpio_defaults[4] gpio_defaults_block_27/gpio_defaults[5]
+ gpio_defaults_block_27/gpio_defaults[6] gpio_defaults_block_27/gpio_defaults[7]
+ gpio_defaults_block_27/gpio_defaults[8] gpio_defaults_block_27/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[33] gpio_control_in_2\[14\]/zero housekeeping/mgmt_gpio_out[33]
+ gpio_control_in_2\[14\]/one padframe/mprj_io_drive_sel[66] padframe/mprj_io_drive_sel[67]
+ padframe/mprj_io_in[33] padframe/mprj_io_inen[33] padframe/mprj_io_out[33] padframe/mprj_io_outen[33]
+ padframe/mprj_io_pd_select[33] padframe/mprj_io_pu_select[33] padframe/mprj_io_schmitt_select[33]
+ padframe/mprj_io_slew_select[33] gpio_control_in_2\[14\]/resetn gpio_control_in_2\[13\]/resetn
+ gpio_control_in_2\[14\]/serial_clock gpio_control_in_2\[13\]/serial_clock gpio_control_in_2\[14\]/serial_data_in
+ gpio_control_in_2\[13\]/serial_data_in gpio_control_in_2\[14\]/serial_load gpio_control_in_2\[13\]/serial_load
+ mprj/io_in[33] mprj/io_oeb[33] mprj/io_out[33] gpio_control_in_2\[14\]/zero gpio_control_block
Xgpio_control_in_1a\[3\] soc/VDD soc/VSS gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[1]
+ gpio_defaults_block_28/gpio_defaults[2] gpio_defaults_block_28/gpio_defaults[3]
+ gpio_defaults_block_28/gpio_defaults[4] gpio_defaults_block_28/gpio_defaults[5]
+ gpio_defaults_block_28/gpio_defaults[6] gpio_defaults_block_28/gpio_defaults[7]
+ gpio_defaults_block_28/gpio_defaults[8] gpio_defaults_block_28/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[5] gpio_control_in_1a\[3\]/zero housekeeping/mgmt_gpio_out[5]
+ gpio_control_in_1a\[3\]/one padframe/mprj_io_drive_sel[11] padframe/mprj_io_drive_sel[10]
+ padframe/mprj_io_in[5] padframe/mprj_io_inen[5] padframe/mprj_io_out[5] padframe/mprj_io_outen[5]
+ padframe/mprj_io_pd_select[5] padframe/mprj_io_pu_select[5] padframe/mprj_io_schmitt_select[5]
+ padframe/mprj_io_slew_select[5] gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[4\]/resetn
+ gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[3\]/serial_data_in
+ gpio_control_in_1a\[4\]/serial_data_in gpio_control_in_1a\[3\]/serial_load gpio_control_in_1a\[4\]/serial_load
+ mprj/io_in[5] mprj/io_oeb[5] mprj/io_out[5] gpio_control_in_1a\[3\]/zero gpio_control_block
Xgpio_control_bidir_2\[0\] soc/VDD soc/VSS gpio_defaults_block_30/gpio_defaults[0]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_oeb[35]
+ housekeeping/mgmt_gpio_out[35] gpio_control_bidir_2\[0\]/one padframe/mprj_io_drive_sel[70]
+ padframe/mprj_io_drive_sel[71] padframe/mprj_io_in[35] padframe/mprj_io_inen[35]
+ padframe/mprj_io_out[35] padframe/mprj_io_outen[35] padframe/mprj_io_pd_select[35]
+ padframe/mprj_io_pu_select[35] padframe/mprj_io_schmitt_select[35] padframe/mprj_io_slew_select[35]
+ gpio_control_bidir_2\[0\]/resetn gpio_control_in_2\[15\]/resetn gpio_control_bidir_2\[0\]/serial_clock
+ gpio_control_in_2\[15\]/serial_clock gpio_control_bidir_2\[0\]/serial_data_in gpio_control_in_2\[15\]/serial_data_in
+ gpio_control_bidir_2\[0\]/serial_load gpio_control_in_2\[15\]/serial_load mprj/io_in[35]
+ mprj/io_oeb[35] mprj/io_out[35] gpio_control_bidir_2\[0\]/zero gpio_control_block
Xsoc soc/VDD soc/VSS soc/core_clk soc/core_rstn soc/debug_in soc/debug_mode soc/debug_oeb
+ soc/debug_out soc/flash_clk soc/flash_csb soc/flash_io0_di soc/flash_io0_do soc/flash_io0_oeb
+ soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb soc/flash_io2_di soc/flash_io2_do
+ soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do soc/flash_io3_oeb soc/gpio_in_pad
+ soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_out_pad soc/gpio_outenb_pad
+ soc/hk_ack_i soc/hk_cyc_o soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11] soc/hk_dat_i[12]
+ soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16] soc/hk_dat_i[17]
+ soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20] soc/hk_dat_i[21]
+ soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25] soc/hk_dat_i[26]
+ soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2] soc/hk_dat_i[30]
+ soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5] soc/hk_dat_i[6]
+ soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] soc/hk_stb_o soc/irq[0] soc/irq[1]
+ soc/irq[2] soc/irq[3] soc/irq[4] soc/irq[5] soc/la_iena[0] soc/la_iena[10] soc/la_iena[11]
+ soc/la_iena[12] soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16]
+ soc/la_iena[17] soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21]
+ soc/la_iena[22] soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26]
+ soc/la_iena[27] soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31]
+ soc/la_iena[32] soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36]
+ soc/la_iena[37] soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41]
+ soc/la_iena[42] soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46]
+ soc/la_iena[47] soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51]
+ soc/la_iena[52] soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56]
+ soc/la_iena[57] soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61]
+ soc/la_iena[62] soc/la_iena[63] soc/la_iena[6] soc/la_iena[7] soc/la_iena[8] soc/la_iena[9]
+ soc/la_input[0] soc/la_input[10] soc/la_input[11] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[6] soc/la_input[7] soc/la_input[8] soc/la_input[9] soc/la_oenb[0] soc/la_oenb[10]
+ soc/la_oenb[11] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14] soc/la_oenb[15]
+ soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19] soc/la_oenb[1] soc/la_oenb[20]
+ soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24] soc/la_oenb[25]
+ soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29] soc/la_oenb[2] soc/la_oenb[30]
+ soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34] soc/la_oenb[35]
+ soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39] soc/la_oenb[3] soc/la_oenb[40]
+ soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44] soc/la_oenb[45]
+ soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49] soc/la_oenb[4] soc/la_oenb[50]
+ soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54] soc/la_oenb[55]
+ soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59] soc/la_oenb[5] soc/la_oenb[60]
+ soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[6] soc/la_oenb[7] soc/la_oenb[8]
+ soc/la_oenb[9] soc/la_output[0] soc/la_output[10] soc/la_output[11] soc/la_output[12]
+ soc/la_output[13] soc/la_output[14] soc/la_output[15] soc/la_output[16] soc/la_output[17]
+ soc/la_output[18] soc/la_output[19] soc/la_output[1] soc/la_output[20] soc/la_output[21]
+ soc/la_output[22] soc/la_output[23] soc/la_output[24] soc/la_output[25] soc/la_output[26]
+ soc/la_output[27] soc/la_output[28] soc/la_output[29] soc/la_output[2] soc/la_output[30]
+ soc/la_output[31] soc/la_output[32] soc/la_output[33] soc/la_output[34] soc/la_output[35]
+ soc/la_output[36] soc/la_output[37] soc/la_output[38] soc/la_output[39] soc/la_output[3]
+ soc/la_output[40] soc/la_output[41] soc/la_output[42] soc/la_output[43] soc/la_output[44]
+ soc/la_output[45] soc/la_output[46] soc/la_output[47] soc/la_output[48] soc/la_output[49]
+ soc/la_output[4] soc/la_output[50] soc/la_output[51] soc/la_output[52] soc/la_output[53]
+ soc/la_output[54] soc/la_output[55] soc/la_output[56] soc/la_output[57] soc/la_output[58]
+ soc/la_output[59] soc/la_output[5] soc/la_output[60] soc/la_output[61] soc/la_output[62]
+ soc/la_output[63] soc/la_output[6] soc/la_output[7] soc/la_output[8] soc/la_output[9]
+ soc/mprj_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12]
+ soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17]
+ soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21]
+ soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26]
+ soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30]
+ soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6]
+ soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/mprj_cyc_o soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12]
+ soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17]
+ soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21]
+ soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26]
+ soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30]
+ soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6]
+ soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/mprj_stb_o soc/mprj_wb_iena soc/mprj_we_o
+ soc/qspi_enabled soc/ser_rx soc/ser_tx soc/spi_csb soc/spi_enabled soc/spi_sck soc/spi_sdi
+ soc/spi_sdo soc/spi_sdoenb soc/trap soc/uart_enabled soc/user_irq_ena[0] soc/user_irq_ena[1]
+ soc/user_irq_ena[2] mgmt_core_wrapper
Xgpio_defaults_block_14 gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[1]
+ gpio_defaults_block_14/gpio_defaults[2] gpio_defaults_block_14/gpio_defaults[3]
+ gpio_defaults_block_14/gpio_defaults[4] gpio_defaults_block_14/gpio_defaults[5]
+ gpio_defaults_block_14/gpio_defaults[6] gpio_defaults_block_14/gpio_defaults[7]
+ gpio_defaults_block_14/gpio_defaults[8] gpio_defaults_block_14/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[9\] soc/VDD soc/VSS gpio_defaults_block_18/gpio_defaults[0] gpio_defaults_block_18/gpio_defaults[1]
+ gpio_defaults_block_18/gpio_defaults[2] gpio_defaults_block_18/gpio_defaults[3]
+ gpio_defaults_block_18/gpio_defaults[4] gpio_defaults_block_18/gpio_defaults[5]
+ gpio_defaults_block_18/gpio_defaults[6] gpio_defaults_block_18/gpio_defaults[7]
+ gpio_defaults_block_18/gpio_defaults[8] gpio_defaults_block_18/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[28] gpio_control_in_2\[9\]/zero housekeeping/mgmt_gpio_out[28]
+ gpio_control_in_2\[9\]/one padframe/mprj_io_drive_sel[56] padframe/mprj_io_drive_sel[57]
+ padframe/mprj_io_in[28] padframe/mprj_io_inen[28] padframe/mprj_io_out[28] padframe/mprj_io_outen[28]
+ padframe/mprj_io_pd_select[28] padframe/mprj_io_pu_select[28] padframe/mprj_io_schmitt_select[28]
+ padframe/mprj_io_slew_select[28] gpio_control_in_2\[9\]/resetn gpio_control_in_2\[8\]/resetn
+ gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[9\]/serial_data_in
+ gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[9\]/serial_load gpio_control_in_2\[8\]/serial_load
+ mprj/io_in[28] mprj/io_oeb[28] mprj/io_out[28] gpio_control_in_2\[9\]/zero gpio_control_block
Xgpio_defaults_block_25 gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[1]
+ gpio_defaults_block_25/gpio_defaults[2] gpio_defaults_block_25/gpio_defaults[3]
+ gpio_defaults_block_25/gpio_defaults[4] gpio_defaults_block_25/gpio_defaults[5]
+ gpio_defaults_block_25/gpio_defaults[6] gpio_defaults_block_25/gpio_defaults[7]
+ gpio_defaults_block_25/gpio_defaults[8] gpio_defaults_block_25/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xsimple_por_0 soc/VDD soc/VSS simple_por_0/porb simple_por_0/por simple_por
Xgpio_control_in_1\[4\] soc/VDD soc/VSS gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[1]
+ gpio_defaults_block_11/gpio_defaults[2] gpio_defaults_block_11/gpio_defaults[3]
+ gpio_defaults_block_11/gpio_defaults[4] gpio_defaults_block_11/gpio_defaults[5]
+ gpio_defaults_block_11/gpio_defaults[6] gpio_defaults_block_11/gpio_defaults[7]
+ gpio_defaults_block_11/gpio_defaults[8] gpio_defaults_block_11/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[12] gpio_control_in_1\[4\]/zero housekeeping/mgmt_gpio_out[12]
+ gpio_control_in_1\[4\]/one padframe/mprj_io_drive_sel[25] padframe/mprj_io_drive_sel[24]
+ padframe/mprj_io_in[12] padframe/mprj_io_inen[12] padframe/mprj_io_out[12] padframe/mprj_io_outen[12]
+ padframe/mprj_io_pd_select[12] padframe/mprj_io_pu_select[12] padframe/mprj_io_schmitt_select[12]
+ padframe/mprj_io_slew_select[12] gpio_control_in_1\[4\]/resetn gpio_control_in_1\[5\]/resetn
+ gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[4\]/serial_data_in
+ gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[4\]/serial_load gpio_control_in_1\[5\]/serial_load
+ mprj/io_in[12] mprj/io_oeb[12] mprj/io_out[12] gpio_control_in_1\[4\]/zero gpio_control_block
Xgpio_defaults_block_15 gpio_defaults_block_15/gpio_defaults[0] gpio_defaults_block_15/gpio_defaults[1]
+ gpio_defaults_block_15/gpio_defaults[2] gpio_defaults_block_15/gpio_defaults[3]
+ gpio_defaults_block_15/gpio_defaults[4] gpio_defaults_block_15/gpio_defaults[5]
+ gpio_defaults_block_15/gpio_defaults[6] gpio_defaults_block_15/gpio_defaults[7]
+ gpio_defaults_block_15/gpio_defaults[8] gpio_defaults_block_15/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_26 gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[1]
+ gpio_defaults_block_26/gpio_defaults[2] gpio_defaults_block_26/gpio_defaults[3]
+ gpio_defaults_block_26/gpio_defaults[4] gpio_defaults_block_26/gpio_defaults[5]
+ gpio_defaults_block_26/gpio_defaults[6] gpio_defaults_block_26/gpio_defaults[7]
+ gpio_defaults_block_26/gpio_defaults[8] gpio_defaults_block_26/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_16 gpio_defaults_block_16/gpio_defaults[0] gpio_defaults_block_16/gpio_defaults[1]
+ gpio_defaults_block_16/gpio_defaults[2] gpio_defaults_block_16/gpio_defaults[3]
+ gpio_defaults_block_16/gpio_defaults[4] gpio_defaults_block_16/gpio_defaults[5]
+ gpio_defaults_block_16/gpio_defaults[6] gpio_defaults_block_16/gpio_defaults[7]
+ gpio_defaults_block_16/gpio_defaults[8] gpio_defaults_block_16/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[12\] soc/VDD soc/VSS gpio_defaults_block_22/gpio_defaults[0] gpio_defaults_block_22/gpio_defaults[1]
+ gpio_defaults_block_22/gpio_defaults[2] gpio_defaults_block_22/gpio_defaults[3]
+ gpio_defaults_block_22/gpio_defaults[4] gpio_defaults_block_22/gpio_defaults[5]
+ gpio_defaults_block_22/gpio_defaults[6] gpio_defaults_block_22/gpio_defaults[7]
+ gpio_defaults_block_22/gpio_defaults[8] gpio_defaults_block_22/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[31] gpio_control_in_2\[12\]/zero housekeeping/mgmt_gpio_out[31]
+ gpio_control_in_2\[12\]/one padframe/mprj_io_drive_sel[62] padframe/mprj_io_drive_sel[63]
+ padframe/mprj_io_in[31] padframe/mprj_io_inen[31] padframe/mprj_io_out[31] padframe/mprj_io_outen[31]
+ padframe/mprj_io_pd_select[31] padframe/mprj_io_pu_select[31] padframe/mprj_io_schmitt_select[31]
+ padframe/mprj_io_slew_select[31] gpio_control_in_2\[12\]/resetn gpio_control_in_2\[11\]/resetn
+ gpio_control_in_2\[12\]/serial_clock gpio_control_in_2\[11\]/serial_clock gpio_control_in_2\[12\]/serial_data_in
+ gpio_control_in_2\[11\]/serial_data_in gpio_control_in_2\[12\]/serial_load gpio_control_in_2\[11\]/serial_load
+ mprj/io_in[31] mprj/io_oeb[31] mprj/io_out[31] gpio_control_in_2\[12\]/zero gpio_control_block
Xgpio_defaults_block_27 gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[1]
+ gpio_defaults_block_27/gpio_defaults[2] gpio_defaults_block_27/gpio_defaults[3]
+ gpio_defaults_block_27/gpio_defaults[4] gpio_defaults_block_27/gpio_defaults[5]
+ gpio_defaults_block_27/gpio_defaults[6] gpio_defaults_block_27/gpio_defaults[7]
+ gpio_defaults_block_27/gpio_defaults[8] gpio_defaults_block_27/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1a\[1\] soc/VDD soc/VSS gpio_control_in_1a\[1\]/gpio_defaults[0]
+ gpio_control_in_1a\[1\]/gpio_defaults[1] gpio_control_in_1a\[1\]/gpio_defaults[2]
+ gpio_control_in_1a\[1\]/gpio_defaults[3] gpio_control_in_1a\[1\]/gpio_defaults[4]
+ gpio_control_in_1a\[1\]/gpio_defaults[5] gpio_control_in_1a\[1\]/gpio_defaults[6]
+ gpio_control_in_1a\[1\]/gpio_defaults[7] gpio_control_in_1a\[1\]/gpio_defaults[8]
+ gpio_control_in_1a\[1\]/gpio_defaults[9] housekeeping/mgmt_gpio_in[3] gpio_control_in_1a\[1\]/zero
+ housekeeping/mgmt_gpio_out[3] gpio_control_in_1a\[1\]/one padframe/mprj_io_drive_sel[7]
+ padframe/mprj_io_drive_sel[6] padframe/mprj_io_in[3] padframe/mprj_io_inen[3] padframe/mprj_io_out[3]
+ padframe/mprj_io_outen[3] padframe/mprj_io_pd_select[3] padframe/mprj_io_pu_select[3]
+ padframe/mprj_io_schmitt_select[3] padframe/mprj_io_slew_select[3] gpio_control_in_1a\[1\]/resetn
+ gpio_control_in_1a\[2\]/resetn gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[2\]/serial_clock
+ gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[1\]/serial_load
+ gpio_control_in_1a\[2\]/serial_load mprj/io_in[3] mprj/io_oeb[3] mprj/io_out[3]
+ gpio_control_in_1a\[1\]/zero gpio_control_block
Xclock_ctrl soc/VDD soc/VSS soc/core_clk pll/osc clock_ctrl/ext_clk_sel housekeeping/reset
+ pll/clockp[1] pll/clockp[0] pll/resetb soc/core_rstn clock_ctrl/sel2[0] clock_ctrl/sel2[1]
+ clock_ctrl/sel2[2] clock_ctrl/sel[0] clock_ctrl/sel[1] clock_ctrl/sel[2] clock_ctrl/user_clk
+ caravel_clocking
Xgpio_control_in_2\[7\] soc/VDD soc/VSS gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[1]
+ gpio_defaults_block_13/gpio_defaults[2] gpio_defaults_block_13/gpio_defaults[3]
+ gpio_defaults_block_13/gpio_defaults[4] gpio_defaults_block_13/gpio_defaults[5]
+ gpio_defaults_block_13/gpio_defaults[6] gpio_defaults_block_13/gpio_defaults[7]
+ gpio_defaults_block_13/gpio_defaults[8] gpio_defaults_block_13/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[26] gpio_control_in_2\[7\]/zero housekeeping/mgmt_gpio_out[26]
+ gpio_control_in_2\[7\]/one padframe/mprj_io_drive_sel[52] padframe/mprj_io_drive_sel[53]
+ padframe/mprj_io_in[26] padframe/mprj_io_inen[26] padframe/mprj_io_out[26] padframe/mprj_io_outen[26]
+ padframe/mprj_io_pd_select[26] padframe/mprj_io_pu_select[26] padframe/mprj_io_schmitt_select[26]
+ padframe/mprj_io_slew_select[26] gpio_control_in_2\[7\]/resetn gpio_control_in_2\[6\]/resetn
+ gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[7\]/serial_data_in
+ gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[7\]/serial_load gpio_control_in_2\[6\]/serial_load
+ mprj/io_in[26] mprj/io_oeb[26] mprj/io_out[26] gpio_control_in_2\[7\]/zero gpio_control_block
Xgpio_defaults_block_17 gpio_defaults_block_17/gpio_defaults[0] gpio_defaults_block_17/gpio_defaults[1]
+ gpio_defaults_block_17/gpio_defaults[2] gpio_defaults_block_17/gpio_defaults[3]
+ gpio_defaults_block_17/gpio_defaults[4] gpio_defaults_block_17/gpio_defaults[5]
+ gpio_defaults_block_17/gpio_defaults[6] gpio_defaults_block_17/gpio_defaults[7]
+ gpio_defaults_block_17/gpio_defaults[8] gpio_defaults_block_17/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_28 gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[1]
+ gpio_defaults_block_28/gpio_defaults[2] gpio_defaults_block_28/gpio_defaults[3]
+ gpio_defaults_block_28/gpio_defaults[4] gpio_defaults_block_28/gpio_defaults[5]
+ gpio_defaults_block_28/gpio_defaults[6] gpio_defaults_block_28/gpio_defaults[7]
+ gpio_defaults_block_28/gpio_defaults[8] gpio_defaults_block_28/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1\[2\] soc/VDD soc/VSS gpio_defaults_block_16/gpio_defaults[0] gpio_defaults_block_16/gpio_defaults[1]
+ gpio_defaults_block_16/gpio_defaults[2] gpio_defaults_block_16/gpio_defaults[3]
+ gpio_defaults_block_16/gpio_defaults[4] gpio_defaults_block_16/gpio_defaults[5]
+ gpio_defaults_block_16/gpio_defaults[6] gpio_defaults_block_16/gpio_defaults[7]
+ gpio_defaults_block_16/gpio_defaults[8] gpio_defaults_block_16/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[10] gpio_control_in_1\[2\]/zero housekeeping/mgmt_gpio_out[10]
+ gpio_control_in_1\[2\]/one padframe/mprj_io_drive_sel[21] padframe/mprj_io_drive_sel[20]
+ padframe/mprj_io_in[10] padframe/mprj_io_inen[10] padframe/mprj_io_out[10] padframe/mprj_io_outen[10]
+ padframe/mprj_io_pd_select[10] padframe/mprj_io_pu_select[10] padframe/mprj_io_schmitt_select[10]
+ padframe/mprj_io_slew_select[10] gpio_control_in_1\[2\]/resetn gpio_control_in_1\[3\]/resetn
+ gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[2\]/serial_data_in
+ gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[2\]/serial_load gpio_control_in_1\[3\]/serial_load
+ mprj/io_in[10] mprj/io_oeb[10] mprj/io_out[10] gpio_control_in_1\[2\]/zero gpio_control_block
Xgpio_defaults_block_18 gpio_defaults_block_18/gpio_defaults[0] gpio_defaults_block_18/gpio_defaults[1]
+ gpio_defaults_block_18/gpio_defaults[2] gpio_defaults_block_18/gpio_defaults[3]
+ gpio_defaults_block_18/gpio_defaults[4] gpio_defaults_block_18/gpio_defaults[5]
+ gpio_defaults_block_18/gpio_defaults[6] gpio_defaults_block_18/gpio_defaults[7]
+ gpio_defaults_block_18/gpio_defaults[8] gpio_defaults_block_18/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_19 gpio_defaults_block_19/gpio_defaults[0] gpio_defaults_block_19/gpio_defaults[1]
+ gpio_defaults_block_19/gpio_defaults[2] gpio_defaults_block_19/gpio_defaults[3]
+ gpio_defaults_block_19/gpio_defaults[4] gpio_defaults_block_19/gpio_defaults[5]
+ gpio_defaults_block_19/gpio_defaults[6] gpio_defaults_block_19/gpio_defaults[7]
+ gpio_defaults_block_19/gpio_defaults[8] gpio_defaults_block_19/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_29 gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[1]
+ gpio_defaults_block_29/gpio_defaults[2] gpio_defaults_block_29/gpio_defaults[3]
+ gpio_defaults_block_29/gpio_defaults[4] gpio_defaults_block_29/gpio_defaults[5]
+ gpio_defaults_block_29/gpio_defaults[6] gpio_defaults_block_29/gpio_defaults[7]
+ gpio_defaults_block_29/gpio_defaults[8] gpio_defaults_block_29/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[10\] soc/VDD soc/VSS gpio_defaults_block_17/gpio_defaults[0] gpio_defaults_block_17/gpio_defaults[1]
+ gpio_defaults_block_17/gpio_defaults[2] gpio_defaults_block_17/gpio_defaults[3]
+ gpio_defaults_block_17/gpio_defaults[4] gpio_defaults_block_17/gpio_defaults[5]
+ gpio_defaults_block_17/gpio_defaults[6] gpio_defaults_block_17/gpio_defaults[7]
+ gpio_defaults_block_17/gpio_defaults[8] gpio_defaults_block_17/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[29] gpio_control_in_2\[10\]/zero housekeeping/mgmt_gpio_out[29]
+ gpio_control_in_2\[10\]/one padframe/mprj_io_drive_sel[58] padframe/mprj_io_drive_sel[59]
+ padframe/mprj_io_in[29] padframe/mprj_io_inen[29] padframe/mprj_io_out[29] padframe/mprj_io_outen[29]
+ padframe/mprj_io_pd_select[29] padframe/mprj_io_pu_select[29] padframe/mprj_io_schmitt_select[29]
+ padframe/mprj_io_slew_select[29] gpio_control_in_2\[10\]/resetn gpio_control_in_2\[9\]/resetn
+ gpio_control_in_2\[10\]/serial_clock gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[10\]/serial_data_in
+ gpio_control_in_2\[9\]/serial_data_in gpio_control_in_2\[10\]/serial_load gpio_control_in_2\[9\]/serial_load
+ mprj/io_in[29] mprj/io_oeb[29] mprj/io_out[29] gpio_control_in_2\[10\]/zero gpio_control_block
Xgpio_defaults_block_0 gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[1]
+ gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3] gpio_defaults_block_0/gpio_defaults[4]
+ gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6] gpio_defaults_block_0/gpio_defaults[7]
+ gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9] gpio_defaults_block_0/VDD
+ gpio_defaults_block_0/VSS gpio_defaults_block
Xgpio_control_in_1\[10\] soc/VDD soc/VSS gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[1]
+ gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3] gpio_defaults_block_4/gpio_defaults[4]
+ gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6] gpio_defaults_block_4/gpio_defaults[7]
+ gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9] housekeeping/mgmt_gpio_in[18]
+ gpio_control_in_1\[10\]/zero housekeeping/mgmt_gpio_out[18] gpio_control_in_1\[10\]/one
+ padframe/mprj_io_drive_sel[36] padframe/mprj_io_drive_sel[37] padframe/mprj_io_in[18]
+ padframe/mprj_io_inen[18] padframe/mprj_io_out[18] padframe/mprj_io_outen[18] padframe/mprj_io_pd_select[18]
+ padframe/mprj_io_pu_select[18] padframe/mprj_io_schmitt_select[18] padframe/mprj_io_slew_select[18]
+ gpio_control_in_1\[10\]/resetn gpio_control_in_1\[10\]/resetn_out gpio_control_in_1\[10\]/serial_clock
+ gpio_control_in_1\[10\]/serial_clock_out gpio_control_in_1\[9\]/serial_data_out
+ gpio_control_in_1\[10\]/serial_data_out gpio_control_in_1\[10\]/serial_load gpio_control_in_1\[10\]/serial_load_out
+ mprj/io_in[18] mprj/io_oeb[18] mprj/io_out[18] gpio_control_in_1\[10\]/zero gpio_control_block
Xgpio_control_in_2\[5\] soc/VDD soc/VSS gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[1]
+ gpio_defaults_block_10/gpio_defaults[2] gpio_defaults_block_10/gpio_defaults[3]
+ gpio_defaults_block_10/gpio_defaults[4] gpio_defaults_block_10/gpio_defaults[5]
+ gpio_defaults_block_10/gpio_defaults[6] gpio_defaults_block_10/gpio_defaults[7]
+ gpio_defaults_block_10/gpio_defaults[8] gpio_defaults_block_10/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[24] gpio_control_in_2\[5\]/zero housekeeping/mgmt_gpio_out[24]
+ gpio_control_in_2\[5\]/one padframe/mprj_io_drive_sel[48] padframe/mprj_io_drive_sel[49]
+ padframe/mprj_io_in[24] padframe/mprj_io_inen[24] padframe/mprj_io_out[24] padframe/mprj_io_outen[24]
+ padframe/mprj_io_pd_select[24] padframe/mprj_io_pu_select[24] padframe/mprj_io_schmitt_select[24]
+ padframe/mprj_io_slew_select[24] gpio_control_in_2\[5\]/resetn gpio_control_in_2\[4\]/resetn
+ gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[4\]/serial_clock gpio_control_in_2\[5\]/serial_data_in
+ gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[5\]/serial_load gpio_control_in_2\[4\]/serial_load
+ mprj/io_in[24] mprj/io_oeb[24] mprj/io_out[24] gpio_control_in_2\[5\]/zero gpio_control_block
Xgpio_control_in_1\[0\] soc/VDD soc/VSS gpio_defaults_block_21/gpio_defaults[0] gpio_defaults_block_21/gpio_defaults[1]
+ gpio_defaults_block_21/gpio_defaults[2] gpio_defaults_block_21/gpio_defaults[3]
+ gpio_defaults_block_21/gpio_defaults[4] gpio_defaults_block_21/gpio_defaults[5]
+ gpio_defaults_block_21/gpio_defaults[6] gpio_defaults_block_21/gpio_defaults[7]
+ gpio_defaults_block_21/gpio_defaults[8] gpio_defaults_block_21/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[8] gpio_control_in_1\[0\]/zero housekeeping/mgmt_gpio_out[8]
+ gpio_control_in_1\[0\]/one padframe/mprj_io_drive_sel[17] padframe/mprj_io_drive_sel[16]
+ padframe/mprj_io_in[8] padframe/mprj_io_inen[8] padframe/mprj_io_out[8] padframe/mprj_io_outen[8]
+ padframe/mprj_io_pd_select[8] padframe/mprj_io_pu_select[8] padframe/mprj_io_schmitt_select[8]
+ padframe/mprj_io_slew_select[8] gpio_control_in_1\[0\]/resetn gpio_control_in_1\[1\]/resetn
+ gpio_control_in_1\[0\]/serial_clock gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[0\]/serial_data_in
+ gpio_control_in_1\[1\]/serial_data_in gpio_control_in_1\[0\]/serial_load gpio_control_in_1\[1\]/serial_load
+ mprj/io_in[8] mprj/io_oeb[8] mprj/io_out[8] gpio_control_in_1\[0\]/zero gpio_control_block
Xgpio_defaults_block_1 gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[1]
+ gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3] gpio_defaults_block_1/gpio_defaults[4]
+ gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6] gpio_defaults_block_1/gpio_defaults[7]
+ gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9] soc/VDD
+ soc/VSS gpio_defaults_block
Xspare_logic\[3\] soc/VDD soc/VSS spare_logic\[3\]/spare_xfq[0] spare_logic\[3\]/spare_xfq[1]
+ spare_logic\[3\]/spare_xi[0] spare_logic\[3\]/spare_xi[1] spare_logic\[3\]/spare_xi[2]
+ spare_logic\[3\]/spare_xi[3] spare_logic\[3\]/spare_xib spare_logic\[3\]/spare_xmx[0]
+ spare_logic\[3\]/spare_xmx[1] spare_logic\[3\]/spare_xna[0] spare_logic\[3\]/spare_xna[1]
+ spare_logic\[3\]/spare_xno[0] spare_logic\[3\]/spare_xno[1] spare_logic\[3\]/spare_xz[0]
+ spare_logic\[3\]/spare_xz[10] spare_logic\[3\]/spare_xz[11] spare_logic\[3\]/spare_xz[12]
+ spare_logic\[3\]/spare_xz[13] spare_logic\[3\]/spare_xz[14] spare_logic\[3\]/spare_xz[15]
+ spare_logic\[3\]/spare_xz[16] spare_logic\[3\]/spare_xz[17] spare_logic\[3\]/spare_xz[18]
+ spare_logic\[3\]/spare_xz[19] spare_logic\[3\]/spare_xz[1] spare_logic\[3\]/spare_xz[20]
+ spare_logic\[3\]/spare_xz[21] spare_logic\[3\]/spare_xz[22] spare_logic\[3\]/spare_xz[23]
+ spare_logic\[3\]/spare_xz[24] spare_logic\[3\]/spare_xz[25] spare_logic\[3\]/spare_xz[26]
+ spare_logic\[3\]/spare_xz[27] spare_logic\[3\]/spare_xz[28] spare_logic\[3\]/spare_xz[29]
+ spare_logic\[3\]/spare_xz[2] spare_logic\[3\]/spare_xz[30] spare_logic\[3\]/spare_xz[3]
+ spare_logic\[3\]/spare_xz[4] spare_logic\[3\]/spare_xz[5] spare_logic\[3\]/spare_xz[6]
+ spare_logic\[3\]/spare_xz[7] spare_logic\[3\]/spare_xz[8] spare_logic\[3\]/spare_xz[9]
+ spare_logic_block
Xuser_id_value user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ user_id_value/VDD user_id_value/VSS user_id_programming
Xgpio_defaults_block_2 gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[1]
+ gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3] gpio_defaults_block_2/gpio_defaults[4]
+ gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6] gpio_defaults_block_2/gpio_defaults[7]
+ gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9] gpio_defaults_block_2/VDD
+ gpio_defaults_block_2/VSS gpio_defaults_block
Xgpio_control_in_2\[3\] soc/VDD soc/VSS gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[1]
+ gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3] gpio_defaults_block_9/gpio_defaults[4]
+ gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6] gpio_defaults_block_9/gpio_defaults[7]
+ gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9] housekeeping/mgmt_gpio_in[22]
+ gpio_control_in_2\[3\]/zero housekeeping/mgmt_gpio_out[22] gpio_control_in_2\[3\]/one
+ padframe/mprj_io_drive_sel[44] padframe/mprj_io_drive_sel[45] padframe/mprj_io_in[22]
+ padframe/mprj_io_inen[22] padframe/mprj_io_out[22] padframe/mprj_io_outen[22] padframe/mprj_io_pd_select[22]
+ padframe/mprj_io_pu_select[22] padframe/mprj_io_schmitt_select[22] padframe/mprj_io_slew_select[22]
+ gpio_control_in_2\[3\]/resetn gpio_control_in_2\[2\]/resetn gpio_control_in_2\[3\]/serial_clock
+ gpio_control_in_2\[2\]/serial_clock gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[2\]/serial_data_in
+ gpio_control_in_2\[3\]/serial_load gpio_control_in_2\[2\]/serial_load mprj/io_in[22]
+ mprj/io_oeb[22] mprj/io_out[22] gpio_control_in_2\[3\]/zero gpio_control_block
Xgpio_defaults_block_3 gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[1]
+ gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3] gpio_defaults_block_3/gpio_defaults[4]
+ gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6] gpio_defaults_block_3/gpio_defaults[7]
+ gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9] gpio_defaults_block_3/VDD
+ gpio_defaults_block_3/VSS gpio_defaults_block
Xgpio_control_bidir_1\[0\] soc/VDD soc/VSS gpio_defaults_block_009_1/gpio_defaults[0]
+ gpio_defaults_block_009_1/gpio_defaults[1] gpio_defaults_block_009_1/gpio_defaults[2]
+ gpio_defaults_block_009_1/gpio_defaults[3] gpio_defaults_block_009_1/gpio_defaults[4]
+ gpio_defaults_block_009_1/gpio_defaults[5] gpio_defaults_block_009_1/gpio_defaults[6]
+ gpio_defaults_block_009_1/gpio_defaults[7] gpio_defaults_block_009_1/gpio_defaults[8]
+ gpio_defaults_block_009_1/gpio_defaults[9] housekeeping/mgmt_gpio_in[0] housekeeping/mgmt_gpio_oeb[0]
+ housekeeping/mgmt_gpio_out[0] gpio_control_bidir_1\[0\]/one padframe/mprj_io_drive_sel[0]
+ padframe/mprj_io_drive_sel[1] padframe/mprj_io_in[0] padframe/mprj_io_inen[0] padframe/mprj_io_out[0]
+ padframe/mprj_io_outen[0] padframe/mprj_io_pd_select[0] padframe/mprj_io_pu_select[0]
+ padframe/mprj_io_schmitt_select[0] padframe/mprj_io_slew_select[0] housekeeping/serial_resetn
+ gpio_control_bidir_1\[1\]/resetn housekeeping/serial_clock gpio_control_bidir_1\[1\]/serial_clock
+ housekeeping/serial_data_1 gpio_control_bidir_1\[1\]/serial_data_in housekeeping/serial_load
+ gpio_control_bidir_1\[1\]/serial_load mprj/io_in[0] mprj/io_oeb[0] mprj/io_out[0]
+ gpio_control_bidir_1\[0\]/zero gpio_control_block
Xgpio_control_in_1\[9\] soc/VDD soc/VSS gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[1]
+ gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3] gpio_defaults_block_3/gpio_defaults[4]
+ gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6] gpio_defaults_block_3/gpio_defaults[7]
+ gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9] housekeeping/mgmt_gpio_in[17]
+ gpio_control_in_1\[9\]/zero housekeeping/mgmt_gpio_out[17] gpio_control_in_1\[9\]/one
+ padframe/mprj_io_drive_sel[34] padframe/mprj_io_drive_sel[35] padframe/mprj_io_in[17]
+ padframe/mprj_io_inen[17] padframe/mprj_io_out[17] padframe/mprj_io_outen[17] padframe/mprj_io_pd_select[17]
+ padframe/mprj_io_pu_select[17] padframe/mprj_io_schmitt_select[17] padframe/mprj_io_slew_select[17]
+ gpio_control_in_1\[9\]/resetn gpio_control_in_1\[10\]/resetn gpio_control_in_1\[9\]/serial_clock
+ gpio_control_in_1\[10\]/serial_clock gpio_control_in_1\[9\]/serial_data_in gpio_control_in_1\[9\]/serial_data_out
+ gpio_control_in_1\[9\]/serial_load gpio_control_in_1\[10\]/serial_load mprj/io_in[17]
+ mprj/io_oeb[17] mprj/io_out[17] gpio_control_in_1\[9\]/zero gpio_control_block
Xgpio_defaults_block_4 gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[1]
+ gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3] gpio_defaults_block_4/gpio_defaults[4]
+ gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6] gpio_defaults_block_4/gpio_defaults[7]
+ gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9] gpio_defaults_block_4/VDD
+ gpio_defaults_block_4/VSS gpio_defaults_block
Xgpio_defaults_block_5 gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[1]
+ gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3] gpio_defaults_block_5/gpio_defaults[4]
+ gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6] gpio_defaults_block_5/gpio_defaults[7]
+ gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9] gpio_defaults_block_5/VDD
+ gpio_defaults_block_5/VSS gpio_defaults_block
Xspare_logic\[1\] soc/VDD soc/VSS spare_logic\[1\]/spare_xfq[0] spare_logic\[1\]/spare_xfq[1]
+ spare_logic\[1\]/spare_xi[0] spare_logic\[1\]/spare_xi[1] spare_logic\[1\]/spare_xi[2]
+ spare_logic\[1\]/spare_xi[3] spare_logic\[1\]/spare_xib spare_logic\[1\]/spare_xmx[0]
+ spare_logic\[1\]/spare_xmx[1] spare_logic\[1\]/spare_xna[0] spare_logic\[1\]/spare_xna[1]
+ spare_logic\[1\]/spare_xno[0] spare_logic\[1\]/spare_xno[1] spare_logic\[1\]/spare_xz[0]
+ spare_logic\[1\]/spare_xz[10] spare_logic\[1\]/spare_xz[11] spare_logic\[1\]/spare_xz[12]
+ spare_logic\[1\]/spare_xz[13] spare_logic\[1\]/spare_xz[14] spare_logic\[1\]/spare_xz[15]
+ spare_logic\[1\]/spare_xz[16] spare_logic\[1\]/spare_xz[17] spare_logic\[1\]/spare_xz[18]
+ spare_logic\[1\]/spare_xz[19] spare_logic\[1\]/spare_xz[1] spare_logic\[1\]/spare_xz[20]
+ spare_logic\[1\]/spare_xz[21] spare_logic\[1\]/spare_xz[22] spare_logic\[1\]/spare_xz[23]
+ spare_logic\[1\]/spare_xz[24] spare_logic\[1\]/spare_xz[25] spare_logic\[1\]/spare_xz[26]
+ spare_logic\[1\]/spare_xz[27] spare_logic\[1\]/spare_xz[28] spare_logic\[1\]/spare_xz[29]
+ spare_logic\[1\]/spare_xz[2] spare_logic\[1\]/spare_xz[30] spare_logic\[1\]/spare_xz[3]
+ spare_logic\[1\]/spare_xz[4] spare_logic\[1\]/spare_xz[5] spare_logic\[1\]/spare_xz[6]
+ spare_logic\[1\]/spare_xz[7] spare_logic\[1\]/spare_xz[8] spare_logic\[1\]/spare_xz[9]
+ spare_logic_block
Xgpio_defaults_block_6 gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[1]
+ gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3] gpio_defaults_block_6/gpio_defaults[4]
+ gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6] gpio_defaults_block_6/gpio_defaults[7]
+ gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9] gpio_defaults_block_6/VDD
+ gpio_defaults_block_6/VSS gpio_defaults_block
Xgpio_control_in_2\[1\] soc/VDD soc/VSS gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[1]
+ gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3] gpio_defaults_block_5/gpio_defaults[4]
+ gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6] gpio_defaults_block_5/gpio_defaults[7]
+ gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9] housekeeping/mgmt_gpio_in[20]
+ gpio_control_in_2\[1\]/zero housekeeping/mgmt_gpio_out[20] gpio_control_in_2\[1\]/one
+ padframe/mprj_io_drive_sel[40] padframe/mprj_io_drive_sel[41] padframe/mprj_io_in[20]
+ padframe/mprj_io_inen[20] padframe/mprj_io_out[20] padframe/mprj_io_outen[20] padframe/mprj_io_pd_select[20]
+ padframe/mprj_io_pu_select[20] padframe/mprj_io_schmitt_select[20] padframe/mprj_io_slew_select[20]
+ gpio_control_in_2\[1\]/resetn gpio_control_in_2\[0\]/resetn gpio_control_in_2\[1\]/serial_clock
+ gpio_control_in_2\[0\]/serial_clock gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[0\]/serial_data_in
+ gpio_control_in_2\[1\]/serial_load gpio_control_in_2\[0\]/serial_load mprj/io_in[20]
+ mprj/io_oeb[20] mprj/io_out[20] gpio_control_in_2\[1\]/zero gpio_control_block
Xgpio_defaults_block_7 gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[1]
+ gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3] gpio_defaults_block_7/gpio_defaults[4]
+ gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6] gpio_defaults_block_7/gpio_defaults[7]
+ gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9] gpio_defaults_block_7/VDD
+ gpio_defaults_block_7/VSS gpio_defaults_block
Xgpio_control_in_1\[7\] soc/VDD soc/VSS gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[1]
+ gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3] gpio_defaults_block_0/gpio_defaults[4]
+ gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6] gpio_defaults_block_0/gpio_defaults[7]
+ gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9] housekeeping/mgmt_gpio_in[15]
+ gpio_control_in_1\[7\]/zero housekeeping/mgmt_gpio_out[15] gpio_control_in_1\[7\]/one
+ padframe/mprj_io_drive_sel[30] padframe/mprj_io_drive_sel[31] padframe/mprj_io_in[15]
+ padframe/mprj_io_inen[15] padframe/mprj_io_out[15] padframe/mprj_io_outen[15] padframe/mprj_io_pd_select[15]
+ padframe/mprj_io_pu_select[15] padframe/mprj_io_schmitt_select[15] padframe/mprj_io_slew_select[15]
+ gpio_control_in_1\[7\]/resetn gpio_control_in_1\[8\]/resetn gpio_control_in_1\[7\]/serial_clock
+ gpio_control_in_1\[8\]/serial_clock gpio_control_in_1\[7\]/serial_data_in gpio_control_in_1\[8\]/serial_data_in
+ gpio_control_in_1\[7\]/serial_load gpio_control_in_1\[8\]/serial_load mprj/io_in[15]
+ mprj/io_oeb[15] mprj/io_out[15] gpio_control_in_1\[7\]/zero gpio_control_block
Xgpio_defaults_block_8 gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[1]
+ gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3] gpio_defaults_block_8/gpio_defaults[4]
+ gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6] gpio_defaults_block_8/gpio_defaults[7]
+ gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9] gpio_defaults_block_8/VDD
+ gpio_defaults_block_8/VSS gpio_defaults_block
Xgpio_control_in_1a\[4\] soc/VDD soc/VSS gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[1]
+ gpio_defaults_block_26/gpio_defaults[2] gpio_defaults_block_26/gpio_defaults[3]
+ gpio_defaults_block_26/gpio_defaults[4] gpio_defaults_block_26/gpio_defaults[5]
+ gpio_defaults_block_26/gpio_defaults[6] gpio_defaults_block_26/gpio_defaults[7]
+ gpio_defaults_block_26/gpio_defaults[8] gpio_defaults_block_26/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[6] gpio_control_in_1a\[4\]/zero housekeeping/mgmt_gpio_out[6]
+ gpio_control_in_1a\[4\]/one padframe/mprj_io_drive_sel[13] padframe/mprj_io_drive_sel[12]
+ padframe/mprj_io_in[6] padframe/mprj_io_inen[6] padframe/mprj_io_out[6] padframe/mprj_io_outen[6]
+ padframe/mprj_io_pd_select[6] padframe/mprj_io_pu_select[6] padframe/mprj_io_schmitt_select[6]
+ padframe/mprj_io_slew_select[6] gpio_control_in_1a\[4\]/resetn gpio_control_in_1a\[5\]/resetn
+ gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1a\[4\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1a\[4\]/serial_load gpio_control_in_1a\[5\]/serial_load
+ mprj/io_in[6] mprj/io_oeb[6] mprj/io_out[6] gpio_control_in_1a\[4\]/zero gpio_control_block
Xmgmt_buffers soc/VDD soc/VSS soc/core_clk clock_ctrl/user_clk soc/core_rstn mprj/la_data_in[0]
+ mprj/la_data_in[10] mprj/la_data_in[11] mprj/la_data_in[12] mprj/la_data_in[13]
+ mprj/la_data_in[14] mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17]
+ mprj/la_data_in[18] mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21]
+ mprj/la_data_in[22] mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25]
+ mprj/la_data_in[26] mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29]
+ mprj/la_data_in[2] mprj/la_data_in[30] mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33]
+ mprj/la_data_in[34] mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37]
+ mprj/la_data_in[38] mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41]
+ mprj/la_data_in[42] mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45]
+ mprj/la_data_in[46] mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49]
+ mprj/la_data_in[4] mprj/la_data_in[50] mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53]
+ mprj/la_data_in[54] mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57]
+ mprj/la_data_in[58] mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61]
+ mprj/la_data_in[62] mprj/la_data_in[63] mprj/la_data_in[6] mprj/la_data_in[7] mprj/la_data_in[8]
+ mprj/la_data_in[9] soc/la_input[0] soc/la_input[10] soc/la_input[11] soc/la_input[12]
+ soc/la_input[13] soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17]
+ soc/la_input[18] soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21]
+ soc/la_input[22] soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26]
+ soc/la_input[27] soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30]
+ soc/la_input[31] soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35]
+ soc/la_input[36] soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3]
+ soc/la_input[40] soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44]
+ soc/la_input[45] soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49]
+ soc/la_input[4] soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53]
+ soc/la_input[54] soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58]
+ soc/la_input[59] soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62]
+ soc/la_input[63] soc/la_input[6] soc/la_input[7] soc/la_input[8] soc/la_input[9]
+ mprj/la_data_out[0] mprj/la_data_out[10] mprj/la_data_out[11] mprj/la_data_out[12]
+ mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16]
+ mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1]
+ mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23]
+ mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27]
+ mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30]
+ mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34]
+ mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38]
+ mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41]
+ mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45]
+ mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49]
+ mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52]
+ mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56]
+ mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5]
+ mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63]
+ mprj/la_data_out[6] mprj/la_data_out[7] mprj/la_data_out[8] mprj/la_data_out[9]
+ soc/la_output[0] soc/la_output[10] soc/la_output[11] soc/la_output[12] soc/la_output[13]
+ soc/la_output[14] soc/la_output[15] soc/la_output[16] soc/la_output[17] soc/la_output[18]
+ soc/la_output[19] soc/la_output[1] soc/la_output[20] soc/la_output[21] soc/la_output[22]
+ soc/la_output[23] soc/la_output[24] soc/la_output[25] soc/la_output[26] soc/la_output[27]
+ soc/la_output[28] soc/la_output[29] soc/la_output[2] soc/la_output[30] soc/la_output[31]
+ soc/la_output[32] soc/la_output[33] soc/la_output[34] soc/la_output[35] soc/la_output[36]
+ soc/la_output[37] soc/la_output[38] soc/la_output[39] soc/la_output[3] soc/la_output[40]
+ soc/la_output[41] soc/la_output[42] soc/la_output[43] soc/la_output[44] soc/la_output[45]
+ soc/la_output[46] soc/la_output[47] soc/la_output[48] soc/la_output[49] soc/la_output[4]
+ soc/la_output[50] soc/la_output[51] soc/la_output[52] soc/la_output[53] soc/la_output[54]
+ soc/la_output[55] soc/la_output[56] soc/la_output[57] soc/la_output[58] soc/la_output[59]
+ soc/la_output[5] soc/la_output[60] soc/la_output[61] soc/la_output[62] soc/la_output[63]
+ soc/la_output[6] soc/la_output[7] soc/la_output[8] soc/la_output[9] soc/la_iena[0]
+ soc/la_iena[10] soc/la_iena[11] soc/la_iena[12] soc/la_iena[13] soc/la_iena[14]
+ soc/la_iena[15] soc/la_iena[16] soc/la_iena[17] soc/la_iena[18] soc/la_iena[19]
+ soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22] soc/la_iena[23] soc/la_iena[24]
+ soc/la_iena[25] soc/la_iena[26] soc/la_iena[27] soc/la_iena[28] soc/la_iena[29]
+ soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32] soc/la_iena[33] soc/la_iena[34]
+ soc/la_iena[35] soc/la_iena[36] soc/la_iena[37] soc/la_iena[38] soc/la_iena[39]
+ soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42] soc/la_iena[43] soc/la_iena[44]
+ soc/la_iena[45] soc/la_iena[46] soc/la_iena[47] soc/la_iena[48] soc/la_iena[49]
+ soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52] soc/la_iena[53] soc/la_iena[54]
+ soc/la_iena[55] soc/la_iena[56] soc/la_iena[57] soc/la_iena[58] soc/la_iena[59]
+ soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62] soc/la_iena[63] soc/la_iena[6]
+ soc/la_iena[7] soc/la_iena[8] soc/la_iena[9] mprj/la_oenb[0] mprj/la_oenb[10] mprj/la_oenb[11]
+ mprj/la_oenb[12] mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16]
+ mprj/la_oenb[17] mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20]
+ mprj/la_oenb[21] mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25]
+ mprj/la_oenb[26] mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2]
+ mprj/la_oenb[30] mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34]
+ mprj/la_oenb[35] mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39]
+ mprj/la_oenb[3] mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43]
+ mprj/la_oenb[44] mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48]
+ mprj/la_oenb[49] mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52]
+ mprj/la_oenb[53] mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57]
+ mprj/la_oenb[58] mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61]
+ mprj/la_oenb[62] mprj/la_oenb[63] mprj/la_oenb[6] mprj/la_oenb[7] mprj/la_oenb[8]
+ mprj/la_oenb[9] soc/la_oenb[0] soc/la_oenb[10] soc/la_oenb[11] soc/la_oenb[12] soc/la_oenb[13]
+ soc/la_oenb[14] soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18]
+ soc/la_oenb[19] soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23]
+ soc/la_oenb[24] soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28]
+ soc/la_oenb[29] soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33]
+ soc/la_oenb[34] soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38]
+ soc/la_oenb[39] soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43]
+ soc/la_oenb[44] soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48]
+ soc/la_oenb[49] soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53]
+ soc/la_oenb[54] soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58]
+ soc/la_oenb[59] soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63]
+ soc/la_oenb[6] soc/la_oenb[7] soc/la_oenb[8] soc/la_oenb[9] soc/mprj_ack_i mprj/wbs_ack_o
+ soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13]
+ soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18]
+ soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22]
+ soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27]
+ soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31]
+ soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7]
+ soc/mprj_adr_o[8] soc/mprj_adr_o[9] mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11]
+ mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16]
+ mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20]
+ mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25]
+ mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2]
+ mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5]
+ mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] soc/mprj_cyc_o
+ mprj/wbs_cyc_i soc/mprj_dat_i[0] soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12]
+ soc/mprj_dat_i[13] soc/mprj_dat_i[14] soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17]
+ soc/mprj_dat_i[18] soc/mprj_dat_i[19] soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21]
+ soc/mprj_dat_i[22] soc/mprj_dat_i[23] soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26]
+ soc/mprj_dat_i[27] soc/mprj_dat_i[28] soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30]
+ soc/mprj_dat_i[31] soc/mprj_dat_i[3] soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6]
+ soc/mprj_dat_i[7] soc/mprj_dat_i[8] soc/mprj_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10]
+ mprj/wbs_dat_o[11] mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15]
+ mprj/wbs_dat_o[16] mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1]
+ mprj/wbs_dat_o[20] mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24]
+ mprj/wbs_dat_o[25] mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29]
+ mprj/wbs_dat_o[2] mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4]
+ mprj/wbs_dat_o[5] mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9]
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11]
+ mprj/wbs_dat_i[12] mprj/wbs_dat_i[13] mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16]
+ mprj/wbs_dat_i[17] mprj/wbs_dat_i[18] mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20]
+ mprj/wbs_dat_i[21] mprj/wbs_dat_i[22] mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25]
+ mprj/wbs_dat_i[26] mprj/wbs_dat_i[27] mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2]
+ mprj/wbs_dat_i[30] mprj/wbs_dat_i[31] mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5]
+ mprj/wbs_dat_i[6] mprj/wbs_dat_i[7] mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] soc/mprj_wb_iena
+ soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] mprj/wbs_sel_i[0]
+ mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] soc/mprj_stb_o mprj/wbs_stb_i
+ soc/mprj_we_o mprj/wbs_we_i mprj/wb_clk_i mprj/user_clock2 soc/irq[0] soc/irq[1]
+ soc/irq[2] mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] soc/user_irq_ena[0]
+ soc/user_irq_ena[1] soc/user_irq_ena[2] mprj/wb_rst_i mgmt_protect
Xgpio_defaults_block_009_0 gpio_defaults_block_009_0/gpio_defaults[0] gpio_defaults_block_009_0/gpio_defaults[1]
+ gpio_defaults_block_009_0/gpio_defaults[2] gpio_defaults_block_009_0/gpio_defaults[3]
+ gpio_defaults_block_009_0/gpio_defaults[4] gpio_defaults_block_009_0/gpio_defaults[5]
+ gpio_defaults_block_009_0/gpio_defaults[6] gpio_defaults_block_009_0/gpio_defaults[7]
+ gpio_defaults_block_009_0/gpio_defaults[8] gpio_defaults_block_009_0/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_009
Xgpio_defaults_block_009_1 gpio_defaults_block_009_1/gpio_defaults[0] gpio_defaults_block_009_1/gpio_defaults[1]
+ gpio_defaults_block_009_1/gpio_defaults[2] gpio_defaults_block_009_1/gpio_defaults[3]
+ gpio_defaults_block_009_1/gpio_defaults[4] gpio_defaults_block_009_1/gpio_defaults[5]
+ gpio_defaults_block_009_1/gpio_defaults[6] gpio_defaults_block_009_1/gpio_defaults[7]
+ gpio_defaults_block_009_1/gpio_defaults[8] gpio_defaults_block_009_1/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_009
Xgpio_defaults_block_9 gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[1]
+ gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3] gpio_defaults_block_9/gpio_defaults[4]
+ gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6] gpio_defaults_block_9/gpio_defaults[7]
+ gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9] gpio_defaults_block_9/VDD
+ gpio_defaults_block_9/VSS gpio_defaults_block
Xgpio_control_in_2\[15\] soc/VDD soc/VSS gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[1]
+ gpio_defaults_block_29/gpio_defaults[2] gpio_defaults_block_29/gpio_defaults[3]
+ gpio_defaults_block_29/gpio_defaults[4] gpio_defaults_block_29/gpio_defaults[5]
+ gpio_defaults_block_29/gpio_defaults[6] gpio_defaults_block_29/gpio_defaults[7]
+ gpio_defaults_block_29/gpio_defaults[8] gpio_defaults_block_29/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[34] gpio_control_in_2\[15\]/zero housekeeping/mgmt_gpio_out[34]
+ gpio_control_in_2\[15\]/one padframe/mprj_io_drive_sel[68] padframe/mprj_io_drive_sel[69]
+ padframe/mprj_io_in[34] padframe/mprj_io_inen[34] padframe/mprj_io_out[34] padframe/mprj_io_outen[34]
+ padframe/mprj_io_pd_select[34] padframe/mprj_io_pu_select[34] padframe/mprj_io_schmitt_select[34]
+ padframe/mprj_io_slew_select[34] gpio_control_in_2\[15\]/resetn gpio_control_in_2\[14\]/resetn
+ gpio_control_in_2\[15\]/serial_clock gpio_control_in_2\[14\]/serial_clock gpio_control_in_2\[15\]/serial_data_in
+ gpio_control_in_2\[14\]/serial_data_in gpio_control_in_2\[15\]/serial_load gpio_control_in_2\[14\]/serial_load
+ mprj/io_in[34] mprj/io_oeb[34] mprj/io_out[34] gpio_control_in_2\[15\]/zero gpio_control_block
Xgpio_control_bidir_2\[1\] soc/VDD soc/VSS gpio_defaults_block_31/gpio_defaults[0]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] housekeeping/mgmt_gpio_in[36] housekeeping/mgmt_gpio_oeb[36]
+ housekeeping/mgmt_gpio_out[36] gpio_control_bidir_2\[1\]/one padframe/mprj_io_drive_sel[72]
+ padframe/mprj_io_drive_sel[73] padframe/mprj_io_in[36] padframe/mprj_io_inen[36]
+ padframe/mprj_io_out[36] padframe/mprj_io_outen[36] padframe/mprj_io_pd_select[36]
+ padframe/mprj_io_pu_select[36] padframe/mprj_io_schmitt_select[36] padframe/mprj_io_slew_select[36]
+ gpio_control_bidir_2\[1\]/resetn gpio_control_bidir_2\[0\]/resetn gpio_control_bidir_2\[1\]/serial_clock
+ gpio_control_bidir_2\[0\]/serial_clock gpio_control_bidir_2\[1\]/serial_data_in
+ gpio_control_bidir_2\[0\]/serial_data_in gpio_control_bidir_2\[1\]/serial_load gpio_control_bidir_2\[0\]/serial_load
+ mprj/io_in[36] mprj/io_oeb[36] mprj/io_out[36] gpio_control_bidir_2\[1\]/zero gpio_control_block
Xgpio_control_in_1\[5\] soc/VDD soc/VSS gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[1]
+ gpio_defaults_block_12/gpio_defaults[2] gpio_defaults_block_12/gpio_defaults[3]
+ gpio_defaults_block_12/gpio_defaults[4] gpio_defaults_block_12/gpio_defaults[5]
+ gpio_defaults_block_12/gpio_defaults[6] gpio_defaults_block_12/gpio_defaults[7]
+ gpio_defaults_block_12/gpio_defaults[8] gpio_defaults_block_12/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[13] gpio_control_in_1\[5\]/zero housekeeping/mgmt_gpio_out[13]
+ gpio_control_in_1\[5\]/one padframe/mprj_io_drive_sel[26] padframe/mprj_io_drive_sel[27]
+ padframe/mprj_io_in[13] padframe/mprj_io_inen[13] padframe/mprj_io_out[13] padframe/mprj_io_outen[13]
+ padframe/mprj_io_pd_select[13] padframe/mprj_io_pu_select[13] padframe/mprj_io_schmitt_select[13]
+ padframe/mprj_io_slew_select[13] gpio_control_in_1\[5\]/resetn gpio_control_in_1\[6\]/resetn
+ gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[6\]/serial_clock gpio_control_in_1\[5\]/serial_data_in
+ gpio_control_in_1\[6\]/serial_data_in gpio_control_in_1\[5\]/serial_load gpio_control_in_1\[6\]/serial_load
+ mprj/io_in[13] mprj/io_oeb[13] mprj/io_out[13] gpio_control_in_1\[5\]/zero gpio_control_block
Xgpio_defaults_block_007_0 gpio_control_in_1a\[2\]/gpio_defaults[0] gpio_control_in_1a\[2\]/gpio_defaults[1]
+ gpio_control_in_1a\[2\]/gpio_defaults[2] gpio_control_in_1a\[2\]/gpio_defaults[3]
+ gpio_control_in_1a\[2\]/gpio_defaults[4] gpio_control_in_1a\[2\]/gpio_defaults[5]
+ gpio_control_in_1a\[2\]/gpio_defaults[6] gpio_control_in_1a\[2\]/gpio_defaults[7]
+ gpio_control_in_1a\[2\]/gpio_defaults[8] gpio_control_in_1a\[2\]/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_007
Xgpio_control_in_2\[13\] soc/VDD soc/VSS gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[1]
+ gpio_defaults_block_25/gpio_defaults[2] gpio_defaults_block_25/gpio_defaults[3]
+ gpio_defaults_block_25/gpio_defaults[4] gpio_defaults_block_25/gpio_defaults[5]
+ gpio_defaults_block_25/gpio_defaults[6] gpio_defaults_block_25/gpio_defaults[7]
+ gpio_defaults_block_25/gpio_defaults[8] gpio_defaults_block_25/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[32] gpio_control_in_2\[13\]/zero housekeeping/mgmt_gpio_out[32]
+ gpio_control_in_2\[13\]/one padframe/mprj_io_drive_sel[64] padframe/mprj_io_drive_sel[65]
+ padframe/mprj_io_in[32] padframe/mprj_io_inen[32] padframe/mprj_io_out[32] padframe/mprj_io_outen[32]
+ padframe/mprj_io_pd_select[32] padframe/mprj_io_pu_select[32] padframe/mprj_io_schmitt_select[32]
+ padframe/mprj_io_slew_select[32] gpio_control_in_2\[13\]/resetn gpio_control_in_2\[12\]/resetn
+ gpio_control_in_2\[13\]/serial_clock gpio_control_in_2\[12\]/serial_clock gpio_control_in_2\[13\]/serial_data_in
+ gpio_control_in_2\[12\]/serial_data_in gpio_control_in_2\[13\]/serial_load gpio_control_in_2\[12\]/serial_load
+ mprj/io_in[32] mprj/io_oeb[32] mprj/io_out[32] gpio_control_in_2\[13\]/zero gpio_control_block
Xgpio_control_in_1a\[2\] soc/VDD soc/VSS gpio_control_in_1a\[2\]/gpio_defaults[0]
+ gpio_control_in_1a\[2\]/gpio_defaults[1] gpio_control_in_1a\[2\]/gpio_defaults[2]
+ gpio_control_in_1a\[2\]/gpio_defaults[3] gpio_control_in_1a\[2\]/gpio_defaults[4]
+ gpio_control_in_1a\[2\]/gpio_defaults[5] gpio_control_in_1a\[2\]/gpio_defaults[6]
+ gpio_control_in_1a\[2\]/gpio_defaults[7] gpio_control_in_1a\[2\]/gpio_defaults[8]
+ gpio_control_in_1a\[2\]/gpio_defaults[9] housekeeping/mgmt_gpio_in[4] gpio_control_in_1a\[2\]/zero
+ housekeeping/mgmt_gpio_out[4] gpio_control_in_1a\[2\]/one padframe/mprj_io_drive_sel[9]
+ padframe/mprj_io_drive_sel[8] padframe/mprj_io_in[4] padframe/mprj_io_inen[4] padframe/mprj_io_out[4]
+ padframe/mprj_io_outen[4] padframe/mprj_io_pd_select[4] padframe/mprj_io_pu_select[4]
+ padframe/mprj_io_schmitt_select[4] padframe/mprj_io_slew_select[4] gpio_control_in_1a\[2\]/resetn
+ gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[3\]/serial_clock
+ gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[3\]/serial_data_in gpio_control_in_1a\[2\]/serial_load
+ gpio_control_in_1a\[3\]/serial_load mprj/io_in[4] mprj/io_oeb[4] mprj/io_out[4]
+ gpio_control_in_1a\[2\]/zero gpio_control_block
Xgpio_defaults_block_007_1 gpio_control_in_1a\[1\]/gpio_defaults[0] gpio_control_in_1a\[1\]/gpio_defaults[1]
+ gpio_control_in_1a\[1\]/gpio_defaults[2] gpio_control_in_1a\[1\]/gpio_defaults[3]
+ gpio_control_in_1a\[1\]/gpio_defaults[4] gpio_control_in_1a\[1\]/gpio_defaults[5]
+ gpio_control_in_1a\[1\]/gpio_defaults[6] gpio_control_in_1a\[1\]/gpio_defaults[7]
+ gpio_control_in_1a\[1\]/gpio_defaults[8] gpio_control_in_1a\[1\]/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_007
Xgpio_control_in_2\[8\] soc/VDD soc/VSS gpio_defaults_block_19/gpio_defaults[0] gpio_defaults_block_19/gpio_defaults[1]
+ gpio_defaults_block_19/gpio_defaults[2] gpio_defaults_block_19/gpio_defaults[3]
+ gpio_defaults_block_19/gpio_defaults[4] gpio_defaults_block_19/gpio_defaults[5]
+ gpio_defaults_block_19/gpio_defaults[6] gpio_defaults_block_19/gpio_defaults[7]
+ gpio_defaults_block_19/gpio_defaults[8] gpio_defaults_block_19/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[27] gpio_control_in_2\[8\]/zero housekeeping/mgmt_gpio_out[27]
+ gpio_control_in_2\[8\]/one padframe/mprj_io_drive_sel[54] padframe/mprj_io_drive_sel[55]
+ padframe/mprj_io_in[27] padframe/mprj_io_inen[27] padframe/mprj_io_out[27] padframe/mprj_io_outen[27]
+ padframe/mprj_io_pd_select[27] padframe/mprj_io_pu_select[27] padframe/mprj_io_schmitt_select[27]
+ padframe/mprj_io_slew_select[27] gpio_control_in_2\[8\]/resetn gpio_control_in_2\[7\]/resetn
+ gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[8\]/serial_data_in
+ gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[8\]/serial_load gpio_control_in_2\[7\]/serial_load
+ mprj/io_in[27] mprj/io_oeb[27] mprj/io_out[27] gpio_control_in_2\[8\]/zero gpio_control_block
Xgpio_defaults_block_007_2 gpio_control_in_1a\[0\]/gpio_defaults[0] gpio_control_in_1a\[0\]/gpio_defaults[1]
+ gpio_control_in_1a\[0\]/gpio_defaults[2] gpio_control_in_1a\[0\]/gpio_defaults[3]
+ gpio_control_in_1a\[0\]/gpio_defaults[4] gpio_control_in_1a\[0\]/gpio_defaults[5]
+ gpio_control_in_1a\[0\]/gpio_defaults[6] gpio_control_in_1a\[0\]/gpio_defaults[7]
+ gpio_control_in_1a\[0\]/gpio_defaults[8] gpio_control_in_1a\[0\]/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_007
Xgpio_control_in_1\[3\] soc/VDD soc/VSS gpio_defaults_block_15/gpio_defaults[0] gpio_defaults_block_15/gpio_defaults[1]
+ gpio_defaults_block_15/gpio_defaults[2] gpio_defaults_block_15/gpio_defaults[3]
+ gpio_defaults_block_15/gpio_defaults[4] gpio_defaults_block_15/gpio_defaults[5]
+ gpio_defaults_block_15/gpio_defaults[6] gpio_defaults_block_15/gpio_defaults[7]
+ gpio_defaults_block_15/gpio_defaults[8] gpio_defaults_block_15/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[11] gpio_control_in_1\[3\]/zero housekeeping/mgmt_gpio_out[11]
+ gpio_control_in_1\[3\]/one padframe/mprj_io_drive_sel[23] padframe/mprj_io_drive_sel[22]
+ padframe/mprj_io_in[11] padframe/mprj_io_inen[11] padframe/mprj_io_out[11] padframe/mprj_io_outen[11]
+ padframe/mprj_io_pd_select[11] padframe/mprj_io_pu_select[11] padframe/mprj_io_schmitt_select[11]
+ padframe/mprj_io_slew_select[11] gpio_control_in_1\[3\]/resetn gpio_control_in_1\[4\]/resetn
+ gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[3\]/serial_data_in
+ gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[3\]/serial_load gpio_control_in_1\[4\]/serial_load
+ mprj/io_in[11] mprj/io_oeb[11] mprj/io_out[11] gpio_control_in_1\[3\]/zero gpio_control_block
Xgpio_control_in_2\[11\] soc/VDD soc/VSS gpio_defaults_block_23/gpio_defaults[0] gpio_defaults_block_23/gpio_defaults[1]
+ gpio_defaults_block_23/gpio_defaults[2] gpio_defaults_block_23/gpio_defaults[3]
+ gpio_defaults_block_23/gpio_defaults[4] gpio_defaults_block_23/gpio_defaults[5]
+ gpio_defaults_block_23/gpio_defaults[6] gpio_defaults_block_23/gpio_defaults[7]
+ gpio_defaults_block_23/gpio_defaults[8] gpio_defaults_block_23/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[30] gpio_control_in_2\[11\]/zero housekeeping/mgmt_gpio_out[30]
+ gpio_control_in_2\[11\]/one padframe/mprj_io_drive_sel[63] padframe/mprj_io_drive_sel[61]
+ padframe/mprj_io_in[30] padframe/mprj_io_inen[30] padframe/mprj_io_out[30] padframe/mprj_io_outen[30]
+ padframe/mprj_io_pd_select[30] padframe/mprj_io_pu_select[30] padframe/mprj_io_schmitt_select[30]
+ padframe/mprj_io_slew_select[30] gpio_control_in_2\[11\]/resetn gpio_control_in_2\[10\]/resetn
+ gpio_control_in_2\[11\]/serial_clock gpio_control_in_2\[10\]/serial_clock gpio_control_in_2\[11\]/serial_data_in
+ gpio_control_in_2\[10\]/serial_data_in gpio_control_in_2\[11\]/serial_load gpio_control_in_2\[10\]/serial_load
+ mprj/io_in[30] mprj/io_oeb[30] mprj/io_out[30] gpio_control_in_2\[11\]/zero gpio_control_block
Xgpio_control_in_1a\[0\] soc/VDD soc/VSS gpio_control_in_1a\[0\]/gpio_defaults[0]
+ gpio_control_in_1a\[0\]/gpio_defaults[1] gpio_control_in_1a\[0\]/gpio_defaults[2]
+ gpio_control_in_1a\[0\]/gpio_defaults[3] gpio_control_in_1a\[0\]/gpio_defaults[4]
+ gpio_control_in_1a\[0\]/gpio_defaults[5] gpio_control_in_1a\[0\]/gpio_defaults[6]
+ gpio_control_in_1a\[0\]/gpio_defaults[7] gpio_control_in_1a\[0\]/gpio_defaults[8]
+ gpio_control_in_1a\[0\]/gpio_defaults[9] housekeeping/mgmt_gpio_in[2] gpio_control_in_1a\[0\]/zero
+ housekeeping/mgmt_gpio_out[2] gpio_control_in_1a\[0\]/one padframe/mprj_io_drive_sel[5]
+ padframe/mprj_io_drive_sel[4] padframe/mprj_io_in[2] padframe/mprj_io_inen[2] padframe/mprj_io_out[2]
+ padframe/mprj_io_outen[2] padframe/mprj_io_pd_select[2] padframe/mprj_io_pu_select[2]
+ padframe/mprj_io_schmitt_select[2] padframe/mprj_io_slew_select[2] gpio_control_in_1a\[0\]/resetn
+ gpio_control_in_1a\[1\]/resetn gpio_control_in_1a\[0\]/serial_clock gpio_control_in_1a\[1\]/serial_clock
+ gpio_control_in_1a\[0\]/serial_data_in gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_load
+ gpio_control_in_1a\[1\]/serial_load mprj/io_in[2] mprj/io_oeb[2] mprj/io_out[2]
+ gpio_control_in_1a\[0\]/zero gpio_control_block
Xgpio_control_in_2\[6\] soc/VDD soc/VSS gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[1]
+ gpio_defaults_block_14/gpio_defaults[2] gpio_defaults_block_14/gpio_defaults[3]
+ gpio_defaults_block_14/gpio_defaults[4] gpio_defaults_block_14/gpio_defaults[5]
+ gpio_defaults_block_14/gpio_defaults[6] gpio_defaults_block_14/gpio_defaults[7]
+ gpio_defaults_block_14/gpio_defaults[8] gpio_defaults_block_14/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[25] gpio_control_in_2\[6\]/zero housekeeping/mgmt_gpio_out[25]
+ gpio_control_in_2\[6\]/one padframe/mprj_io_drive_sel[525] padframe/mprj_io_drive_sel[51]
+ padframe/mprj_io_in[25] padframe/mprj_io_inen[25] padframe/mprj_io_out[25] padframe/mprj_io_outen[25]
+ padframe/mprj_io_pd_select[25] padframe/mprj_io_pu_select[25] padframe/mprj_io_schmitt_select[25]
+ padframe/mprj_io_slew_select[25] gpio_control_in_2\[6\]/resetn gpio_control_in_2\[5\]/resetn
+ gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[6\]/serial_data_in
+ gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[6\]/serial_load gpio_control_in_2\[5\]/serial_load
+ mprj/io_in[25] mprj/io_oeb[25] mprj/io_out[25] gpio_control_in_2\[6\]/zero gpio_control_block
Xgpio_control_in_1\[1\] soc/VDD soc/VSS gpio_defaults_block_20/gpio_defaults[0] gpio_defaults_block_20/gpio_defaults[1]
+ gpio_defaults_block_20/gpio_defaults[2] gpio_defaults_block_20/gpio_defaults[3]
+ gpio_defaults_block_20/gpio_defaults[4] gpio_defaults_block_20/gpio_defaults[5]
+ gpio_defaults_block_20/gpio_defaults[6] gpio_defaults_block_20/gpio_defaults[7]
+ gpio_defaults_block_20/gpio_defaults[8] gpio_defaults_block_20/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[9] gpio_control_in_1\[1\]/zero housekeeping/mgmt_gpio_out[9]
+ gpio_control_in_1\[1\]/one padframe/mprj_io_drive_sel[19] padframe/mprj_io_drive_sel[18]
+ padframe/mprj_io_in[9] padframe/mprj_io_inen[9] padframe/mprj_io_out[9] padframe/mprj_io_outen[9]
+ padframe/mprj_io_pd_select[9] padframe/mprj_io_pu_select[9] padframe/mprj_io_schmitt_select[9]
+ padframe/mprj_io_slew_select[9] gpio_control_in_1\[1\]/resetn gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[1\]/serial_data_in
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[1\]/serial_load gpio_control_in_1\[2\]/serial_load
+ mprj/io_in[9] mprj/io_oeb[9] mprj/io_out[9] gpio_control_in_1\[1\]/zero gpio_control_block
Xmprj mprj/io_in[0] mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13] mprj/io_in[14]
+ mprj/io_in[15] mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19] mprj/io_in[1]
+ mprj/io_in[20] mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24] mprj/io_in[25]
+ mprj/io_in[26] mprj/io_in[27] mprj/io_in[28] mprj/io_in[29] mprj/io_in[2] mprj/io_in[30]
+ mprj/io_in[31] mprj/io_in[32] mprj/io_in[33] mprj/io_in[34] mprj/io_in[35] mprj/io_in[36]
+ mprj/io_in[37] mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6] mprj/io_in[7]
+ mprj/io_in[8] mprj/io_in[9] mprj/io_oeb[0] mprj/io_oeb[10] mprj/io_oeb[11] mprj/io_oeb[12]
+ mprj/io_oeb[13] mprj/io_oeb[14] mprj/io_oeb[15] mprj/io_oeb[16] mprj/io_oeb[17]
+ mprj/io_oeb[18] mprj/io_oeb[19] mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21] mprj/io_oeb[22]
+ mprj/io_oeb[23] mprj/io_oeb[24] mprj/io_oeb[25] mprj/io_oeb[26] mprj/io_oeb[27]
+ mprj/io_oeb[28] mprj/io_oeb[29] mprj/io_oeb[2] mprj/io_oeb[30] mprj/io_oeb[31] mprj/io_oeb[32]
+ mprj/io_oeb[33] mprj/io_oeb[34] mprj/io_oeb[35] mprj/io_oeb[36] mprj/io_oeb[37]
+ mprj/io_oeb[3] mprj/io_oeb[4] mprj/io_oeb[5] mprj/io_oeb[6] mprj/io_oeb[7] mprj/io_oeb[8]
+ mprj/io_oeb[9] mprj/io_out[0] mprj/io_out[10] mprj/io_out[11] mprj/io_out[12] mprj/io_out[13]
+ mprj/io_out[14] mprj/io_out[15] mprj/io_out[16] mprj/io_out[17] mprj/io_out[18]
+ mprj/io_out[19] mprj/io_out[1] mprj/io_out[20] mprj/io_out[21] mprj/io_out[22] mprj/io_out[23]
+ mprj/io_out[24] mprj/io_out[25] mprj/io_out[26] mprj/io_out[27] mprj/io_out[28]
+ mprj/io_out[29] mprj/io_out[2] mprj/io_out[30] mprj/io_out[31] mprj/io_out[32] mprj/io_out[33]
+ mprj/io_out[34] mprj/io_out[35] mprj/io_out[36] mprj/io_out[37] mprj/io_out[3] mprj/io_out[4]
+ mprj/io_out[5] mprj/io_out[6] mprj/io_out[7] mprj/io_out[8] mprj/io_out[9] mprj/la_data_in[0]
+ mprj/la_data_in[10] mprj/la_data_in[11] mprj/la_data_in[12] mprj/la_data_in[13]
+ mprj/la_data_in[14] mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17]
+ mprj/la_data_in[18] mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21]
+ mprj/la_data_in[22] mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25]
+ mprj/la_data_in[26] mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29]
+ mprj/la_data_in[2] mprj/la_data_in[30] mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33]
+ mprj/la_data_in[34] mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37]
+ mprj/la_data_in[38] mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41]
+ mprj/la_data_in[42] mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45]
+ mprj/la_data_in[46] mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49]
+ mprj/la_data_in[4] mprj/la_data_in[50] mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53]
+ mprj/la_data_in[54] mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57]
+ mprj/la_data_in[58] mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61]
+ mprj/la_data_in[62] mprj/la_data_in[63] mprj/la_data_in[6] mprj/la_data_in[7] mprj/la_data_in[8]
+ mprj/la_data_in[9] mprj/la_data_out[0] mprj/la_data_out[10] mprj/la_data_out[11]
+ mprj/la_data_out[12] mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15]
+ mprj/la_data_out[16] mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19]
+ mprj/la_data_out[1] mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22]
+ mprj/la_data_out[23] mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26]
+ mprj/la_data_out[27] mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2]
+ mprj/la_data_out[30] mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33]
+ mprj/la_data_out[34] mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37]
+ mprj/la_data_out[38] mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40]
+ mprj/la_data_out[41] mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44]
+ mprj/la_data_out[45] mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48]
+ mprj/la_data_out[49] mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51]
+ mprj/la_data_out[52] mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55]
+ mprj/la_data_out[56] mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59]
+ mprj/la_data_out[5] mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62]
+ mprj/la_data_out[63] mprj/la_data_out[6] mprj/la_data_out[7] mprj/la_data_out[8]
+ mprj/la_data_out[9] mprj/la_oenb[0] mprj/la_oenb[10] mprj/la_oenb[11] mprj/la_oenb[12]
+ mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17]
+ mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21]
+ mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26]
+ mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30]
+ mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35]
+ mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3]
+ mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44]
+ mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49]
+ mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53]
+ mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58]
+ mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62]
+ mprj/la_oenb[63] mprj/la_oenb[6] mprj/la_oenb[7] mprj/la_oenb[8] mprj/la_oenb[9]
+ mprj/user_clock2 mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] soc/VDD soc/VSS
+ mprj/wb_clk_i mprj/wb_rst_i mprj/wbs_ack_o mprj/wbs_adr_i[0] mprj/wbs_adr_i[10]
+ mprj/wbs_adr_i[11] mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15]
+ mprj/wbs_adr_i[16] mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1]
+ mprj/wbs_adr_i[20] mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24]
+ mprj/wbs_adr_i[25] mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29]
+ mprj/wbs_adr_i[2] mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4]
+ mprj/wbs_adr_i[5] mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9]
+ mprj/wbs_cyc_i mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12]
+ mprj/wbs_dat_i[13] mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17]
+ mprj/wbs_dat_i[18] mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21]
+ mprj/wbs_dat_i[22] mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26]
+ mprj/wbs_dat_i[27] mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30]
+ mprj/wbs_dat_i[31] mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6]
+ mprj/wbs_dat_i[7] mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10]
+ mprj/wbs_dat_o[11] mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15]
+ mprj/wbs_dat_o[16] mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1]
+ mprj/wbs_dat_o[20] mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24]
+ mprj/wbs_dat_o[25] mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29]
+ mprj/wbs_dat_o[2] mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4]
+ mprj/wbs_dat_o[5] mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9]
+ mprj/wbs_sel_i[0] mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i
+ mprj/wbs_we_i user_project_wrapper
Xgpio_control_in_2\[4\] soc/VDD soc/VSS gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[1]
+ gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3] gpio_defaults_block_8/gpio_defaults[4]
+ gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6] gpio_defaults_block_8/gpio_defaults[7]
+ gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9] housekeeping/mgmt_gpio_in[23]
+ gpio_control_in_2\[4\]/zero housekeeping/mgmt_gpio_out[23] gpio_control_in_2\[4\]/one
+ padframe/mprj_io_drive_sel[46] padframe/mprj_io_drive_sel[47] padframe/mprj_io_in[23]
+ padframe/mprj_io_inen[23] padframe/mprj_io_out[23] padframe/mprj_io_outen[23] padframe/mprj_io_pd_select[23]
+ padframe/mprj_io_pu_select[23] padframe/mprj_io_schmitt_select[23] padframe/mprj_io_slew_select[23]
+ gpio_control_in_2\[4\]/resetn gpio_control_in_2\[3\]/resetn gpio_control_in_2\[4\]/serial_clock
+ gpio_control_in_2\[3\]/serial_clock gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[3\]/serial_data_in
+ gpio_control_in_2\[4\]/serial_load gpio_control_in_2\[3\]/serial_load mprj/io_in[23]
+ mprj/io_oeb[23] mprj/io_out[23] gpio_control_in_2\[4\]/zero gpio_control_block
Xgpio_control_bidir_1\[1\] soc/VDD soc/VSS gpio_defaults_block_009_0/gpio_defaults[0]
+ gpio_defaults_block_009_0/gpio_defaults[1] gpio_defaults_block_009_0/gpio_defaults[2]
+ gpio_defaults_block_009_0/gpio_defaults[3] gpio_defaults_block_009_0/gpio_defaults[4]
+ gpio_defaults_block_009_0/gpio_defaults[5] gpio_defaults_block_009_0/gpio_defaults[6]
+ gpio_defaults_block_009_0/gpio_defaults[7] gpio_defaults_block_009_0/gpio_defaults[8]
+ gpio_defaults_block_009_0/gpio_defaults[9] housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_oeb[1]
+ housekeeping/mgmt_gpio_out[1] gpio_control_bidir_1\[1\]/one padframe/mprj_io_drive_sel[2]
+ padframe/mprj_io_drive_sel[3] padframe/mprj_io_in[1] padframe/mprj_io_inen[1] padframe/mprj_io_out[1]
+ padframe/mprj_io_outen[1] padframe/mprj_io_pd_select[1] padframe/mprj_io_pu_select[1]
+ padframe/mprj_io_schmitt_select[1] padframe/mprj_io_slew_select[1] gpio_control_bidir_1\[1\]/resetn
+ gpio_control_in_1a\[0\]/resetn gpio_control_bidir_1\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_clock
+ gpio_control_bidir_1\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_data_in
+ gpio_control_bidir_1\[1\]/serial_load gpio_control_in_1a\[0\]/serial_load mprj/io_in[1]
+ mprj/io_oeb[1] mprj/io_out[1] gpio_control_bidir_1\[1\]/zero gpio_control_block
Xspare_logic\[2\] soc/VDD soc/VSS spare_logic\[2\]/spare_xfq[0] spare_logic\[2\]/spare_xfq[1]
+ spare_logic\[2\]/spare_xi[0] spare_logic\[2\]/spare_xi[1] spare_logic\[2\]/spare_xi[2]
+ spare_logic\[2\]/spare_xi[3] spare_logic\[2\]/spare_xib spare_logic\[2\]/spare_xmx[0]
+ spare_logic\[2\]/spare_xmx[1] spare_logic\[2\]/spare_xna[0] spare_logic\[2\]/spare_xna[1]
+ spare_logic\[2\]/spare_xno[0] spare_logic\[2\]/spare_xno[1] spare_logic\[2\]/spare_xz[0]
+ spare_logic\[2\]/spare_xz[10] spare_logic\[2\]/spare_xz[11] spare_logic\[2\]/spare_xz[12]
+ spare_logic\[2\]/spare_xz[13] spare_logic\[2\]/spare_xz[14] spare_logic\[2\]/spare_xz[15]
+ spare_logic\[2\]/spare_xz[16] spare_logic\[2\]/spare_xz[17] spare_logic\[2\]/spare_xz[18]
+ spare_logic\[2\]/spare_xz[19] spare_logic\[2\]/spare_xz[1] spare_logic\[2\]/spare_xz[20]
+ spare_logic\[2\]/spare_xz[21] spare_logic\[2\]/spare_xz[22] spare_logic\[2\]/spare_xz[23]
+ spare_logic\[2\]/spare_xz[24] spare_logic\[2\]/spare_xz[25] spare_logic\[2\]/spare_xz[26]
+ spare_logic\[2\]/spare_xz[27] spare_logic\[2\]/spare_xz[28] spare_logic\[2\]/spare_xz[29]
+ spare_logic\[2\]/spare_xz[2] spare_logic\[2\]/spare_xz[30] spare_logic\[2\]/spare_xz[3]
+ spare_logic\[2\]/spare_xz[4] spare_logic\[2\]/spare_xz[5] spare_logic\[2\]/spare_xz[6]
+ spare_logic\[2\]/spare_xz[7] spare_logic\[2\]/spare_xz[8] spare_logic\[2\]/spare_xz[9]
+ spare_logic_block
Xhousekeeping soc/VDD soc/VSS soc/debug_in soc/debug_mode soc/debug_oeb soc/debug_out
+ soc/irq[3] soc/irq[4] soc/irq[5] user_id_value/mask_rev[0] user_id_value/mask_rev[10]
+ user_id_value/mask_rev[11] user_id_value/mask_rev[12] user_id_value/mask_rev[13]
+ user_id_value/mask_rev[14] user_id_value/mask_rev[15] user_id_value/mask_rev[16]
+ user_id_value/mask_rev[17] user_id_value/mask_rev[18] user_id_value/mask_rev[19]
+ user_id_value/mask_rev[1] user_id_value/mask_rev[20] user_id_value/mask_rev[21]
+ user_id_value/mask_rev[22] user_id_value/mask_rev[23] user_id_value/mask_rev[24]
+ user_id_value/mask_rev[25] user_id_value/mask_rev[26] user_id_value/mask_rev[27]
+ user_id_value/mask_rev[28] user_id_value/mask_rev[29] user_id_value/mask_rev[2]
+ user_id_value/mask_rev[30] user_id_value/mask_rev[31] user_id_value/mask_rev[3]
+ user_id_value/mask_rev[4] user_id_value/mask_rev[5] user_id_value/mask_rev[6] user_id_value/mask_rev[7]
+ user_id_value/mask_rev[8] user_id_value/mask_rev[9] housekeeping/mgmt_gpio_in[0]
+ housekeeping/mgmt_gpio_in[10] housekeeping/mgmt_gpio_in[11] housekeeping/mgmt_gpio_in[12]
+ housekeeping/mgmt_gpio_in[13] housekeeping/mgmt_gpio_in[14] housekeeping/mgmt_gpio_in[15]
+ housekeeping/mgmt_gpio_in[16] housekeeping/mgmt_gpio_in[17] housekeeping/mgmt_gpio_in[18]
+ housekeeping/mgmt_gpio_in[19] housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_in[20]
+ housekeeping/mgmt_gpio_in[21] housekeeping/mgmt_gpio_in[22] housekeeping/mgmt_gpio_in[23]
+ housekeeping/mgmt_gpio_in[24] housekeeping/mgmt_gpio_in[25] housekeeping/mgmt_gpio_in[26]
+ housekeeping/mgmt_gpio_in[27] housekeeping/mgmt_gpio_in[28] housekeeping/mgmt_gpio_in[29]
+ housekeeping/mgmt_gpio_in[2] housekeeping/mgmt_gpio_in[30] housekeeping/mgmt_gpio_in[31]
+ housekeeping/mgmt_gpio_in[32] housekeeping/mgmt_gpio_in[33] housekeeping/mgmt_gpio_in[34]
+ housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_in[36] housekeeping/mgmt_gpio_in[37]
+ housekeeping/mgmt_gpio_in[3] housekeeping/mgmt_gpio_in[4] housekeeping/mgmt_gpio_in[5]
+ housekeeping/mgmt_gpio_in[6] housekeeping/mgmt_gpio_in[7] housekeeping/mgmt_gpio_in[8]
+ housekeeping/mgmt_gpio_in[9] housekeeping/mgmt_gpio_oeb[0] housekeeping/mgmt_gpio_oeb[10]
+ housekeeping/mgmt_gpio_oeb[11] housekeeping/mgmt_gpio_oeb[12] housekeeping/mgmt_gpio_oeb[13]
+ housekeeping/mgmt_gpio_oeb[14] housekeeping/mgmt_gpio_oeb[15] housekeeping/mgmt_gpio_oeb[16]
+ housekeeping/mgmt_gpio_oeb[17] housekeeping/mgmt_gpio_oeb[18] housekeeping/mgmt_gpio_oeb[19]
+ housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_oeb[20] housekeeping/mgmt_gpio_oeb[21]
+ housekeeping/mgmt_gpio_oeb[22] housekeeping/mgmt_gpio_oeb[23] housekeeping/mgmt_gpio_oeb[24]
+ housekeeping/mgmt_gpio_oeb[25] housekeeping/mgmt_gpio_oeb[26] housekeeping/mgmt_gpio_oeb[27]
+ housekeeping/mgmt_gpio_oeb[28] housekeeping/mgmt_gpio_oeb[29] housekeeping/mgmt_gpio_oeb[2]
+ housekeeping/mgmt_gpio_oeb[30] housekeeping/mgmt_gpio_oeb[31] housekeeping/mgmt_gpio_oeb[32]
+ housekeeping/mgmt_gpio_oeb[33] housekeeping/mgmt_gpio_oeb[34] housekeeping/mgmt_gpio_oeb[35]
+ housekeeping/mgmt_gpio_oeb[36] housekeeping/mgmt_gpio_oeb[37] housekeeping/mgmt_gpio_oeb[3]
+ housekeeping/mgmt_gpio_oeb[4] housekeeping/mgmt_gpio_oeb[5] housekeeping/mgmt_gpio_oeb[6]
+ housekeeping/mgmt_gpio_oeb[7] housekeeping/mgmt_gpio_oeb[8] housekeeping/mgmt_gpio_oeb[9]
+ housekeeping/mgmt_gpio_out[0] housekeeping/mgmt_gpio_out[10] housekeeping/mgmt_gpio_out[11]
+ housekeeping/mgmt_gpio_out[12] housekeeping/mgmt_gpio_out[13] housekeeping/mgmt_gpio_out[14]
+ housekeeping/mgmt_gpio_out[15] housekeeping/mgmt_gpio_out[16] housekeeping/mgmt_gpio_out[17]
+ housekeeping/mgmt_gpio_out[18] housekeeping/mgmt_gpio_out[19] housekeeping/mgmt_gpio_out[1]
+ housekeeping/mgmt_gpio_out[20] housekeeping/mgmt_gpio_out[21] housekeeping/mgmt_gpio_out[22]
+ housekeeping/mgmt_gpio_out[23] housekeeping/mgmt_gpio_out[24] housekeeping/mgmt_gpio_out[25]
+ housekeeping/mgmt_gpio_out[26] housekeeping/mgmt_gpio_out[27] housekeeping/mgmt_gpio_out[28]
+ housekeeping/mgmt_gpio_out[29] housekeeping/mgmt_gpio_out[2] housekeeping/mgmt_gpio_out[30]
+ housekeeping/mgmt_gpio_out[31] housekeeping/mgmt_gpio_out[32] housekeeping/mgmt_gpio_out[33]
+ housekeeping/mgmt_gpio_out[34] housekeeping/mgmt_gpio_out[35] housekeeping/mgmt_gpio_out[36]
+ housekeeping/mgmt_gpio_out[37] housekeeping/mgmt_gpio_out[3] housekeeping/mgmt_gpio_out[4]
+ housekeeping/mgmt_gpio_out[5] housekeeping/mgmt_gpio_out[6] housekeeping/mgmt_gpio_out[7]
+ housekeeping/mgmt_gpio_out[8] housekeeping/mgmt_gpio_out[9] padframe/flash_clk_core
+ padframe/flash_clk_oe_core padframe/flash_csb_core padframe/flash_csb_oe_core padframe/flash_io0_di_core
+ padframe/flash_io0_do_core padframe/flash_io0_ie_core padframe/flash_io0_oe_core
+ padframe/flash_io1_di_core padframe/flash_io1_do_core padframe/flash_io1_ie_core
+ padframe/flash_io1_oe_core clock_ctrl/sel2[0] clock_ctrl/sel2[1] clock_ctrl/sel2[2]
+ clock_ctrl/ext_clk_sel pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3] pll/div[4]
+ pll/enable clock_ctrl/sel[0] clock_ctrl/sel[1] clock_ctrl/sel[2] pll/ext_trim[0]
+ pll/ext_trim[10] pll/ext_trim[11] pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14]
+ pll/ext_trim[15] pll/ext_trim[16] pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19]
+ pll/ext_trim[1] pll/ext_trim[20] pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23]
+ pll/ext_trim[24] pll/ext_trim[25] pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4]
+ pll/ext_trim[5] pll/ext_trim[6] pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9]
+ simple_por_0/porb housekeeping/pwr_ctrl_out soc/qspi_enabled housekeeping/reset
+ soc/ser_rx soc/ser_tx housekeeping/serial_clock housekeeping/serial_data_1 housekeeping/serial_data_2
+ housekeeping/serial_load housekeeping/serial_resetn soc/spi_csb soc/spi_enabled
+ soc/spi_sck soc/spi_sdi soc/spi_sdo soc/spi_sdoenb soc/flash_clk soc/flash_csb soc/flash_io0_di
+ soc/flash_io0_do soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb
+ soc/flash_io2_di soc/flash_io2_do soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do
+ soc/flash_io3_oeb soc/trap soc/uart_enabled clock_ctrl/user_clk soc/hk_ack_i soc/mprj_adr_o[0]
+ soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14]
+ soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19]
+ soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23]
+ soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28]
+ soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3]
+ soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8]
+ soc/mprj_adr_o[9] soc/core_clk soc/hk_cyc_o soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11] soc/hk_dat_i[12] soc/hk_dat_i[13]
+ soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16] soc/hk_dat_i[17] soc/hk_dat_i[18]
+ soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20] soc/hk_dat_i[21] soc/hk_dat_i[22]
+ soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25] soc/hk_dat_i[26] soc/hk_dat_i[27]
+ soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2] soc/hk_dat_i[30] soc/hk_dat_i[31]
+ soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5] soc/hk_dat_i[6] soc/hk_dat_i[7]
+ soc/hk_dat_i[8] soc/hk_dat_i[9] soc/core_rstn soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/hk_stb_o soc/mprj_we_o housekeeping
Xgpio_control_in_2\[2\] soc/VDD soc/VSS gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[1]
+ gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3] gpio_defaults_block_7/gpio_defaults[4]
+ gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6] gpio_defaults_block_7/gpio_defaults[7]
+ gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9] housekeeping/mgmt_gpio_in[21]
+ gpio_control_in_2\[2\]/zero housekeeping/mgmt_gpio_out[21] gpio_control_in_2\[2\]/one
+ padframe/mprj_io_drive_sel[42] padframe/mprj_io_drive_sel[43] padframe/mprj_io_in[21]
+ padframe/mprj_io_inen[21] padframe/mprj_io_out[21] padframe/mprj_io_outen[21] padframe/mprj_io_pd_select[21]
+ padframe/mprj_io_pu_select[21] padframe/mprj_io_schmitt_select[21] padframe/mprj_io_slew_select[21]
+ gpio_control_in_2\[2\]/resetn gpio_control_in_2\[1\]/resetn gpio_control_in_2\[2\]/serial_clock
+ gpio_control_in_2\[1\]/serial_clock gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[1\]/serial_data_in
+ gpio_control_in_2\[2\]/serial_load gpio_control_in_2\[1\]/serial_load mprj/io_in[21]
+ mprj/io_oeb[21] mprj/io_out[21] gpio_control_in_2\[2\]/zero gpio_control_block
Xgpio_control_in_1\[8\] soc/VDD soc/VSS gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[1]
+ gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3] gpio_defaults_block_2/gpio_defaults[4]
+ gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6] gpio_defaults_block_2/gpio_defaults[7]
+ gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9] housekeeping/mgmt_gpio_in[16]
+ gpio_control_in_1\[8\]/zero housekeeping/mgmt_gpio_out[16] gpio_control_in_1\[8\]/one
+ padframe/mprj_io_drive_sel[32] padframe/mprj_io_drive_sel[33] padframe/mprj_io_in[16]
+ padframe/mprj_io_inen[16] padframe/mprj_io_out[16] padframe/mprj_io_outen[16] padframe/mprj_io_pd_select[16]
+ padframe/mprj_io_pu_select[16] padframe/mprj_io_schmitt_select[16] padframe/mprj_io_slew_select[16]
+ gpio_control_in_1\[8\]/resetn gpio_control_in_1\[9\]/resetn gpio_control_in_1\[8\]/serial_clock
+ gpio_control_in_1\[9\]/serial_clock gpio_control_in_1\[8\]/serial_data_in gpio_control_in_1\[9\]/serial_data_in
+ gpio_control_in_1\[8\]/serial_load gpio_control_in_1\[9\]/serial_load mprj/io_in[16]
+ mprj/io_oeb[16] mprj/io_out[16] gpio_control_in_1\[8\]/zero gpio_control_block
Xspare_logic\[0\] soc/VDD soc/VSS spare_logic\[0\]/spare_xfq[0] spare_logic\[0\]/spare_xfq[1]
+ spare_logic\[0\]/spare_xi[0] spare_logic\[0\]/spare_xi[1] spare_logic\[0\]/spare_xi[2]
+ spare_logic\[0\]/spare_xi[3] spare_logic\[0\]/spare_xib spare_logic\[0\]/spare_xmx[0]
+ spare_logic\[0\]/spare_xmx[1] spare_logic\[0\]/spare_xna[0] spare_logic\[0\]/spare_xna[1]
+ spare_logic\[0\]/spare_xno[0] spare_logic\[0\]/spare_xno[1] spare_logic\[0\]/spare_xz[0]
+ spare_logic\[0\]/spare_xz[10] spare_logic\[0\]/spare_xz[11] spare_logic\[0\]/spare_xz[12]
+ spare_logic\[0\]/spare_xz[13] spare_logic\[0\]/spare_xz[14] spare_logic\[0\]/spare_xz[15]
+ spare_logic\[0\]/spare_xz[16] spare_logic\[0\]/spare_xz[17] spare_logic\[0\]/spare_xz[18]
+ spare_logic\[0\]/spare_xz[19] spare_logic\[0\]/spare_xz[1] spare_logic\[0\]/spare_xz[20]
+ spare_logic\[0\]/spare_xz[21] spare_logic\[0\]/spare_xz[22] spare_logic\[0\]/spare_xz[23]
+ spare_logic\[0\]/spare_xz[24] spare_logic\[0\]/spare_xz[25] spare_logic\[0\]/spare_xz[26]
+ spare_logic\[0\]/spare_xz[27] spare_logic\[0\]/spare_xz[28] spare_logic\[0\]/spare_xz[29]
+ spare_logic\[0\]/spare_xz[2] spare_logic\[0\]/spare_xz[30] spare_logic\[0\]/spare_xz[3]
+ spare_logic\[0\]/spare_xz[4] spare_logic\[0\]/spare_xz[5] spare_logic\[0\]/spare_xz[6]
+ spare_logic\[0\]/spare_xz[7] spare_logic\[0\]/spare_xz[8] spare_logic\[0\]/spare_xz[9]
+ spare_logic_block
Xgpio_defaults_block_30 gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[1]
+ gpio_defaults_block_30/gpio_defaults[2] gpio_defaults_block_30/gpio_defaults[3]
+ gpio_defaults_block_30/gpio_defaults[4] gpio_defaults_block_30/gpio_defaults[5]
+ gpio_defaults_block_30/gpio_defaults[6] gpio_defaults_block_30/gpio_defaults[7]
+ gpio_defaults_block_30/gpio_defaults[8] gpio_defaults_block_30/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_10 gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[1]
+ gpio_defaults_block_10/gpio_defaults[2] gpio_defaults_block_10/gpio_defaults[3]
+ gpio_defaults_block_10/gpio_defaults[4] gpio_defaults_block_10/gpio_defaults[5]
+ gpio_defaults_block_10/gpio_defaults[6] gpio_defaults_block_10/gpio_defaults[7]
+ gpio_defaults_block_10/gpio_defaults[8] gpio_defaults_block_10/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_20 gpio_defaults_block_20/gpio_defaults[0] gpio_defaults_block_20/gpio_defaults[1]
+ gpio_defaults_block_20/gpio_defaults[2] gpio_defaults_block_20/gpio_defaults[3]
+ gpio_defaults_block_20/gpio_defaults[4] gpio_defaults_block_20/gpio_defaults[5]
+ gpio_defaults_block_20/gpio_defaults[6] gpio_defaults_block_20/gpio_defaults[7]
+ gpio_defaults_block_20/gpio_defaults[8] gpio_defaults_block_20/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_21 gpio_defaults_block_21/gpio_defaults[0] gpio_defaults_block_21/gpio_defaults[1]
+ gpio_defaults_block_21/gpio_defaults[2] gpio_defaults_block_21/gpio_defaults[3]
+ gpio_defaults_block_21/gpio_defaults[4] gpio_defaults_block_21/gpio_defaults[5]
+ gpio_defaults_block_21/gpio_defaults[6] gpio_defaults_block_21/gpio_defaults[7]
+ gpio_defaults_block_21/gpio_defaults[8] gpio_defaults_block_21/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1a\[5\] soc/VDD soc/VSS gpio_defaults_block_24/gpio_defaults[0] gpio_defaults_block_24/gpio_defaults[1]
+ gpio_defaults_block_24/gpio_defaults[2] gpio_defaults_block_24/gpio_defaults[3]
+ gpio_defaults_block_24/gpio_defaults[4] gpio_defaults_block_24/gpio_defaults[5]
+ gpio_defaults_block_24/gpio_defaults[6] gpio_defaults_block_24/gpio_defaults[7]
+ gpio_defaults_block_24/gpio_defaults[8] gpio_defaults_block_24/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[7] gpio_control_in_1a\[5\]/zero housekeeping/mgmt_gpio_out[7]
+ gpio_control_in_1a\[5\]/one padframe/mprj_io_drive_sel[15] padframe/mprj_io_drive_sel[14]
+ padframe/mprj_io_in[7] padframe/mprj_io_inen[7] padframe/mprj_io_out[7] padframe/mprj_io_outen[7]
+ padframe/mprj_io_pd_select[7] padframe/mprj_io_pu_select[7] padframe/mprj_io_schmitt_select[7]
+ padframe/mprj_io_slew_select[7] gpio_control_in_1a\[5\]/resetn gpio_control_in_1\[0\]/resetn
+ gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1\[0\]/serial_clock gpio_control_in_1a\[5\]/serial_data_in
+ gpio_control_in_1\[0\]/serial_data_in gpio_control_in_1a\[5\]/serial_load gpio_control_in_1\[0\]/serial_load
+ mprj/io_in[7] mprj/io_oeb[7] mprj/io_out[7] gpio_control_in_1a\[5\]/zero gpio_control_block
Xgpio_defaults_block_31 gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[1]
+ gpio_defaults_block_31/gpio_defaults[2] gpio_defaults_block_31/gpio_defaults[3]
+ gpio_defaults_block_31/gpio_defaults[4] gpio_defaults_block_31/gpio_defaults[5]
+ gpio_defaults_block_31/gpio_defaults[6] gpio_defaults_block_31/gpio_defaults[7]
+ gpio_defaults_block_31/gpio_defaults[8] gpio_defaults_block_31/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_32 gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[1]
+ gpio_defaults_block_32/gpio_defaults[2] gpio_defaults_block_32/gpio_defaults[3]
+ gpio_defaults_block_32/gpio_defaults[4] gpio_defaults_block_32/gpio_defaults[5]
+ gpio_defaults_block_32/gpio_defaults[6] gpio_defaults_block_32/gpio_defaults[7]
+ gpio_defaults_block_32/gpio_defaults[8] gpio_defaults_block_32/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_bidir_2\[2\] soc/VDD soc/VSS gpio_defaults_block_32/gpio_defaults[0]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] housekeeping/mgmt_gpio_in[37] housekeeping/mgmt_gpio_oeb[37]
+ housekeeping/mgmt_gpio_out[37] gpio_control_bidir_2\[2\]/one padframe/mprj_io_drive_sel[74]
+ padframe/mprj_io_drive_sel[75] padframe/mprj_io_in[37] padframe/mprj_io_inen[37]
+ padframe/mprj_io_out[37] padframe/mprj_io_outen[37] padframe/mprj_io_pd_select[37]
+ padframe/mprj_io_pu_select[37] padframe/mprj_io_schmitt_select[37] padframe/mprj_io_slew_select[37]
+ housekeeping/serial_resetn gpio_control_bidir_2\[1\]/resetn housekeeping/serial_clock
+ gpio_control_bidir_2\[1\]/serial_clock housekeeping/serial_data_2 gpio_control_bidir_2\[1\]/serial_data_in
+ housekeeping/serial_load gpio_control_bidir_2\[1\]/serial_load mprj/io_in[37] mprj/io_oeb[37]
+ mprj/io_out[37] gpio_control_bidir_2\[2\]/zero gpio_control_block
.ends

