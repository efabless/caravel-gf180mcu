VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_core
  CLASS BLOCK ;
  FOREIGN caravel_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 3170.000 BY 4360.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 14.080 17.440 24.080 4341.600 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.080 17.440 3154.960 27.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.080 4331.600 3154.960 4341.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3144.960 17.440 3154.960 4341.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.080 5.440 109.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.080 4275.080 109.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 186.080 5.440 189.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 186.080 4275.080 189.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 266.080 5.440 269.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 266.080 4275.080 269.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 346.080 5.440 349.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 346.080 4275.080 349.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.080 5.440 429.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.080 4275.080 429.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.080 5.440 509.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.080 4275.080 509.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.080 5.440 589.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.080 4275.080 589.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 666.080 5.440 669.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 666.080 4275.080 669.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 746.080 5.440 749.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 746.080 4275.080 749.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 826.080 5.440 829.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 826.080 4275.080 829.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.080 5.440 909.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.080 4275.080 909.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.080 5.440 989.080 66.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.080 545.520 989.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.080 4275.080 989.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1066.080 5.440 1069.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1066.080 4275.080 1069.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1146.080 5.440 1149.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1146.080 4275.080 1149.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1226.080 5.440 1229.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1226.080 4275.080 1229.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1306.080 5.440 1309.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1306.080 4275.080 1309.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1386.080 5.440 1389.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1386.080 4275.080 1389.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1466.080 5.440 1469.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1466.080 4275.080 1469.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 5.440 1549.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 4275.080 1549.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1626.080 5.440 1629.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1626.080 4275.080 1629.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1706.080 5.440 1709.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1706.080 4275.080 1709.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1786.080 5.440 1789.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1786.080 4275.080 1789.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1866.080 5.440 1869.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1866.080 4275.080 1869.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1946.080 5.440 1949.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1946.080 4275.080 1949.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2026.080 5.440 2029.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2026.080 4275.080 2029.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2106.080 5.440 2109.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2106.080 4275.080 2109.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2186.080 5.440 2189.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2186.080 4275.080 2189.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2266.080 5.440 2269.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2266.080 4275.080 2269.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2346.080 5.440 2349.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2346.080 4275.080 2349.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2426.080 5.440 2429.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2426.080 999.280 2429.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2426.080 4275.080 2429.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.080 5.440 2509.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.080 999.280 2509.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.080 4275.080 2509.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.080 5.440 2589.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.080 999.280 2589.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.080 4275.080 2589.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 5.440 2669.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 999.280 2669.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 4275.080 2669.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.080 5.440 2749.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.080 999.280 2749.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.080 4275.080 2749.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.080 5.440 2829.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.080 999.280 2829.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.080 4275.080 2829.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 5.440 2909.080 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 144.725 2909.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 999.280 2909.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 4275.080 2909.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.080 5.440 2989.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.080 999.280 2989.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.080 4275.080 2989.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3099.080 5.440 3102.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3126.620 5.440 3129.620 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 36.080 5.440 39.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.940 5.440 63.940 4353.600 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 56.590 3166.960 59.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 116.590 2896.355 119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 176.590 3166.960 179.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 236.590 2432.720 239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 296.590 2432.720 299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 356.590 2432.720 359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 416.590 2432.720 419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 476.590 2432.720 479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 536.590 2432.720 539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 596.590 2432.720 599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 656.590 2432.720 659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 716.590 2432.720 719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 776.590 2432.720 779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 836.590 2432.720 839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 896.590 601.540 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 956.590 601.540 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1016.590 3166.960 1019.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1076.590 1561.540 1079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1136.590 3166.960 1139.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1196.590 3166.960 1199.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1256.590 3166.960 1259.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1316.590 94.615 1319.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1376.590 94.615 1379.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1436.590 94.615 1439.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1496.590 94.615 1499.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1556.590 94.615 1559.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1616.590 94.615 1619.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1676.590 94.615 1679.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1736.590 94.615 1739.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1796.590 94.615 1799.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1856.590 94.615 1859.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1916.590 94.615 1919.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1976.590 94.615 1979.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2036.590 94.615 2039.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2096.590 94.615 2099.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2156.590 94.615 2159.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2216.590 94.615 2219.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2276.590 94.615 2279.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2336.590 94.615 2339.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2396.590 94.615 2399.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2456.590 94.615 2459.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2516.590 94.615 2519.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2576.590 94.615 2579.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2636.590 94.615 2639.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2696.590 94.615 2699.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2756.590 94.615 2759.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2816.590 94.615 2819.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2876.590 94.615 2879.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2936.590 94.615 2939.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2996.590 94.615 2999.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3056.590 94.615 3059.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3116.590 94.615 3119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3176.590 94.615 3179.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3236.590 94.615 3239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3296.590 94.615 3299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3356.590 94.615 3359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3416.590 94.615 3419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3476.590 94.615 3479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3536.590 94.615 3539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3596.590 94.615 3599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3656.590 94.615 3659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3716.590 94.615 3719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3776.590 94.615 3779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3836.590 94.615 3839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3896.590 94.615 3899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3956.590 94.615 3959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4016.590 94.615 4019.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4076.590 94.615 4079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4136.590 94.615 4139.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4196.590 94.615 4199.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4256.590 94.615 4259.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4316.590 3166.960 4319.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 677.460 896.590 1081.540 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 677.460 956.590 1081.540 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1157.460 896.590 2432.720 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1157.460 956.590 2432.720 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1637.460 1076.590 2121.040 1079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2196.960 1076.590 3166.960 1079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2966.995 116.590 3166.960 119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 236.590 3166.960 239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 296.590 3166.960 299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 356.590 3166.960 359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 416.590 3166.960 419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 476.590 3166.960 479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 536.590 3166.960 539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 596.590 3166.960 599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 656.590 3166.960 659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 716.590 3166.960 719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 776.590 3166.960 779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 836.590 3166.960 839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 896.590 3166.960 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 956.590 3166.960 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1316.590 3166.960 1319.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1376.590 3166.960 1379.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1436.590 3166.960 1439.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1496.590 3166.960 1499.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1556.590 3166.960 1559.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1616.590 3166.960 1619.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1676.590 3166.960 1679.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1736.590 3166.960 1739.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1796.590 3166.960 1799.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1856.590 3166.960 1859.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1916.590 3166.960 1919.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1976.590 3166.960 1979.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2036.590 3166.960 2039.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2096.590 3166.960 2099.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2156.590 3166.960 2159.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2216.590 3166.960 2219.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2276.590 3166.960 2279.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2336.590 3166.960 2339.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2396.590 3166.960 2399.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2456.590 3166.960 2459.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2516.590 3166.960 2519.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2576.590 3166.960 2579.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2636.590 3166.960 2639.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2696.590 3166.960 2699.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2756.590 3166.960 2759.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2816.590 3166.960 2819.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2876.590 3166.960 2879.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2936.590 3166.960 2939.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2996.590 3166.960 2999.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3056.590 3166.960 3059.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3116.590 3166.960 3119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3176.590 3166.960 3179.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3236.590 3166.960 3239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3296.590 3166.960 3299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3356.590 3166.960 3359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3416.590 3166.960 3419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3476.590 3166.960 3479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3536.590 3166.960 3539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3596.590 3166.960 3599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3656.590 3166.960 3659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3716.590 3166.960 3719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3776.590 3166.960 3779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3836.590 3166.960 3839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3896.590 3166.960 3899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3956.590 3166.960 3959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4016.590 3166.960 4019.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4076.590 3166.960 4079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4136.590 3166.960 4139.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4196.590 3166.960 4199.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4256.590 3166.960 4259.590 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2331.080 5.440 2334.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2331.080 4275.080 2334.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2880.580 5.440 2883.580 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2880.580 999.280 2883.580 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2880.580 4275.080 2883.580 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2163.080 5.440 2166.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2163.080 4275.080 2166.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1916.380 5.440 1919.380 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1916.380 4275.080 1919.380 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1359.380 5.440 1362.380 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1359.380 4275.080 1362.380 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1116.480 5.440 1119.480 899.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1116.480 967.380 1119.480 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1116.480 4275.080 1119.480 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 864.780 5.440 867.780 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 864.780 4275.080 867.780 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 556.280 5.440 559.280 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 556.280 4275.080 559.280 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 306.580 5.440 309.580 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 306.580 4275.080 309.580 4353.600 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 2.080 5.440 12.080 4353.600 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 5.440 3166.960 15.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4343.600 3166.960 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3156.960 5.440 3166.960 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.080 5.440 131.080 66.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.080 545.520 131.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.080 4275.080 131.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.080 5.440 211.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.080 4275.080 211.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 288.080 5.440 291.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 288.080 4275.080 291.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.080 5.440 371.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.080 4275.080 371.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.080 5.440 451.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.080 4275.080 451.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 528.080 5.440 531.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 528.080 4275.080 531.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 608.080 5.440 611.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 608.080 4275.080 611.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 688.080 5.440 691.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 688.080 4275.080 691.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 768.080 5.440 771.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 768.080 4275.080 771.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 848.080 5.440 851.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 848.080 4275.080 851.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 928.080 5.440 931.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 928.080 4275.080 931.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1008.080 5.440 1011.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1008.080 4275.080 1011.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.080 5.440 1091.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.080 4275.080 1091.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1168.080 5.440 1171.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1168.080 4275.080 1171.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1248.080 5.440 1251.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1248.080 4275.080 1251.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1328.080 5.440 1331.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1328.080 4275.080 1331.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1408.080 5.440 1411.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1408.080 4275.080 1411.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1488.080 5.440 1491.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1488.080 4275.080 1491.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1568.080 5.440 1571.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1568.080 4275.080 1571.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1648.080 5.440 1651.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1648.080 4275.080 1651.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1728.080 5.440 1731.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1728.080 4275.080 1731.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1808.080 5.440 1811.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1808.080 4275.080 1811.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1888.080 5.440 1891.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1888.080 4275.080 1891.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.080 5.440 1971.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.080 4275.080 1971.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2048.080 5.440 2051.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2048.080 4275.080 2051.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2128.080 5.440 2131.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2128.080 4275.080 2131.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2208.080 5.440 2211.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2208.080 4275.080 2211.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2288.080 5.440 2291.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2288.080 4275.080 2291.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2368.080 5.440 2371.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2368.080 4275.080 2371.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.080 5.440 2451.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.080 999.280 2451.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.080 4275.080 2451.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2528.080 5.440 2531.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2528.080 999.280 2531.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2528.080 4275.080 2531.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2608.080 5.440 2611.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2608.080 999.280 2611.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2608.080 4275.080 2611.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 5.440 2691.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 999.280 2691.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 4275.080 2691.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2768.080 5.440 2771.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2768.080 999.280 2771.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2768.080 4275.080 2771.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2848.080 5.440 2851.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2848.080 999.280 2851.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2848.080 4275.080 2851.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 5.440 2931.080 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 144.725 2931.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 999.280 2931.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 4275.080 2931.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3008.080 5.440 3011.080 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3008.080 999.280 3011.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3008.080 4275.080 3011.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3108.080 5.440 3111.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3135.620 5.440 3138.620 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 45.080 5.440 48.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 69.940 5.440 72.940 4353.600 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 86.590 2896.855 89.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 146.590 2896.355 149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 206.590 2432.720 209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 266.590 2432.720 269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 326.590 2432.720 329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 386.590 2432.720 389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 446.590 2432.720 449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 506.590 2432.720 509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 566.590 2432.720 569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 626.590 2432.720 629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 686.590 2432.720 689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 746.590 2432.720 749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 806.590 2432.720 809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 866.590 2432.720 869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 926.590 601.540 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 986.590 2432.720 989.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1046.590 1561.540 1049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1106.590 1561.540 1109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1166.590 3166.960 1169.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1226.590 3166.960 1229.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1286.590 94.615 1289.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1346.590 94.615 1349.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1406.590 94.615 1409.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1466.590 94.615 1469.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1526.590 94.615 1529.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1586.590 94.615 1589.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1646.590 94.615 1649.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1706.590 94.615 1709.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1766.590 94.615 1769.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1826.590 94.615 1829.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1886.590 94.615 1889.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1946.590 94.615 1949.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2006.590 94.615 2009.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2066.590 94.615 2069.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2126.590 94.615 2129.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2186.590 94.615 2189.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2246.590 94.615 2249.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2306.590 94.615 2309.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2366.590 94.615 2369.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2426.590 94.615 2429.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2486.590 94.615 2489.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2546.590 94.615 2549.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2606.590 94.615 2609.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2666.590 94.615 2669.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2726.590 94.615 2729.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2786.590 94.615 2789.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2846.590 94.615 2849.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2906.590 94.615 2909.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2966.590 94.615 2969.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3026.590 94.615 3029.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3086.590 94.615 3089.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3146.590 94.615 3149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3206.590 94.615 3209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3266.590 94.615 3269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3326.590 94.615 3329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3386.590 94.615 3389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3446.590 94.615 3449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3506.590 94.615 3509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3566.590 94.615 3569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3626.590 94.615 3629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3686.590 94.615 3689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3746.590 94.615 3749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3806.590 94.615 3809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3866.590 94.615 3869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3926.590 94.615 3929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3986.590 94.615 3989.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4046.590 94.615 4049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4106.590 94.615 4109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4166.590 94.615 4169.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4226.590 94.615 4229.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4286.590 3166.960 4289.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 677.460 926.590 1081.540 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1157.460 926.590 2432.720 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1637.460 1046.590 2121.040 1049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1637.460 1106.590 2121.040 1109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2196.960 1046.590 3166.960 1049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2196.960 1106.590 3166.960 1109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2966.995 86.590 3166.960 89.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2966.995 146.590 3166.960 149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 206.590 3166.960 209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 266.590 3166.960 269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 326.590 3166.960 329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 386.590 3166.960 389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 446.590 3166.960 449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 506.590 3166.960 509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 566.590 3166.960 569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 626.590 3166.960 629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 686.590 3166.960 689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 746.590 3166.960 749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 806.590 3166.960 809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 866.590 3166.960 869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 926.590 3166.960 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3051.280 986.590 3166.960 989.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1286.590 3166.960 1289.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1346.590 3166.960 1349.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1406.590 3166.960 1409.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1466.590 3166.960 1469.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1526.590 3166.960 1529.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1586.590 3166.960 1589.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1646.590 3166.960 1649.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1706.590 3166.960 1709.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1766.590 3166.960 1769.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1826.590 3166.960 1829.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1886.590 3166.960 1889.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 1946.590 3166.960 1949.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2006.590 3166.960 2009.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2066.590 3166.960 2069.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2126.590 3166.960 2129.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2186.590 3166.960 2189.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2246.590 3166.960 2249.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2306.590 3166.960 2309.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2366.590 3166.960 2369.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2426.590 3166.960 2429.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2486.590 3166.960 2489.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2546.590 3166.960 2549.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2606.590 3166.960 2609.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2666.590 3166.960 2669.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2726.590 3166.960 2729.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2786.590 3166.960 2789.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2846.590 3166.960 2849.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2906.590 3166.960 2909.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 2966.590 3166.960 2969.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3026.590 3166.960 3029.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3086.590 3166.960 3089.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3146.590 3166.960 3149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3206.590 3166.960 3209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3266.590 3166.960 3269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3326.590 3166.960 3329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3386.590 3166.960 3389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3446.590 3166.960 3449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3506.590 3166.960 3509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3566.590 3166.960 3569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3626.590 3166.960 3629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3686.590 3166.960 3689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3746.590 3166.960 3749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3806.590 3166.960 3809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3866.590 3166.960 3869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3926.590 3166.960 3929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 3986.590 3166.960 3989.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4046.590 3166.960 4049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4106.590 3166.960 4109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4166.590 3166.960 4169.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3075.235 4226.590 3166.960 4229.590 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2353.080 5.440 2356.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2353.080 4275.080 2356.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2892.580 5.440 2895.580 202.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2892.580 999.280 2895.580 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2892.580 4275.080 2895.580 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2170.080 5.440 2173.080 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2170.080 4275.080 2173.080 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1923.380 5.440 1926.380 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1923.380 4275.080 1926.380 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1366.380 5.440 1369.380 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1366.380 4275.080 1369.380 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1123.480 5.440 1126.480 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1123.480 4275.080 1126.480 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 871.780 5.440 874.780 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 871.780 4275.080 874.780 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.280 5.440 566.280 66.400 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.280 545.520 566.280 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.280 4275.080 566.280 4353.600 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.580 5.440 316.580 1260.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.580 4275.080 316.580 4353.600 ;
    END
  END VSS
  PIN clock_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 790.860 -4.000 791.240 4.000 ;
    END
  END clock_core
  PIN const_one[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.965 -4.000 451.345 4.000 ;
    END
  END const_one[0]
  PIN const_one[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1275.965 -4.220 1276.345 4.000 ;
    END
  END const_one[1]
  PIN const_zero[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2163.670 -4.010 2164.050 4.000 ;
    END
  END const_zero[0]
  PIN const_zero[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1888.670 -4.010 1889.050 4.000 ;
    END
  END const_zero[1]
  PIN const_zero[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1613.670 -4.010 1614.050 4.000 ;
    END
  END const_zero[2]
  PIN const_zero[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1338.665 -4.000 1339.055 4.000 ;
    END
  END const_zero[3]
  PIN const_zero[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.965 -4.050 726.345 4.000 ;
    END
  END const_zero[4]
  PIN const_zero[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 455.330 -4.000 455.710 4.000 ;
    END
  END const_zero[5]
  PIN const_zero[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2373.360 -4.010 2373.740 4.000 ;
    END
  END const_zero[6]
  PIN const_zero[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2375.965 -4.010 2376.345 4.000 ;
    END
  END const_zero[7]
  PIN const_zero[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2380.330 -4.010 2380.710 4.000 ;
    END
  END const_zero[8]
  PIN const_zero[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2438.670 -4.010 2439.050 4.000 ;
    END
  END const_zero[9]
  PIN flash_clk_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1614.400 -4.000 1614.780 4.000 ;
    END
  END flash_clk_frame
  PIN flash_clk_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1615.130 -4.000 1615.510 4.000 ;
    END
  END flash_clk_oe
  PIN flash_csb_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1339.400 -4.000 1339.780 4.000 ;
    END
  END flash_csb_frame
  PIN flash_csb_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1340.130 -4.000 1340.510 4.000 ;
    END
  END flash_csb_oe
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1890.855 -4.000 1891.235 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1889.400 -4.000 1889.780 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1831.385 -4.000 1831.765 4.000 ;
    END
  END flash_io0_ie
  PIN flash_io0_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1890.130 -4.000 1890.510 4.000 ;
    END
  END flash_io0_oe
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2165.860 -4.000 2166.240 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2164.400 -4.000 2164.780 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2106.385 -4.000 2106.765 4.000 ;
    END
  END flash_io1_ie
  PIN flash_io1_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2165.130 -4.000 2165.510 4.000 ;
    END
  END flash_io1_oe
  PIN gpio_drive_select_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2377.110 -4.000 2377.490 4.000 ;
    END
  END gpio_drive_select_core[0]
  PIN gpio_drive_select_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2377.820 -4.500 2378.200 4.000 ;
    END
  END gpio_drive_select_core[1]
  PIN gpio_in_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2440.860 -4.000 2441.240 4.000 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2381.385 -4.000 2381.765 4.000 ;
    END
  END gpio_inenb_core
  PIN gpio_out_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2439.400 -4.000 2439.780 4.000 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2440.130 -4.000 2440.510 4.000 ;
    END
  END gpio_outenb_core
  PIN mprj_io_drive_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 97.110 3174.000 97.490 ;
    END
  END mprj_io_drive_sel[0]
  PIN mprj_io_drive_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 1172.110 3174.000 1172.490 ;
    END
  END mprj_io_drive_sel[10]
  PIN mprj_io_drive_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 1172.820 3174.000 1173.200 ;
    END
  END mprj_io_drive_sel[11]
  PIN mprj_io_drive_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 1387.110 3174.000 1387.490 ;
    END
  END mprj_io_drive_sel[12]
  PIN mprj_io_drive_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 1387.820 3174.000 1388.200 ;
    END
  END mprj_io_drive_sel[13]
  PIN mprj_io_drive_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2247.110 3174.000 2247.490 ;
    END
  END mprj_io_drive_sel[14]
  PIN mprj_io_drive_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2247.820 3174.000 2248.200 ;
    END
  END mprj_io_drive_sel[15]
  PIN mprj_io_drive_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2462.110 3174.000 2462.490 ;
    END
  END mprj_io_drive_sel[16]
  PIN mprj_io_drive_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2462.820 3174.000 2463.200 ;
    END
  END mprj_io_drive_sel[17]
  PIN mprj_io_drive_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2677.110 3174.000 2677.490 ;
    END
  END mprj_io_drive_sel[18]
  PIN mprj_io_drive_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2677.820 3174.000 2678.200 ;
    END
  END mprj_io_drive_sel[19]
  PIN mprj_io_drive_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 97.820 3174.000 98.200 ;
    END
  END mprj_io_drive_sel[1]
  PIN mprj_io_drive_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2892.110 3174.000 2892.490 ;
    END
  END mprj_io_drive_sel[20]
  PIN mprj_io_drive_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2892.820 3174.000 2893.200 ;
    END
  END mprj_io_drive_sel[21]
  PIN mprj_io_drive_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 3107.110 3174.000 3107.490 ;
    END
  END mprj_io_drive_sel[22]
  PIN mprj_io_drive_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 3107.820 3174.000 3108.200 ;
    END
  END mprj_io_drive_sel[23]
  PIN mprj_io_drive_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 3322.110 3174.000 3322.490 ;
    END
  END mprj_io_drive_sel[24]
  PIN mprj_io_drive_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 3322.820 3174.000 3323.200 ;
    END
  END mprj_io_drive_sel[25]
  PIN mprj_io_drive_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 3752.110 3174.000 3752.490 ;
    END
  END mprj_io_drive_sel[26]
  PIN mprj_io_drive_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 3752.820 3174.000 3753.200 ;
    END
  END mprj_io_drive_sel[27]
  PIN mprj_io_drive_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 4182.110 3174.000 4182.490 ;
    END
  END mprj_io_drive_sel[28]
  PIN mprj_io_drive_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 4182.820 3174.000 4183.200 ;
    END
  END mprj_io_drive_sel[29]
  PIN mprj_io_drive_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 312.110 3174.000 312.490 ;
    END
  END mprj_io_drive_sel[2]
  PIN mprj_io_drive_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2982.510 4356.000 2982.890 4364.000 ;
    END
  END mprj_io_drive_sel[30]
  PIN mprj_io_drive_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2981.800 4356.000 2982.180 4364.000 ;
    END
  END mprj_io_drive_sel[31]
  PIN mprj_io_drive_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2432.510 4356.000 2432.890 4364.000 ;
    END
  END mprj_io_drive_sel[32]
  PIN mprj_io_drive_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2431.800 4356.000 2432.180 4364.000 ;
    END
  END mprj_io_drive_sel[33]
  PIN mprj_io_drive_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2157.510 4356.000 2157.890 4364.000 ;
    END
  END mprj_io_drive_sel[34]
  PIN mprj_io_drive_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2156.800 4356.000 2157.180 4364.000 ;
    END
  END mprj_io_drive_sel[35]
  PIN mprj_io_drive_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1882.510 4356.000 1882.890 4364.000 ;
    END
  END mprj_io_drive_sel[36]
  PIN mprj_io_drive_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1881.800 4356.000 1882.180 4364.000 ;
    END
  END mprj_io_drive_sel[37]
  PIN mprj_io_drive_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1332.510 4356.000 1332.890 4364.000 ;
    END
  END mprj_io_drive_sel[38]
  PIN mprj_io_drive_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1331.800 4356.000 1332.180 4364.000 ;
    END
  END mprj_io_drive_sel[39]
  PIN mprj_io_drive_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 312.820 3174.000 313.200 ;
    END
  END mprj_io_drive_sel[3]
  PIN mprj_io_drive_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1057.510 4356.000 1057.890 4364.000 ;
    END
  END mprj_io_drive_sel[40]
  PIN mprj_io_drive_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.800 4356.000 1057.180 4364.000 ;
    END
  END mprj_io_drive_sel[41]
  PIN mprj_io_drive_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.510 4356.000 782.890 4364.000 ;
    END
  END mprj_io_drive_sel[42]
  PIN mprj_io_drive_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 781.800 4356.000 782.180 4364.000 ;
    END
  END mprj_io_drive_sel[43]
  PIN mprj_io_drive_sel[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.510 4356.000 507.890 4364.000 ;
    END
  END mprj_io_drive_sel[44]
  PIN mprj_io_drive_sel[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.800 4356.000 507.180 4364.000 ;
    END
  END mprj_io_drive_sel[45]
  PIN mprj_io_drive_sel[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.510 4356.000 232.890 4364.000 ;
    END
  END mprj_io_drive_sel[46]
  PIN mprj_io_drive_sel[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.800 4356.000 232.180 4364.000 ;
    END
  END mprj_io_drive_sel[47]
  PIN mprj_io_drive_sel[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4237.510 6.500 4237.890 ;
    END
  END mprj_io_drive_sel[48]
  PIN mprj_io_drive_sel[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4236.800 9.000 4237.180 ;
    END
  END mprj_io_drive_sel[49]
  PIN mprj_io_drive_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 527.110 3174.000 527.490 ;
    END
  END mprj_io_drive_sel[4]
  PIN mprj_io_drive_sel[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3417.510 6.500 3417.890 ;
    END
  END mprj_io_drive_sel[50]
  PIN mprj_io_drive_sel[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3416.800 9.000 3417.180 ;
    END
  END mprj_io_drive_sel[51]
  PIN mprj_io_drive_sel[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3212.510 6.500 3212.890 ;
    END
  END mprj_io_drive_sel[52]
  PIN mprj_io_drive_sel[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3211.800 9.000 3212.180 ;
    END
  END mprj_io_drive_sel[53]
  PIN mprj_io_drive_sel[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3007.510 6.500 3007.890 ;
    END
  END mprj_io_drive_sel[54]
  PIN mprj_io_drive_sel[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3006.800 9.000 3007.180 ;
    END
  END mprj_io_drive_sel[55]
  PIN mprj_io_drive_sel[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2802.510 6.500 2802.890 ;
    END
  END mprj_io_drive_sel[56]
  PIN mprj_io_drive_sel[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2801.800 9.000 2802.180 ;
    END
  END mprj_io_drive_sel[57]
  PIN mprj_io_drive_sel[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2597.510 6.500 2597.890 ;
    END
  END mprj_io_drive_sel[58]
  PIN mprj_io_drive_sel[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2596.800 9.000 2597.180 ;
    END
  END mprj_io_drive_sel[59]
  PIN mprj_io_drive_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 527.820 3174.000 528.200 ;
    END
  END mprj_io_drive_sel[5]
  PIN mprj_io_drive_sel[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2392.510 6.500 2392.890 ;
    END
  END mprj_io_drive_sel[60]
  PIN mprj_io_drive_sel[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2391.800 9.000 2392.180 ;
    END
  END mprj_io_drive_sel[61]
  PIN mprj_io_drive_sel[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2187.510 6.500 2187.890 ;
    END
  END mprj_io_drive_sel[62]
  PIN mprj_io_drive_sel[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2186.800 9.000 2187.180 ;
    END
  END mprj_io_drive_sel[63]
  PIN mprj_io_drive_sel[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1572.510 6.500 1572.890 ;
    END
  END mprj_io_drive_sel[64]
  PIN mprj_io_drive_sel[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1571.800 9.000 1572.180 ;
    END
  END mprj_io_drive_sel[65]
  PIN mprj_io_drive_sel[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1367.510 6.500 1367.890 ;
    END
  END mprj_io_drive_sel[66]
  PIN mprj_io_drive_sel[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1366.800 9.000 1367.180 ;
    END
  END mprj_io_drive_sel[67]
  PIN mprj_io_drive_sel[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1162.510 6.500 1162.890 ;
    END
  END mprj_io_drive_sel[68]
  PIN mprj_io_drive_sel[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1161.800 9.000 1162.180 ;
    END
  END mprj_io_drive_sel[69]
  PIN mprj_io_drive_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 742.110 3174.000 742.490 ;
    END
  END mprj_io_drive_sel[6]
  PIN mprj_io_drive_sel[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 957.510 6.500 957.890 ;
    END
  END mprj_io_drive_sel[70]
  PIN mprj_io_drive_sel[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 956.800 9.000 957.180 ;
    END
  END mprj_io_drive_sel[71]
  PIN mprj_io_drive_sel[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 752.510 6.500 752.890 ;
    END
  END mprj_io_drive_sel[72]
  PIN mprj_io_drive_sel[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 751.800 9.000 752.180 ;
    END
  END mprj_io_drive_sel[73]
  PIN mprj_io_drive_sel[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 547.510 6.500 547.890 ;
    END
  END mprj_io_drive_sel[74]
  PIN mprj_io_drive_sel[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 546.800 9.000 547.180 ;
    END
  END mprj_io_drive_sel[75]
  PIN mprj_io_drive_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 742.820 3174.000 743.200 ;
    END
  END mprj_io_drive_sel[7]
  PIN mprj_io_drive_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 957.110 3174.000 957.490 ;
    END
  END mprj_io_drive_sel[8]
  PIN mprj_io_drive_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 957.820 3174.000 958.200 ;
    END
  END mprj_io_drive_sel[9]
  PIN mprj_io_ie[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 101.385 3174.000 101.765 ;
    END
  END mprj_io_ie[0]
  PIN mprj_io_ie[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 2896.385 3174.000 2896.765 ;
    END
  END mprj_io_ie[10]
  PIN mprj_io_ie[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 3111.385 3174.000 3111.765 ;
    END
  END mprj_io_ie[11]
  PIN mprj_io_ie[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 3326.385 3174.000 3326.765 ;
    END
  END mprj_io_ie[12]
  PIN mprj_io_ie[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 3756.385 3174.000 3756.765 ;
    END
  END mprj_io_ie[13]
  PIN mprj_io_ie[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 4186.385 3174.000 4186.765 ;
    END
  END mprj_io_ie[14]
  PIN mprj_io_ie[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2978.235 4356.000 2978.615 4364.000 ;
    END
  END mprj_io_ie[15]
  PIN mprj_io_ie[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2428.235 4356.000 2428.615 4364.000 ;
    END
  END mprj_io_ie[16]
  PIN mprj_io_ie[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2153.235 4356.000 2153.615 4364.000 ;
    END
  END mprj_io_ie[17]
  PIN mprj_io_ie[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1878.235 4356.000 1878.615 4364.000 ;
    END
  END mprj_io_ie[18]
  PIN mprj_io_ie[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1328.235 4356.000 1328.615 4364.000 ;
    END
  END mprj_io_ie[19]
  PIN mprj_io_ie[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 316.385 3174.000 316.765 ;
    END
  END mprj_io_ie[1]
  PIN mprj_io_ie[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1053.235 4356.000 1053.615 4364.000 ;
    END
  END mprj_io_ie[20]
  PIN mprj_io_ie[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 778.235 4356.000 778.615 4364.000 ;
    END
  END mprj_io_ie[21]
  PIN mprj_io_ie[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.235 4356.000 503.615 4364.000 ;
    END
  END mprj_io_ie[22]
  PIN mprj_io_ie[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.235 4356.000 228.615 4364.000 ;
    END
  END mprj_io_ie[23]
  PIN mprj_io_ie[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4233.235 14.000 4233.615 ;
    END
  END mprj_io_ie[24]
  PIN mprj_io_ie[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3413.235 14.000 3413.615 ;
    END
  END mprj_io_ie[25]
  PIN mprj_io_ie[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3208.235 14.000 3208.615 ;
    END
  END mprj_io_ie[26]
  PIN mprj_io_ie[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3003.235 14.000 3003.615 ;
    END
  END mprj_io_ie[27]
  PIN mprj_io_ie[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2798.235 14.000 2798.615 ;
    END
  END mprj_io_ie[28]
  PIN mprj_io_ie[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2593.235 14.000 2593.615 ;
    END
  END mprj_io_ie[29]
  PIN mprj_io_ie[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 531.385 3174.000 531.765 ;
    END
  END mprj_io_ie[2]
  PIN mprj_io_ie[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2388.235 14.000 2388.615 ;
    END
  END mprj_io_ie[30]
  PIN mprj_io_ie[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2183.235 14.000 2183.615 ;
    END
  END mprj_io_ie[31]
  PIN mprj_io_ie[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1568.235 14.000 1568.615 ;
    END
  END mprj_io_ie[32]
  PIN mprj_io_ie[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1363.235 14.000 1363.615 ;
    END
  END mprj_io_ie[33]
  PIN mprj_io_ie[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1158.235 14.000 1158.615 ;
    END
  END mprj_io_ie[34]
  PIN mprj_io_ie[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 953.235 14.000 953.615 ;
    END
  END mprj_io_ie[35]
  PIN mprj_io_ie[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 748.235 14.000 748.615 ;
    END
  END mprj_io_ie[36]
  PIN mprj_io_ie[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 543.235 14.000 543.615 ;
    END
  END mprj_io_ie[37]
  PIN mprj_io_ie[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 746.385 3174.000 746.765 ;
    END
  END mprj_io_ie[3]
  PIN mprj_io_ie[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 961.385 3174.000 961.765 ;
    END
  END mprj_io_ie[4]
  PIN mprj_io_ie[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 1176.385 3174.000 1176.765 ;
    END
  END mprj_io_ie[5]
  PIN mprj_io_ie[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 1391.385 3174.000 1391.765 ;
    END
  END mprj_io_ie[6]
  PIN mprj_io_ie[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 2251.385 3174.000 2251.765 ;
    END
  END mprj_io_ie[7]
  PIN mprj_io_ie[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 2466.385 3174.000 2466.765 ;
    END
  END mprj_io_ie[8]
  PIN mprj_io_ie[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3156.000 2681.385 3174.000 2681.765 ;
    END
  END mprj_io_ie[9]
  PIN mprj_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 160.860 3174.000 161.240 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2955.860 3174.000 2956.240 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 3170.860 3174.000 3171.240 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 3385.860 3174.000 3386.240 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 3815.860 3174.000 3816.240 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 4245.860 3174.000 4246.240 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2918.760 4356.000 2919.140 4364.000 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2368.760 4356.000 2369.140 4364.000 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2093.760 4356.000 2094.140 4364.000 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1818.760 4356.000 1819.140 4364.000 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1268.760 4356.000 1269.140 4364.000 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 375.860 3174.000 376.240 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 993.760 4356.000 994.140 4364.000 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 718.760 4356.000 719.140 4364.000 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.760 4356.000 444.140 4364.000 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.760 4356.000 169.140 4364.000 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4173.760 9.000 4174.140 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3353.760 9.000 3354.140 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3148.760 9.000 3149.140 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2943.760 9.000 2944.140 ;
    END
  END mprj_io_in[27]
  PIN mprj_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2738.760 9.000 2739.140 ;
    END
  END mprj_io_in[28]
  PIN mprj_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2533.760 9.000 2534.140 ;
    END
  END mprj_io_in[29]
  PIN mprj_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 590.860 3174.000 591.240 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2328.760 9.000 2329.140 ;
    END
  END mprj_io_in[30]
  PIN mprj_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2123.760 9.000 2124.140 ;
    END
  END mprj_io_in[31]
  PIN mprj_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1508.760 9.000 1509.140 ;
    END
  END mprj_io_in[32]
  PIN mprj_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1303.760 9.000 1304.140 ;
    END
  END mprj_io_in[33]
  PIN mprj_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1098.760 9.000 1099.140 ;
    END
  END mprj_io_in[34]
  PIN mprj_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 893.760 9.000 894.140 ;
    END
  END mprj_io_in[35]
  PIN mprj_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 688.760 9.000 689.140 ;
    END
  END mprj_io_in[36]
  PIN mprj_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 483.760 9.000 484.140 ;
    END
  END mprj_io_in[37]
  PIN mprj_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 805.860 3174.000 806.240 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 1020.860 3174.000 1021.240 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 1235.860 3174.000 1236.240 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 1450.860 3174.000 1451.240 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2310.860 3174.000 2311.240 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2525.860 3174.000 2526.240 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3161.000 2740.860 3174.000 2741.240 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 160.130 3174.000 160.510 ;
    END
  END mprj_io_oe[0]
  PIN mprj_io_oe[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2955.130 3174.000 2955.510 ;
    END
  END mprj_io_oe[10]
  PIN mprj_io_oe[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 3170.130 3174.000 3170.510 ;
    END
  END mprj_io_oe[11]
  PIN mprj_io_oe[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 3385.130 3174.000 3385.510 ;
    END
  END mprj_io_oe[12]
  PIN mprj_io_oe[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 3815.130 3174.000 3815.510 ;
    END
  END mprj_io_oe[13]
  PIN mprj_io_oe[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 4245.130 3174.000 4245.510 ;
    END
  END mprj_io_oe[14]
  PIN mprj_io_oe[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2919.490 4356.000 2919.870 4364.000 ;
    END
  END mprj_io_oe[15]
  PIN mprj_io_oe[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2369.490 4356.000 2369.870 4364.000 ;
    END
  END mprj_io_oe[16]
  PIN mprj_io_oe[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2094.490 4356.000 2094.870 4364.000 ;
    END
  END mprj_io_oe[17]
  PIN mprj_io_oe[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1819.490 4356.000 1819.870 4364.000 ;
    END
  END mprj_io_oe[18]
  PIN mprj_io_oe[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1269.490 4356.000 1269.870 4364.000 ;
    END
  END mprj_io_oe[19]
  PIN mprj_io_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 375.130 3174.000 375.510 ;
    END
  END mprj_io_oe[1]
  PIN mprj_io_oe[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.490 4356.000 994.870 4364.000 ;
    END
  END mprj_io_oe[20]
  PIN mprj_io_oe[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.490 4356.000 719.870 4364.000 ;
    END
  END mprj_io_oe[21]
  PIN mprj_io_oe[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.490 4356.000 444.870 4364.000 ;
    END
  END mprj_io_oe[22]
  PIN mprj_io_oe[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.490 4356.000 169.870 4364.000 ;
    END
  END mprj_io_oe[23]
  PIN mprj_io_oe[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4174.490 6.500 4174.870 ;
    END
  END mprj_io_oe[24]
  PIN mprj_io_oe[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3354.490 6.500 3354.870 ;
    END
  END mprj_io_oe[25]
  PIN mprj_io_oe[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3149.490 6.500 3149.870 ;
    END
  END mprj_io_oe[26]
  PIN mprj_io_oe[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2944.490 6.500 2944.870 ;
    END
  END mprj_io_oe[27]
  PIN mprj_io_oe[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2739.490 6.500 2739.870 ;
    END
  END mprj_io_oe[28]
  PIN mprj_io_oe[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2534.490 6.500 2534.870 ;
    END
  END mprj_io_oe[29]
  PIN mprj_io_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 590.130 3174.000 590.510 ;
    END
  END mprj_io_oe[2]
  PIN mprj_io_oe[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2329.490 6.500 2329.870 ;
    END
  END mprj_io_oe[30]
  PIN mprj_io_oe[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2124.490 6.500 2124.870 ;
    END
  END mprj_io_oe[31]
  PIN mprj_io_oe[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1509.490 6.500 1509.870 ;
    END
  END mprj_io_oe[32]
  PIN mprj_io_oe[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1304.490 6.500 1304.870 ;
    END
  END mprj_io_oe[33]
  PIN mprj_io_oe[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1099.490 6.500 1099.870 ;
    END
  END mprj_io_oe[34]
  PIN mprj_io_oe[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 894.490 6.500 894.870 ;
    END
  END mprj_io_oe[35]
  PIN mprj_io_oe[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 689.490 6.500 689.870 ;
    END
  END mprj_io_oe[36]
  PIN mprj_io_oe[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 484.490 6.500 484.870 ;
    END
  END mprj_io_oe[37]
  PIN mprj_io_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 805.130 3174.000 805.510 ;
    END
  END mprj_io_oe[3]
  PIN mprj_io_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 1020.130 3174.000 1020.510 ;
    END
  END mprj_io_oe[4]
  PIN mprj_io_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 1235.130 3174.000 1235.510 ;
    END
  END mprj_io_oe[5]
  PIN mprj_io_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 1450.130 3174.000 1450.510 ;
    END
  END mprj_io_oe[6]
  PIN mprj_io_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2310.130 3174.000 2310.510 ;
    END
  END mprj_io_oe[7]
  PIN mprj_io_oe[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2525.130 3174.000 2525.510 ;
    END
  END mprj_io_oe[8]
  PIN mprj_io_oe[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3163.500 2740.130 3174.000 2740.510 ;
    END
  END mprj_io_oe[9]
  PIN mprj_io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 159.400 3174.000 159.780 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2954.400 3174.000 2954.780 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 3169.400 3174.000 3169.780 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 3384.400 3174.000 3384.780 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 3814.400 3174.000 3814.780 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 4244.400 3174.000 4244.780 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2920.220 4356.000 2920.600 4364.000 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2370.220 4356.000 2370.600 4364.000 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2095.220 4356.000 2095.600 4364.000 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1820.220 4356.000 1820.600 4364.000 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1270.220 4356.000 1270.600 4364.000 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 374.400 3174.000 374.780 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 995.220 4356.000 995.600 4364.000 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.220 4356.000 720.600 4364.000 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.220 4356.000 445.600 4364.000 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.220 4356.000 170.600 4364.000 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4175.220 4.000 4175.600 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3355.220 4.000 3355.600 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3150.220 4.000 3150.600 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2945.220 4.000 2945.600 ;
    END
  END mprj_io_out[27]
  PIN mprj_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2740.220 4.000 2740.600 ;
    END
  END mprj_io_out[28]
  PIN mprj_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2535.220 4.000 2535.600 ;
    END
  END mprj_io_out[29]
  PIN mprj_io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 589.400 3174.000 589.780 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2330.220 4.000 2330.600 ;
    END
  END mprj_io_out[30]
  PIN mprj_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2125.220 4.000 2125.600 ;
    END
  END mprj_io_out[31]
  PIN mprj_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1510.220 4.000 1510.600 ;
    END
  END mprj_io_out[32]
  PIN mprj_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1305.220 4.000 1305.600 ;
    END
  END mprj_io_out[33]
  PIN mprj_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1100.220 4.000 1100.600 ;
    END
  END mprj_io_out[34]
  PIN mprj_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 895.220 4.000 895.600 ;
    END
  END mprj_io_out[35]
  PIN mprj_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 690.220 4.000 690.600 ;
    END
  END mprj_io_out[36]
  PIN mprj_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 485.220 4.000 485.600 ;
    END
  END mprj_io_out[37]
  PIN mprj_io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 804.400 3174.000 804.780 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 1019.400 3174.000 1019.780 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 1234.400 3174.000 1234.780 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 1449.400 3174.000 1449.780 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2309.400 3174.000 2309.780 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2524.400 3174.000 2524.780 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2739.400 3174.000 2739.780 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_pulldown_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 100.330 3174.000 100.710 ;
    END
  END mprj_io_pulldown_sel[0]
  PIN mprj_io_pulldown_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 2895.330 3174.000 2895.710 ;
    END
  END mprj_io_pulldown_sel[10]
  PIN mprj_io_pulldown_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 3110.330 3174.000 3110.710 ;
    END
  END mprj_io_pulldown_sel[11]
  PIN mprj_io_pulldown_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 3325.330 3174.000 3325.710 ;
    END
  END mprj_io_pulldown_sel[12]
  PIN mprj_io_pulldown_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 3755.330 3174.000 3755.710 ;
    END
  END mprj_io_pulldown_sel[13]
  PIN mprj_io_pulldown_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 4185.330 3174.000 4185.710 ;
    END
  END mprj_io_pulldown_sel[14]
  PIN mprj_io_pulldown_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2979.290 4356.000 2979.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[15]
  PIN mprj_io_pulldown_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2429.290 4356.000 2429.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[16]
  PIN mprj_io_pulldown_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2154.290 4356.000 2154.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[17]
  PIN mprj_io_pulldown_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1879.290 4356.000 1879.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[18]
  PIN mprj_io_pulldown_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1329.290 4356.000 1329.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[19]
  PIN mprj_io_pulldown_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 315.330 3174.000 315.710 ;
    END
  END mprj_io_pulldown_sel[1]
  PIN mprj_io_pulldown_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1054.290 4356.000 1054.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[20]
  PIN mprj_io_pulldown_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.290 4356.000 779.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[21]
  PIN mprj_io_pulldown_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.290 4356.000 504.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[22]
  PIN mprj_io_pulldown_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.290 4356.000 229.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[23]
  PIN mprj_io_pulldown_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4234.290 11.500 4234.670 ;
    END
  END mprj_io_pulldown_sel[24]
  PIN mprj_io_pulldown_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3414.290 11.500 3414.670 ;
    END
  END mprj_io_pulldown_sel[25]
  PIN mprj_io_pulldown_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3209.290 11.500 3209.670 ;
    END
  END mprj_io_pulldown_sel[26]
  PIN mprj_io_pulldown_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3004.290 11.500 3004.670 ;
    END
  END mprj_io_pulldown_sel[27]
  PIN mprj_io_pulldown_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2799.290 11.500 2799.670 ;
    END
  END mprj_io_pulldown_sel[28]
  PIN mprj_io_pulldown_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2594.290 11.500 2594.670 ;
    END
  END mprj_io_pulldown_sel[29]
  PIN mprj_io_pulldown_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 530.330 3174.000 530.710 ;
    END
  END mprj_io_pulldown_sel[2]
  PIN mprj_io_pulldown_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2389.290 11.500 2389.670 ;
    END
  END mprj_io_pulldown_sel[30]
  PIN mprj_io_pulldown_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2184.290 11.500 2184.670 ;
    END
  END mprj_io_pulldown_sel[31]
  PIN mprj_io_pulldown_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1569.290 11.500 1569.670 ;
    END
  END mprj_io_pulldown_sel[32]
  PIN mprj_io_pulldown_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1364.290 11.500 1364.670 ;
    END
  END mprj_io_pulldown_sel[33]
  PIN mprj_io_pulldown_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1159.290 11.500 1159.670 ;
    END
  END mprj_io_pulldown_sel[34]
  PIN mprj_io_pulldown_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 954.290 11.500 954.670 ;
    END
  END mprj_io_pulldown_sel[35]
  PIN mprj_io_pulldown_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 749.290 11.500 749.670 ;
    END
  END mprj_io_pulldown_sel[36]
  PIN mprj_io_pulldown_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 544.290 11.500 544.670 ;
    END
  END mprj_io_pulldown_sel[37]
  PIN mprj_io_pulldown_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 745.330 3174.000 745.710 ;
    END
  END mprj_io_pulldown_sel[3]
  PIN mprj_io_pulldown_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 960.330 3174.000 960.710 ;
    END
  END mprj_io_pulldown_sel[4]
  PIN mprj_io_pulldown_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 1175.330 3174.000 1175.710 ;
    END
  END mprj_io_pulldown_sel[5]
  PIN mprj_io_pulldown_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 1390.330 3174.000 1390.710 ;
    END
  END mprj_io_pulldown_sel[6]
  PIN mprj_io_pulldown_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 2250.330 3174.000 2250.710 ;
    END
  END mprj_io_pulldown_sel[7]
  PIN mprj_io_pulldown_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 2465.330 3174.000 2465.710 ;
    END
  END mprj_io_pulldown_sel[8]
  PIN mprj_io_pulldown_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3158.500 2680.330 3174.000 2680.710 ;
    END
  END mprj_io_pulldown_sel[9]
  PIN mprj_io_pullup_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 95.965 3174.000 96.345 ;
    END
  END mprj_io_pullup_sel[0]
  PIN mprj_io_pullup_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2890.965 3174.000 2891.345 ;
    END
  END mprj_io_pullup_sel[10]
  PIN mprj_io_pullup_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 3105.965 3174.000 3106.345 ;
    END
  END mprj_io_pullup_sel[11]
  PIN mprj_io_pullup_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 3320.965 3174.000 3321.345 ;
    END
  END mprj_io_pullup_sel[12]
  PIN mprj_io_pullup_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 3750.965 3174.000 3751.345 ;
    END
  END mprj_io_pullup_sel[13]
  PIN mprj_io_pullup_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 4180.965 3174.000 4181.345 ;
    END
  END mprj_io_pullup_sel[14]
  PIN mprj_io_pullup_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2983.655 4356.000 2984.035 4364.000 ;
    END
  END mprj_io_pullup_sel[15]
  PIN mprj_io_pullup_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2433.655 4356.000 2434.035 4364.000 ;
    END
  END mprj_io_pullup_sel[16]
  PIN mprj_io_pullup_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2158.655 4356.000 2159.035 4364.000 ;
    END
  END mprj_io_pullup_sel[17]
  PIN mprj_io_pullup_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1883.655 4356.000 1884.035 4364.000 ;
    END
  END mprj_io_pullup_sel[18]
  PIN mprj_io_pullup_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1333.655 4356.000 1334.035 4364.000 ;
    END
  END mprj_io_pullup_sel[19]
  PIN mprj_io_pullup_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 310.965 3174.000 311.345 ;
    END
  END mprj_io_pullup_sel[1]
  PIN mprj_io_pullup_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1058.655 4356.000 1059.035 4364.000 ;
    END
  END mprj_io_pullup_sel[20]
  PIN mprj_io_pullup_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 783.655 4356.000 784.035 4364.000 ;
    END
  END mprj_io_pullup_sel[21]
  PIN mprj_io_pullup_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.655 4356.000 509.035 4364.000 ;
    END
  END mprj_io_pullup_sel[22]
  PIN mprj_io_pullup_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 233.655 4356.000 234.035 4364.000 ;
    END
  END mprj_io_pullup_sel[23]
  PIN mprj_io_pullup_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4238.655 4.000 4239.035 ;
    END
  END mprj_io_pullup_sel[24]
  PIN mprj_io_pullup_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3418.655 4.000 3419.035 ;
    END
  END mprj_io_pullup_sel[25]
  PIN mprj_io_pullup_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3213.655 4.000 3214.035 ;
    END
  END mprj_io_pullup_sel[26]
  PIN mprj_io_pullup_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3008.655 4.000 3009.035 ;
    END
  END mprj_io_pullup_sel[27]
  PIN mprj_io_pullup_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2803.655 4.000 2804.035 ;
    END
  END mprj_io_pullup_sel[28]
  PIN mprj_io_pullup_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2598.655 4.000 2599.035 ;
    END
  END mprj_io_pullup_sel[29]
  PIN mprj_io_pullup_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 525.965 3174.000 526.345 ;
    END
  END mprj_io_pullup_sel[2]
  PIN mprj_io_pullup_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2393.655 4.000 2394.035 ;
    END
  END mprj_io_pullup_sel[30]
  PIN mprj_io_pullup_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2188.655 4.000 2189.035 ;
    END
  END mprj_io_pullup_sel[31]
  PIN mprj_io_pullup_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1573.655 4.000 1574.035 ;
    END
  END mprj_io_pullup_sel[32]
  PIN mprj_io_pullup_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1368.655 4.000 1369.035 ;
    END
  END mprj_io_pullup_sel[33]
  PIN mprj_io_pullup_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1163.655 4.000 1164.035 ;
    END
  END mprj_io_pullup_sel[34]
  PIN mprj_io_pullup_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 958.655 4.000 959.035 ;
    END
  END mprj_io_pullup_sel[35]
  PIN mprj_io_pullup_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 753.655 4.000 754.035 ;
    END
  END mprj_io_pullup_sel[36]
  PIN mprj_io_pullup_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 548.655 4.000 549.035 ;
    END
  END mprj_io_pullup_sel[37]
  PIN mprj_io_pullup_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 740.965 3174.000 741.345 ;
    END
  END mprj_io_pullup_sel[3]
  PIN mprj_io_pullup_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 955.965 3174.000 956.345 ;
    END
  END mprj_io_pullup_sel[4]
  PIN mprj_io_pullup_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 1170.965 3174.000 1171.345 ;
    END
  END mprj_io_pullup_sel[5]
  PIN mprj_io_pullup_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 1385.965 3174.000 1386.345 ;
    END
  END mprj_io_pullup_sel[6]
  PIN mprj_io_pullup_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2245.965 3174.000 2246.345 ;
    END
  END mprj_io_pullup_sel[7]
  PIN mprj_io_pullup_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2460.965 3174.000 2461.345 ;
    END
  END mprj_io_pullup_sel[8]
  PIN mprj_io_pullup_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3166.000 2675.965 3174.000 2676.345 ;
    END
  END mprj_io_pullup_sel[9]
  PIN mprj_io_schmitt_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 93.360 3174.000 93.740 ;
    END
  END mprj_io_schmitt_sel[0]
  PIN mprj_io_schmitt_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2888.360 3174.000 2888.740 ;
    END
  END mprj_io_schmitt_sel[10]
  PIN mprj_io_schmitt_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 3103.360 3174.000 3103.740 ;
    END
  END mprj_io_schmitt_sel[11]
  PIN mprj_io_schmitt_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 3318.360 3174.000 3318.740 ;
    END
  END mprj_io_schmitt_sel[12]
  PIN mprj_io_schmitt_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 3748.360 3174.000 3748.740 ;
    END
  END mprj_io_schmitt_sel[13]
  PIN mprj_io_schmitt_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 4178.360 3174.000 4178.740 ;
    END
  END mprj_io_schmitt_sel[14]
  PIN mprj_io_schmitt_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2986.260 4356.000 2986.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[15]
  PIN mprj_io_schmitt_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2436.260 4356.000 2436.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[16]
  PIN mprj_io_schmitt_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2161.260 4356.000 2161.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[17]
  PIN mprj_io_schmitt_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1886.260 4356.000 1886.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[18]
  PIN mprj_io_schmitt_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1336.260 4356.000 1336.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[19]
  PIN mprj_io_schmitt_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 308.360 3174.000 308.740 ;
    END
  END mprj_io_schmitt_sel[1]
  PIN mprj_io_schmitt_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1061.260 4356.000 1061.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[20]
  PIN mprj_io_schmitt_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.260 4356.000 786.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[21]
  PIN mprj_io_schmitt_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.260 4356.000 511.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[22]
  PIN mprj_io_schmitt_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.260 4356.000 236.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[23]
  PIN mprj_io_schmitt_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4241.260 1.500 4241.640 ;
    END
  END mprj_io_schmitt_sel[24]
  PIN mprj_io_schmitt_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3421.260 1.500 3421.640 ;
    END
  END mprj_io_schmitt_sel[25]
  PIN mprj_io_schmitt_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3216.260 1.500 3216.640 ;
    END
  END mprj_io_schmitt_sel[26]
  PIN mprj_io_schmitt_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3011.260 1.500 3011.640 ;
    END
  END mprj_io_schmitt_sel[27]
  PIN mprj_io_schmitt_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2806.260 1.500 2806.640 ;
    END
  END mprj_io_schmitt_sel[28]
  PIN mprj_io_schmitt_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2601.260 1.500 2601.640 ;
    END
  END mprj_io_schmitt_sel[29]
  PIN mprj_io_schmitt_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 523.360 3174.000 523.740 ;
    END
  END mprj_io_schmitt_sel[2]
  PIN mprj_io_schmitt_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2396.260 1.500 2396.640 ;
    END
  END mprj_io_schmitt_sel[30]
  PIN mprj_io_schmitt_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2191.260 1.500 2191.640 ;
    END
  END mprj_io_schmitt_sel[31]
  PIN mprj_io_schmitt_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1576.260 1.500 1576.640 ;
    END
  END mprj_io_schmitt_sel[32]
  PIN mprj_io_schmitt_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1371.260 1.500 1371.640 ;
    END
  END mprj_io_schmitt_sel[33]
  PIN mprj_io_schmitt_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1166.260 1.500 1166.640 ;
    END
  END mprj_io_schmitt_sel[34]
  PIN mprj_io_schmitt_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 961.260 1.500 961.640 ;
    END
  END mprj_io_schmitt_sel[35]
  PIN mprj_io_schmitt_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 756.260 1.500 756.640 ;
    END
  END mprj_io_schmitt_sel[36]
  PIN mprj_io_schmitt_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 551.260 1.500 551.640 ;
    END
  END mprj_io_schmitt_sel[37]
  PIN mprj_io_schmitt_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 738.360 3174.000 738.740 ;
    END
  END mprj_io_schmitt_sel[3]
  PIN mprj_io_schmitt_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 953.360 3174.000 953.740 ;
    END
  END mprj_io_schmitt_sel[4]
  PIN mprj_io_schmitt_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 1168.360 3174.000 1168.740 ;
    END
  END mprj_io_schmitt_sel[5]
  PIN mprj_io_schmitt_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 1383.360 3174.000 1383.740 ;
    END
  END mprj_io_schmitt_sel[6]
  PIN mprj_io_schmitt_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2243.360 3174.000 2243.740 ;
    END
  END mprj_io_schmitt_sel[7]
  PIN mprj_io_schmitt_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2458.360 3174.000 2458.740 ;
    END
  END mprj_io_schmitt_sel[8]
  PIN mprj_io_schmitt_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2673.360 3174.000 2673.740 ;
    END
  END mprj_io_schmitt_sel[9]
  PIN mprj_io_slew_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 158.670 3174.000 159.050 ;
    END
  END mprj_io_slew_sel[0]
  PIN mprj_io_slew_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2953.670 3174.000 2954.050 ;
    END
  END mprj_io_slew_sel[10]
  PIN mprj_io_slew_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 3168.670 3174.000 3169.050 ;
    END
  END mprj_io_slew_sel[11]
  PIN mprj_io_slew_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 3383.670 3174.000 3384.050 ;
    END
  END mprj_io_slew_sel[12]
  PIN mprj_io_slew_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 3813.670 3174.000 3814.050 ;
    END
  END mprj_io_slew_sel[13]
  PIN mprj_io_slew_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 4243.670 3174.000 4244.050 ;
    END
  END mprj_io_slew_sel[14]
  PIN mprj_io_slew_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2920.950 4356.000 2921.330 4364.000 ;
    END
  END mprj_io_slew_sel[15]
  PIN mprj_io_slew_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2370.950 4356.000 2371.330 4364.000 ;
    END
  END mprj_io_slew_sel[16]
  PIN mprj_io_slew_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2095.950 4356.000 2096.330 4364.000 ;
    END
  END mprj_io_slew_sel[17]
  PIN mprj_io_slew_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1820.950 4356.000 1821.330 4364.000 ;
    END
  END mprj_io_slew_sel[18]
  PIN mprj_io_slew_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1270.950 4356.000 1271.330 4364.000 ;
    END
  END mprj_io_slew_sel[19]
  PIN mprj_io_slew_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 373.670 3174.000 374.050 ;
    END
  END mprj_io_slew_sel[1]
  PIN mprj_io_slew_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 995.950 4356.000 996.330 4364.000 ;
    END
  END mprj_io_slew_sel[20]
  PIN mprj_io_slew_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.950 4356.000 721.330 4364.000 ;
    END
  END mprj_io_slew_sel[21]
  PIN mprj_io_slew_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.950 4356.000 446.330 4364.000 ;
    END
  END mprj_io_slew_sel[22]
  PIN mprj_io_slew_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.950 4356.000 171.330 4364.000 ;
    END
  END mprj_io_slew_sel[23]
  PIN mprj_io_slew_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 4175.950 1.500 4176.330 ;
    END
  END mprj_io_slew_sel[24]
  PIN mprj_io_slew_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3355.950 1.500 3356.330 ;
    END
  END mprj_io_slew_sel[25]
  PIN mprj_io_slew_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 3150.950 1.500 3151.330 ;
    END
  END mprj_io_slew_sel[26]
  PIN mprj_io_slew_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2945.950 1.500 2946.330 ;
    END
  END mprj_io_slew_sel[27]
  PIN mprj_io_slew_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2740.950 1.500 2741.330 ;
    END
  END mprj_io_slew_sel[28]
  PIN mprj_io_slew_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2535.950 1.500 2536.330 ;
    END
  END mprj_io_slew_sel[29]
  PIN mprj_io_slew_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 588.670 3174.000 589.050 ;
    END
  END mprj_io_slew_sel[2]
  PIN mprj_io_slew_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2330.950 1.500 2331.330 ;
    END
  END mprj_io_slew_sel[30]
  PIN mprj_io_slew_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 2125.950 1.500 2126.330 ;
    END
  END mprj_io_slew_sel[31]
  PIN mprj_io_slew_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1510.950 1.500 1511.330 ;
    END
  END mprj_io_slew_sel[32]
  PIN mprj_io_slew_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1305.950 1.500 1306.330 ;
    END
  END mprj_io_slew_sel[33]
  PIN mprj_io_slew_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 1100.950 1.500 1101.330 ;
    END
  END mprj_io_slew_sel[34]
  PIN mprj_io_slew_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 895.950 1.500 896.330 ;
    END
  END mprj_io_slew_sel[35]
  PIN mprj_io_slew_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 690.950 1.500 691.330 ;
    END
  END mprj_io_slew_sel[36]
  PIN mprj_io_slew_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -4.000 485.950 1.500 486.330 ;
    END
  END mprj_io_slew_sel[37]
  PIN mprj_io_slew_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 803.670 3174.000 804.050 ;
    END
  END mprj_io_slew_sel[3]
  PIN mprj_io_slew_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 1018.670 3174.000 1019.050 ;
    END
  END mprj_io_slew_sel[4]
  PIN mprj_io_slew_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 1233.670 3174.000 1234.050 ;
    END
  END mprj_io_slew_sel[5]
  PIN mprj_io_slew_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 1448.670 3174.000 1449.050 ;
    END
  END mprj_io_slew_sel[6]
  PIN mprj_io_slew_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2308.670 3174.000 2309.050 ;
    END
  END mprj_io_slew_sel[7]
  PIN mprj_io_slew_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2523.670 3174.000 2524.050 ;
    END
  END mprj_io_slew_sel[8]
  PIN mprj_io_slew_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3168.500 2738.670 3174.000 2739.050 ;
    END
  END mprj_io_slew_sel[9]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 515.860 -4.000 516.240 4.000 ;
    END
  END rstb
  OBS
      LAYER Metal1 ;
        RECT 2.890 25.350 3169.510 4354.410 ;
      LAYER Metal2 ;
        RECT 1.260 4355.700 168.460 4356.660 ;
        RECT 171.630 4355.700 227.935 4356.660 ;
        RECT 228.915 4355.700 228.990 4356.660 ;
        RECT 229.970 4355.700 231.500 4356.660 ;
        RECT 233.190 4355.700 233.355 4356.660 ;
        RECT 234.335 4355.700 235.960 4356.660 ;
        RECT 236.940 4355.700 443.460 4356.660 ;
        RECT 446.630 4355.700 502.935 4356.660 ;
        RECT 503.915 4355.700 503.990 4356.660 ;
        RECT 504.970 4355.700 506.500 4356.660 ;
        RECT 508.190 4355.700 508.355 4356.660 ;
        RECT 509.335 4355.700 510.960 4356.660 ;
        RECT 511.940 4355.700 718.460 4356.660 ;
        RECT 721.630 4355.700 777.935 4356.660 ;
        RECT 778.915 4355.700 778.990 4356.660 ;
        RECT 779.970 4355.700 781.500 4356.660 ;
        RECT 783.190 4355.700 783.355 4356.660 ;
        RECT 784.335 4355.700 785.960 4356.660 ;
        RECT 786.940 4355.700 993.460 4356.660 ;
        RECT 996.630 4355.700 1052.935 4356.660 ;
        RECT 1053.915 4355.700 1053.990 4356.660 ;
        RECT 1054.970 4355.700 1056.500 4356.660 ;
        RECT 1058.190 4355.700 1058.355 4356.660 ;
        RECT 1059.335 4355.700 1060.960 4356.660 ;
        RECT 1061.940 4355.700 1268.460 4356.660 ;
        RECT 1271.630 4355.700 1327.935 4356.660 ;
        RECT 1328.915 4355.700 1328.990 4356.660 ;
        RECT 1329.970 4355.700 1331.500 4356.660 ;
        RECT 1333.190 4355.700 1333.355 4356.660 ;
        RECT 1334.335 4355.700 1335.960 4356.660 ;
        RECT 1336.940 4355.700 1818.460 4356.660 ;
        RECT 1821.630 4355.700 1877.935 4356.660 ;
        RECT 1878.915 4355.700 1878.990 4356.660 ;
        RECT 1879.970 4355.700 1881.500 4356.660 ;
        RECT 1883.190 4355.700 1883.355 4356.660 ;
        RECT 1884.335 4355.700 1885.960 4356.660 ;
        RECT 1886.940 4355.700 2093.460 4356.660 ;
        RECT 2096.630 4355.700 2152.935 4356.660 ;
        RECT 2153.915 4355.700 2153.990 4356.660 ;
        RECT 2154.970 4355.700 2156.500 4356.660 ;
        RECT 2158.190 4355.700 2158.355 4356.660 ;
        RECT 2159.335 4355.700 2160.960 4356.660 ;
        RECT 2161.940 4355.700 2368.460 4356.660 ;
        RECT 2371.630 4355.700 2427.935 4356.660 ;
        RECT 2428.915 4355.700 2428.990 4356.660 ;
        RECT 2429.970 4355.700 2431.500 4356.660 ;
        RECT 2433.190 4355.700 2433.355 4356.660 ;
        RECT 2434.335 4355.700 2435.960 4356.660 ;
        RECT 2436.940 4355.700 2918.460 4356.660 ;
        RECT 2921.630 4355.700 2977.935 4356.660 ;
        RECT 2978.915 4355.700 2978.990 4356.660 ;
        RECT 2979.970 4355.700 2981.500 4356.660 ;
        RECT 2983.190 4355.700 2983.355 4356.660 ;
        RECT 2984.335 4355.700 2985.960 4356.660 ;
        RECT 2986.940 4355.700 3169.460 4356.660 ;
        RECT 1.260 4246.540 3169.460 4355.700 ;
        RECT 1.260 4245.560 3160.700 4246.540 ;
        RECT 1.260 4244.830 3163.200 4245.560 ;
        RECT 1.260 4244.100 3165.700 4244.830 ;
        RECT 1.260 4243.370 3168.200 4244.100 ;
        RECT 1.260 4241.940 3169.460 4243.370 ;
        RECT 1.800 4240.960 3169.460 4241.940 ;
        RECT 1.260 4239.335 3169.460 4240.960 ;
        RECT 4.300 4238.355 3169.460 4239.335 ;
        RECT 1.260 4238.190 3169.460 4238.355 ;
        RECT 6.800 4237.480 3169.460 4238.190 ;
        RECT 9.300 4236.500 3169.460 4237.480 ;
        RECT 1.260 4234.970 3169.460 4236.500 ;
        RECT 11.800 4233.990 3169.460 4234.970 ;
        RECT 1.260 4233.915 3169.460 4233.990 ;
        RECT 14.300 4232.935 3169.460 4233.915 ;
        RECT 1.260 4187.065 3169.460 4232.935 ;
        RECT 1.260 4186.085 3155.700 4187.065 ;
        RECT 1.260 4186.010 3169.460 4186.085 ;
        RECT 1.260 4185.030 3158.200 4186.010 ;
        RECT 1.260 4183.500 3169.460 4185.030 ;
        RECT 1.260 4182.520 3160.700 4183.500 ;
        RECT 1.260 4181.810 3163.200 4182.520 ;
        RECT 1.260 4181.645 3169.460 4181.810 ;
        RECT 1.260 4180.665 3165.700 4181.645 ;
        RECT 1.260 4179.040 3169.460 4180.665 ;
        RECT 1.260 4178.060 3168.200 4179.040 ;
        RECT 1.260 4176.630 3169.460 4178.060 ;
        RECT 1.800 4175.900 3169.460 4176.630 ;
        RECT 4.300 4175.170 3169.460 4175.900 ;
        RECT 6.800 4174.440 3169.460 4175.170 ;
        RECT 9.300 4173.460 3169.460 4174.440 ;
        RECT 1.260 3816.540 3169.460 4173.460 ;
        RECT 1.260 3815.560 3160.700 3816.540 ;
        RECT 1.260 3814.830 3163.200 3815.560 ;
        RECT 1.260 3814.100 3165.700 3814.830 ;
        RECT 1.260 3813.370 3168.200 3814.100 ;
        RECT 1.260 3757.065 3169.460 3813.370 ;
        RECT 1.260 3756.085 3155.700 3757.065 ;
        RECT 1.260 3756.010 3169.460 3756.085 ;
        RECT 1.260 3755.030 3158.200 3756.010 ;
        RECT 1.260 3753.500 3169.460 3755.030 ;
        RECT 1.260 3752.520 3160.700 3753.500 ;
        RECT 1.260 3751.810 3163.200 3752.520 ;
        RECT 1.260 3751.645 3169.460 3751.810 ;
        RECT 1.260 3750.665 3165.700 3751.645 ;
        RECT 1.260 3749.040 3169.460 3750.665 ;
        RECT 1.260 3748.060 3168.200 3749.040 ;
        RECT 1.260 3421.940 3169.460 3748.060 ;
        RECT 1.800 3420.960 3169.460 3421.940 ;
        RECT 1.260 3419.335 3169.460 3420.960 ;
        RECT 4.300 3418.355 3169.460 3419.335 ;
        RECT 1.260 3418.190 3169.460 3418.355 ;
        RECT 6.800 3417.480 3169.460 3418.190 ;
        RECT 9.300 3416.500 3169.460 3417.480 ;
        RECT 1.260 3414.970 3169.460 3416.500 ;
        RECT 11.800 3413.990 3169.460 3414.970 ;
        RECT 1.260 3413.915 3169.460 3413.990 ;
        RECT 14.300 3412.935 3169.460 3413.915 ;
        RECT 1.260 3386.540 3169.460 3412.935 ;
        RECT 1.260 3385.560 3160.700 3386.540 ;
        RECT 1.260 3384.830 3163.200 3385.560 ;
        RECT 1.260 3384.100 3165.700 3384.830 ;
        RECT 1.260 3383.370 3168.200 3384.100 ;
        RECT 1.260 3356.630 3169.460 3383.370 ;
        RECT 1.800 3355.900 3169.460 3356.630 ;
        RECT 4.300 3355.170 3169.460 3355.900 ;
        RECT 6.800 3354.440 3169.460 3355.170 ;
        RECT 9.300 3353.460 3169.460 3354.440 ;
        RECT 1.260 3327.065 3169.460 3353.460 ;
        RECT 1.260 3326.085 3155.700 3327.065 ;
        RECT 1.260 3326.010 3169.460 3326.085 ;
        RECT 1.260 3325.030 3158.200 3326.010 ;
        RECT 1.260 3323.500 3169.460 3325.030 ;
        RECT 1.260 3322.520 3160.700 3323.500 ;
        RECT 1.260 3321.810 3163.200 3322.520 ;
        RECT 1.260 3321.645 3169.460 3321.810 ;
        RECT 1.260 3320.665 3165.700 3321.645 ;
        RECT 1.260 3319.040 3169.460 3320.665 ;
        RECT 1.260 3318.060 3168.200 3319.040 ;
        RECT 1.260 3216.940 3169.460 3318.060 ;
        RECT 1.800 3215.960 3169.460 3216.940 ;
        RECT 1.260 3214.335 3169.460 3215.960 ;
        RECT 4.300 3213.355 3169.460 3214.335 ;
        RECT 1.260 3213.190 3169.460 3213.355 ;
        RECT 6.800 3212.480 3169.460 3213.190 ;
        RECT 9.300 3211.500 3169.460 3212.480 ;
        RECT 1.260 3209.970 3169.460 3211.500 ;
        RECT 11.800 3208.990 3169.460 3209.970 ;
        RECT 1.260 3208.915 3169.460 3208.990 ;
        RECT 14.300 3207.935 3169.460 3208.915 ;
        RECT 1.260 3171.540 3169.460 3207.935 ;
        RECT 1.260 3170.560 3160.700 3171.540 ;
        RECT 1.260 3169.830 3163.200 3170.560 ;
        RECT 1.260 3169.100 3165.700 3169.830 ;
        RECT 1.260 3168.370 3168.200 3169.100 ;
        RECT 1.260 3151.630 3169.460 3168.370 ;
        RECT 1.800 3150.900 3169.460 3151.630 ;
        RECT 4.300 3150.170 3169.460 3150.900 ;
        RECT 6.800 3149.440 3169.460 3150.170 ;
        RECT 9.300 3148.460 3169.460 3149.440 ;
        RECT 1.260 3112.065 3169.460 3148.460 ;
        RECT 1.260 3111.085 3155.700 3112.065 ;
        RECT 1.260 3111.010 3169.460 3111.085 ;
        RECT 1.260 3110.030 3158.200 3111.010 ;
        RECT 1.260 3108.500 3169.460 3110.030 ;
        RECT 1.260 3107.520 3160.700 3108.500 ;
        RECT 1.260 3106.810 3163.200 3107.520 ;
        RECT 1.260 3106.645 3169.460 3106.810 ;
        RECT 1.260 3105.665 3165.700 3106.645 ;
        RECT 1.260 3104.040 3169.460 3105.665 ;
        RECT 1.260 3103.060 3168.200 3104.040 ;
        RECT 1.260 3011.940 3169.460 3103.060 ;
        RECT 1.800 3010.960 3169.460 3011.940 ;
        RECT 1.260 3009.335 3169.460 3010.960 ;
        RECT 4.300 3008.355 3169.460 3009.335 ;
        RECT 1.260 3008.190 3169.460 3008.355 ;
        RECT 6.800 3007.480 3169.460 3008.190 ;
        RECT 9.300 3006.500 3169.460 3007.480 ;
        RECT 1.260 3004.970 3169.460 3006.500 ;
        RECT 11.800 3003.990 3169.460 3004.970 ;
        RECT 1.260 3003.915 3169.460 3003.990 ;
        RECT 14.300 3002.935 3169.460 3003.915 ;
        RECT 1.260 2956.540 3169.460 3002.935 ;
        RECT 1.260 2955.560 3160.700 2956.540 ;
        RECT 1.260 2954.830 3163.200 2955.560 ;
        RECT 1.260 2954.100 3165.700 2954.830 ;
        RECT 1.260 2953.370 3168.200 2954.100 ;
        RECT 1.260 2946.630 3169.460 2953.370 ;
        RECT 1.800 2945.900 3169.460 2946.630 ;
        RECT 4.300 2945.170 3169.460 2945.900 ;
        RECT 6.800 2944.440 3169.460 2945.170 ;
        RECT 9.300 2943.460 3169.460 2944.440 ;
        RECT 1.260 2897.065 3169.460 2943.460 ;
        RECT 1.260 2896.085 3155.700 2897.065 ;
        RECT 1.260 2896.010 3169.460 2896.085 ;
        RECT 1.260 2895.030 3158.200 2896.010 ;
        RECT 1.260 2893.500 3169.460 2895.030 ;
        RECT 1.260 2892.520 3160.700 2893.500 ;
        RECT 1.260 2891.810 3163.200 2892.520 ;
        RECT 1.260 2891.645 3169.460 2891.810 ;
        RECT 1.260 2890.665 3165.700 2891.645 ;
        RECT 1.260 2889.040 3169.460 2890.665 ;
        RECT 1.260 2888.060 3168.200 2889.040 ;
        RECT 1.260 2806.940 3169.460 2888.060 ;
        RECT 1.800 2805.960 3169.460 2806.940 ;
        RECT 1.260 2804.335 3169.460 2805.960 ;
        RECT 4.300 2803.355 3169.460 2804.335 ;
        RECT 1.260 2803.190 3169.460 2803.355 ;
        RECT 6.800 2802.480 3169.460 2803.190 ;
        RECT 9.300 2801.500 3169.460 2802.480 ;
        RECT 1.260 2799.970 3169.460 2801.500 ;
        RECT 11.800 2798.990 3169.460 2799.970 ;
        RECT 1.260 2798.915 3169.460 2798.990 ;
        RECT 14.300 2797.935 3169.460 2798.915 ;
        RECT 1.260 2741.630 3169.460 2797.935 ;
        RECT 1.800 2741.540 3169.460 2741.630 ;
        RECT 1.800 2740.900 3160.700 2741.540 ;
        RECT 4.300 2740.560 3160.700 2740.900 ;
        RECT 4.300 2740.170 3163.200 2740.560 ;
        RECT 6.800 2739.830 3163.200 2740.170 ;
        RECT 6.800 2739.440 3165.700 2739.830 ;
        RECT 9.300 2739.100 3165.700 2739.440 ;
        RECT 9.300 2738.460 3168.200 2739.100 ;
        RECT 1.260 2738.370 3168.200 2738.460 ;
        RECT 1.260 2682.065 3169.460 2738.370 ;
        RECT 1.260 2681.085 3155.700 2682.065 ;
        RECT 1.260 2681.010 3169.460 2681.085 ;
        RECT 1.260 2680.030 3158.200 2681.010 ;
        RECT 1.260 2678.500 3169.460 2680.030 ;
        RECT 1.260 2677.520 3160.700 2678.500 ;
        RECT 1.260 2676.810 3163.200 2677.520 ;
        RECT 1.260 2676.645 3169.460 2676.810 ;
        RECT 1.260 2675.665 3165.700 2676.645 ;
        RECT 1.260 2674.040 3169.460 2675.665 ;
        RECT 1.260 2673.060 3168.200 2674.040 ;
        RECT 1.260 2601.940 3169.460 2673.060 ;
        RECT 1.800 2600.960 3169.460 2601.940 ;
        RECT 1.260 2599.335 3169.460 2600.960 ;
        RECT 4.300 2598.355 3169.460 2599.335 ;
        RECT 1.260 2598.190 3169.460 2598.355 ;
        RECT 6.800 2597.480 3169.460 2598.190 ;
        RECT 9.300 2596.500 3169.460 2597.480 ;
        RECT 1.260 2594.970 3169.460 2596.500 ;
        RECT 11.800 2593.990 3169.460 2594.970 ;
        RECT 1.260 2593.915 3169.460 2593.990 ;
        RECT 14.300 2592.935 3169.460 2593.915 ;
        RECT 1.260 2536.630 3169.460 2592.935 ;
        RECT 1.800 2535.900 3169.460 2536.630 ;
        RECT 4.300 2535.170 3169.460 2535.900 ;
        RECT 6.800 2534.440 3169.460 2535.170 ;
        RECT 9.300 2533.460 3169.460 2534.440 ;
        RECT 1.260 2526.540 3169.460 2533.460 ;
        RECT 1.260 2525.560 3160.700 2526.540 ;
        RECT 1.260 2524.830 3163.200 2525.560 ;
        RECT 1.260 2524.100 3165.700 2524.830 ;
        RECT 1.260 2523.370 3168.200 2524.100 ;
        RECT 1.260 2467.065 3169.460 2523.370 ;
        RECT 1.260 2466.085 3155.700 2467.065 ;
        RECT 1.260 2466.010 3169.460 2466.085 ;
        RECT 1.260 2465.030 3158.200 2466.010 ;
        RECT 1.260 2463.500 3169.460 2465.030 ;
        RECT 1.260 2462.520 3160.700 2463.500 ;
        RECT 1.260 2461.810 3163.200 2462.520 ;
        RECT 1.260 2461.645 3169.460 2461.810 ;
        RECT 1.260 2460.665 3165.700 2461.645 ;
        RECT 1.260 2459.040 3169.460 2460.665 ;
        RECT 1.260 2458.060 3168.200 2459.040 ;
        RECT 1.260 2396.940 3169.460 2458.060 ;
        RECT 1.800 2395.960 3169.460 2396.940 ;
        RECT 1.260 2394.335 3169.460 2395.960 ;
        RECT 4.300 2393.355 3169.460 2394.335 ;
        RECT 1.260 2393.190 3169.460 2393.355 ;
        RECT 6.800 2392.480 3169.460 2393.190 ;
        RECT 9.300 2391.500 3169.460 2392.480 ;
        RECT 1.260 2389.970 3169.460 2391.500 ;
        RECT 11.800 2388.990 3169.460 2389.970 ;
        RECT 1.260 2388.915 3169.460 2388.990 ;
        RECT 14.300 2387.935 3169.460 2388.915 ;
        RECT 1.260 2331.630 3169.460 2387.935 ;
        RECT 1.800 2330.900 3169.460 2331.630 ;
        RECT 4.300 2330.170 3169.460 2330.900 ;
        RECT 6.800 2329.440 3169.460 2330.170 ;
        RECT 9.300 2328.460 3169.460 2329.440 ;
        RECT 1.260 2311.540 3169.460 2328.460 ;
        RECT 1.260 2310.560 3160.700 2311.540 ;
        RECT 1.260 2309.830 3163.200 2310.560 ;
        RECT 1.260 2309.100 3165.700 2309.830 ;
        RECT 1.260 2308.370 3168.200 2309.100 ;
        RECT 1.260 2252.065 3169.460 2308.370 ;
        RECT 1.260 2251.085 3155.700 2252.065 ;
        RECT 1.260 2251.010 3169.460 2251.085 ;
        RECT 1.260 2250.030 3158.200 2251.010 ;
        RECT 1.260 2248.500 3169.460 2250.030 ;
        RECT 1.260 2247.520 3160.700 2248.500 ;
        RECT 1.260 2246.810 3163.200 2247.520 ;
        RECT 1.260 2246.645 3169.460 2246.810 ;
        RECT 1.260 2245.665 3165.700 2246.645 ;
        RECT 1.260 2244.040 3169.460 2245.665 ;
        RECT 1.260 2243.060 3168.200 2244.040 ;
        RECT 1.260 2191.940 3169.460 2243.060 ;
        RECT 1.800 2190.960 3169.460 2191.940 ;
        RECT 1.260 2189.335 3169.460 2190.960 ;
        RECT 4.300 2188.355 3169.460 2189.335 ;
        RECT 1.260 2188.190 3169.460 2188.355 ;
        RECT 6.800 2187.480 3169.460 2188.190 ;
        RECT 9.300 2186.500 3169.460 2187.480 ;
        RECT 1.260 2184.970 3169.460 2186.500 ;
        RECT 11.800 2183.990 3169.460 2184.970 ;
        RECT 1.260 2183.915 3169.460 2183.990 ;
        RECT 14.300 2182.935 3169.460 2183.915 ;
        RECT 1.260 2126.630 3169.460 2182.935 ;
        RECT 1.800 2125.900 3169.460 2126.630 ;
        RECT 4.300 2125.170 3169.460 2125.900 ;
        RECT 6.800 2124.440 3169.460 2125.170 ;
        RECT 9.300 2123.460 3169.460 2124.440 ;
        RECT 1.260 1576.940 3169.460 2123.460 ;
        RECT 1.800 1575.960 3169.460 1576.940 ;
        RECT 1.260 1574.335 3169.460 1575.960 ;
        RECT 4.300 1573.355 3169.460 1574.335 ;
        RECT 1.260 1573.190 3169.460 1573.355 ;
        RECT 6.800 1572.480 3169.460 1573.190 ;
        RECT 9.300 1571.500 3169.460 1572.480 ;
        RECT 1.260 1569.970 3169.460 1571.500 ;
        RECT 11.800 1568.990 3169.460 1569.970 ;
        RECT 1.260 1568.915 3169.460 1568.990 ;
        RECT 14.300 1567.935 3169.460 1568.915 ;
        RECT 1.260 1511.630 3169.460 1567.935 ;
        RECT 1.800 1510.900 3169.460 1511.630 ;
        RECT 4.300 1510.170 3169.460 1510.900 ;
        RECT 6.800 1509.440 3169.460 1510.170 ;
        RECT 9.300 1508.460 3169.460 1509.440 ;
        RECT 1.260 1451.540 3169.460 1508.460 ;
        RECT 1.260 1450.560 3160.700 1451.540 ;
        RECT 1.260 1449.830 3163.200 1450.560 ;
        RECT 1.260 1449.100 3165.700 1449.830 ;
        RECT 1.260 1448.370 3168.200 1449.100 ;
        RECT 1.260 1392.065 3169.460 1448.370 ;
        RECT 1.260 1391.085 3155.700 1392.065 ;
        RECT 1.260 1391.010 3169.460 1391.085 ;
        RECT 1.260 1390.030 3158.200 1391.010 ;
        RECT 1.260 1388.500 3169.460 1390.030 ;
        RECT 1.260 1387.520 3160.700 1388.500 ;
        RECT 1.260 1386.810 3163.200 1387.520 ;
        RECT 1.260 1386.645 3169.460 1386.810 ;
        RECT 1.260 1385.665 3165.700 1386.645 ;
        RECT 1.260 1384.040 3169.460 1385.665 ;
        RECT 1.260 1383.060 3168.200 1384.040 ;
        RECT 1.260 1371.940 3169.460 1383.060 ;
        RECT 1.800 1370.960 3169.460 1371.940 ;
        RECT 1.260 1369.335 3169.460 1370.960 ;
        RECT 4.300 1368.355 3169.460 1369.335 ;
        RECT 1.260 1368.190 3169.460 1368.355 ;
        RECT 6.800 1367.480 3169.460 1368.190 ;
        RECT 9.300 1366.500 3169.460 1367.480 ;
        RECT 1.260 1364.970 3169.460 1366.500 ;
        RECT 11.800 1363.990 3169.460 1364.970 ;
        RECT 1.260 1363.915 3169.460 1363.990 ;
        RECT 14.300 1362.935 3169.460 1363.915 ;
        RECT 1.260 1306.630 3169.460 1362.935 ;
        RECT 1.800 1305.900 3169.460 1306.630 ;
        RECT 4.300 1305.170 3169.460 1305.900 ;
        RECT 6.800 1304.440 3169.460 1305.170 ;
        RECT 9.300 1303.460 3169.460 1304.440 ;
        RECT 1.260 1236.540 3169.460 1303.460 ;
        RECT 1.260 1235.560 3160.700 1236.540 ;
        RECT 1.260 1234.830 3163.200 1235.560 ;
        RECT 1.260 1234.100 3165.700 1234.830 ;
        RECT 1.260 1233.370 3168.200 1234.100 ;
        RECT 1.260 1177.065 3169.460 1233.370 ;
        RECT 1.260 1176.085 3155.700 1177.065 ;
        RECT 1.260 1176.010 3169.460 1176.085 ;
        RECT 1.260 1175.030 3158.200 1176.010 ;
        RECT 1.260 1173.500 3169.460 1175.030 ;
        RECT 1.260 1172.520 3160.700 1173.500 ;
        RECT 1.260 1171.810 3163.200 1172.520 ;
        RECT 1.260 1171.645 3169.460 1171.810 ;
        RECT 1.260 1170.665 3165.700 1171.645 ;
        RECT 1.260 1169.040 3169.460 1170.665 ;
        RECT 1.260 1168.060 3168.200 1169.040 ;
        RECT 1.260 1166.940 3169.460 1168.060 ;
        RECT 1.800 1165.960 3169.460 1166.940 ;
        RECT 1.260 1164.335 3169.460 1165.960 ;
        RECT 4.300 1163.355 3169.460 1164.335 ;
        RECT 1.260 1163.190 3169.460 1163.355 ;
        RECT 6.800 1162.480 3169.460 1163.190 ;
        RECT 9.300 1161.500 3169.460 1162.480 ;
        RECT 1.260 1159.970 3169.460 1161.500 ;
        RECT 11.800 1158.990 3169.460 1159.970 ;
        RECT 1.260 1158.915 3169.460 1158.990 ;
        RECT 14.300 1157.935 3169.460 1158.915 ;
        RECT 1.260 1101.630 3169.460 1157.935 ;
        RECT 1.800 1100.900 3169.460 1101.630 ;
        RECT 4.300 1100.170 3169.460 1100.900 ;
        RECT 6.800 1099.440 3169.460 1100.170 ;
        RECT 9.300 1098.460 3169.460 1099.440 ;
        RECT 1.260 1021.540 3169.460 1098.460 ;
        RECT 1.260 1020.560 3160.700 1021.540 ;
        RECT 1.260 1019.830 3163.200 1020.560 ;
        RECT 1.260 1019.100 3165.700 1019.830 ;
        RECT 1.260 1018.370 3168.200 1019.100 ;
        RECT 1.260 962.065 3169.460 1018.370 ;
        RECT 1.260 961.940 3155.700 962.065 ;
        RECT 1.800 961.085 3155.700 961.940 ;
        RECT 1.800 961.010 3169.460 961.085 ;
        RECT 1.800 960.960 3158.200 961.010 ;
        RECT 1.260 960.030 3158.200 960.960 ;
        RECT 1.260 959.335 3169.460 960.030 ;
        RECT 4.300 958.500 3169.460 959.335 ;
        RECT 4.300 958.355 3160.700 958.500 ;
        RECT 1.260 958.190 3160.700 958.355 ;
        RECT 6.800 957.520 3160.700 958.190 ;
        RECT 6.800 957.480 3163.200 957.520 ;
        RECT 9.300 956.810 3163.200 957.480 ;
        RECT 9.300 956.645 3169.460 956.810 ;
        RECT 9.300 956.500 3165.700 956.645 ;
        RECT 1.260 955.665 3165.700 956.500 ;
        RECT 1.260 954.970 3169.460 955.665 ;
        RECT 11.800 954.040 3169.460 954.970 ;
        RECT 11.800 953.990 3168.200 954.040 ;
        RECT 1.260 953.915 3168.200 953.990 ;
        RECT 14.300 953.060 3168.200 953.915 ;
        RECT 14.300 952.935 3169.460 953.060 ;
        RECT 1.260 896.630 3169.460 952.935 ;
        RECT 1.800 895.900 3169.460 896.630 ;
        RECT 4.300 895.170 3169.460 895.900 ;
        RECT 6.800 894.440 3169.460 895.170 ;
        RECT 9.300 893.460 3169.460 894.440 ;
        RECT 1.260 806.540 3169.460 893.460 ;
        RECT 1.260 805.560 3160.700 806.540 ;
        RECT 1.260 804.830 3163.200 805.560 ;
        RECT 1.260 804.100 3165.700 804.830 ;
        RECT 1.260 803.370 3168.200 804.100 ;
        RECT 1.260 756.940 3169.460 803.370 ;
        RECT 1.800 755.960 3169.460 756.940 ;
        RECT 1.260 754.335 3169.460 755.960 ;
        RECT 4.300 753.355 3169.460 754.335 ;
        RECT 1.260 753.190 3169.460 753.355 ;
        RECT 6.800 752.480 3169.460 753.190 ;
        RECT 9.300 751.500 3169.460 752.480 ;
        RECT 1.260 749.970 3169.460 751.500 ;
        RECT 11.800 748.990 3169.460 749.970 ;
        RECT 1.260 748.915 3169.460 748.990 ;
        RECT 14.300 747.935 3169.460 748.915 ;
        RECT 1.260 747.065 3169.460 747.935 ;
        RECT 1.260 746.085 3155.700 747.065 ;
        RECT 1.260 746.010 3169.460 746.085 ;
        RECT 1.260 745.030 3158.200 746.010 ;
        RECT 1.260 743.500 3169.460 745.030 ;
        RECT 1.260 742.520 3160.700 743.500 ;
        RECT 1.260 741.810 3163.200 742.520 ;
        RECT 1.260 741.645 3169.460 741.810 ;
        RECT 1.260 740.665 3165.700 741.645 ;
        RECT 1.260 739.040 3169.460 740.665 ;
        RECT 1.260 738.060 3168.200 739.040 ;
        RECT 1.260 691.630 3169.460 738.060 ;
        RECT 1.800 690.900 3169.460 691.630 ;
        RECT 4.300 690.170 3169.460 690.900 ;
        RECT 6.800 689.440 3169.460 690.170 ;
        RECT 9.300 688.460 3169.460 689.440 ;
        RECT 1.260 591.540 3169.460 688.460 ;
        RECT 1.260 590.560 3160.700 591.540 ;
        RECT 1.260 589.830 3163.200 590.560 ;
        RECT 1.260 589.100 3165.700 589.830 ;
        RECT 1.260 588.370 3168.200 589.100 ;
        RECT 1.260 551.940 3169.460 588.370 ;
        RECT 1.800 550.960 3169.460 551.940 ;
        RECT 1.260 549.335 3169.460 550.960 ;
        RECT 4.300 548.355 3169.460 549.335 ;
        RECT 1.260 548.190 3169.460 548.355 ;
        RECT 6.800 547.480 3169.460 548.190 ;
        RECT 9.300 546.500 3169.460 547.480 ;
        RECT 1.260 544.970 3169.460 546.500 ;
        RECT 11.800 543.990 3169.460 544.970 ;
        RECT 1.260 543.915 3169.460 543.990 ;
        RECT 14.300 542.935 3169.460 543.915 ;
        RECT 1.260 532.065 3169.460 542.935 ;
        RECT 1.260 531.085 3155.700 532.065 ;
        RECT 1.260 531.010 3169.460 531.085 ;
        RECT 1.260 530.030 3158.200 531.010 ;
        RECT 1.260 528.500 3169.460 530.030 ;
        RECT 1.260 527.520 3160.700 528.500 ;
        RECT 1.260 526.810 3163.200 527.520 ;
        RECT 1.260 526.645 3169.460 526.810 ;
        RECT 1.260 525.665 3165.700 526.645 ;
        RECT 1.260 524.040 3169.460 525.665 ;
        RECT 1.260 523.060 3168.200 524.040 ;
        RECT 1.260 486.630 3169.460 523.060 ;
        RECT 1.800 485.900 3169.460 486.630 ;
        RECT 4.300 485.170 3169.460 485.900 ;
        RECT 6.800 484.440 3169.460 485.170 ;
        RECT 9.300 483.460 3169.460 484.440 ;
        RECT 1.260 376.540 3169.460 483.460 ;
        RECT 1.260 375.560 3160.700 376.540 ;
        RECT 1.260 374.830 3163.200 375.560 ;
        RECT 1.260 374.100 3165.700 374.830 ;
        RECT 1.260 373.370 3168.200 374.100 ;
        RECT 1.260 317.065 3169.460 373.370 ;
        RECT 1.260 316.085 3155.700 317.065 ;
        RECT 1.260 316.010 3169.460 316.085 ;
        RECT 1.260 315.030 3158.200 316.010 ;
        RECT 1.260 313.500 3169.460 315.030 ;
        RECT 1.260 312.520 3160.700 313.500 ;
        RECT 1.260 311.810 3163.200 312.520 ;
        RECT 1.260 311.645 3169.460 311.810 ;
        RECT 1.260 310.665 3165.700 311.645 ;
        RECT 1.260 309.040 3169.460 310.665 ;
        RECT 1.260 308.060 3168.200 309.040 ;
        RECT 1.260 161.540 3169.460 308.060 ;
        RECT 1.260 160.560 3160.700 161.540 ;
        RECT 1.260 159.830 3163.200 160.560 ;
        RECT 1.260 159.100 3165.700 159.830 ;
        RECT 1.260 158.370 3168.200 159.100 ;
        RECT 1.260 102.065 3169.460 158.370 ;
        RECT 1.260 101.085 3155.700 102.065 ;
        RECT 1.260 101.010 3169.460 101.085 ;
        RECT 1.260 100.030 3158.200 101.010 ;
        RECT 1.260 98.500 3169.460 100.030 ;
        RECT 1.260 97.520 3160.700 98.500 ;
        RECT 1.260 96.810 3163.200 97.520 ;
        RECT 1.260 96.645 3169.460 96.810 ;
        RECT 1.260 95.665 3165.700 96.645 ;
        RECT 1.260 94.040 3169.460 95.665 ;
        RECT 1.260 93.060 3168.200 94.040 ;
        RECT 1.260 4.300 3169.460 93.060 ;
        RECT 1.260 3.500 450.665 4.300 ;
        RECT 451.645 3.500 455.030 4.300 ;
        RECT 456.010 3.500 515.560 4.300 ;
        RECT 516.540 3.500 725.665 4.300 ;
        RECT 726.645 3.500 790.560 4.300 ;
        RECT 791.540 3.500 1275.665 4.300 ;
        RECT 1276.645 3.500 1338.365 4.300 ;
        RECT 1340.810 3.500 1613.370 4.300 ;
        RECT 1615.810 3.500 1831.085 4.300 ;
        RECT 1832.065 3.500 1888.370 4.300 ;
        RECT 1891.535 3.500 2106.085 4.300 ;
        RECT 2107.065 3.500 2163.370 4.300 ;
        RECT 2166.540 3.500 2373.060 4.300 ;
        RECT 2374.040 3.500 2375.665 4.300 ;
        RECT 2376.645 3.500 2376.810 4.300 ;
        RECT 2378.500 3.500 2380.030 4.300 ;
        RECT 2381.010 3.500 2381.085 4.300 ;
        RECT 2382.065 3.500 2438.370 4.300 ;
        RECT 2441.540 3.500 3169.460 4.300 ;
      LAYER Metal3 ;
        RECT 1.210 5.740 3169.510 4354.980 ;
      LAYER Metal4 ;
        RECT 26.460 26.410 35.780 4329.270 ;
        RECT 39.380 26.410 44.780 4329.270 ;
        RECT 48.380 26.410 60.640 4329.270 ;
        RECT 64.240 26.410 69.640 4329.270 ;
        RECT 73.240 4274.780 105.780 4329.270 ;
        RECT 109.380 4274.780 127.780 4329.270 ;
        RECT 131.380 4274.780 185.780 4329.270 ;
        RECT 189.380 4274.780 207.780 4329.270 ;
        RECT 211.380 4274.780 265.780 4329.270 ;
        RECT 269.380 4274.780 287.780 4329.270 ;
        RECT 291.380 4274.780 306.280 4329.270 ;
        RECT 309.880 4274.780 313.280 4329.270 ;
        RECT 316.880 4274.780 345.780 4329.270 ;
        RECT 349.380 4274.780 367.780 4329.270 ;
        RECT 371.380 4274.780 425.780 4329.270 ;
        RECT 429.380 4274.780 447.780 4329.270 ;
        RECT 451.380 4274.780 505.780 4329.270 ;
        RECT 509.380 4274.780 527.780 4329.270 ;
        RECT 531.380 4274.780 555.980 4329.270 ;
        RECT 559.580 4274.780 562.980 4329.270 ;
        RECT 566.580 4274.780 585.780 4329.270 ;
        RECT 589.380 4274.780 607.780 4329.270 ;
        RECT 611.380 4274.780 665.780 4329.270 ;
        RECT 669.380 4274.780 687.780 4329.270 ;
        RECT 691.380 4274.780 745.780 4329.270 ;
        RECT 749.380 4274.780 767.780 4329.270 ;
        RECT 771.380 4274.780 825.780 4329.270 ;
        RECT 829.380 4274.780 847.780 4329.270 ;
        RECT 851.380 4274.780 864.480 4329.270 ;
        RECT 868.080 4274.780 871.480 4329.270 ;
        RECT 875.080 4274.780 905.780 4329.270 ;
        RECT 909.380 4274.780 927.780 4329.270 ;
        RECT 931.380 4274.780 985.780 4329.270 ;
        RECT 989.380 4274.780 1007.780 4329.270 ;
        RECT 1011.380 4274.780 1065.780 4329.270 ;
        RECT 1069.380 4274.780 1087.780 4329.270 ;
        RECT 1091.380 4274.780 1116.180 4329.270 ;
        RECT 1119.780 4274.780 1123.180 4329.270 ;
        RECT 1126.780 4274.780 1145.780 4329.270 ;
        RECT 1149.380 4274.780 1167.780 4329.270 ;
        RECT 1171.380 4274.780 1225.780 4329.270 ;
        RECT 1229.380 4274.780 1247.780 4329.270 ;
        RECT 1251.380 4274.780 1305.780 4329.270 ;
        RECT 1309.380 4274.780 1327.780 4329.270 ;
        RECT 1331.380 4274.780 1359.080 4329.270 ;
        RECT 1362.680 4274.780 1366.080 4329.270 ;
        RECT 1369.680 4274.780 1385.780 4329.270 ;
        RECT 1389.380 4274.780 1407.780 4329.270 ;
        RECT 1411.380 4274.780 1465.780 4329.270 ;
        RECT 1469.380 4274.780 1487.780 4329.270 ;
        RECT 1491.380 4274.780 1545.780 4329.270 ;
        RECT 1549.380 4274.780 1567.780 4329.270 ;
        RECT 1571.380 4274.780 1625.780 4329.270 ;
        RECT 1629.380 4274.780 1647.780 4329.270 ;
        RECT 1651.380 4274.780 1705.780 4329.270 ;
        RECT 1709.380 4274.780 1727.780 4329.270 ;
        RECT 1731.380 4274.780 1785.780 4329.270 ;
        RECT 1789.380 4274.780 1807.780 4329.270 ;
        RECT 1811.380 4274.780 1865.780 4329.270 ;
        RECT 1869.380 4274.780 1887.780 4329.270 ;
        RECT 1891.380 4274.780 1916.080 4329.270 ;
        RECT 1919.680 4274.780 1923.080 4329.270 ;
        RECT 1926.680 4274.780 1945.780 4329.270 ;
        RECT 1949.380 4274.780 1967.780 4329.270 ;
        RECT 1971.380 4274.780 2025.780 4329.270 ;
        RECT 2029.380 4274.780 2047.780 4329.270 ;
        RECT 2051.380 4274.780 2105.780 4329.270 ;
        RECT 2109.380 4274.780 2127.780 4329.270 ;
        RECT 2131.380 4274.780 2162.780 4329.270 ;
        RECT 2166.380 4274.780 2169.780 4329.270 ;
        RECT 2173.380 4274.780 2185.780 4329.270 ;
        RECT 2189.380 4274.780 2207.780 4329.270 ;
        RECT 2211.380 4274.780 2265.780 4329.270 ;
        RECT 2269.380 4274.780 2287.780 4329.270 ;
        RECT 2291.380 4274.780 2330.780 4329.270 ;
        RECT 2334.380 4274.780 2345.780 4329.270 ;
        RECT 2349.380 4274.780 2352.780 4329.270 ;
        RECT 2356.380 4274.780 2367.780 4329.270 ;
        RECT 2371.380 4274.780 2425.780 4329.270 ;
        RECT 2429.380 4274.780 2447.780 4329.270 ;
        RECT 2451.380 4274.780 2505.780 4329.270 ;
        RECT 2509.380 4274.780 2527.780 4329.270 ;
        RECT 2531.380 4274.780 2585.780 4329.270 ;
        RECT 2589.380 4274.780 2607.780 4329.270 ;
        RECT 2611.380 4274.780 2665.780 4329.270 ;
        RECT 2669.380 4274.780 2687.780 4329.270 ;
        RECT 2691.380 4274.780 2745.780 4329.270 ;
        RECT 2749.380 4274.780 2767.780 4329.270 ;
        RECT 2771.380 4274.780 2825.780 4329.270 ;
        RECT 2829.380 4274.780 2847.780 4329.270 ;
        RECT 2851.380 4274.780 2880.280 4329.270 ;
        RECT 2883.880 4274.780 2892.280 4329.270 ;
        RECT 2895.880 4274.780 2905.780 4329.270 ;
        RECT 2909.380 4274.780 2927.780 4329.270 ;
        RECT 2931.380 4274.780 2985.780 4329.270 ;
        RECT 2989.380 4274.780 3007.780 4329.270 ;
        RECT 3011.380 4274.780 3098.780 4329.270 ;
        RECT 73.240 1260.620 3098.780 4274.780 ;
        RECT 73.240 26.410 105.780 1260.620 ;
        RECT 109.380 545.220 127.780 1260.620 ;
        RECT 131.380 545.220 185.780 1260.620 ;
        RECT 109.380 66.700 185.780 545.220 ;
        RECT 109.380 26.410 127.780 66.700 ;
        RECT 131.380 26.410 185.780 66.700 ;
        RECT 189.380 26.410 207.780 1260.620 ;
        RECT 211.380 26.410 265.780 1260.620 ;
        RECT 269.380 26.410 287.780 1260.620 ;
        RECT 291.380 26.410 306.280 1260.620 ;
        RECT 309.880 26.410 313.280 1260.620 ;
        RECT 316.880 26.410 345.780 1260.620 ;
        RECT 349.380 26.410 367.780 1260.620 ;
        RECT 371.380 26.410 425.780 1260.620 ;
        RECT 429.380 26.410 447.780 1260.620 ;
        RECT 451.380 26.410 505.780 1260.620 ;
        RECT 509.380 26.410 527.780 1260.620 ;
        RECT 531.380 26.410 555.980 1260.620 ;
        RECT 559.580 545.220 562.980 1260.620 ;
        RECT 566.580 545.220 585.780 1260.620 ;
        RECT 559.580 66.700 585.780 545.220 ;
        RECT 559.580 26.410 562.980 66.700 ;
        RECT 566.580 26.410 585.780 66.700 ;
        RECT 589.380 26.410 607.780 1260.620 ;
        RECT 611.380 26.410 665.780 1260.620 ;
        RECT 669.380 26.410 687.780 1260.620 ;
        RECT 691.380 26.410 745.780 1260.620 ;
        RECT 749.380 26.410 767.780 1260.620 ;
        RECT 771.380 26.410 825.780 1260.620 ;
        RECT 829.380 26.410 847.780 1260.620 ;
        RECT 851.380 26.410 864.480 1260.620 ;
        RECT 868.080 26.410 871.480 1260.620 ;
        RECT 875.080 26.410 905.780 1260.620 ;
        RECT 909.380 26.410 927.780 1260.620 ;
        RECT 931.380 545.220 985.780 1260.620 ;
        RECT 989.380 545.220 1007.780 1260.620 ;
        RECT 931.380 66.700 1007.780 545.220 ;
        RECT 931.380 26.410 985.780 66.700 ;
        RECT 989.380 26.410 1007.780 66.700 ;
        RECT 1011.380 26.410 1065.780 1260.620 ;
        RECT 1069.380 26.410 1087.780 1260.620 ;
        RECT 1091.380 967.080 1116.180 1260.620 ;
        RECT 1119.780 967.080 1123.180 1260.620 ;
        RECT 1091.380 899.560 1123.180 967.080 ;
        RECT 1091.380 26.410 1116.180 899.560 ;
        RECT 1119.780 26.410 1123.180 899.560 ;
        RECT 1126.780 26.410 1145.780 1260.620 ;
        RECT 1149.380 26.410 1167.780 1260.620 ;
        RECT 1171.380 26.410 1225.780 1260.620 ;
        RECT 1229.380 26.410 1247.780 1260.620 ;
        RECT 1251.380 26.410 1305.780 1260.620 ;
        RECT 1309.380 26.410 1327.780 1260.620 ;
        RECT 1331.380 26.410 1359.080 1260.620 ;
        RECT 1362.680 26.410 1366.080 1260.620 ;
        RECT 1369.680 26.410 1385.780 1260.620 ;
        RECT 1389.380 26.410 1407.780 1260.620 ;
        RECT 1411.380 26.410 1465.780 1260.620 ;
        RECT 1469.380 26.410 1487.780 1260.620 ;
        RECT 1491.380 26.410 1545.780 1260.620 ;
        RECT 1549.380 26.410 1567.780 1260.620 ;
        RECT 1571.380 26.410 1625.780 1260.620 ;
        RECT 1629.380 26.410 1647.780 1260.620 ;
        RECT 1651.380 26.410 1705.780 1260.620 ;
        RECT 1709.380 26.410 1727.780 1260.620 ;
        RECT 1731.380 26.410 1785.780 1260.620 ;
        RECT 1789.380 26.410 1807.780 1260.620 ;
        RECT 1811.380 26.410 1865.780 1260.620 ;
        RECT 1869.380 26.410 1887.780 1260.620 ;
        RECT 1891.380 26.410 1916.080 1260.620 ;
        RECT 1919.680 26.410 1923.080 1260.620 ;
        RECT 1926.680 26.410 1945.780 1260.620 ;
        RECT 1949.380 26.410 1967.780 1260.620 ;
        RECT 1971.380 26.410 2025.780 1260.620 ;
        RECT 2029.380 26.410 2047.780 1260.620 ;
        RECT 2051.380 26.410 2105.780 1260.620 ;
        RECT 2109.380 26.410 2127.780 1260.620 ;
        RECT 2131.380 26.410 2162.780 1260.620 ;
        RECT 2166.380 26.410 2169.780 1260.620 ;
        RECT 2173.380 26.410 2185.780 1260.620 ;
        RECT 2189.380 26.410 2207.780 1260.620 ;
        RECT 2211.380 26.410 2265.780 1260.620 ;
        RECT 2269.380 26.410 2287.780 1260.620 ;
        RECT 2291.380 26.410 2330.780 1260.620 ;
        RECT 2334.380 26.410 2345.780 1260.620 ;
        RECT 2349.380 26.410 2352.780 1260.620 ;
        RECT 2356.380 26.410 2367.780 1260.620 ;
        RECT 2371.380 998.980 2425.780 1260.620 ;
        RECT 2429.380 998.980 2447.780 1260.620 ;
        RECT 2451.380 998.980 2505.780 1260.620 ;
        RECT 2509.380 998.980 2527.780 1260.620 ;
        RECT 2531.380 998.980 2585.780 1260.620 ;
        RECT 2589.380 998.980 2607.780 1260.620 ;
        RECT 2611.380 998.980 2665.780 1260.620 ;
        RECT 2669.380 998.980 2687.780 1260.620 ;
        RECT 2691.380 998.980 2745.780 1260.620 ;
        RECT 2749.380 998.980 2767.780 1260.620 ;
        RECT 2771.380 998.980 2825.780 1260.620 ;
        RECT 2829.380 998.980 2847.780 1260.620 ;
        RECT 2851.380 998.980 2880.280 1260.620 ;
        RECT 2883.880 998.980 2892.280 1260.620 ;
        RECT 2895.880 998.980 2905.780 1260.620 ;
        RECT 2909.380 998.980 2927.780 1260.620 ;
        RECT 2931.380 998.980 2985.780 1260.620 ;
        RECT 2989.380 998.980 3007.780 1260.620 ;
        RECT 3011.380 998.980 3098.780 1260.620 ;
        RECT 2371.380 203.020 3098.780 998.980 ;
        RECT 2371.380 26.410 2425.780 203.020 ;
        RECT 2429.380 26.410 2447.780 203.020 ;
        RECT 2451.380 26.410 2505.780 203.020 ;
        RECT 2509.380 26.410 2527.780 203.020 ;
        RECT 2531.380 26.410 2585.780 203.020 ;
        RECT 2589.380 26.410 2607.780 203.020 ;
        RECT 2611.380 26.410 2665.780 203.020 ;
        RECT 2669.380 26.410 2687.780 203.020 ;
        RECT 2691.380 26.410 2745.780 203.020 ;
        RECT 2749.380 26.410 2767.780 203.020 ;
        RECT 2771.380 26.410 2825.780 203.020 ;
        RECT 2829.380 26.410 2847.780 203.020 ;
        RECT 2851.380 26.410 2880.280 203.020 ;
        RECT 2883.880 26.410 2892.280 203.020 ;
        RECT 2895.880 144.425 2905.780 203.020 ;
        RECT 2909.380 144.425 2927.780 203.020 ;
        RECT 2931.380 144.425 2985.780 203.020 ;
        RECT 2895.880 87.030 2985.780 144.425 ;
        RECT 2895.880 26.410 2905.780 87.030 ;
        RECT 2909.380 26.410 2927.780 87.030 ;
        RECT 2931.380 26.410 2985.780 87.030 ;
        RECT 2989.380 26.410 3007.780 203.020 ;
        RECT 3011.380 26.410 3098.780 203.020 ;
        RECT 3102.380 26.410 3107.780 4329.270 ;
        RECT 3111.380 26.410 3126.320 4329.270 ;
        RECT 3129.920 26.410 3135.320 4329.270 ;
        RECT 3138.920 26.410 3144.660 4329.270 ;
        RECT 3155.260 26.410 3156.660 4329.270 ;
        RECT 3167.260 26.410 3167.780 4329.270 ;
      LAYER Metal5 ;
        RECT 84.995 4260.090 3167.860 4278.900 ;
        RECT 95.115 4256.090 3074.735 4260.090 ;
        RECT 3167.460 4256.090 3167.860 4260.090 ;
        RECT 84.995 4230.090 3167.860 4256.090 ;
        RECT 95.115 4226.090 3074.735 4230.090 ;
        RECT 3167.460 4226.090 3167.860 4230.090 ;
        RECT 84.995 4200.090 3167.860 4226.090 ;
        RECT 95.115 4196.090 3074.735 4200.090 ;
        RECT 3167.460 4196.090 3167.860 4200.090 ;
        RECT 84.995 4170.090 3167.860 4196.090 ;
        RECT 95.115 4166.090 3074.735 4170.090 ;
        RECT 3167.460 4166.090 3167.860 4170.090 ;
        RECT 84.995 4140.090 3167.860 4166.090 ;
        RECT 95.115 4136.090 3074.735 4140.090 ;
        RECT 3167.460 4136.090 3167.860 4140.090 ;
        RECT 84.995 4110.090 3167.860 4136.090 ;
        RECT 95.115 4106.090 3074.735 4110.090 ;
        RECT 3167.460 4106.090 3167.860 4110.090 ;
        RECT 84.995 4080.090 3167.860 4106.090 ;
        RECT 95.115 4076.090 3074.735 4080.090 ;
        RECT 3167.460 4076.090 3167.860 4080.090 ;
        RECT 84.995 4050.090 3167.860 4076.090 ;
        RECT 95.115 4046.090 3074.735 4050.090 ;
        RECT 3167.460 4046.090 3167.860 4050.090 ;
        RECT 84.995 4020.090 3167.860 4046.090 ;
        RECT 95.115 4016.090 3074.735 4020.090 ;
        RECT 3167.460 4016.090 3167.860 4020.090 ;
        RECT 84.995 3990.090 3167.860 4016.090 ;
        RECT 95.115 3986.090 3074.735 3990.090 ;
        RECT 3167.460 3986.090 3167.860 3990.090 ;
        RECT 84.995 3960.090 3167.860 3986.090 ;
        RECT 95.115 3956.090 3074.735 3960.090 ;
        RECT 3167.460 3956.090 3167.860 3960.090 ;
        RECT 84.995 3930.090 3167.860 3956.090 ;
        RECT 95.115 3926.090 3074.735 3930.090 ;
        RECT 3167.460 3926.090 3167.860 3930.090 ;
        RECT 84.995 3900.090 3167.860 3926.090 ;
        RECT 95.115 3896.090 3074.735 3900.090 ;
        RECT 3167.460 3896.090 3167.860 3900.090 ;
        RECT 84.995 3870.090 3167.860 3896.090 ;
        RECT 95.115 3866.090 3074.735 3870.090 ;
        RECT 3167.460 3866.090 3167.860 3870.090 ;
        RECT 84.995 3840.090 3167.860 3866.090 ;
        RECT 95.115 3836.090 3074.735 3840.090 ;
        RECT 3167.460 3836.090 3167.860 3840.090 ;
        RECT 84.995 3810.090 3167.860 3836.090 ;
        RECT 95.115 3806.090 3074.735 3810.090 ;
        RECT 3167.460 3806.090 3167.860 3810.090 ;
        RECT 84.995 3780.090 3167.860 3806.090 ;
        RECT 95.115 3776.090 3074.735 3780.090 ;
        RECT 3167.460 3776.090 3167.860 3780.090 ;
        RECT 84.995 3750.090 3167.860 3776.090 ;
        RECT 95.115 3746.090 3074.735 3750.090 ;
        RECT 3167.460 3746.090 3167.860 3750.090 ;
        RECT 84.995 3720.090 3167.860 3746.090 ;
        RECT 95.115 3716.090 3074.735 3720.090 ;
        RECT 3167.460 3716.090 3167.860 3720.090 ;
        RECT 84.995 3690.090 3167.860 3716.090 ;
        RECT 95.115 3686.090 3074.735 3690.090 ;
        RECT 3167.460 3686.090 3167.860 3690.090 ;
        RECT 84.995 3660.090 3167.860 3686.090 ;
        RECT 95.115 3656.090 3074.735 3660.090 ;
        RECT 3167.460 3656.090 3167.860 3660.090 ;
        RECT 84.995 3630.090 3167.860 3656.090 ;
        RECT 95.115 3626.090 3074.735 3630.090 ;
        RECT 3167.460 3626.090 3167.860 3630.090 ;
        RECT 84.995 3600.090 3167.860 3626.090 ;
        RECT 95.115 3596.090 3074.735 3600.090 ;
        RECT 3167.460 3596.090 3167.860 3600.090 ;
        RECT 84.995 3570.090 3167.860 3596.090 ;
        RECT 95.115 3566.090 3074.735 3570.090 ;
        RECT 3167.460 3566.090 3167.860 3570.090 ;
        RECT 84.995 3540.090 3167.860 3566.090 ;
        RECT 95.115 3536.090 3074.735 3540.090 ;
        RECT 3167.460 3536.090 3167.860 3540.090 ;
        RECT 84.995 3510.090 3167.860 3536.090 ;
        RECT 95.115 3506.090 3074.735 3510.090 ;
        RECT 3167.460 3506.090 3167.860 3510.090 ;
        RECT 84.995 3480.090 3167.860 3506.090 ;
        RECT 95.115 3476.090 3074.735 3480.090 ;
        RECT 3167.460 3476.090 3167.860 3480.090 ;
        RECT 84.995 3450.090 3167.860 3476.090 ;
        RECT 95.115 3446.090 3074.735 3450.090 ;
        RECT 3167.460 3446.090 3167.860 3450.090 ;
        RECT 84.995 3420.090 3167.860 3446.090 ;
        RECT 95.115 3416.090 3074.735 3420.090 ;
        RECT 3167.460 3416.090 3167.860 3420.090 ;
        RECT 84.995 3390.090 3167.860 3416.090 ;
        RECT 95.115 3386.090 3074.735 3390.090 ;
        RECT 3167.460 3386.090 3167.860 3390.090 ;
        RECT 84.995 3360.090 3167.860 3386.090 ;
        RECT 95.115 3356.090 3074.735 3360.090 ;
        RECT 3167.460 3356.090 3167.860 3360.090 ;
        RECT 84.995 3330.090 3167.860 3356.090 ;
        RECT 95.115 3326.090 3074.735 3330.090 ;
        RECT 3167.460 3326.090 3167.860 3330.090 ;
        RECT 84.995 3300.090 3167.860 3326.090 ;
        RECT 95.115 3296.090 3074.735 3300.090 ;
        RECT 3167.460 3296.090 3167.860 3300.090 ;
        RECT 84.995 3270.090 3167.860 3296.090 ;
        RECT 95.115 3266.090 3074.735 3270.090 ;
        RECT 3167.460 3266.090 3167.860 3270.090 ;
        RECT 84.995 3240.090 3167.860 3266.090 ;
        RECT 95.115 3236.090 3074.735 3240.090 ;
        RECT 3167.460 3236.090 3167.860 3240.090 ;
        RECT 84.995 3210.090 3167.860 3236.090 ;
        RECT 95.115 3206.090 3074.735 3210.090 ;
        RECT 3167.460 3206.090 3167.860 3210.090 ;
        RECT 84.995 3180.090 3167.860 3206.090 ;
        RECT 95.115 3176.090 3074.735 3180.090 ;
        RECT 3167.460 3176.090 3167.860 3180.090 ;
        RECT 84.995 3150.090 3167.860 3176.090 ;
        RECT 95.115 3146.090 3074.735 3150.090 ;
        RECT 3167.460 3146.090 3167.860 3150.090 ;
        RECT 84.995 3120.090 3167.860 3146.090 ;
        RECT 95.115 3116.090 3074.735 3120.090 ;
        RECT 3167.460 3116.090 3167.860 3120.090 ;
        RECT 84.995 3090.090 3167.860 3116.090 ;
        RECT 95.115 3086.090 3074.735 3090.090 ;
        RECT 3167.460 3086.090 3167.860 3090.090 ;
        RECT 84.995 3060.090 3167.860 3086.090 ;
        RECT 95.115 3056.090 3074.735 3060.090 ;
        RECT 3167.460 3056.090 3167.860 3060.090 ;
        RECT 84.995 3030.090 3167.860 3056.090 ;
        RECT 95.115 3026.090 3074.735 3030.090 ;
        RECT 3167.460 3026.090 3167.860 3030.090 ;
        RECT 84.995 3000.090 3167.860 3026.090 ;
        RECT 95.115 2996.090 3074.735 3000.090 ;
        RECT 3167.460 2996.090 3167.860 3000.090 ;
        RECT 84.995 2970.090 3167.860 2996.090 ;
        RECT 95.115 2966.090 3074.735 2970.090 ;
        RECT 3167.460 2966.090 3167.860 2970.090 ;
        RECT 84.995 2940.090 3167.860 2966.090 ;
        RECT 95.115 2936.090 3074.735 2940.090 ;
        RECT 3167.460 2936.090 3167.860 2940.090 ;
        RECT 84.995 2910.090 3167.860 2936.090 ;
        RECT 95.115 2906.090 3074.735 2910.090 ;
        RECT 3167.460 2906.090 3167.860 2910.090 ;
        RECT 84.995 2880.090 3167.860 2906.090 ;
        RECT 95.115 2876.090 3074.735 2880.090 ;
        RECT 3167.460 2876.090 3167.860 2880.090 ;
        RECT 84.995 2850.090 3167.860 2876.090 ;
        RECT 95.115 2846.090 3074.735 2850.090 ;
        RECT 3167.460 2846.090 3167.860 2850.090 ;
        RECT 84.995 2820.090 3167.860 2846.090 ;
        RECT 95.115 2816.090 3074.735 2820.090 ;
        RECT 3167.460 2816.090 3167.860 2820.090 ;
        RECT 84.995 2790.090 3167.860 2816.090 ;
        RECT 95.115 2786.090 3074.735 2790.090 ;
        RECT 3167.460 2786.090 3167.860 2790.090 ;
        RECT 84.995 2760.090 3167.860 2786.090 ;
        RECT 95.115 2756.090 3074.735 2760.090 ;
        RECT 3167.460 2756.090 3167.860 2760.090 ;
        RECT 84.995 2730.090 3167.860 2756.090 ;
        RECT 95.115 2726.090 3074.735 2730.090 ;
        RECT 3167.460 2726.090 3167.860 2730.090 ;
        RECT 84.995 2700.090 3167.860 2726.090 ;
        RECT 95.115 2696.090 3074.735 2700.090 ;
        RECT 3167.460 2696.090 3167.860 2700.090 ;
        RECT 84.995 2670.090 3167.860 2696.090 ;
        RECT 95.115 2666.090 3074.735 2670.090 ;
        RECT 3167.460 2666.090 3167.860 2670.090 ;
        RECT 84.995 2640.090 3167.860 2666.090 ;
        RECT 95.115 2636.090 3074.735 2640.090 ;
        RECT 3167.460 2636.090 3167.860 2640.090 ;
        RECT 84.995 2610.090 3167.860 2636.090 ;
        RECT 95.115 2606.090 3074.735 2610.090 ;
        RECT 3167.460 2606.090 3167.860 2610.090 ;
        RECT 84.995 2580.090 3167.860 2606.090 ;
        RECT 95.115 2576.090 3074.735 2580.090 ;
        RECT 3167.460 2576.090 3167.860 2580.090 ;
        RECT 84.995 2550.090 3167.860 2576.090 ;
        RECT 95.115 2546.090 3074.735 2550.090 ;
        RECT 3167.460 2546.090 3167.860 2550.090 ;
        RECT 84.995 2520.090 3167.860 2546.090 ;
        RECT 95.115 2516.090 3074.735 2520.090 ;
        RECT 3167.460 2516.090 3167.860 2520.090 ;
        RECT 84.995 2490.090 3167.860 2516.090 ;
        RECT 95.115 2486.090 3074.735 2490.090 ;
        RECT 3167.460 2486.090 3167.860 2490.090 ;
        RECT 84.995 2460.090 3167.860 2486.090 ;
        RECT 95.115 2456.090 3074.735 2460.090 ;
        RECT 3167.460 2456.090 3167.860 2460.090 ;
        RECT 84.995 2430.090 3167.860 2456.090 ;
        RECT 95.115 2426.090 3074.735 2430.090 ;
        RECT 3167.460 2426.090 3167.860 2430.090 ;
        RECT 84.995 2400.090 3167.860 2426.090 ;
        RECT 95.115 2396.090 3074.735 2400.090 ;
        RECT 3167.460 2396.090 3167.860 2400.090 ;
        RECT 84.995 2370.090 3167.860 2396.090 ;
        RECT 95.115 2366.090 3074.735 2370.090 ;
        RECT 3167.460 2366.090 3167.860 2370.090 ;
        RECT 84.995 2340.090 3167.860 2366.090 ;
        RECT 95.115 2336.090 3074.735 2340.090 ;
        RECT 3167.460 2336.090 3167.860 2340.090 ;
        RECT 84.995 2310.090 3167.860 2336.090 ;
        RECT 95.115 2306.090 3074.735 2310.090 ;
        RECT 3167.460 2306.090 3167.860 2310.090 ;
        RECT 84.995 2280.090 3167.860 2306.090 ;
        RECT 95.115 2276.090 3074.735 2280.090 ;
        RECT 3167.460 2276.090 3167.860 2280.090 ;
        RECT 84.995 2250.090 3167.860 2276.090 ;
        RECT 95.115 2246.090 3074.735 2250.090 ;
        RECT 3167.460 2246.090 3167.860 2250.090 ;
        RECT 84.995 2220.090 3167.860 2246.090 ;
        RECT 95.115 2216.090 3074.735 2220.090 ;
        RECT 3167.460 2216.090 3167.860 2220.090 ;
        RECT 84.995 2190.090 3167.860 2216.090 ;
        RECT 95.115 2186.090 3074.735 2190.090 ;
        RECT 3167.460 2186.090 3167.860 2190.090 ;
        RECT 84.995 2160.090 3167.860 2186.090 ;
        RECT 95.115 2156.090 3074.735 2160.090 ;
        RECT 3167.460 2156.090 3167.860 2160.090 ;
        RECT 84.995 2130.090 3167.860 2156.090 ;
        RECT 95.115 2126.090 3074.735 2130.090 ;
        RECT 3167.460 2126.090 3167.860 2130.090 ;
        RECT 84.995 2100.090 3167.860 2126.090 ;
        RECT 95.115 2096.090 3074.735 2100.090 ;
        RECT 3167.460 2096.090 3167.860 2100.090 ;
        RECT 84.995 2070.090 3167.860 2096.090 ;
        RECT 95.115 2066.090 3074.735 2070.090 ;
        RECT 3167.460 2066.090 3167.860 2070.090 ;
        RECT 84.995 2040.090 3167.860 2066.090 ;
        RECT 95.115 2036.090 3074.735 2040.090 ;
        RECT 3167.460 2036.090 3167.860 2040.090 ;
        RECT 84.995 2010.090 3167.860 2036.090 ;
        RECT 95.115 2006.090 3074.735 2010.090 ;
        RECT 3167.460 2006.090 3167.860 2010.090 ;
        RECT 84.995 1980.090 3167.860 2006.090 ;
        RECT 95.115 1976.090 3074.735 1980.090 ;
        RECT 3167.460 1976.090 3167.860 1980.090 ;
        RECT 84.995 1950.090 3167.860 1976.090 ;
        RECT 95.115 1946.090 3074.735 1950.090 ;
        RECT 3167.460 1946.090 3167.860 1950.090 ;
        RECT 84.995 1920.090 3167.860 1946.090 ;
        RECT 95.115 1916.090 3074.735 1920.090 ;
        RECT 3167.460 1916.090 3167.860 1920.090 ;
        RECT 84.995 1890.090 3167.860 1916.090 ;
        RECT 95.115 1886.090 3074.735 1890.090 ;
        RECT 3167.460 1886.090 3167.860 1890.090 ;
        RECT 84.995 1860.090 3167.860 1886.090 ;
        RECT 95.115 1856.090 3074.735 1860.090 ;
        RECT 3167.460 1856.090 3167.860 1860.090 ;
        RECT 84.995 1830.090 3167.860 1856.090 ;
        RECT 95.115 1826.090 3074.735 1830.090 ;
        RECT 3167.460 1826.090 3167.860 1830.090 ;
        RECT 84.995 1800.090 3167.860 1826.090 ;
        RECT 95.115 1796.090 3074.735 1800.090 ;
        RECT 3167.460 1796.090 3167.860 1800.090 ;
        RECT 84.995 1770.090 3167.860 1796.090 ;
        RECT 95.115 1766.090 3074.735 1770.090 ;
        RECT 3167.460 1766.090 3167.860 1770.090 ;
        RECT 84.995 1740.090 3167.860 1766.090 ;
        RECT 95.115 1736.090 3074.735 1740.090 ;
        RECT 3167.460 1736.090 3167.860 1740.090 ;
        RECT 84.995 1710.090 3167.860 1736.090 ;
        RECT 95.115 1706.090 3074.735 1710.090 ;
        RECT 3167.460 1706.090 3167.860 1710.090 ;
        RECT 84.995 1680.090 3167.860 1706.090 ;
        RECT 95.115 1676.090 3074.735 1680.090 ;
        RECT 3167.460 1676.090 3167.860 1680.090 ;
        RECT 84.995 1650.090 3167.860 1676.090 ;
        RECT 95.115 1646.090 3074.735 1650.090 ;
        RECT 3167.460 1646.090 3167.860 1650.090 ;
        RECT 84.995 1620.090 3167.860 1646.090 ;
        RECT 95.115 1616.090 3074.735 1620.090 ;
        RECT 3167.460 1616.090 3167.860 1620.090 ;
        RECT 84.995 1590.090 3167.860 1616.090 ;
        RECT 95.115 1586.090 3074.735 1590.090 ;
        RECT 3167.460 1586.090 3167.860 1590.090 ;
        RECT 84.995 1560.090 3167.860 1586.090 ;
        RECT 95.115 1556.090 3074.735 1560.090 ;
        RECT 3167.460 1556.090 3167.860 1560.090 ;
        RECT 84.995 1530.090 3167.860 1556.090 ;
        RECT 95.115 1526.090 3074.735 1530.090 ;
        RECT 3167.460 1526.090 3167.860 1530.090 ;
        RECT 84.995 1500.090 3167.860 1526.090 ;
        RECT 95.115 1496.090 3074.735 1500.090 ;
        RECT 3167.460 1496.090 3167.860 1500.090 ;
        RECT 84.995 1470.090 3167.860 1496.090 ;
        RECT 95.115 1466.090 3074.735 1470.090 ;
        RECT 3167.460 1466.090 3167.860 1470.090 ;
        RECT 84.995 1440.090 3167.860 1466.090 ;
        RECT 95.115 1436.090 3074.735 1440.090 ;
        RECT 3167.460 1436.090 3167.860 1440.090 ;
        RECT 84.995 1410.090 3167.860 1436.090 ;
        RECT 95.115 1406.090 3074.735 1410.090 ;
        RECT 3167.460 1406.090 3167.860 1410.090 ;
        RECT 84.995 1380.090 3167.860 1406.090 ;
        RECT 95.115 1376.090 3074.735 1380.090 ;
        RECT 3167.460 1376.090 3167.860 1380.090 ;
        RECT 84.995 1350.090 3167.860 1376.090 ;
        RECT 95.115 1346.090 3074.735 1350.090 ;
        RECT 3167.460 1346.090 3167.860 1350.090 ;
        RECT 84.995 1320.090 3167.860 1346.090 ;
        RECT 95.115 1316.090 3074.735 1320.090 ;
        RECT 3167.460 1316.090 3167.860 1320.090 ;
        RECT 84.995 1290.090 3167.860 1316.090 ;
        RECT 95.115 1286.090 3074.735 1290.090 ;
        RECT 3167.460 1286.090 3167.860 1290.090 ;
        RECT 84.995 1260.090 3167.860 1286.090 ;
        RECT 3167.460 1256.090 3167.860 1260.090 ;
        RECT 84.995 1230.090 3167.860 1256.090 ;
        RECT 3167.460 1226.090 3167.860 1230.090 ;
        RECT 84.995 1200.090 3167.860 1226.090 ;
        RECT 3167.460 1196.090 3167.860 1200.090 ;
        RECT 84.995 1170.090 3167.860 1196.090 ;
        RECT 3167.460 1166.090 3167.860 1170.090 ;
        RECT 84.995 1140.090 3167.860 1166.090 ;
        RECT 3167.460 1136.090 3167.860 1140.090 ;
        RECT 84.995 1110.090 3167.860 1136.090 ;
        RECT 1562.040 1106.090 1636.960 1110.090 ;
        RECT 2121.540 1106.090 2196.460 1110.090 ;
        RECT 3167.460 1106.090 3167.860 1110.090 ;
        RECT 84.995 1080.090 3167.860 1106.090 ;
        RECT 1562.040 1076.090 1636.960 1080.090 ;
        RECT 2121.540 1076.090 2196.460 1080.090 ;
        RECT 3167.460 1076.090 3167.860 1080.090 ;
        RECT 84.995 1050.090 3167.860 1076.090 ;
        RECT 1562.040 1046.090 1636.960 1050.090 ;
        RECT 2121.540 1046.090 2196.460 1050.090 ;
        RECT 3167.460 1046.090 3167.860 1050.090 ;
        RECT 84.995 1020.090 3167.860 1046.090 ;
        RECT 3167.460 1016.090 3167.860 1020.090 ;
        RECT 84.995 990.090 3167.860 1016.090 ;
        RECT 2433.220 986.090 3050.780 990.090 ;
        RECT 3167.460 986.090 3167.860 990.090 ;
        RECT 84.995 960.090 3167.860 986.090 ;
        RECT 602.040 956.090 676.960 960.090 ;
        RECT 1082.040 956.090 1156.960 960.090 ;
        RECT 2433.220 956.090 3050.780 960.090 ;
        RECT 3167.460 956.090 3167.860 960.090 ;
        RECT 84.995 930.090 3167.860 956.090 ;
        RECT 602.040 926.090 676.960 930.090 ;
        RECT 1082.040 926.090 1156.960 930.090 ;
        RECT 2433.220 926.090 3050.780 930.090 ;
        RECT 3167.460 926.090 3167.860 930.090 ;
        RECT 84.995 900.090 3167.860 926.090 ;
        RECT 602.040 896.090 676.960 900.090 ;
        RECT 1082.040 896.090 1156.960 900.090 ;
        RECT 2433.220 896.090 3050.780 900.090 ;
        RECT 3167.460 896.090 3167.860 900.090 ;
        RECT 84.995 870.090 3167.860 896.090 ;
        RECT 2433.220 866.090 3050.780 870.090 ;
        RECT 3167.460 866.090 3167.860 870.090 ;
        RECT 84.995 840.090 3167.860 866.090 ;
        RECT 2433.220 836.090 3050.780 840.090 ;
        RECT 3167.460 836.090 3167.860 840.090 ;
        RECT 84.995 810.090 3167.860 836.090 ;
        RECT 2433.220 806.090 3050.780 810.090 ;
        RECT 3167.460 806.090 3167.860 810.090 ;
        RECT 84.995 780.090 3167.860 806.090 ;
        RECT 2433.220 776.090 3050.780 780.090 ;
        RECT 3167.460 776.090 3167.860 780.090 ;
        RECT 84.995 750.090 3167.860 776.090 ;
        RECT 2433.220 746.090 3050.780 750.090 ;
        RECT 3167.460 746.090 3167.860 750.090 ;
        RECT 84.995 720.090 3167.860 746.090 ;
        RECT 2433.220 716.090 3050.780 720.090 ;
        RECT 3167.460 716.090 3167.860 720.090 ;
        RECT 84.995 690.090 3167.860 716.090 ;
        RECT 2433.220 686.090 3050.780 690.090 ;
        RECT 3167.460 686.090 3167.860 690.090 ;
        RECT 84.995 660.090 3167.860 686.090 ;
        RECT 2433.220 656.090 3050.780 660.090 ;
        RECT 3167.460 656.090 3167.860 660.090 ;
        RECT 84.995 630.090 3167.860 656.090 ;
        RECT 2433.220 626.090 3050.780 630.090 ;
        RECT 3167.460 626.090 3167.860 630.090 ;
        RECT 84.995 600.090 3167.860 626.090 ;
        RECT 2433.220 596.090 3050.780 600.090 ;
        RECT 3167.460 596.090 3167.860 600.090 ;
        RECT 84.995 570.090 3167.860 596.090 ;
        RECT 2433.220 566.090 3050.780 570.090 ;
        RECT 3167.460 566.090 3167.860 570.090 ;
        RECT 84.995 540.090 3167.860 566.090 ;
        RECT 2433.220 536.090 3050.780 540.090 ;
        RECT 3167.460 536.090 3167.860 540.090 ;
        RECT 84.995 510.090 3167.860 536.090 ;
        RECT 2433.220 506.090 3050.780 510.090 ;
        RECT 3167.460 506.090 3167.860 510.090 ;
        RECT 84.995 480.090 3167.860 506.090 ;
        RECT 2433.220 476.090 3050.780 480.090 ;
        RECT 3167.460 476.090 3167.860 480.090 ;
        RECT 84.995 450.090 3167.860 476.090 ;
        RECT 2433.220 446.090 3050.780 450.090 ;
        RECT 3167.460 446.090 3167.860 450.090 ;
        RECT 84.995 420.090 3167.860 446.090 ;
        RECT 2433.220 416.090 3050.780 420.090 ;
        RECT 3167.460 416.090 3167.860 420.090 ;
        RECT 84.995 390.090 3167.860 416.090 ;
        RECT 2433.220 386.090 3050.780 390.090 ;
        RECT 3167.460 386.090 3167.860 390.090 ;
        RECT 84.995 360.090 3167.860 386.090 ;
        RECT 2433.220 356.090 3050.780 360.090 ;
        RECT 3167.460 356.090 3167.860 360.090 ;
        RECT 84.995 330.090 3167.860 356.090 ;
        RECT 2433.220 326.090 3050.780 330.090 ;
        RECT 3167.460 326.090 3167.860 330.090 ;
        RECT 84.995 300.090 3167.860 326.090 ;
        RECT 2433.220 296.090 3050.780 300.090 ;
        RECT 3167.460 296.090 3167.860 300.090 ;
        RECT 84.995 270.090 3167.860 296.090 ;
        RECT 2433.220 266.090 3050.780 270.090 ;
        RECT 3167.460 266.090 3167.860 270.090 ;
        RECT 84.995 240.090 3167.860 266.090 ;
        RECT 2433.220 236.090 3050.780 240.090 ;
        RECT 3167.460 236.090 3167.860 240.090 ;
        RECT 84.995 210.090 3167.860 236.090 ;
        RECT 2433.220 206.090 3050.780 210.090 ;
        RECT 3167.460 206.090 3167.860 210.090 ;
        RECT 84.995 180.090 3167.860 206.090 ;
        RECT 3167.460 176.090 3167.860 180.090 ;
        RECT 84.995 150.090 3167.860 176.090 ;
        RECT 2896.855 146.090 2966.495 150.090 ;
        RECT 3167.460 146.090 3167.860 150.090 ;
        RECT 84.995 120.090 3167.860 146.090 ;
        RECT 2896.855 116.090 2966.495 120.090 ;
        RECT 3167.460 116.090 3167.860 120.090 ;
        RECT 84.995 90.090 3167.860 116.090 ;
        RECT 2897.355 86.090 2966.495 90.090 ;
        RECT 3167.460 86.090 3167.860 90.090 ;
        RECT 84.995 60.090 3167.860 86.090 ;
        RECT 3167.460 56.090 3167.860 60.090 ;
        RECT 84.995 45.980 3167.860 56.090 ;
  END
END caravel_core
END LIBRARY

