magic
tech gf180mcuC
magscale 1 10
timestamp 1655473255
<< checkpaint >>
rect -2000 -2000 23672 4313
<< obsm1 >>
rect 889 528 20825 2216
<< metal2 >>
rect 0 0 56 1076
rect 672 0 728 899
rect 1456 0 1512 766
rect 2128 0 2184 608
rect 2800 0 2856 618
rect 3472 0 3528 899
rect 4144 0 4200 722
rect 4928 0 4984 899
rect 5600 0 5656 659
rect 6272 0 6328 899
rect 6944 0 7000 1909
rect 7728 0 7784 900
rect 8400 0 8456 1909
rect 9072 0 9128 899
rect 9744 0 9800 1909
rect 10416 0 10472 899
rect 11200 0 11256 1909
rect 11872 0 11928 899
rect 12544 0 12600 1909
rect 13216 0 13272 878
rect 14000 0 14056 609
rect 14672 0 14728 899
rect 15344 0 15400 709
rect 16016 0 16072 899
rect 16688 0 16744 717
rect 17472 0 17528 899
rect 18144 0 18200 774
rect 18816 0 18872 731
rect 19488 0 19544 779
rect 20272 0 20328 767
rect 20944 0 21000 769
rect 21616 0 21672 899
<< obsm2 >>
rect 56 1969 21616 2313
rect 56 1136 6884 1969
rect 116 959 6884 1136
rect 116 425 612 959
rect 788 826 3412 959
rect 788 425 1396 826
rect 1572 678 3412 826
rect 1572 668 2740 678
rect 1572 425 2068 668
rect 2244 425 2740 668
rect 2916 425 3412 678
rect 3588 782 4868 959
rect 3588 425 4084 782
rect 4260 425 4868 782
rect 5044 719 6212 959
rect 5044 425 5540 719
rect 5716 425 6212 719
rect 6388 425 6884 959
rect 7060 960 8340 1969
rect 7060 425 7668 960
rect 7844 425 8340 960
rect 8516 959 9684 1969
rect 8516 425 9012 959
rect 9188 425 9684 959
rect 9860 959 11140 1969
rect 9860 425 10356 959
rect 10532 425 11140 959
rect 11316 959 12484 1969
rect 11316 425 11812 959
rect 11988 425 12484 959
rect 12660 959 21616 1969
rect 12660 938 14612 959
rect 12660 425 13156 938
rect 13332 669 14612 938
rect 13332 425 13940 669
rect 14116 425 14612 669
rect 14788 769 15956 959
rect 14788 425 15284 769
rect 15460 425 15956 769
rect 16132 777 17412 959
rect 16132 425 16628 777
rect 16804 425 17412 777
rect 17588 839 21556 959
rect 17588 834 19428 839
rect 17588 425 18084 834
rect 18260 791 19428 834
rect 18260 425 18756 791
rect 18932 425 19428 791
rect 19604 829 21556 839
rect 19604 827 20884 829
rect 19604 425 20212 827
rect 20388 425 20884 827
rect 21060 425 21556 829
<< obsm3 >>
rect 1696 425 20014 2313
<< obsm4 >>
rect 1696 425 20013 2313
<< metal5 >>
rect 741 1225 6209 1545
rect 741 425 1709 745
<< obsm5 >>
rect 741 1645 20916 2313
rect 6309 1125 20916 1645
rect 741 845 20916 1125
rect 1809 425 20916 845
<< labels >>
rlabel metal2 s 0 0 56 1076 6 mask_rev[0]
port 1 nsew
rlabel metal2 s 6944 0 7000 1909 6 mask_rev[10]
port 2 nsew
rlabel metal2 s 7728 0 7784 900 6 mask_rev[11]
port 3 nsew
rlabel metal2 s 8400 0 8456 1909 6 mask_rev[12]
port 4 nsew
rlabel metal2 s 9072 0 9128 899 6 mask_rev[13]
port 5 nsew
rlabel metal2 s 9744 0 9800 1909 6 mask_rev[14]
port 6 nsew
rlabel metal2 s 10416 0 10472 899 6 mask_rev[15]
port 7 nsew
rlabel metal2 s 11200 0 11256 1909 6 mask_rev[16]
port 8 nsew
rlabel metal2 s 11872 0 11928 899 6 mask_rev[17]
port 9 nsew
rlabel metal2 s 12544 0 12600 1909 6 mask_rev[18]
port 10 nsew
rlabel metal2 s 13216 0 13272 878 6 mask_rev[19]
port 11 nsew
rlabel metal2 s 672 0 728 899 6 mask_rev[1]
port 12 nsew
rlabel metal2 s 14000 0 14056 609 6 mask_rev[20]
port 13 nsew
rlabel metal2 s 14672 0 14728 899 6 mask_rev[21]
port 14 nsew
rlabel metal2 s 15344 0 15400 709 6 mask_rev[22]
port 15 nsew
rlabel metal2 s 16016 0 16072 899 6 mask_rev[23]
port 16 nsew
rlabel metal2 s 16688 0 16744 717 6 mask_rev[24]
port 17 nsew
rlabel metal2 s 17472 0 17528 899 6 mask_rev[25]
port 18 nsew
rlabel metal2 s 18144 0 18200 774 6 mask_rev[26]
port 19 nsew
rlabel metal2 s 18816 0 18872 731 6 mask_rev[27]
port 20 nsew
rlabel metal2 s 19488 0 19544 779 6 mask_rev[28]
port 21 nsew
rlabel metal2 s 20272 0 20328 767 6 mask_rev[29]
port 22 nsew
rlabel metal2 s 1456 0 1512 766 6 mask_rev[2]
port 23 nsew
rlabel metal2 s 20944 0 21000 769 6 mask_rev[30]
port 24 nsew
rlabel metal2 s 21616 0 21672 899 6 mask_rev[31]
port 25 nsew
rlabel metal2 s 2128 0 2184 608 6 mask_rev[3]
port 26 nsew
rlabel metal2 s 2800 0 2856 618 6 mask_rev[4]
port 27 nsew
rlabel metal2 s 3472 0 3528 899 6 mask_rev[5]
port 28 nsew
rlabel metal2 s 4144 0 4200 722 6 mask_rev[6]
port 29 nsew
rlabel metal2 s 4928 0 4984 899 6 mask_rev[7]
port 30 nsew
rlabel metal2 s 5600 0 5656 659 6 mask_rev[8]
port 31 nsew
rlabel metal2 s 6272 0 6328 899 6 mask_rev[9]
port 32 nsew
rlabel metal5 s 741 1225 6209 1545 6 VDD
port 33 nsew power default
rlabel metal5 s 741 425 1709 745 6 VSS
port 34 nsew ground default
<< properties >>
string FIXED_BBOX 0 0 21672 2313
string GDS_END 66360
string GDS_FILE ../gds/user_id_programming.gds
string GDS_START 9860
string LEFclass BLOCK
string LEFview TRUE
<< end >>
