VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_gf180_pdn
  CLASS BLOCK ;
  FOREIGN caravel_gf180_pdn ;
  ORIGIN 0 0 ;
  SIZE 3192.000 BY 4402.000 ;
  OBS
      LAYER Metal2 ;
        RECT 1906.360 4749.000 1915.860 4751.000 ;
        RECT 1918.760 4749.000 1929.010 4751.000 ;
        RECT 1930.610 4749.000 1940.860 4751.000 ;
        RECT 1944.140 4749.000 1954.390 4751.000 ;
        RECT 1955.990 4749.000 1966.240 4751.000 ;
        RECT 1969.140 4749.000 1978.640 4751.000 ;
        RECT 3006.360 4749.000 3015.860 4751.000 ;
        RECT 3018.760 4749.000 3029.010 4751.000 ;
        RECT 3030.610 4749.000 3040.860 4751.000 ;
        RECT 3044.140 4749.000 3054.390 4751.000 ;
        RECT 3055.990 4749.000 3066.240 4751.000 ;
        RECT 3069.140 4749.000 3078.640 4751.000 ;
        RECT 349.000 4414.140 351.000 4423.640 ;
        RECT 349.000 4400.990 351.000 4411.240 ;
        RECT 3539.000 4409.140 3541.000 4418.640 ;
        RECT 349.000 4389.140 351.000 4399.390 ;
        RECT 3539.000 4395.990 3541.000 4406.240 ;
        RECT 349.000 4375.610 351.000 4385.860 ;
        RECT 3539.000 4384.140 3541.000 4394.390 ;
        RECT 349.000 4363.760 351.000 4374.010 ;
        RECT 3539.000 4370.610 3541.000 4380.860 ;
        RECT 349.000 4351.360 351.000 4360.860 ;
        RECT 3539.000 4358.760 3541.000 4369.010 ;
        RECT 3539.000 4346.360 3541.000 4355.860 ;
        RECT 349.000 4209.140 351.000 4218.640 ;
        RECT 349.000 4195.990 351.000 4206.240 ;
        RECT 349.000 4184.140 351.000 4194.390 ;
        RECT 349.000 4170.610 351.000 4180.860 ;
        RECT 349.000 4158.760 351.000 4169.010 ;
        RECT 349.000 4146.360 351.000 4155.860 ;
        RECT 349.000 4004.140 351.000 4013.640 ;
        RECT 349.000 3990.990 351.000 4001.240 ;
        RECT 349.000 3979.140 351.000 3989.390 ;
        RECT 3539.000 3979.140 3541.000 3988.640 ;
        RECT 349.000 3965.610 351.000 3975.860 ;
        RECT 3539.000 3965.990 3541.000 3976.240 ;
        RECT 349.000 3953.760 351.000 3964.010 ;
        RECT 3539.000 3954.140 3541.000 3964.390 ;
        RECT 349.000 3941.360 351.000 3950.860 ;
        RECT 3539.000 3940.610 3541.000 3950.860 ;
        RECT 3539.000 3928.760 3541.000 3939.010 ;
        RECT 3539.000 3916.360 3541.000 3925.860 ;
        RECT 3539.000 2474.140 3541.000 2483.640 ;
        RECT 3539.000 2460.990 3541.000 2471.240 ;
        RECT 3539.000 2449.140 3541.000 2459.390 ;
        RECT 3539.000 2435.610 3541.000 2445.860 ;
        RECT 3539.000 2423.760 3541.000 2434.010 ;
        RECT 3539.000 2411.360 3541.000 2420.860 ;
        RECT 349.000 2364.140 351.000 2373.640 ;
        RECT 349.000 2350.990 351.000 2361.240 ;
        RECT 349.000 2339.140 351.000 2349.390 ;
        RECT 349.000 2325.610 351.000 2335.860 ;
        RECT 349.000 2313.760 351.000 2324.010 ;
        RECT 349.000 2301.360 351.000 2310.860 ;
        RECT 3539.000 2259.140 3541.000 2268.640 ;
        RECT 3539.000 2245.990 3541.000 2256.240 ;
        RECT 3539.000 2234.140 3541.000 2244.390 ;
        RECT 3539.000 2220.610 3541.000 2230.860 ;
        RECT 3539.000 2208.760 3541.000 2219.010 ;
        RECT 3539.000 2196.360 3541.000 2205.860 ;
        RECT 349.000 2159.140 351.000 2168.640 ;
        RECT 349.000 2145.990 351.000 2156.240 ;
        RECT 349.000 2134.140 351.000 2144.390 ;
        RECT 349.000 2120.610 351.000 2130.860 ;
        RECT 349.000 2108.760 351.000 2119.010 ;
        RECT 349.000 2096.360 351.000 2105.860 ;
        RECT 3539.000 2044.140 3541.000 2053.640 ;
        RECT 3539.000 2030.990 3541.000 2041.240 ;
        RECT 3539.000 2019.140 3541.000 2029.390 ;
        RECT 3539.000 2005.610 3541.000 2015.860 ;
        RECT 3539.000 1993.760 3541.000 2004.010 ;
        RECT 3539.000 1981.360 3541.000 1990.860 ;
        RECT 349.000 724.140 351.000 733.640 ;
        RECT 349.000 710.990 351.000 721.240 ;
        RECT 349.000 699.140 351.000 709.390 ;
        RECT 349.000 685.610 351.000 695.860 ;
        RECT 349.000 673.760 351.000 684.010 ;
        RECT 349.000 661.360 351.000 670.860 ;
        RECT 349.000 519.140 351.000 528.640 ;
        RECT 349.000 505.990 351.000 516.240 ;
        RECT 349.000 494.140 351.000 504.390 ;
        RECT 349.000 480.610 351.000 490.860 ;
        RECT 349.000 468.760 351.000 479.010 ;
        RECT 349.000 456.360 351.000 465.860 ;
        RECT 536.360 349.000 545.860 351.000 ;
        RECT 548.760 349.000 559.010 351.000 ;
        RECT 560.610 349.000 570.860 351.000 ;
        RECT 574.140 349.000 584.390 351.000 ;
        RECT 585.990 349.000 596.240 351.000 ;
        RECT 599.140 349.000 608.640 351.000 ;
        RECT 1361.360 349.000 1370.860 351.000 ;
        RECT 1373.760 349.000 1384.010 351.000 ;
        RECT 1385.610 349.000 1395.860 351.000 ;
        RECT 1399.140 349.000 1409.390 351.000 ;
        RECT 1410.990 349.000 1421.240 351.000 ;
        RECT 1424.140 349.000 1433.640 351.000 ;
        RECT 3011.360 349.000 3020.860 351.000 ;
        RECT 3023.760 349.000 3034.010 351.000 ;
        RECT 3035.610 349.000 3045.860 351.000 ;
        RECT 3049.140 349.000 3059.390 351.000 ;
        RECT 3060.990 349.000 3071.240 351.000 ;
        RECT 3074.140 349.000 3083.640 351.000 ;
        RECT 3286.360 349.000 3295.860 351.000 ;
        RECT 3298.760 349.000 3309.010 351.000 ;
        RECT 3310.610 349.000 3320.860 351.000 ;
        RECT 3324.140 349.000 3334.390 351.000 ;
        RECT 3335.990 349.000 3346.240 351.000 ;
        RECT 3349.140 349.000 3358.640 351.000 ;
      LAYER VIA2 ;
        RECT 1906.710 4749.350 1906.990 4749.630 ;
        RECT 1907.330 4749.350 1907.610 4749.630 ;
        RECT 1907.950 4749.350 1908.230 4749.630 ;
        RECT 1908.570 4749.350 1908.850 4749.630 ;
        RECT 1909.190 4749.350 1909.470 4749.630 ;
        RECT 1909.810 4749.350 1910.090 4749.630 ;
        RECT 1910.430 4749.350 1910.710 4749.630 ;
        RECT 1911.050 4749.350 1911.330 4749.630 ;
        RECT 1911.670 4749.350 1911.950 4749.630 ;
        RECT 1912.290 4749.350 1912.570 4749.630 ;
        RECT 1912.910 4749.350 1913.190 4749.630 ;
        RECT 1913.530 4749.350 1913.810 4749.630 ;
        RECT 1914.150 4749.350 1914.430 4749.630 ;
        RECT 1914.770 4749.350 1915.050 4749.630 ;
        RECT 1915.390 4749.350 1915.670 4749.630 ;
        RECT 1919.110 4749.350 1919.390 4749.630 ;
        RECT 1919.730 4749.350 1920.010 4749.630 ;
        RECT 1920.350 4749.350 1920.630 4749.630 ;
        RECT 1920.970 4749.350 1921.250 4749.630 ;
        RECT 1921.590 4749.350 1921.870 4749.630 ;
        RECT 1922.210 4749.350 1922.490 4749.630 ;
        RECT 1922.830 4749.350 1923.110 4749.630 ;
        RECT 1923.450 4749.350 1923.730 4749.630 ;
        RECT 1924.070 4749.350 1924.350 4749.630 ;
        RECT 1924.690 4749.350 1924.970 4749.630 ;
        RECT 1925.310 4749.350 1925.590 4749.630 ;
        RECT 1925.930 4749.350 1926.210 4749.630 ;
        RECT 1926.550 4749.350 1926.830 4749.630 ;
        RECT 1927.170 4749.350 1927.450 4749.630 ;
        RECT 1927.790 4749.350 1928.070 4749.630 ;
        RECT 1928.410 4749.350 1928.690 4749.630 ;
        RECT 1930.960 4749.350 1931.240 4749.630 ;
        RECT 1931.580 4749.350 1931.860 4749.630 ;
        RECT 1932.200 4749.350 1932.480 4749.630 ;
        RECT 1932.820 4749.350 1933.100 4749.630 ;
        RECT 1933.440 4749.350 1933.720 4749.630 ;
        RECT 1934.060 4749.350 1934.340 4749.630 ;
        RECT 1934.680 4749.350 1934.960 4749.630 ;
        RECT 1935.300 4749.350 1935.580 4749.630 ;
        RECT 1935.920 4749.350 1936.200 4749.630 ;
        RECT 1936.540 4749.350 1936.820 4749.630 ;
        RECT 1937.160 4749.350 1937.440 4749.630 ;
        RECT 1937.780 4749.350 1938.060 4749.630 ;
        RECT 1938.400 4749.350 1938.680 4749.630 ;
        RECT 1939.020 4749.350 1939.300 4749.630 ;
        RECT 1939.640 4749.350 1939.920 4749.630 ;
        RECT 1940.260 4749.350 1940.540 4749.630 ;
        RECT 1944.460 4749.350 1944.740 4749.630 ;
        RECT 1945.080 4749.350 1945.360 4749.630 ;
        RECT 1945.700 4749.350 1945.980 4749.630 ;
        RECT 1946.320 4749.350 1946.600 4749.630 ;
        RECT 1946.940 4749.350 1947.220 4749.630 ;
        RECT 1947.560 4749.350 1947.840 4749.630 ;
        RECT 1948.180 4749.350 1948.460 4749.630 ;
        RECT 1948.800 4749.350 1949.080 4749.630 ;
        RECT 1949.420 4749.350 1949.700 4749.630 ;
        RECT 1950.040 4749.350 1950.320 4749.630 ;
        RECT 1950.660 4749.350 1950.940 4749.630 ;
        RECT 1951.280 4749.350 1951.560 4749.630 ;
        RECT 1951.900 4749.350 1952.180 4749.630 ;
        RECT 1952.520 4749.350 1952.800 4749.630 ;
        RECT 1953.140 4749.350 1953.420 4749.630 ;
        RECT 1953.760 4749.350 1954.040 4749.630 ;
        RECT 1956.310 4749.350 1956.590 4749.630 ;
        RECT 1956.930 4749.350 1957.210 4749.630 ;
        RECT 1957.550 4749.350 1957.830 4749.630 ;
        RECT 1958.170 4749.350 1958.450 4749.630 ;
        RECT 1958.790 4749.350 1959.070 4749.630 ;
        RECT 1959.410 4749.350 1959.690 4749.630 ;
        RECT 1960.030 4749.350 1960.310 4749.630 ;
        RECT 1960.650 4749.350 1960.930 4749.630 ;
        RECT 1961.270 4749.350 1961.550 4749.630 ;
        RECT 1961.890 4749.350 1962.170 4749.630 ;
        RECT 1962.510 4749.350 1962.790 4749.630 ;
        RECT 1963.130 4749.350 1963.410 4749.630 ;
        RECT 1963.750 4749.350 1964.030 4749.630 ;
        RECT 1964.370 4749.350 1964.650 4749.630 ;
        RECT 1964.990 4749.350 1965.270 4749.630 ;
        RECT 1965.610 4749.350 1965.890 4749.630 ;
        RECT 1969.330 4749.350 1969.610 4749.630 ;
        RECT 1969.950 4749.350 1970.230 4749.630 ;
        RECT 1970.570 4749.350 1970.850 4749.630 ;
        RECT 1971.190 4749.350 1971.470 4749.630 ;
        RECT 1971.810 4749.350 1972.090 4749.630 ;
        RECT 1972.430 4749.350 1972.710 4749.630 ;
        RECT 1973.050 4749.350 1973.330 4749.630 ;
        RECT 1973.670 4749.350 1973.950 4749.630 ;
        RECT 1974.290 4749.350 1974.570 4749.630 ;
        RECT 1974.910 4749.350 1975.190 4749.630 ;
        RECT 1975.530 4749.350 1975.810 4749.630 ;
        RECT 1976.150 4749.350 1976.430 4749.630 ;
        RECT 1976.770 4749.350 1977.050 4749.630 ;
        RECT 1977.390 4749.350 1977.670 4749.630 ;
        RECT 1978.010 4749.350 1978.290 4749.630 ;
        RECT 3006.710 4749.350 3006.990 4749.630 ;
        RECT 3007.330 4749.350 3007.610 4749.630 ;
        RECT 3007.950 4749.350 3008.230 4749.630 ;
        RECT 3008.570 4749.350 3008.850 4749.630 ;
        RECT 3009.190 4749.350 3009.470 4749.630 ;
        RECT 3009.810 4749.350 3010.090 4749.630 ;
        RECT 3010.430 4749.350 3010.710 4749.630 ;
        RECT 3011.050 4749.350 3011.330 4749.630 ;
        RECT 3011.670 4749.350 3011.950 4749.630 ;
        RECT 3012.290 4749.350 3012.570 4749.630 ;
        RECT 3012.910 4749.350 3013.190 4749.630 ;
        RECT 3013.530 4749.350 3013.810 4749.630 ;
        RECT 3014.150 4749.350 3014.430 4749.630 ;
        RECT 3014.770 4749.350 3015.050 4749.630 ;
        RECT 3015.390 4749.350 3015.670 4749.630 ;
        RECT 3019.110 4749.350 3019.390 4749.630 ;
        RECT 3019.730 4749.350 3020.010 4749.630 ;
        RECT 3020.350 4749.350 3020.630 4749.630 ;
        RECT 3020.970 4749.350 3021.250 4749.630 ;
        RECT 3021.590 4749.350 3021.870 4749.630 ;
        RECT 3022.210 4749.350 3022.490 4749.630 ;
        RECT 3022.830 4749.350 3023.110 4749.630 ;
        RECT 3023.450 4749.350 3023.730 4749.630 ;
        RECT 3024.070 4749.350 3024.350 4749.630 ;
        RECT 3024.690 4749.350 3024.970 4749.630 ;
        RECT 3025.310 4749.350 3025.590 4749.630 ;
        RECT 3025.930 4749.350 3026.210 4749.630 ;
        RECT 3026.550 4749.350 3026.830 4749.630 ;
        RECT 3027.170 4749.350 3027.450 4749.630 ;
        RECT 3027.790 4749.350 3028.070 4749.630 ;
        RECT 3028.410 4749.350 3028.690 4749.630 ;
        RECT 3030.960 4749.350 3031.240 4749.630 ;
        RECT 3031.580 4749.350 3031.860 4749.630 ;
        RECT 3032.200 4749.350 3032.480 4749.630 ;
        RECT 3032.820 4749.350 3033.100 4749.630 ;
        RECT 3033.440 4749.350 3033.720 4749.630 ;
        RECT 3034.060 4749.350 3034.340 4749.630 ;
        RECT 3034.680 4749.350 3034.960 4749.630 ;
        RECT 3035.300 4749.350 3035.580 4749.630 ;
        RECT 3035.920 4749.350 3036.200 4749.630 ;
        RECT 3036.540 4749.350 3036.820 4749.630 ;
        RECT 3037.160 4749.350 3037.440 4749.630 ;
        RECT 3037.780 4749.350 3038.060 4749.630 ;
        RECT 3038.400 4749.350 3038.680 4749.630 ;
        RECT 3039.020 4749.350 3039.300 4749.630 ;
        RECT 3039.640 4749.350 3039.920 4749.630 ;
        RECT 3040.260 4749.350 3040.540 4749.630 ;
        RECT 3044.460 4749.350 3044.740 4749.630 ;
        RECT 3045.080 4749.350 3045.360 4749.630 ;
        RECT 3045.700 4749.350 3045.980 4749.630 ;
        RECT 3046.320 4749.350 3046.600 4749.630 ;
        RECT 3046.940 4749.350 3047.220 4749.630 ;
        RECT 3047.560 4749.350 3047.840 4749.630 ;
        RECT 3048.180 4749.350 3048.460 4749.630 ;
        RECT 3048.800 4749.350 3049.080 4749.630 ;
        RECT 3049.420 4749.350 3049.700 4749.630 ;
        RECT 3050.040 4749.350 3050.320 4749.630 ;
        RECT 3050.660 4749.350 3050.940 4749.630 ;
        RECT 3051.280 4749.350 3051.560 4749.630 ;
        RECT 3051.900 4749.350 3052.180 4749.630 ;
        RECT 3052.520 4749.350 3052.800 4749.630 ;
        RECT 3053.140 4749.350 3053.420 4749.630 ;
        RECT 3053.760 4749.350 3054.040 4749.630 ;
        RECT 3056.310 4749.350 3056.590 4749.630 ;
        RECT 3056.930 4749.350 3057.210 4749.630 ;
        RECT 3057.550 4749.350 3057.830 4749.630 ;
        RECT 3058.170 4749.350 3058.450 4749.630 ;
        RECT 3058.790 4749.350 3059.070 4749.630 ;
        RECT 3059.410 4749.350 3059.690 4749.630 ;
        RECT 3060.030 4749.350 3060.310 4749.630 ;
        RECT 3060.650 4749.350 3060.930 4749.630 ;
        RECT 3061.270 4749.350 3061.550 4749.630 ;
        RECT 3061.890 4749.350 3062.170 4749.630 ;
        RECT 3062.510 4749.350 3062.790 4749.630 ;
        RECT 3063.130 4749.350 3063.410 4749.630 ;
        RECT 3063.750 4749.350 3064.030 4749.630 ;
        RECT 3064.370 4749.350 3064.650 4749.630 ;
        RECT 3064.990 4749.350 3065.270 4749.630 ;
        RECT 3065.610 4749.350 3065.890 4749.630 ;
        RECT 3069.330 4749.350 3069.610 4749.630 ;
        RECT 3069.950 4749.350 3070.230 4749.630 ;
        RECT 3070.570 4749.350 3070.850 4749.630 ;
        RECT 3071.190 4749.350 3071.470 4749.630 ;
        RECT 3071.810 4749.350 3072.090 4749.630 ;
        RECT 3072.430 4749.350 3072.710 4749.630 ;
        RECT 3073.050 4749.350 3073.330 4749.630 ;
        RECT 3073.670 4749.350 3073.950 4749.630 ;
        RECT 3074.290 4749.350 3074.570 4749.630 ;
        RECT 3074.910 4749.350 3075.190 4749.630 ;
        RECT 3075.530 4749.350 3075.810 4749.630 ;
        RECT 3076.150 4749.350 3076.430 4749.630 ;
        RECT 3076.770 4749.350 3077.050 4749.630 ;
        RECT 3077.390 4749.350 3077.670 4749.630 ;
        RECT 3078.010 4749.350 3078.290 4749.630 ;
        RECT 350.370 4423.010 350.650 4423.290 ;
        RECT 350.370 4422.390 350.650 4422.670 ;
        RECT 350.370 4421.770 350.650 4422.050 ;
        RECT 350.370 4421.150 350.650 4421.430 ;
        RECT 350.370 4420.530 350.650 4420.810 ;
        RECT 350.370 4419.910 350.650 4420.190 ;
        RECT 350.370 4419.290 350.650 4419.570 ;
        RECT 350.370 4418.670 350.650 4418.950 ;
        RECT 350.370 4418.050 350.650 4418.330 ;
        RECT 350.370 4417.430 350.650 4417.710 ;
        RECT 350.370 4416.810 350.650 4417.090 ;
        RECT 350.370 4416.190 350.650 4416.470 ;
        RECT 350.370 4415.570 350.650 4415.850 ;
        RECT 350.370 4414.950 350.650 4415.230 ;
        RECT 350.370 4414.330 350.650 4414.610 ;
        RECT 3539.350 4418.010 3539.630 4418.290 ;
        RECT 3539.350 4417.390 3539.630 4417.670 ;
        RECT 3539.350 4416.770 3539.630 4417.050 ;
        RECT 3539.350 4416.150 3539.630 4416.430 ;
        RECT 3539.350 4415.530 3539.630 4415.810 ;
        RECT 3539.350 4414.910 3539.630 4415.190 ;
        RECT 3539.350 4414.290 3539.630 4414.570 ;
        RECT 3539.350 4413.670 3539.630 4413.950 ;
        RECT 3539.350 4413.050 3539.630 4413.330 ;
        RECT 3539.350 4412.430 3539.630 4412.710 ;
        RECT 3539.350 4411.810 3539.630 4412.090 ;
        RECT 350.370 4410.640 350.650 4410.920 ;
        RECT 350.370 4410.020 350.650 4410.300 ;
        RECT 350.370 4409.400 350.650 4409.680 ;
        RECT 3539.350 4411.190 3539.630 4411.470 ;
        RECT 3539.350 4410.570 3539.630 4410.850 ;
        RECT 3539.350 4409.950 3539.630 4410.230 ;
        RECT 3539.350 4409.330 3539.630 4409.610 ;
        RECT 350.370 4408.780 350.650 4409.060 ;
        RECT 350.370 4408.160 350.650 4408.440 ;
        RECT 350.370 4407.540 350.650 4407.820 ;
        RECT 350.370 4406.920 350.650 4407.200 ;
        RECT 350.370 4406.300 350.650 4406.580 ;
        RECT 350.370 4405.680 350.650 4405.960 ;
        RECT 350.370 4405.060 350.650 4405.340 ;
        RECT 350.370 4404.440 350.650 4404.720 ;
        RECT 350.370 4403.820 350.650 4404.100 ;
        RECT 350.370 4403.200 350.650 4403.480 ;
        RECT 350.370 4402.580 350.650 4402.860 ;
        RECT 350.370 4401.960 350.650 4402.240 ;
        RECT 350.370 4401.340 350.650 4401.620 ;
        RECT 3539.350 4405.610 3539.630 4405.890 ;
        RECT 3539.350 4404.990 3539.630 4405.270 ;
        RECT 3539.350 4404.370 3539.630 4404.650 ;
        RECT 3539.350 4403.750 3539.630 4404.030 ;
        RECT 3539.350 4403.130 3539.630 4403.410 ;
        RECT 3539.350 4402.510 3539.630 4402.790 ;
        RECT 3539.350 4401.890 3539.630 4402.170 ;
        RECT 3539.350 4401.270 3539.630 4401.550 ;
        RECT 3539.350 4400.650 3539.630 4400.930 ;
        RECT 3539.350 4400.030 3539.630 4400.310 ;
        RECT 3539.350 4399.410 3539.630 4399.690 ;
        RECT 350.370 4398.790 350.650 4399.070 ;
        RECT 350.370 4398.170 350.650 4398.450 ;
        RECT 350.370 4397.550 350.650 4397.830 ;
        RECT 350.370 4396.930 350.650 4397.210 ;
        RECT 350.370 4396.310 350.650 4396.590 ;
        RECT 3539.350 4398.790 3539.630 4399.070 ;
        RECT 3539.350 4398.170 3539.630 4398.450 ;
        RECT 3539.350 4397.550 3539.630 4397.830 ;
        RECT 3539.350 4396.930 3539.630 4397.210 ;
        RECT 3539.350 4396.310 3539.630 4396.590 ;
        RECT 350.370 4395.690 350.650 4395.970 ;
        RECT 350.370 4395.070 350.650 4395.350 ;
        RECT 350.370 4394.450 350.650 4394.730 ;
        RECT 350.370 4393.830 350.650 4394.110 ;
        RECT 350.370 4393.210 350.650 4393.490 ;
        RECT 350.370 4392.590 350.650 4392.870 ;
        RECT 350.370 4391.970 350.650 4392.250 ;
        RECT 350.370 4391.350 350.650 4391.630 ;
        RECT 350.370 4390.730 350.650 4391.010 ;
        RECT 350.370 4390.110 350.650 4390.390 ;
        RECT 350.370 4389.490 350.650 4389.770 ;
        RECT 3539.350 4393.760 3539.630 4394.040 ;
        RECT 3539.350 4393.140 3539.630 4393.420 ;
        RECT 3539.350 4392.520 3539.630 4392.800 ;
        RECT 3539.350 4391.900 3539.630 4392.180 ;
        RECT 3539.350 4391.280 3539.630 4391.560 ;
        RECT 3539.350 4390.660 3539.630 4390.940 ;
        RECT 3539.350 4390.040 3539.630 4390.320 ;
        RECT 3539.350 4389.420 3539.630 4389.700 ;
        RECT 3539.350 4388.800 3539.630 4389.080 ;
        RECT 3539.350 4388.180 3539.630 4388.460 ;
        RECT 3539.350 4387.560 3539.630 4387.840 ;
        RECT 3539.350 4386.940 3539.630 4387.220 ;
        RECT 3539.350 4386.320 3539.630 4386.600 ;
        RECT 350.370 4385.260 350.650 4385.540 ;
        RECT 350.370 4384.640 350.650 4384.920 ;
        RECT 350.370 4384.020 350.650 4384.300 ;
        RECT 3539.350 4385.700 3539.630 4385.980 ;
        RECT 3539.350 4385.080 3539.630 4385.360 ;
        RECT 3539.350 4384.460 3539.630 4384.740 ;
        RECT 350.370 4383.400 350.650 4383.680 ;
        RECT 350.370 4382.780 350.650 4383.060 ;
        RECT 350.370 4382.160 350.650 4382.440 ;
        RECT 350.370 4381.540 350.650 4381.820 ;
        RECT 350.370 4380.920 350.650 4381.200 ;
        RECT 350.370 4380.300 350.650 4380.580 ;
        RECT 350.370 4379.680 350.650 4379.960 ;
        RECT 350.370 4379.060 350.650 4379.340 ;
        RECT 350.370 4378.440 350.650 4378.720 ;
        RECT 350.370 4377.820 350.650 4378.100 ;
        RECT 350.370 4377.200 350.650 4377.480 ;
        RECT 350.370 4376.580 350.650 4376.860 ;
        RECT 350.370 4375.960 350.650 4376.240 ;
        RECT 3539.350 4380.230 3539.630 4380.510 ;
        RECT 3539.350 4379.610 3539.630 4379.890 ;
        RECT 3539.350 4378.990 3539.630 4379.270 ;
        RECT 3539.350 4378.370 3539.630 4378.650 ;
        RECT 3539.350 4377.750 3539.630 4378.030 ;
        RECT 3539.350 4377.130 3539.630 4377.410 ;
        RECT 3539.350 4376.510 3539.630 4376.790 ;
        RECT 3539.350 4375.890 3539.630 4376.170 ;
        RECT 3539.350 4375.270 3539.630 4375.550 ;
        RECT 3539.350 4374.650 3539.630 4374.930 ;
        RECT 3539.350 4374.030 3539.630 4374.310 ;
        RECT 350.370 4373.410 350.650 4373.690 ;
        RECT 350.370 4372.790 350.650 4373.070 ;
        RECT 350.370 4372.170 350.650 4372.450 ;
        RECT 350.370 4371.550 350.650 4371.830 ;
        RECT 350.370 4370.930 350.650 4371.210 ;
        RECT 3539.350 4373.410 3539.630 4373.690 ;
        RECT 3539.350 4372.790 3539.630 4373.070 ;
        RECT 3539.350 4372.170 3539.630 4372.450 ;
        RECT 3539.350 4371.550 3539.630 4371.830 ;
        RECT 3539.350 4370.930 3539.630 4371.210 ;
        RECT 350.370 4370.310 350.650 4370.590 ;
        RECT 350.370 4369.690 350.650 4369.970 ;
        RECT 350.370 4369.070 350.650 4369.350 ;
        RECT 350.370 4368.450 350.650 4368.730 ;
        RECT 350.370 4367.830 350.650 4368.110 ;
        RECT 350.370 4367.210 350.650 4367.490 ;
        RECT 350.370 4366.590 350.650 4366.870 ;
        RECT 350.370 4365.970 350.650 4366.250 ;
        RECT 350.370 4365.350 350.650 4365.630 ;
        RECT 350.370 4364.730 350.650 4365.010 ;
        RECT 350.370 4364.110 350.650 4364.390 ;
        RECT 3539.350 4368.380 3539.630 4368.660 ;
        RECT 3539.350 4367.760 3539.630 4368.040 ;
        RECT 3539.350 4367.140 3539.630 4367.420 ;
        RECT 3539.350 4366.520 3539.630 4366.800 ;
        RECT 3539.350 4365.900 3539.630 4366.180 ;
        RECT 3539.350 4365.280 3539.630 4365.560 ;
        RECT 3539.350 4364.660 3539.630 4364.940 ;
        RECT 3539.350 4364.040 3539.630 4364.320 ;
        RECT 3539.350 4363.420 3539.630 4363.700 ;
        RECT 3539.350 4362.800 3539.630 4363.080 ;
        RECT 3539.350 4362.180 3539.630 4362.460 ;
        RECT 3539.350 4361.560 3539.630 4361.840 ;
        RECT 3539.350 4360.940 3539.630 4361.220 ;
        RECT 350.370 4360.390 350.650 4360.670 ;
        RECT 350.370 4359.770 350.650 4360.050 ;
        RECT 350.370 4359.150 350.650 4359.430 ;
        RECT 350.370 4358.530 350.650 4358.810 ;
        RECT 3539.350 4360.320 3539.630 4360.600 ;
        RECT 3539.350 4359.700 3539.630 4359.980 ;
        RECT 3539.350 4359.080 3539.630 4359.360 ;
        RECT 350.370 4357.910 350.650 4358.190 ;
        RECT 350.370 4357.290 350.650 4357.570 ;
        RECT 350.370 4356.670 350.650 4356.950 ;
        RECT 350.370 4356.050 350.650 4356.330 ;
        RECT 350.370 4355.430 350.650 4355.710 ;
        RECT 350.370 4354.810 350.650 4355.090 ;
        RECT 350.370 4354.190 350.650 4354.470 ;
        RECT 350.370 4353.570 350.650 4353.850 ;
        RECT 350.370 4352.950 350.650 4353.230 ;
        RECT 350.370 4352.330 350.650 4352.610 ;
        RECT 350.370 4351.710 350.650 4351.990 ;
        RECT 3539.350 4355.390 3539.630 4355.670 ;
        RECT 3539.350 4354.770 3539.630 4355.050 ;
        RECT 3539.350 4354.150 3539.630 4354.430 ;
        RECT 3539.350 4353.530 3539.630 4353.810 ;
        RECT 3539.350 4352.910 3539.630 4353.190 ;
        RECT 3539.350 4352.290 3539.630 4352.570 ;
        RECT 3539.350 4351.670 3539.630 4351.950 ;
        RECT 3539.350 4351.050 3539.630 4351.330 ;
        RECT 3539.350 4350.430 3539.630 4350.710 ;
        RECT 3539.350 4349.810 3539.630 4350.090 ;
        RECT 3539.350 4349.190 3539.630 4349.470 ;
        RECT 3539.350 4348.570 3539.630 4348.850 ;
        RECT 3539.350 4347.950 3539.630 4348.230 ;
        RECT 3539.350 4347.330 3539.630 4347.610 ;
        RECT 3539.350 4346.710 3539.630 4346.990 ;
        RECT 350.370 4218.010 350.650 4218.290 ;
        RECT 350.370 4217.390 350.650 4217.670 ;
        RECT 350.370 4216.770 350.650 4217.050 ;
        RECT 350.370 4216.150 350.650 4216.430 ;
        RECT 350.370 4215.530 350.650 4215.810 ;
        RECT 350.370 4214.910 350.650 4215.190 ;
        RECT 350.370 4214.290 350.650 4214.570 ;
        RECT 350.370 4213.670 350.650 4213.950 ;
        RECT 350.370 4213.050 350.650 4213.330 ;
        RECT 350.370 4212.430 350.650 4212.710 ;
        RECT 350.370 4211.810 350.650 4212.090 ;
        RECT 350.370 4211.190 350.650 4211.470 ;
        RECT 350.370 4210.570 350.650 4210.850 ;
        RECT 350.370 4209.950 350.650 4210.230 ;
        RECT 350.370 4209.330 350.650 4209.610 ;
        RECT 350.370 4205.640 350.650 4205.920 ;
        RECT 350.370 4205.020 350.650 4205.300 ;
        RECT 350.370 4204.400 350.650 4204.680 ;
        RECT 350.370 4203.780 350.650 4204.060 ;
        RECT 350.370 4203.160 350.650 4203.440 ;
        RECT 350.370 4202.540 350.650 4202.820 ;
        RECT 350.370 4201.920 350.650 4202.200 ;
        RECT 350.370 4201.300 350.650 4201.580 ;
        RECT 350.370 4200.680 350.650 4200.960 ;
        RECT 350.370 4200.060 350.650 4200.340 ;
        RECT 350.370 4199.440 350.650 4199.720 ;
        RECT 350.370 4198.820 350.650 4199.100 ;
        RECT 350.370 4198.200 350.650 4198.480 ;
        RECT 350.370 4197.580 350.650 4197.860 ;
        RECT 350.370 4196.960 350.650 4197.240 ;
        RECT 350.370 4196.340 350.650 4196.620 ;
        RECT 350.370 4193.790 350.650 4194.070 ;
        RECT 350.370 4193.170 350.650 4193.450 ;
        RECT 350.370 4192.550 350.650 4192.830 ;
        RECT 350.370 4191.930 350.650 4192.210 ;
        RECT 350.370 4191.310 350.650 4191.590 ;
        RECT 350.370 4190.690 350.650 4190.970 ;
        RECT 350.370 4190.070 350.650 4190.350 ;
        RECT 350.370 4189.450 350.650 4189.730 ;
        RECT 350.370 4188.830 350.650 4189.110 ;
        RECT 350.370 4188.210 350.650 4188.490 ;
        RECT 350.370 4187.590 350.650 4187.870 ;
        RECT 350.370 4186.970 350.650 4187.250 ;
        RECT 350.370 4186.350 350.650 4186.630 ;
        RECT 350.370 4185.730 350.650 4186.010 ;
        RECT 350.370 4185.110 350.650 4185.390 ;
        RECT 350.370 4184.490 350.650 4184.770 ;
        RECT 350.370 4180.260 350.650 4180.540 ;
        RECT 350.370 4179.640 350.650 4179.920 ;
        RECT 350.370 4179.020 350.650 4179.300 ;
        RECT 350.370 4178.400 350.650 4178.680 ;
        RECT 350.370 4177.780 350.650 4178.060 ;
        RECT 350.370 4177.160 350.650 4177.440 ;
        RECT 350.370 4176.540 350.650 4176.820 ;
        RECT 350.370 4175.920 350.650 4176.200 ;
        RECT 350.370 4175.300 350.650 4175.580 ;
        RECT 350.370 4174.680 350.650 4174.960 ;
        RECT 350.370 4174.060 350.650 4174.340 ;
        RECT 350.370 4173.440 350.650 4173.720 ;
        RECT 350.370 4172.820 350.650 4173.100 ;
        RECT 350.370 4172.200 350.650 4172.480 ;
        RECT 350.370 4171.580 350.650 4171.860 ;
        RECT 350.370 4170.960 350.650 4171.240 ;
        RECT 350.370 4168.410 350.650 4168.690 ;
        RECT 350.370 4167.790 350.650 4168.070 ;
        RECT 350.370 4167.170 350.650 4167.450 ;
        RECT 350.370 4166.550 350.650 4166.830 ;
        RECT 350.370 4165.930 350.650 4166.210 ;
        RECT 350.370 4165.310 350.650 4165.590 ;
        RECT 350.370 4164.690 350.650 4164.970 ;
        RECT 350.370 4164.070 350.650 4164.350 ;
        RECT 350.370 4163.450 350.650 4163.730 ;
        RECT 350.370 4162.830 350.650 4163.110 ;
        RECT 350.370 4162.210 350.650 4162.490 ;
        RECT 350.370 4161.590 350.650 4161.870 ;
        RECT 350.370 4160.970 350.650 4161.250 ;
        RECT 350.370 4160.350 350.650 4160.630 ;
        RECT 350.370 4159.730 350.650 4160.010 ;
        RECT 350.370 4159.110 350.650 4159.390 ;
        RECT 350.370 4155.390 350.650 4155.670 ;
        RECT 350.370 4154.770 350.650 4155.050 ;
        RECT 350.370 4154.150 350.650 4154.430 ;
        RECT 350.370 4153.530 350.650 4153.810 ;
        RECT 350.370 4152.910 350.650 4153.190 ;
        RECT 350.370 4152.290 350.650 4152.570 ;
        RECT 350.370 4151.670 350.650 4151.950 ;
        RECT 350.370 4151.050 350.650 4151.330 ;
        RECT 350.370 4150.430 350.650 4150.710 ;
        RECT 350.370 4149.810 350.650 4150.090 ;
        RECT 350.370 4149.190 350.650 4149.470 ;
        RECT 350.370 4148.570 350.650 4148.850 ;
        RECT 350.370 4147.950 350.650 4148.230 ;
        RECT 350.370 4147.330 350.650 4147.610 ;
        RECT 350.370 4146.710 350.650 4146.990 ;
        RECT 350.370 4013.010 350.650 4013.290 ;
        RECT 350.370 4012.390 350.650 4012.670 ;
        RECT 350.370 4011.770 350.650 4012.050 ;
        RECT 350.370 4011.150 350.650 4011.430 ;
        RECT 350.370 4010.530 350.650 4010.810 ;
        RECT 350.370 4009.910 350.650 4010.190 ;
        RECT 350.370 4009.290 350.650 4009.570 ;
        RECT 350.370 4008.670 350.650 4008.950 ;
        RECT 350.370 4008.050 350.650 4008.330 ;
        RECT 350.370 4007.430 350.650 4007.710 ;
        RECT 350.370 4006.810 350.650 4007.090 ;
        RECT 350.370 4006.190 350.650 4006.470 ;
        RECT 350.370 4005.570 350.650 4005.850 ;
        RECT 350.370 4004.950 350.650 4005.230 ;
        RECT 350.370 4004.330 350.650 4004.610 ;
        RECT 350.370 4000.640 350.650 4000.920 ;
        RECT 350.370 4000.020 350.650 4000.300 ;
        RECT 350.370 3999.400 350.650 3999.680 ;
        RECT 350.370 3998.780 350.650 3999.060 ;
        RECT 350.370 3998.160 350.650 3998.440 ;
        RECT 350.370 3997.540 350.650 3997.820 ;
        RECT 350.370 3996.920 350.650 3997.200 ;
        RECT 350.370 3996.300 350.650 3996.580 ;
        RECT 350.370 3995.680 350.650 3995.960 ;
        RECT 350.370 3995.060 350.650 3995.340 ;
        RECT 350.370 3994.440 350.650 3994.720 ;
        RECT 350.370 3993.820 350.650 3994.100 ;
        RECT 350.370 3993.200 350.650 3993.480 ;
        RECT 350.370 3992.580 350.650 3992.860 ;
        RECT 350.370 3991.960 350.650 3992.240 ;
        RECT 350.370 3991.340 350.650 3991.620 ;
        RECT 350.370 3988.790 350.650 3989.070 ;
        RECT 350.370 3988.170 350.650 3988.450 ;
        RECT 350.370 3987.550 350.650 3987.830 ;
        RECT 350.370 3986.930 350.650 3987.210 ;
        RECT 350.370 3986.310 350.650 3986.590 ;
        RECT 350.370 3985.690 350.650 3985.970 ;
        RECT 350.370 3985.070 350.650 3985.350 ;
        RECT 350.370 3984.450 350.650 3984.730 ;
        RECT 350.370 3983.830 350.650 3984.110 ;
        RECT 350.370 3983.210 350.650 3983.490 ;
        RECT 350.370 3982.590 350.650 3982.870 ;
        RECT 350.370 3981.970 350.650 3982.250 ;
        RECT 350.370 3981.350 350.650 3981.630 ;
        RECT 350.370 3980.730 350.650 3981.010 ;
        RECT 350.370 3980.110 350.650 3980.390 ;
        RECT 350.370 3979.490 350.650 3979.770 ;
        RECT 3539.350 3988.010 3539.630 3988.290 ;
        RECT 3539.350 3987.390 3539.630 3987.670 ;
        RECT 3539.350 3986.770 3539.630 3987.050 ;
        RECT 3539.350 3986.150 3539.630 3986.430 ;
        RECT 3539.350 3985.530 3539.630 3985.810 ;
        RECT 3539.350 3984.910 3539.630 3985.190 ;
        RECT 3539.350 3984.290 3539.630 3984.570 ;
        RECT 3539.350 3983.670 3539.630 3983.950 ;
        RECT 3539.350 3983.050 3539.630 3983.330 ;
        RECT 3539.350 3982.430 3539.630 3982.710 ;
        RECT 3539.350 3981.810 3539.630 3982.090 ;
        RECT 3539.350 3981.190 3539.630 3981.470 ;
        RECT 3539.350 3980.570 3539.630 3980.850 ;
        RECT 3539.350 3979.950 3539.630 3980.230 ;
        RECT 3539.350 3979.330 3539.630 3979.610 ;
        RECT 350.370 3975.260 350.650 3975.540 ;
        RECT 350.370 3974.640 350.650 3974.920 ;
        RECT 350.370 3974.020 350.650 3974.300 ;
        RECT 350.370 3973.400 350.650 3973.680 ;
        RECT 350.370 3972.780 350.650 3973.060 ;
        RECT 350.370 3972.160 350.650 3972.440 ;
        RECT 350.370 3971.540 350.650 3971.820 ;
        RECT 350.370 3970.920 350.650 3971.200 ;
        RECT 350.370 3970.300 350.650 3970.580 ;
        RECT 350.370 3969.680 350.650 3969.960 ;
        RECT 350.370 3969.060 350.650 3969.340 ;
        RECT 350.370 3968.440 350.650 3968.720 ;
        RECT 350.370 3967.820 350.650 3968.100 ;
        RECT 350.370 3967.200 350.650 3967.480 ;
        RECT 350.370 3966.580 350.650 3966.860 ;
        RECT 350.370 3965.960 350.650 3966.240 ;
        RECT 3539.350 3975.610 3539.630 3975.890 ;
        RECT 3539.350 3974.990 3539.630 3975.270 ;
        RECT 3539.350 3974.370 3539.630 3974.650 ;
        RECT 3539.350 3973.750 3539.630 3974.030 ;
        RECT 3539.350 3973.130 3539.630 3973.410 ;
        RECT 3539.350 3972.510 3539.630 3972.790 ;
        RECT 3539.350 3971.890 3539.630 3972.170 ;
        RECT 3539.350 3971.270 3539.630 3971.550 ;
        RECT 3539.350 3970.650 3539.630 3970.930 ;
        RECT 3539.350 3970.030 3539.630 3970.310 ;
        RECT 3539.350 3969.410 3539.630 3969.690 ;
        RECT 3539.350 3968.790 3539.630 3969.070 ;
        RECT 3539.350 3968.170 3539.630 3968.450 ;
        RECT 3539.350 3967.550 3539.630 3967.830 ;
        RECT 3539.350 3966.930 3539.630 3967.210 ;
        RECT 3539.350 3966.310 3539.630 3966.590 ;
        RECT 350.370 3963.410 350.650 3963.690 ;
        RECT 350.370 3962.790 350.650 3963.070 ;
        RECT 350.370 3962.170 350.650 3962.450 ;
        RECT 350.370 3961.550 350.650 3961.830 ;
        RECT 350.370 3960.930 350.650 3961.210 ;
        RECT 350.370 3960.310 350.650 3960.590 ;
        RECT 350.370 3959.690 350.650 3959.970 ;
        RECT 350.370 3959.070 350.650 3959.350 ;
        RECT 350.370 3958.450 350.650 3958.730 ;
        RECT 350.370 3957.830 350.650 3958.110 ;
        RECT 350.370 3957.210 350.650 3957.490 ;
        RECT 350.370 3956.590 350.650 3956.870 ;
        RECT 350.370 3955.970 350.650 3956.250 ;
        RECT 350.370 3955.350 350.650 3955.630 ;
        RECT 350.370 3954.730 350.650 3955.010 ;
        RECT 350.370 3954.110 350.650 3954.390 ;
        RECT 3539.350 3963.760 3539.630 3964.040 ;
        RECT 3539.350 3963.140 3539.630 3963.420 ;
        RECT 3539.350 3962.520 3539.630 3962.800 ;
        RECT 3539.350 3961.900 3539.630 3962.180 ;
        RECT 3539.350 3961.280 3539.630 3961.560 ;
        RECT 3539.350 3960.660 3539.630 3960.940 ;
        RECT 3539.350 3960.040 3539.630 3960.320 ;
        RECT 3539.350 3959.420 3539.630 3959.700 ;
        RECT 3539.350 3958.800 3539.630 3959.080 ;
        RECT 3539.350 3958.180 3539.630 3958.460 ;
        RECT 3539.350 3957.560 3539.630 3957.840 ;
        RECT 3539.350 3956.940 3539.630 3957.220 ;
        RECT 3539.350 3956.320 3539.630 3956.600 ;
        RECT 3539.350 3955.700 3539.630 3955.980 ;
        RECT 3539.350 3955.080 3539.630 3955.360 ;
        RECT 3539.350 3954.460 3539.630 3954.740 ;
        RECT 350.370 3950.390 350.650 3950.670 ;
        RECT 350.370 3949.770 350.650 3950.050 ;
        RECT 350.370 3949.150 350.650 3949.430 ;
        RECT 350.370 3948.530 350.650 3948.810 ;
        RECT 350.370 3947.910 350.650 3948.190 ;
        RECT 350.370 3947.290 350.650 3947.570 ;
        RECT 350.370 3946.670 350.650 3946.950 ;
        RECT 350.370 3946.050 350.650 3946.330 ;
        RECT 350.370 3945.430 350.650 3945.710 ;
        RECT 350.370 3944.810 350.650 3945.090 ;
        RECT 350.370 3944.190 350.650 3944.470 ;
        RECT 350.370 3943.570 350.650 3943.850 ;
        RECT 350.370 3942.950 350.650 3943.230 ;
        RECT 350.370 3942.330 350.650 3942.610 ;
        RECT 350.370 3941.710 350.650 3941.990 ;
        RECT 3539.350 3950.230 3539.630 3950.510 ;
        RECT 3539.350 3949.610 3539.630 3949.890 ;
        RECT 3539.350 3948.990 3539.630 3949.270 ;
        RECT 3539.350 3948.370 3539.630 3948.650 ;
        RECT 3539.350 3947.750 3539.630 3948.030 ;
        RECT 3539.350 3947.130 3539.630 3947.410 ;
        RECT 3539.350 3946.510 3539.630 3946.790 ;
        RECT 3539.350 3945.890 3539.630 3946.170 ;
        RECT 3539.350 3945.270 3539.630 3945.550 ;
        RECT 3539.350 3944.650 3539.630 3944.930 ;
        RECT 3539.350 3944.030 3539.630 3944.310 ;
        RECT 3539.350 3943.410 3539.630 3943.690 ;
        RECT 3539.350 3942.790 3539.630 3943.070 ;
        RECT 3539.350 3942.170 3539.630 3942.450 ;
        RECT 3539.350 3941.550 3539.630 3941.830 ;
        RECT 3539.350 3940.930 3539.630 3941.210 ;
        RECT 3539.350 3938.380 3539.630 3938.660 ;
        RECT 3539.350 3937.760 3539.630 3938.040 ;
        RECT 3539.350 3937.140 3539.630 3937.420 ;
        RECT 3539.350 3936.520 3539.630 3936.800 ;
        RECT 3539.350 3935.900 3539.630 3936.180 ;
        RECT 3539.350 3935.280 3539.630 3935.560 ;
        RECT 3539.350 3934.660 3539.630 3934.940 ;
        RECT 3539.350 3934.040 3539.630 3934.320 ;
        RECT 3539.350 3933.420 3539.630 3933.700 ;
        RECT 3539.350 3932.800 3539.630 3933.080 ;
        RECT 3539.350 3932.180 3539.630 3932.460 ;
        RECT 3539.350 3931.560 3539.630 3931.840 ;
        RECT 3539.350 3930.940 3539.630 3931.220 ;
        RECT 3539.350 3930.320 3539.630 3930.600 ;
        RECT 3539.350 3929.700 3539.630 3929.980 ;
        RECT 3539.350 3929.080 3539.630 3929.360 ;
        RECT 3539.350 3925.390 3539.630 3925.670 ;
        RECT 3539.350 3924.770 3539.630 3925.050 ;
        RECT 3539.350 3924.150 3539.630 3924.430 ;
        RECT 3539.350 3923.530 3539.630 3923.810 ;
        RECT 3539.350 3922.910 3539.630 3923.190 ;
        RECT 3539.350 3922.290 3539.630 3922.570 ;
        RECT 3539.350 3921.670 3539.630 3921.950 ;
        RECT 3539.350 3921.050 3539.630 3921.330 ;
        RECT 3539.350 3920.430 3539.630 3920.710 ;
        RECT 3539.350 3919.810 3539.630 3920.090 ;
        RECT 3539.350 3919.190 3539.630 3919.470 ;
        RECT 3539.350 3918.570 3539.630 3918.850 ;
        RECT 3539.350 3917.950 3539.630 3918.230 ;
        RECT 3539.350 3917.330 3539.630 3917.610 ;
        RECT 3539.350 3916.710 3539.630 3916.990 ;
        RECT 3539.350 2483.010 3539.630 2483.290 ;
        RECT 3539.350 2482.390 3539.630 2482.670 ;
        RECT 3539.350 2481.770 3539.630 2482.050 ;
        RECT 3539.350 2481.150 3539.630 2481.430 ;
        RECT 3539.350 2480.530 3539.630 2480.810 ;
        RECT 3539.350 2479.910 3539.630 2480.190 ;
        RECT 3539.350 2479.290 3539.630 2479.570 ;
        RECT 3539.350 2478.670 3539.630 2478.950 ;
        RECT 3539.350 2478.050 3539.630 2478.330 ;
        RECT 3539.350 2477.430 3539.630 2477.710 ;
        RECT 3539.350 2476.810 3539.630 2477.090 ;
        RECT 3539.350 2476.190 3539.630 2476.470 ;
        RECT 3539.350 2475.570 3539.630 2475.850 ;
        RECT 3539.350 2474.950 3539.630 2475.230 ;
        RECT 3539.350 2474.330 3539.630 2474.610 ;
        RECT 3539.350 2470.610 3539.630 2470.890 ;
        RECT 3539.350 2469.990 3539.630 2470.270 ;
        RECT 3539.350 2469.370 3539.630 2469.650 ;
        RECT 3539.350 2468.750 3539.630 2469.030 ;
        RECT 3539.350 2468.130 3539.630 2468.410 ;
        RECT 3539.350 2467.510 3539.630 2467.790 ;
        RECT 3539.350 2466.890 3539.630 2467.170 ;
        RECT 3539.350 2466.270 3539.630 2466.550 ;
        RECT 3539.350 2465.650 3539.630 2465.930 ;
        RECT 3539.350 2465.030 3539.630 2465.310 ;
        RECT 3539.350 2464.410 3539.630 2464.690 ;
        RECT 3539.350 2463.790 3539.630 2464.070 ;
        RECT 3539.350 2463.170 3539.630 2463.450 ;
        RECT 3539.350 2462.550 3539.630 2462.830 ;
        RECT 3539.350 2461.930 3539.630 2462.210 ;
        RECT 3539.350 2461.310 3539.630 2461.590 ;
        RECT 3539.350 2458.760 3539.630 2459.040 ;
        RECT 3539.350 2458.140 3539.630 2458.420 ;
        RECT 3539.350 2457.520 3539.630 2457.800 ;
        RECT 3539.350 2456.900 3539.630 2457.180 ;
        RECT 3539.350 2456.280 3539.630 2456.560 ;
        RECT 3539.350 2455.660 3539.630 2455.940 ;
        RECT 3539.350 2455.040 3539.630 2455.320 ;
        RECT 3539.350 2454.420 3539.630 2454.700 ;
        RECT 3539.350 2453.800 3539.630 2454.080 ;
        RECT 3539.350 2453.180 3539.630 2453.460 ;
        RECT 3539.350 2452.560 3539.630 2452.840 ;
        RECT 3539.350 2451.940 3539.630 2452.220 ;
        RECT 3539.350 2451.320 3539.630 2451.600 ;
        RECT 3539.350 2450.700 3539.630 2450.980 ;
        RECT 3539.350 2450.080 3539.630 2450.360 ;
        RECT 3539.350 2449.460 3539.630 2449.740 ;
        RECT 3539.350 2445.230 3539.630 2445.510 ;
        RECT 3539.350 2444.610 3539.630 2444.890 ;
        RECT 3539.350 2443.990 3539.630 2444.270 ;
        RECT 3539.350 2443.370 3539.630 2443.650 ;
        RECT 3539.350 2442.750 3539.630 2443.030 ;
        RECT 3539.350 2442.130 3539.630 2442.410 ;
        RECT 3539.350 2441.510 3539.630 2441.790 ;
        RECT 3539.350 2440.890 3539.630 2441.170 ;
        RECT 3539.350 2440.270 3539.630 2440.550 ;
        RECT 3539.350 2439.650 3539.630 2439.930 ;
        RECT 3539.350 2439.030 3539.630 2439.310 ;
        RECT 3539.350 2438.410 3539.630 2438.690 ;
        RECT 3539.350 2437.790 3539.630 2438.070 ;
        RECT 3539.350 2437.170 3539.630 2437.450 ;
        RECT 3539.350 2436.550 3539.630 2436.830 ;
        RECT 3539.350 2435.930 3539.630 2436.210 ;
        RECT 3539.350 2433.380 3539.630 2433.660 ;
        RECT 3539.350 2432.760 3539.630 2433.040 ;
        RECT 3539.350 2432.140 3539.630 2432.420 ;
        RECT 3539.350 2431.520 3539.630 2431.800 ;
        RECT 3539.350 2430.900 3539.630 2431.180 ;
        RECT 3539.350 2430.280 3539.630 2430.560 ;
        RECT 3539.350 2429.660 3539.630 2429.940 ;
        RECT 3539.350 2429.040 3539.630 2429.320 ;
        RECT 3539.350 2428.420 3539.630 2428.700 ;
        RECT 3539.350 2427.800 3539.630 2428.080 ;
        RECT 3539.350 2427.180 3539.630 2427.460 ;
        RECT 3539.350 2426.560 3539.630 2426.840 ;
        RECT 3539.350 2425.940 3539.630 2426.220 ;
        RECT 3539.350 2425.320 3539.630 2425.600 ;
        RECT 3539.350 2424.700 3539.630 2424.980 ;
        RECT 3539.350 2424.080 3539.630 2424.360 ;
        RECT 3539.350 2420.390 3539.630 2420.670 ;
        RECT 3539.350 2419.770 3539.630 2420.050 ;
        RECT 3539.350 2419.150 3539.630 2419.430 ;
        RECT 3539.350 2418.530 3539.630 2418.810 ;
        RECT 3539.350 2417.910 3539.630 2418.190 ;
        RECT 3539.350 2417.290 3539.630 2417.570 ;
        RECT 3539.350 2416.670 3539.630 2416.950 ;
        RECT 3539.350 2416.050 3539.630 2416.330 ;
        RECT 3539.350 2415.430 3539.630 2415.710 ;
        RECT 3539.350 2414.810 3539.630 2415.090 ;
        RECT 3539.350 2414.190 3539.630 2414.470 ;
        RECT 3539.350 2413.570 3539.630 2413.850 ;
        RECT 3539.350 2412.950 3539.630 2413.230 ;
        RECT 3539.350 2412.330 3539.630 2412.610 ;
        RECT 3539.350 2411.710 3539.630 2411.990 ;
        RECT 350.370 2373.010 350.650 2373.290 ;
        RECT 350.370 2372.390 350.650 2372.670 ;
        RECT 350.370 2371.770 350.650 2372.050 ;
        RECT 350.370 2371.150 350.650 2371.430 ;
        RECT 350.370 2370.530 350.650 2370.810 ;
        RECT 350.370 2369.910 350.650 2370.190 ;
        RECT 350.370 2369.290 350.650 2369.570 ;
        RECT 350.370 2368.670 350.650 2368.950 ;
        RECT 350.370 2368.050 350.650 2368.330 ;
        RECT 350.370 2367.430 350.650 2367.710 ;
        RECT 350.370 2366.810 350.650 2367.090 ;
        RECT 350.370 2366.190 350.650 2366.470 ;
        RECT 350.370 2365.570 350.650 2365.850 ;
        RECT 350.370 2364.950 350.650 2365.230 ;
        RECT 350.370 2364.330 350.650 2364.610 ;
        RECT 350.370 2360.640 350.650 2360.920 ;
        RECT 350.370 2360.020 350.650 2360.300 ;
        RECT 350.370 2359.400 350.650 2359.680 ;
        RECT 350.370 2358.780 350.650 2359.060 ;
        RECT 350.370 2358.160 350.650 2358.440 ;
        RECT 350.370 2357.540 350.650 2357.820 ;
        RECT 350.370 2356.920 350.650 2357.200 ;
        RECT 350.370 2356.300 350.650 2356.580 ;
        RECT 350.370 2355.680 350.650 2355.960 ;
        RECT 350.370 2355.060 350.650 2355.340 ;
        RECT 350.370 2354.440 350.650 2354.720 ;
        RECT 350.370 2353.820 350.650 2354.100 ;
        RECT 350.370 2353.200 350.650 2353.480 ;
        RECT 350.370 2352.580 350.650 2352.860 ;
        RECT 350.370 2351.960 350.650 2352.240 ;
        RECT 350.370 2351.340 350.650 2351.620 ;
        RECT 350.370 2348.790 350.650 2349.070 ;
        RECT 350.370 2348.170 350.650 2348.450 ;
        RECT 350.370 2347.550 350.650 2347.830 ;
        RECT 350.370 2346.930 350.650 2347.210 ;
        RECT 350.370 2346.310 350.650 2346.590 ;
        RECT 350.370 2345.690 350.650 2345.970 ;
        RECT 350.370 2345.070 350.650 2345.350 ;
        RECT 350.370 2344.450 350.650 2344.730 ;
        RECT 350.370 2343.830 350.650 2344.110 ;
        RECT 350.370 2343.210 350.650 2343.490 ;
        RECT 350.370 2342.590 350.650 2342.870 ;
        RECT 350.370 2341.970 350.650 2342.250 ;
        RECT 350.370 2341.350 350.650 2341.630 ;
        RECT 350.370 2340.730 350.650 2341.010 ;
        RECT 350.370 2340.110 350.650 2340.390 ;
        RECT 350.370 2339.490 350.650 2339.770 ;
        RECT 350.370 2335.260 350.650 2335.540 ;
        RECT 350.370 2334.640 350.650 2334.920 ;
        RECT 350.370 2334.020 350.650 2334.300 ;
        RECT 350.370 2333.400 350.650 2333.680 ;
        RECT 350.370 2332.780 350.650 2333.060 ;
        RECT 350.370 2332.160 350.650 2332.440 ;
        RECT 350.370 2331.540 350.650 2331.820 ;
        RECT 350.370 2330.920 350.650 2331.200 ;
        RECT 350.370 2330.300 350.650 2330.580 ;
        RECT 350.370 2329.680 350.650 2329.960 ;
        RECT 350.370 2329.060 350.650 2329.340 ;
        RECT 350.370 2328.440 350.650 2328.720 ;
        RECT 350.370 2327.820 350.650 2328.100 ;
        RECT 350.370 2327.200 350.650 2327.480 ;
        RECT 350.370 2326.580 350.650 2326.860 ;
        RECT 350.370 2325.960 350.650 2326.240 ;
        RECT 350.370 2323.410 350.650 2323.690 ;
        RECT 350.370 2322.790 350.650 2323.070 ;
        RECT 350.370 2322.170 350.650 2322.450 ;
        RECT 350.370 2321.550 350.650 2321.830 ;
        RECT 350.370 2320.930 350.650 2321.210 ;
        RECT 350.370 2320.310 350.650 2320.590 ;
        RECT 350.370 2319.690 350.650 2319.970 ;
        RECT 350.370 2319.070 350.650 2319.350 ;
        RECT 350.370 2318.450 350.650 2318.730 ;
        RECT 350.370 2317.830 350.650 2318.110 ;
        RECT 350.370 2317.210 350.650 2317.490 ;
        RECT 350.370 2316.590 350.650 2316.870 ;
        RECT 350.370 2315.970 350.650 2316.250 ;
        RECT 350.370 2315.350 350.650 2315.630 ;
        RECT 350.370 2314.730 350.650 2315.010 ;
        RECT 350.370 2314.110 350.650 2314.390 ;
        RECT 350.370 2310.390 350.650 2310.670 ;
        RECT 350.370 2309.770 350.650 2310.050 ;
        RECT 350.370 2309.150 350.650 2309.430 ;
        RECT 350.370 2308.530 350.650 2308.810 ;
        RECT 350.370 2307.910 350.650 2308.190 ;
        RECT 350.370 2307.290 350.650 2307.570 ;
        RECT 350.370 2306.670 350.650 2306.950 ;
        RECT 350.370 2306.050 350.650 2306.330 ;
        RECT 350.370 2305.430 350.650 2305.710 ;
        RECT 350.370 2304.810 350.650 2305.090 ;
        RECT 350.370 2304.190 350.650 2304.470 ;
        RECT 350.370 2303.570 350.650 2303.850 ;
        RECT 350.370 2302.950 350.650 2303.230 ;
        RECT 350.370 2302.330 350.650 2302.610 ;
        RECT 350.370 2301.710 350.650 2301.990 ;
        RECT 3539.350 2268.010 3539.630 2268.290 ;
        RECT 3539.350 2267.390 3539.630 2267.670 ;
        RECT 3539.350 2266.770 3539.630 2267.050 ;
        RECT 3539.350 2266.150 3539.630 2266.430 ;
        RECT 3539.350 2265.530 3539.630 2265.810 ;
        RECT 3539.350 2264.910 3539.630 2265.190 ;
        RECT 3539.350 2264.290 3539.630 2264.570 ;
        RECT 3539.350 2263.670 3539.630 2263.950 ;
        RECT 3539.350 2263.050 3539.630 2263.330 ;
        RECT 3539.350 2262.430 3539.630 2262.710 ;
        RECT 3539.350 2261.810 3539.630 2262.090 ;
        RECT 3539.350 2261.190 3539.630 2261.470 ;
        RECT 3539.350 2260.570 3539.630 2260.850 ;
        RECT 3539.350 2259.950 3539.630 2260.230 ;
        RECT 3539.350 2259.330 3539.630 2259.610 ;
        RECT 3539.350 2255.610 3539.630 2255.890 ;
        RECT 3539.350 2254.990 3539.630 2255.270 ;
        RECT 3539.350 2254.370 3539.630 2254.650 ;
        RECT 3539.350 2253.750 3539.630 2254.030 ;
        RECT 3539.350 2253.130 3539.630 2253.410 ;
        RECT 3539.350 2252.510 3539.630 2252.790 ;
        RECT 3539.350 2251.890 3539.630 2252.170 ;
        RECT 3539.350 2251.270 3539.630 2251.550 ;
        RECT 3539.350 2250.650 3539.630 2250.930 ;
        RECT 3539.350 2250.030 3539.630 2250.310 ;
        RECT 3539.350 2249.410 3539.630 2249.690 ;
        RECT 3539.350 2248.790 3539.630 2249.070 ;
        RECT 3539.350 2248.170 3539.630 2248.450 ;
        RECT 3539.350 2247.550 3539.630 2247.830 ;
        RECT 3539.350 2246.930 3539.630 2247.210 ;
        RECT 3539.350 2246.310 3539.630 2246.590 ;
        RECT 3539.350 2243.760 3539.630 2244.040 ;
        RECT 3539.350 2243.140 3539.630 2243.420 ;
        RECT 3539.350 2242.520 3539.630 2242.800 ;
        RECT 3539.350 2241.900 3539.630 2242.180 ;
        RECT 3539.350 2241.280 3539.630 2241.560 ;
        RECT 3539.350 2240.660 3539.630 2240.940 ;
        RECT 3539.350 2240.040 3539.630 2240.320 ;
        RECT 3539.350 2239.420 3539.630 2239.700 ;
        RECT 3539.350 2238.800 3539.630 2239.080 ;
        RECT 3539.350 2238.180 3539.630 2238.460 ;
        RECT 3539.350 2237.560 3539.630 2237.840 ;
        RECT 3539.350 2236.940 3539.630 2237.220 ;
        RECT 3539.350 2236.320 3539.630 2236.600 ;
        RECT 3539.350 2235.700 3539.630 2235.980 ;
        RECT 3539.350 2235.080 3539.630 2235.360 ;
        RECT 3539.350 2234.460 3539.630 2234.740 ;
        RECT 3539.350 2230.230 3539.630 2230.510 ;
        RECT 3539.350 2229.610 3539.630 2229.890 ;
        RECT 3539.350 2228.990 3539.630 2229.270 ;
        RECT 3539.350 2228.370 3539.630 2228.650 ;
        RECT 3539.350 2227.750 3539.630 2228.030 ;
        RECT 3539.350 2227.130 3539.630 2227.410 ;
        RECT 3539.350 2226.510 3539.630 2226.790 ;
        RECT 3539.350 2225.890 3539.630 2226.170 ;
        RECT 3539.350 2225.270 3539.630 2225.550 ;
        RECT 3539.350 2224.650 3539.630 2224.930 ;
        RECT 3539.350 2224.030 3539.630 2224.310 ;
        RECT 3539.350 2223.410 3539.630 2223.690 ;
        RECT 3539.350 2222.790 3539.630 2223.070 ;
        RECT 3539.350 2222.170 3539.630 2222.450 ;
        RECT 3539.350 2221.550 3539.630 2221.830 ;
        RECT 3539.350 2220.930 3539.630 2221.210 ;
        RECT 3539.350 2218.380 3539.630 2218.660 ;
        RECT 3539.350 2217.760 3539.630 2218.040 ;
        RECT 3539.350 2217.140 3539.630 2217.420 ;
        RECT 3539.350 2216.520 3539.630 2216.800 ;
        RECT 3539.350 2215.900 3539.630 2216.180 ;
        RECT 3539.350 2215.280 3539.630 2215.560 ;
        RECT 3539.350 2214.660 3539.630 2214.940 ;
        RECT 3539.350 2214.040 3539.630 2214.320 ;
        RECT 3539.350 2213.420 3539.630 2213.700 ;
        RECT 3539.350 2212.800 3539.630 2213.080 ;
        RECT 3539.350 2212.180 3539.630 2212.460 ;
        RECT 3539.350 2211.560 3539.630 2211.840 ;
        RECT 3539.350 2210.940 3539.630 2211.220 ;
        RECT 3539.350 2210.320 3539.630 2210.600 ;
        RECT 3539.350 2209.700 3539.630 2209.980 ;
        RECT 3539.350 2209.080 3539.630 2209.360 ;
        RECT 3539.350 2205.390 3539.630 2205.670 ;
        RECT 3539.350 2204.770 3539.630 2205.050 ;
        RECT 3539.350 2204.150 3539.630 2204.430 ;
        RECT 3539.350 2203.530 3539.630 2203.810 ;
        RECT 3539.350 2202.910 3539.630 2203.190 ;
        RECT 3539.350 2202.290 3539.630 2202.570 ;
        RECT 3539.350 2201.670 3539.630 2201.950 ;
        RECT 3539.350 2201.050 3539.630 2201.330 ;
        RECT 3539.350 2200.430 3539.630 2200.710 ;
        RECT 3539.350 2199.810 3539.630 2200.090 ;
        RECT 3539.350 2199.190 3539.630 2199.470 ;
        RECT 3539.350 2198.570 3539.630 2198.850 ;
        RECT 3539.350 2197.950 3539.630 2198.230 ;
        RECT 3539.350 2197.330 3539.630 2197.610 ;
        RECT 3539.350 2196.710 3539.630 2196.990 ;
        RECT 350.370 2168.010 350.650 2168.290 ;
        RECT 350.370 2167.390 350.650 2167.670 ;
        RECT 350.370 2166.770 350.650 2167.050 ;
        RECT 350.370 2166.150 350.650 2166.430 ;
        RECT 350.370 2165.530 350.650 2165.810 ;
        RECT 350.370 2164.910 350.650 2165.190 ;
        RECT 350.370 2164.290 350.650 2164.570 ;
        RECT 350.370 2163.670 350.650 2163.950 ;
        RECT 350.370 2163.050 350.650 2163.330 ;
        RECT 350.370 2162.430 350.650 2162.710 ;
        RECT 350.370 2161.810 350.650 2162.090 ;
        RECT 350.370 2161.190 350.650 2161.470 ;
        RECT 350.370 2160.570 350.650 2160.850 ;
        RECT 350.370 2159.950 350.650 2160.230 ;
        RECT 350.370 2159.330 350.650 2159.610 ;
        RECT 350.370 2155.640 350.650 2155.920 ;
        RECT 350.370 2155.020 350.650 2155.300 ;
        RECT 350.370 2154.400 350.650 2154.680 ;
        RECT 350.370 2153.780 350.650 2154.060 ;
        RECT 350.370 2153.160 350.650 2153.440 ;
        RECT 350.370 2152.540 350.650 2152.820 ;
        RECT 350.370 2151.920 350.650 2152.200 ;
        RECT 350.370 2151.300 350.650 2151.580 ;
        RECT 350.370 2150.680 350.650 2150.960 ;
        RECT 350.370 2150.060 350.650 2150.340 ;
        RECT 350.370 2149.440 350.650 2149.720 ;
        RECT 350.370 2148.820 350.650 2149.100 ;
        RECT 350.370 2148.200 350.650 2148.480 ;
        RECT 350.370 2147.580 350.650 2147.860 ;
        RECT 350.370 2146.960 350.650 2147.240 ;
        RECT 350.370 2146.340 350.650 2146.620 ;
        RECT 350.370 2143.790 350.650 2144.070 ;
        RECT 350.370 2143.170 350.650 2143.450 ;
        RECT 350.370 2142.550 350.650 2142.830 ;
        RECT 350.370 2141.930 350.650 2142.210 ;
        RECT 350.370 2141.310 350.650 2141.590 ;
        RECT 350.370 2140.690 350.650 2140.970 ;
        RECT 350.370 2140.070 350.650 2140.350 ;
        RECT 350.370 2139.450 350.650 2139.730 ;
        RECT 350.370 2138.830 350.650 2139.110 ;
        RECT 350.370 2138.210 350.650 2138.490 ;
        RECT 350.370 2137.590 350.650 2137.870 ;
        RECT 350.370 2136.970 350.650 2137.250 ;
        RECT 350.370 2136.350 350.650 2136.630 ;
        RECT 350.370 2135.730 350.650 2136.010 ;
        RECT 350.370 2135.110 350.650 2135.390 ;
        RECT 350.370 2134.490 350.650 2134.770 ;
        RECT 350.370 2130.260 350.650 2130.540 ;
        RECT 350.370 2129.640 350.650 2129.920 ;
        RECT 350.370 2129.020 350.650 2129.300 ;
        RECT 350.370 2128.400 350.650 2128.680 ;
        RECT 350.370 2127.780 350.650 2128.060 ;
        RECT 350.370 2127.160 350.650 2127.440 ;
        RECT 350.370 2126.540 350.650 2126.820 ;
        RECT 350.370 2125.920 350.650 2126.200 ;
        RECT 350.370 2125.300 350.650 2125.580 ;
        RECT 350.370 2124.680 350.650 2124.960 ;
        RECT 350.370 2124.060 350.650 2124.340 ;
        RECT 350.370 2123.440 350.650 2123.720 ;
        RECT 350.370 2122.820 350.650 2123.100 ;
        RECT 350.370 2122.200 350.650 2122.480 ;
        RECT 350.370 2121.580 350.650 2121.860 ;
        RECT 350.370 2120.960 350.650 2121.240 ;
        RECT 350.370 2118.410 350.650 2118.690 ;
        RECT 350.370 2117.790 350.650 2118.070 ;
        RECT 350.370 2117.170 350.650 2117.450 ;
        RECT 350.370 2116.550 350.650 2116.830 ;
        RECT 350.370 2115.930 350.650 2116.210 ;
        RECT 350.370 2115.310 350.650 2115.590 ;
        RECT 350.370 2114.690 350.650 2114.970 ;
        RECT 350.370 2114.070 350.650 2114.350 ;
        RECT 350.370 2113.450 350.650 2113.730 ;
        RECT 350.370 2112.830 350.650 2113.110 ;
        RECT 350.370 2112.210 350.650 2112.490 ;
        RECT 350.370 2111.590 350.650 2111.870 ;
        RECT 350.370 2110.970 350.650 2111.250 ;
        RECT 350.370 2110.350 350.650 2110.630 ;
        RECT 350.370 2109.730 350.650 2110.010 ;
        RECT 350.370 2109.110 350.650 2109.390 ;
        RECT 350.370 2105.390 350.650 2105.670 ;
        RECT 350.370 2104.770 350.650 2105.050 ;
        RECT 350.370 2104.150 350.650 2104.430 ;
        RECT 350.370 2103.530 350.650 2103.810 ;
        RECT 350.370 2102.910 350.650 2103.190 ;
        RECT 350.370 2102.290 350.650 2102.570 ;
        RECT 350.370 2101.670 350.650 2101.950 ;
        RECT 350.370 2101.050 350.650 2101.330 ;
        RECT 350.370 2100.430 350.650 2100.710 ;
        RECT 350.370 2099.810 350.650 2100.090 ;
        RECT 350.370 2099.190 350.650 2099.470 ;
        RECT 350.370 2098.570 350.650 2098.850 ;
        RECT 350.370 2097.950 350.650 2098.230 ;
        RECT 350.370 2097.330 350.650 2097.610 ;
        RECT 350.370 2096.710 350.650 2096.990 ;
        RECT 3539.350 2053.010 3539.630 2053.290 ;
        RECT 3539.350 2052.390 3539.630 2052.670 ;
        RECT 3539.350 2051.770 3539.630 2052.050 ;
        RECT 3539.350 2051.150 3539.630 2051.430 ;
        RECT 3539.350 2050.530 3539.630 2050.810 ;
        RECT 3539.350 2049.910 3539.630 2050.190 ;
        RECT 3539.350 2049.290 3539.630 2049.570 ;
        RECT 3539.350 2048.670 3539.630 2048.950 ;
        RECT 3539.350 2048.050 3539.630 2048.330 ;
        RECT 3539.350 2047.430 3539.630 2047.710 ;
        RECT 3539.350 2046.810 3539.630 2047.090 ;
        RECT 3539.350 2046.190 3539.630 2046.470 ;
        RECT 3539.350 2045.570 3539.630 2045.850 ;
        RECT 3539.350 2044.950 3539.630 2045.230 ;
        RECT 3539.350 2044.330 3539.630 2044.610 ;
        RECT 3539.350 2040.610 3539.630 2040.890 ;
        RECT 3539.350 2039.990 3539.630 2040.270 ;
        RECT 3539.350 2039.370 3539.630 2039.650 ;
        RECT 3539.350 2038.750 3539.630 2039.030 ;
        RECT 3539.350 2038.130 3539.630 2038.410 ;
        RECT 3539.350 2037.510 3539.630 2037.790 ;
        RECT 3539.350 2036.890 3539.630 2037.170 ;
        RECT 3539.350 2036.270 3539.630 2036.550 ;
        RECT 3539.350 2035.650 3539.630 2035.930 ;
        RECT 3539.350 2035.030 3539.630 2035.310 ;
        RECT 3539.350 2034.410 3539.630 2034.690 ;
        RECT 3539.350 2033.790 3539.630 2034.070 ;
        RECT 3539.350 2033.170 3539.630 2033.450 ;
        RECT 3539.350 2032.550 3539.630 2032.830 ;
        RECT 3539.350 2031.930 3539.630 2032.210 ;
        RECT 3539.350 2031.310 3539.630 2031.590 ;
        RECT 3539.350 2028.760 3539.630 2029.040 ;
        RECT 3539.350 2028.140 3539.630 2028.420 ;
        RECT 3539.350 2027.520 3539.630 2027.800 ;
        RECT 3539.350 2026.900 3539.630 2027.180 ;
        RECT 3539.350 2026.280 3539.630 2026.560 ;
        RECT 3539.350 2025.660 3539.630 2025.940 ;
        RECT 3539.350 2025.040 3539.630 2025.320 ;
        RECT 3539.350 2024.420 3539.630 2024.700 ;
        RECT 3539.350 2023.800 3539.630 2024.080 ;
        RECT 3539.350 2023.180 3539.630 2023.460 ;
        RECT 3539.350 2022.560 3539.630 2022.840 ;
        RECT 3539.350 2021.940 3539.630 2022.220 ;
        RECT 3539.350 2021.320 3539.630 2021.600 ;
        RECT 3539.350 2020.700 3539.630 2020.980 ;
        RECT 3539.350 2020.080 3539.630 2020.360 ;
        RECT 3539.350 2019.460 3539.630 2019.740 ;
        RECT 3539.350 2015.230 3539.630 2015.510 ;
        RECT 3539.350 2014.610 3539.630 2014.890 ;
        RECT 3539.350 2013.990 3539.630 2014.270 ;
        RECT 3539.350 2013.370 3539.630 2013.650 ;
        RECT 3539.350 2012.750 3539.630 2013.030 ;
        RECT 3539.350 2012.130 3539.630 2012.410 ;
        RECT 3539.350 2011.510 3539.630 2011.790 ;
        RECT 3539.350 2010.890 3539.630 2011.170 ;
        RECT 3539.350 2010.270 3539.630 2010.550 ;
        RECT 3539.350 2009.650 3539.630 2009.930 ;
        RECT 3539.350 2009.030 3539.630 2009.310 ;
        RECT 3539.350 2008.410 3539.630 2008.690 ;
        RECT 3539.350 2007.790 3539.630 2008.070 ;
        RECT 3539.350 2007.170 3539.630 2007.450 ;
        RECT 3539.350 2006.550 3539.630 2006.830 ;
        RECT 3539.350 2005.930 3539.630 2006.210 ;
        RECT 3539.350 2003.380 3539.630 2003.660 ;
        RECT 3539.350 2002.760 3539.630 2003.040 ;
        RECT 3539.350 2002.140 3539.630 2002.420 ;
        RECT 3539.350 2001.520 3539.630 2001.800 ;
        RECT 3539.350 2000.900 3539.630 2001.180 ;
        RECT 3539.350 2000.280 3539.630 2000.560 ;
        RECT 3539.350 1999.660 3539.630 1999.940 ;
        RECT 3539.350 1999.040 3539.630 1999.320 ;
        RECT 3539.350 1998.420 3539.630 1998.700 ;
        RECT 3539.350 1997.800 3539.630 1998.080 ;
        RECT 3539.350 1997.180 3539.630 1997.460 ;
        RECT 3539.350 1996.560 3539.630 1996.840 ;
        RECT 3539.350 1995.940 3539.630 1996.220 ;
        RECT 3539.350 1995.320 3539.630 1995.600 ;
        RECT 3539.350 1994.700 3539.630 1994.980 ;
        RECT 3539.350 1994.080 3539.630 1994.360 ;
        RECT 3539.350 1990.390 3539.630 1990.670 ;
        RECT 3539.350 1989.770 3539.630 1990.050 ;
        RECT 3539.350 1989.150 3539.630 1989.430 ;
        RECT 3539.350 1988.530 3539.630 1988.810 ;
        RECT 3539.350 1987.910 3539.630 1988.190 ;
        RECT 3539.350 1987.290 3539.630 1987.570 ;
        RECT 3539.350 1986.670 3539.630 1986.950 ;
        RECT 3539.350 1986.050 3539.630 1986.330 ;
        RECT 3539.350 1985.430 3539.630 1985.710 ;
        RECT 3539.350 1984.810 3539.630 1985.090 ;
        RECT 3539.350 1984.190 3539.630 1984.470 ;
        RECT 3539.350 1983.570 3539.630 1983.850 ;
        RECT 3539.350 1982.950 3539.630 1983.230 ;
        RECT 3539.350 1982.330 3539.630 1982.610 ;
        RECT 3539.350 1981.710 3539.630 1981.990 ;
        RECT 350.370 733.010 350.650 733.290 ;
        RECT 350.370 732.390 350.650 732.670 ;
        RECT 350.370 731.770 350.650 732.050 ;
        RECT 350.370 731.150 350.650 731.430 ;
        RECT 350.370 730.530 350.650 730.810 ;
        RECT 350.370 729.910 350.650 730.190 ;
        RECT 350.370 729.290 350.650 729.570 ;
        RECT 350.370 728.670 350.650 728.950 ;
        RECT 350.370 728.050 350.650 728.330 ;
        RECT 350.370 727.430 350.650 727.710 ;
        RECT 350.370 726.810 350.650 727.090 ;
        RECT 350.370 726.190 350.650 726.470 ;
        RECT 350.370 725.570 350.650 725.850 ;
        RECT 350.370 724.950 350.650 725.230 ;
        RECT 350.370 724.330 350.650 724.610 ;
        RECT 350.370 720.640 350.650 720.920 ;
        RECT 350.370 720.020 350.650 720.300 ;
        RECT 350.370 719.400 350.650 719.680 ;
        RECT 350.370 718.780 350.650 719.060 ;
        RECT 350.370 718.160 350.650 718.440 ;
        RECT 350.370 717.540 350.650 717.820 ;
        RECT 350.370 716.920 350.650 717.200 ;
        RECT 350.370 716.300 350.650 716.580 ;
        RECT 350.370 715.680 350.650 715.960 ;
        RECT 350.370 715.060 350.650 715.340 ;
        RECT 350.370 714.440 350.650 714.720 ;
        RECT 350.370 713.820 350.650 714.100 ;
        RECT 350.370 713.200 350.650 713.480 ;
        RECT 350.370 712.580 350.650 712.860 ;
        RECT 350.370 711.960 350.650 712.240 ;
        RECT 350.370 711.340 350.650 711.620 ;
        RECT 350.370 708.790 350.650 709.070 ;
        RECT 350.370 708.170 350.650 708.450 ;
        RECT 350.370 707.550 350.650 707.830 ;
        RECT 350.370 706.930 350.650 707.210 ;
        RECT 350.370 706.310 350.650 706.590 ;
        RECT 350.370 705.690 350.650 705.970 ;
        RECT 350.370 705.070 350.650 705.350 ;
        RECT 350.370 704.450 350.650 704.730 ;
        RECT 350.370 703.830 350.650 704.110 ;
        RECT 350.370 703.210 350.650 703.490 ;
        RECT 350.370 702.590 350.650 702.870 ;
        RECT 350.370 701.970 350.650 702.250 ;
        RECT 350.370 701.350 350.650 701.630 ;
        RECT 350.370 700.730 350.650 701.010 ;
        RECT 350.370 700.110 350.650 700.390 ;
        RECT 350.370 699.490 350.650 699.770 ;
        RECT 350.370 695.260 350.650 695.540 ;
        RECT 350.370 694.640 350.650 694.920 ;
        RECT 350.370 694.020 350.650 694.300 ;
        RECT 350.370 693.400 350.650 693.680 ;
        RECT 350.370 692.780 350.650 693.060 ;
        RECT 350.370 692.160 350.650 692.440 ;
        RECT 350.370 691.540 350.650 691.820 ;
        RECT 350.370 690.920 350.650 691.200 ;
        RECT 350.370 690.300 350.650 690.580 ;
        RECT 350.370 689.680 350.650 689.960 ;
        RECT 350.370 689.060 350.650 689.340 ;
        RECT 350.370 688.440 350.650 688.720 ;
        RECT 350.370 687.820 350.650 688.100 ;
        RECT 350.370 687.200 350.650 687.480 ;
        RECT 350.370 686.580 350.650 686.860 ;
        RECT 350.370 685.960 350.650 686.240 ;
        RECT 350.370 683.410 350.650 683.690 ;
        RECT 350.370 682.790 350.650 683.070 ;
        RECT 350.370 682.170 350.650 682.450 ;
        RECT 350.370 681.550 350.650 681.830 ;
        RECT 350.370 680.930 350.650 681.210 ;
        RECT 350.370 680.310 350.650 680.590 ;
        RECT 350.370 679.690 350.650 679.970 ;
        RECT 350.370 679.070 350.650 679.350 ;
        RECT 350.370 678.450 350.650 678.730 ;
        RECT 350.370 677.830 350.650 678.110 ;
        RECT 350.370 677.210 350.650 677.490 ;
        RECT 350.370 676.590 350.650 676.870 ;
        RECT 350.370 675.970 350.650 676.250 ;
        RECT 350.370 675.350 350.650 675.630 ;
        RECT 350.370 674.730 350.650 675.010 ;
        RECT 350.370 674.110 350.650 674.390 ;
        RECT 350.370 670.390 350.650 670.670 ;
        RECT 350.370 669.770 350.650 670.050 ;
        RECT 350.370 669.150 350.650 669.430 ;
        RECT 350.370 668.530 350.650 668.810 ;
        RECT 350.370 667.910 350.650 668.190 ;
        RECT 350.370 667.290 350.650 667.570 ;
        RECT 350.370 666.670 350.650 666.950 ;
        RECT 350.370 666.050 350.650 666.330 ;
        RECT 350.370 665.430 350.650 665.710 ;
        RECT 350.370 664.810 350.650 665.090 ;
        RECT 350.370 664.190 350.650 664.470 ;
        RECT 350.370 663.570 350.650 663.850 ;
        RECT 350.370 662.950 350.650 663.230 ;
        RECT 350.370 662.330 350.650 662.610 ;
        RECT 350.370 661.710 350.650 661.990 ;
        RECT 350.370 528.010 350.650 528.290 ;
        RECT 350.370 527.390 350.650 527.670 ;
        RECT 350.370 526.770 350.650 527.050 ;
        RECT 350.370 526.150 350.650 526.430 ;
        RECT 350.370 525.530 350.650 525.810 ;
        RECT 350.370 524.910 350.650 525.190 ;
        RECT 350.370 524.290 350.650 524.570 ;
        RECT 350.370 523.670 350.650 523.950 ;
        RECT 350.370 523.050 350.650 523.330 ;
        RECT 350.370 522.430 350.650 522.710 ;
        RECT 350.370 521.810 350.650 522.090 ;
        RECT 350.370 521.190 350.650 521.470 ;
        RECT 350.370 520.570 350.650 520.850 ;
        RECT 350.370 519.950 350.650 520.230 ;
        RECT 350.370 519.330 350.650 519.610 ;
        RECT 350.370 515.640 350.650 515.920 ;
        RECT 350.370 515.020 350.650 515.300 ;
        RECT 350.370 514.400 350.650 514.680 ;
        RECT 350.370 513.780 350.650 514.060 ;
        RECT 350.370 513.160 350.650 513.440 ;
        RECT 350.370 512.540 350.650 512.820 ;
        RECT 350.370 511.920 350.650 512.200 ;
        RECT 350.370 511.300 350.650 511.580 ;
        RECT 350.370 510.680 350.650 510.960 ;
        RECT 350.370 510.060 350.650 510.340 ;
        RECT 350.370 509.440 350.650 509.720 ;
        RECT 350.370 508.820 350.650 509.100 ;
        RECT 350.370 508.200 350.650 508.480 ;
        RECT 350.370 507.580 350.650 507.860 ;
        RECT 350.370 506.960 350.650 507.240 ;
        RECT 350.370 506.340 350.650 506.620 ;
        RECT 350.370 503.790 350.650 504.070 ;
        RECT 350.370 503.170 350.650 503.450 ;
        RECT 350.370 502.550 350.650 502.830 ;
        RECT 350.370 501.930 350.650 502.210 ;
        RECT 350.370 501.310 350.650 501.590 ;
        RECT 350.370 500.690 350.650 500.970 ;
        RECT 350.370 500.070 350.650 500.350 ;
        RECT 350.370 499.450 350.650 499.730 ;
        RECT 350.370 498.830 350.650 499.110 ;
        RECT 350.370 498.210 350.650 498.490 ;
        RECT 350.370 497.590 350.650 497.870 ;
        RECT 350.370 496.970 350.650 497.250 ;
        RECT 350.370 496.350 350.650 496.630 ;
        RECT 350.370 495.730 350.650 496.010 ;
        RECT 350.370 495.110 350.650 495.390 ;
        RECT 350.370 494.490 350.650 494.770 ;
        RECT 350.370 490.260 350.650 490.540 ;
        RECT 350.370 489.640 350.650 489.920 ;
        RECT 350.370 489.020 350.650 489.300 ;
        RECT 350.370 488.400 350.650 488.680 ;
        RECT 350.370 487.780 350.650 488.060 ;
        RECT 350.370 487.160 350.650 487.440 ;
        RECT 350.370 486.540 350.650 486.820 ;
        RECT 350.370 485.920 350.650 486.200 ;
        RECT 350.370 485.300 350.650 485.580 ;
        RECT 350.370 484.680 350.650 484.960 ;
        RECT 350.370 484.060 350.650 484.340 ;
        RECT 350.370 483.440 350.650 483.720 ;
        RECT 350.370 482.820 350.650 483.100 ;
        RECT 350.370 482.200 350.650 482.480 ;
        RECT 350.370 481.580 350.650 481.860 ;
        RECT 350.370 480.960 350.650 481.240 ;
        RECT 350.370 478.410 350.650 478.690 ;
        RECT 350.370 477.790 350.650 478.070 ;
        RECT 350.370 477.170 350.650 477.450 ;
        RECT 350.370 476.550 350.650 476.830 ;
        RECT 350.370 475.930 350.650 476.210 ;
        RECT 350.370 475.310 350.650 475.590 ;
        RECT 350.370 474.690 350.650 474.970 ;
        RECT 350.370 474.070 350.650 474.350 ;
        RECT 350.370 473.450 350.650 473.730 ;
        RECT 350.370 472.830 350.650 473.110 ;
        RECT 350.370 472.210 350.650 472.490 ;
        RECT 350.370 471.590 350.650 471.870 ;
        RECT 350.370 470.970 350.650 471.250 ;
        RECT 350.370 470.350 350.650 470.630 ;
        RECT 350.370 469.730 350.650 470.010 ;
        RECT 350.370 469.110 350.650 469.390 ;
        RECT 350.370 465.390 350.650 465.670 ;
        RECT 350.370 464.770 350.650 465.050 ;
        RECT 350.370 464.150 350.650 464.430 ;
        RECT 350.370 463.530 350.650 463.810 ;
        RECT 350.370 462.910 350.650 463.190 ;
        RECT 350.370 462.290 350.650 462.570 ;
        RECT 350.370 461.670 350.650 461.950 ;
        RECT 350.370 461.050 350.650 461.330 ;
        RECT 350.370 460.430 350.650 460.710 ;
        RECT 350.370 459.810 350.650 460.090 ;
        RECT 350.370 459.190 350.650 459.470 ;
        RECT 350.370 458.570 350.650 458.850 ;
        RECT 350.370 457.950 350.650 458.230 ;
        RECT 350.370 457.330 350.650 457.610 ;
        RECT 350.370 456.710 350.650 456.990 ;
        RECT 536.710 350.370 536.990 350.650 ;
        RECT 537.330 350.370 537.610 350.650 ;
        RECT 537.950 350.370 538.230 350.650 ;
        RECT 538.570 350.370 538.850 350.650 ;
        RECT 539.190 350.370 539.470 350.650 ;
        RECT 539.810 350.370 540.090 350.650 ;
        RECT 540.430 350.370 540.710 350.650 ;
        RECT 541.050 350.370 541.330 350.650 ;
        RECT 541.670 350.370 541.950 350.650 ;
        RECT 542.290 350.370 542.570 350.650 ;
        RECT 542.910 350.370 543.190 350.650 ;
        RECT 543.530 350.370 543.810 350.650 ;
        RECT 544.150 350.370 544.430 350.650 ;
        RECT 544.770 350.370 545.050 350.650 ;
        RECT 545.390 350.370 545.670 350.650 ;
        RECT 549.110 350.370 549.390 350.650 ;
        RECT 549.730 350.370 550.010 350.650 ;
        RECT 550.350 350.370 550.630 350.650 ;
        RECT 550.970 350.370 551.250 350.650 ;
        RECT 551.590 350.370 551.870 350.650 ;
        RECT 552.210 350.370 552.490 350.650 ;
        RECT 552.830 350.370 553.110 350.650 ;
        RECT 553.450 350.370 553.730 350.650 ;
        RECT 554.070 350.370 554.350 350.650 ;
        RECT 554.690 350.370 554.970 350.650 ;
        RECT 555.310 350.370 555.590 350.650 ;
        RECT 555.930 350.370 556.210 350.650 ;
        RECT 556.550 350.370 556.830 350.650 ;
        RECT 557.170 350.370 557.450 350.650 ;
        RECT 557.790 350.370 558.070 350.650 ;
        RECT 558.410 350.370 558.690 350.650 ;
        RECT 560.960 350.370 561.240 350.650 ;
        RECT 561.580 350.370 561.860 350.650 ;
        RECT 562.200 350.370 562.480 350.650 ;
        RECT 562.820 350.370 563.100 350.650 ;
        RECT 563.440 350.370 563.720 350.650 ;
        RECT 564.060 350.370 564.340 350.650 ;
        RECT 564.680 350.370 564.960 350.650 ;
        RECT 565.300 350.370 565.580 350.650 ;
        RECT 565.920 350.370 566.200 350.650 ;
        RECT 566.540 350.370 566.820 350.650 ;
        RECT 567.160 350.370 567.440 350.650 ;
        RECT 567.780 350.370 568.060 350.650 ;
        RECT 568.400 350.370 568.680 350.650 ;
        RECT 569.020 350.370 569.300 350.650 ;
        RECT 569.640 350.370 569.920 350.650 ;
        RECT 570.260 350.370 570.540 350.650 ;
        RECT 574.460 350.370 574.740 350.650 ;
        RECT 575.080 350.370 575.360 350.650 ;
        RECT 575.700 350.370 575.980 350.650 ;
        RECT 576.320 350.370 576.600 350.650 ;
        RECT 576.940 350.370 577.220 350.650 ;
        RECT 577.560 350.370 577.840 350.650 ;
        RECT 578.180 350.370 578.460 350.650 ;
        RECT 578.800 350.370 579.080 350.650 ;
        RECT 579.420 350.370 579.700 350.650 ;
        RECT 580.040 350.370 580.320 350.650 ;
        RECT 580.660 350.370 580.940 350.650 ;
        RECT 581.280 350.370 581.560 350.650 ;
        RECT 581.900 350.370 582.180 350.650 ;
        RECT 582.520 350.370 582.800 350.650 ;
        RECT 583.140 350.370 583.420 350.650 ;
        RECT 583.760 350.370 584.040 350.650 ;
        RECT 586.310 350.370 586.590 350.650 ;
        RECT 586.930 350.370 587.210 350.650 ;
        RECT 587.550 350.370 587.830 350.650 ;
        RECT 588.170 350.370 588.450 350.650 ;
        RECT 588.790 350.370 589.070 350.650 ;
        RECT 589.410 350.370 589.690 350.650 ;
        RECT 590.030 350.370 590.310 350.650 ;
        RECT 590.650 350.370 590.930 350.650 ;
        RECT 591.270 350.370 591.550 350.650 ;
        RECT 591.890 350.370 592.170 350.650 ;
        RECT 592.510 350.370 592.790 350.650 ;
        RECT 593.130 350.370 593.410 350.650 ;
        RECT 593.750 350.370 594.030 350.650 ;
        RECT 594.370 350.370 594.650 350.650 ;
        RECT 594.990 350.370 595.270 350.650 ;
        RECT 595.610 350.370 595.890 350.650 ;
        RECT 599.330 350.370 599.610 350.650 ;
        RECT 599.950 350.370 600.230 350.650 ;
        RECT 600.570 350.370 600.850 350.650 ;
        RECT 601.190 350.370 601.470 350.650 ;
        RECT 601.810 350.370 602.090 350.650 ;
        RECT 602.430 350.370 602.710 350.650 ;
        RECT 603.050 350.370 603.330 350.650 ;
        RECT 603.670 350.370 603.950 350.650 ;
        RECT 604.290 350.370 604.570 350.650 ;
        RECT 604.910 350.370 605.190 350.650 ;
        RECT 605.530 350.370 605.810 350.650 ;
        RECT 606.150 350.370 606.430 350.650 ;
        RECT 606.770 350.370 607.050 350.650 ;
        RECT 607.390 350.370 607.670 350.650 ;
        RECT 608.010 350.370 608.290 350.650 ;
        RECT 1361.710 350.370 1361.990 350.650 ;
        RECT 1362.330 350.370 1362.610 350.650 ;
        RECT 1362.950 350.370 1363.230 350.650 ;
        RECT 1363.570 350.370 1363.850 350.650 ;
        RECT 1364.190 350.370 1364.470 350.650 ;
        RECT 1364.810 350.370 1365.090 350.650 ;
        RECT 1365.430 350.370 1365.710 350.650 ;
        RECT 1366.050 350.370 1366.330 350.650 ;
        RECT 1366.670 350.370 1366.950 350.650 ;
        RECT 1367.290 350.370 1367.570 350.650 ;
        RECT 1367.910 350.370 1368.190 350.650 ;
        RECT 1368.530 350.370 1368.810 350.650 ;
        RECT 1369.150 350.370 1369.430 350.650 ;
        RECT 1369.770 350.370 1370.050 350.650 ;
        RECT 1370.390 350.370 1370.670 350.650 ;
        RECT 1374.110 350.370 1374.390 350.650 ;
        RECT 1374.730 350.370 1375.010 350.650 ;
        RECT 1375.350 350.370 1375.630 350.650 ;
        RECT 1375.970 350.370 1376.250 350.650 ;
        RECT 1376.590 350.370 1376.870 350.650 ;
        RECT 1377.210 350.370 1377.490 350.650 ;
        RECT 1377.830 350.370 1378.110 350.650 ;
        RECT 1378.450 350.370 1378.730 350.650 ;
        RECT 1379.070 350.370 1379.350 350.650 ;
        RECT 1379.690 350.370 1379.970 350.650 ;
        RECT 1380.310 350.370 1380.590 350.650 ;
        RECT 1380.930 350.370 1381.210 350.650 ;
        RECT 1381.550 350.370 1381.830 350.650 ;
        RECT 1382.170 350.370 1382.450 350.650 ;
        RECT 1382.790 350.370 1383.070 350.650 ;
        RECT 1383.410 350.370 1383.690 350.650 ;
        RECT 1385.960 350.370 1386.240 350.650 ;
        RECT 1386.580 350.370 1386.860 350.650 ;
        RECT 1387.200 350.370 1387.480 350.650 ;
        RECT 1387.820 350.370 1388.100 350.650 ;
        RECT 1388.440 350.370 1388.720 350.650 ;
        RECT 1389.060 350.370 1389.340 350.650 ;
        RECT 1389.680 350.370 1389.960 350.650 ;
        RECT 1390.300 350.370 1390.580 350.650 ;
        RECT 1390.920 350.370 1391.200 350.650 ;
        RECT 1391.540 350.370 1391.820 350.650 ;
        RECT 1392.160 350.370 1392.440 350.650 ;
        RECT 1392.780 350.370 1393.060 350.650 ;
        RECT 1393.400 350.370 1393.680 350.650 ;
        RECT 1394.020 350.370 1394.300 350.650 ;
        RECT 1394.640 350.370 1394.920 350.650 ;
        RECT 1395.260 350.370 1395.540 350.650 ;
        RECT 1399.460 350.370 1399.740 350.650 ;
        RECT 1400.080 350.370 1400.360 350.650 ;
        RECT 1400.700 350.370 1400.980 350.650 ;
        RECT 1401.320 350.370 1401.600 350.650 ;
        RECT 1401.940 350.370 1402.220 350.650 ;
        RECT 1402.560 350.370 1402.840 350.650 ;
        RECT 1403.180 350.370 1403.460 350.650 ;
        RECT 1403.800 350.370 1404.080 350.650 ;
        RECT 1404.420 350.370 1404.700 350.650 ;
        RECT 1405.040 350.370 1405.320 350.650 ;
        RECT 1405.660 350.370 1405.940 350.650 ;
        RECT 1406.280 350.370 1406.560 350.650 ;
        RECT 1406.900 350.370 1407.180 350.650 ;
        RECT 1407.520 350.370 1407.800 350.650 ;
        RECT 1408.140 350.370 1408.420 350.650 ;
        RECT 1408.760 350.370 1409.040 350.650 ;
        RECT 1411.310 350.370 1411.590 350.650 ;
        RECT 1411.930 350.370 1412.210 350.650 ;
        RECT 1412.550 350.370 1412.830 350.650 ;
        RECT 1413.170 350.370 1413.450 350.650 ;
        RECT 1413.790 350.370 1414.070 350.650 ;
        RECT 1414.410 350.370 1414.690 350.650 ;
        RECT 1415.030 350.370 1415.310 350.650 ;
        RECT 1415.650 350.370 1415.930 350.650 ;
        RECT 1416.270 350.370 1416.550 350.650 ;
        RECT 1416.890 350.370 1417.170 350.650 ;
        RECT 1417.510 350.370 1417.790 350.650 ;
        RECT 1418.130 350.370 1418.410 350.650 ;
        RECT 1418.750 350.370 1419.030 350.650 ;
        RECT 1419.370 350.370 1419.650 350.650 ;
        RECT 1419.990 350.370 1420.270 350.650 ;
        RECT 1420.610 350.370 1420.890 350.650 ;
        RECT 1424.330 350.370 1424.610 350.650 ;
        RECT 1424.950 350.370 1425.230 350.650 ;
        RECT 1425.570 350.370 1425.850 350.650 ;
        RECT 1426.190 350.370 1426.470 350.650 ;
        RECT 1426.810 350.370 1427.090 350.650 ;
        RECT 1427.430 350.370 1427.710 350.650 ;
        RECT 1428.050 350.370 1428.330 350.650 ;
        RECT 1428.670 350.370 1428.950 350.650 ;
        RECT 1429.290 350.370 1429.570 350.650 ;
        RECT 1429.910 350.370 1430.190 350.650 ;
        RECT 1430.530 350.370 1430.810 350.650 ;
        RECT 1431.150 350.370 1431.430 350.650 ;
        RECT 1431.770 350.370 1432.050 350.650 ;
        RECT 1432.390 350.370 1432.670 350.650 ;
        RECT 1433.010 350.370 1433.290 350.650 ;
        RECT 3011.710 350.370 3011.990 350.650 ;
        RECT 3012.330 350.370 3012.610 350.650 ;
        RECT 3012.950 350.370 3013.230 350.650 ;
        RECT 3013.570 350.370 3013.850 350.650 ;
        RECT 3014.190 350.370 3014.470 350.650 ;
        RECT 3014.810 350.370 3015.090 350.650 ;
        RECT 3015.430 350.370 3015.710 350.650 ;
        RECT 3016.050 350.370 3016.330 350.650 ;
        RECT 3016.670 350.370 3016.950 350.650 ;
        RECT 3017.290 350.370 3017.570 350.650 ;
        RECT 3017.910 350.370 3018.190 350.650 ;
        RECT 3018.530 350.370 3018.810 350.650 ;
        RECT 3019.150 350.370 3019.430 350.650 ;
        RECT 3019.770 350.370 3020.050 350.650 ;
        RECT 3020.390 350.370 3020.670 350.650 ;
        RECT 3024.110 350.370 3024.390 350.650 ;
        RECT 3024.730 350.370 3025.010 350.650 ;
        RECT 3025.350 350.370 3025.630 350.650 ;
        RECT 3025.970 350.370 3026.250 350.650 ;
        RECT 3026.590 350.370 3026.870 350.650 ;
        RECT 3027.210 350.370 3027.490 350.650 ;
        RECT 3027.830 350.370 3028.110 350.650 ;
        RECT 3028.450 350.370 3028.730 350.650 ;
        RECT 3029.070 350.370 3029.350 350.650 ;
        RECT 3029.690 350.370 3029.970 350.650 ;
        RECT 3030.310 350.370 3030.590 350.650 ;
        RECT 3030.930 350.370 3031.210 350.650 ;
        RECT 3031.550 350.370 3031.830 350.650 ;
        RECT 3032.170 350.370 3032.450 350.650 ;
        RECT 3032.790 350.370 3033.070 350.650 ;
        RECT 3033.410 350.370 3033.690 350.650 ;
        RECT 3035.960 350.370 3036.240 350.650 ;
        RECT 3036.580 350.370 3036.860 350.650 ;
        RECT 3037.200 350.370 3037.480 350.650 ;
        RECT 3037.820 350.370 3038.100 350.650 ;
        RECT 3038.440 350.370 3038.720 350.650 ;
        RECT 3039.060 350.370 3039.340 350.650 ;
        RECT 3039.680 350.370 3039.960 350.650 ;
        RECT 3040.300 350.370 3040.580 350.650 ;
        RECT 3040.920 350.370 3041.200 350.650 ;
        RECT 3041.540 350.370 3041.820 350.650 ;
        RECT 3042.160 350.370 3042.440 350.650 ;
        RECT 3042.780 350.370 3043.060 350.650 ;
        RECT 3043.400 350.370 3043.680 350.650 ;
        RECT 3044.020 350.370 3044.300 350.650 ;
        RECT 3044.640 350.370 3044.920 350.650 ;
        RECT 3045.260 350.370 3045.540 350.650 ;
        RECT 3049.460 350.370 3049.740 350.650 ;
        RECT 3050.080 350.370 3050.360 350.650 ;
        RECT 3050.700 350.370 3050.980 350.650 ;
        RECT 3051.320 350.370 3051.600 350.650 ;
        RECT 3051.940 350.370 3052.220 350.650 ;
        RECT 3052.560 350.370 3052.840 350.650 ;
        RECT 3053.180 350.370 3053.460 350.650 ;
        RECT 3053.800 350.370 3054.080 350.650 ;
        RECT 3054.420 350.370 3054.700 350.650 ;
        RECT 3055.040 350.370 3055.320 350.650 ;
        RECT 3055.660 350.370 3055.940 350.650 ;
        RECT 3056.280 350.370 3056.560 350.650 ;
        RECT 3056.900 350.370 3057.180 350.650 ;
        RECT 3057.520 350.370 3057.800 350.650 ;
        RECT 3058.140 350.370 3058.420 350.650 ;
        RECT 3058.760 350.370 3059.040 350.650 ;
        RECT 3061.310 350.370 3061.590 350.650 ;
        RECT 3061.930 350.370 3062.210 350.650 ;
        RECT 3062.550 350.370 3062.830 350.650 ;
        RECT 3063.170 350.370 3063.450 350.650 ;
        RECT 3063.790 350.370 3064.070 350.650 ;
        RECT 3064.410 350.370 3064.690 350.650 ;
        RECT 3065.030 350.370 3065.310 350.650 ;
        RECT 3065.650 350.370 3065.930 350.650 ;
        RECT 3066.270 350.370 3066.550 350.650 ;
        RECT 3066.890 350.370 3067.170 350.650 ;
        RECT 3067.510 350.370 3067.790 350.650 ;
        RECT 3068.130 350.370 3068.410 350.650 ;
        RECT 3068.750 350.370 3069.030 350.650 ;
        RECT 3069.370 350.370 3069.650 350.650 ;
        RECT 3069.990 350.370 3070.270 350.650 ;
        RECT 3070.610 350.370 3070.890 350.650 ;
        RECT 3074.330 350.370 3074.610 350.650 ;
        RECT 3074.950 350.370 3075.230 350.650 ;
        RECT 3075.570 350.370 3075.850 350.650 ;
        RECT 3076.190 350.370 3076.470 350.650 ;
        RECT 3076.810 350.370 3077.090 350.650 ;
        RECT 3077.430 350.370 3077.710 350.650 ;
        RECT 3078.050 350.370 3078.330 350.650 ;
        RECT 3078.670 350.370 3078.950 350.650 ;
        RECT 3079.290 350.370 3079.570 350.650 ;
        RECT 3079.910 350.370 3080.190 350.650 ;
        RECT 3080.530 350.370 3080.810 350.650 ;
        RECT 3081.150 350.370 3081.430 350.650 ;
        RECT 3081.770 350.370 3082.050 350.650 ;
        RECT 3082.390 350.370 3082.670 350.650 ;
        RECT 3083.010 350.370 3083.290 350.650 ;
        RECT 3286.710 350.370 3286.990 350.650 ;
        RECT 3287.330 350.370 3287.610 350.650 ;
        RECT 3287.950 350.370 3288.230 350.650 ;
        RECT 3288.570 350.370 3288.850 350.650 ;
        RECT 3289.190 350.370 3289.470 350.650 ;
        RECT 3289.810 350.370 3290.090 350.650 ;
        RECT 3290.430 350.370 3290.710 350.650 ;
        RECT 3291.050 350.370 3291.330 350.650 ;
        RECT 3291.670 350.370 3291.950 350.650 ;
        RECT 3292.290 350.370 3292.570 350.650 ;
        RECT 3292.910 350.370 3293.190 350.650 ;
        RECT 3293.530 350.370 3293.810 350.650 ;
        RECT 3294.150 350.370 3294.430 350.650 ;
        RECT 3294.770 350.370 3295.050 350.650 ;
        RECT 3295.390 350.370 3295.670 350.650 ;
        RECT 3299.110 350.370 3299.390 350.650 ;
        RECT 3299.730 350.370 3300.010 350.650 ;
        RECT 3300.350 350.370 3300.630 350.650 ;
        RECT 3300.970 350.370 3301.250 350.650 ;
        RECT 3301.590 350.370 3301.870 350.650 ;
        RECT 3302.210 350.370 3302.490 350.650 ;
        RECT 3302.830 350.370 3303.110 350.650 ;
        RECT 3303.450 350.370 3303.730 350.650 ;
        RECT 3304.070 350.370 3304.350 350.650 ;
        RECT 3304.690 350.370 3304.970 350.650 ;
        RECT 3305.310 350.370 3305.590 350.650 ;
        RECT 3305.930 350.370 3306.210 350.650 ;
        RECT 3306.550 350.370 3306.830 350.650 ;
        RECT 3307.170 350.370 3307.450 350.650 ;
        RECT 3307.790 350.370 3308.070 350.650 ;
        RECT 3308.410 350.370 3308.690 350.650 ;
        RECT 3310.960 350.370 3311.240 350.650 ;
        RECT 3311.580 350.370 3311.860 350.650 ;
        RECT 3312.200 350.370 3312.480 350.650 ;
        RECT 3312.820 350.370 3313.100 350.650 ;
        RECT 3313.440 350.370 3313.720 350.650 ;
        RECT 3314.060 350.370 3314.340 350.650 ;
        RECT 3314.680 350.370 3314.960 350.650 ;
        RECT 3315.300 350.370 3315.580 350.650 ;
        RECT 3315.920 350.370 3316.200 350.650 ;
        RECT 3316.540 350.370 3316.820 350.650 ;
        RECT 3317.160 350.370 3317.440 350.650 ;
        RECT 3317.780 350.370 3318.060 350.650 ;
        RECT 3318.400 350.370 3318.680 350.650 ;
        RECT 3319.020 350.370 3319.300 350.650 ;
        RECT 3319.640 350.370 3319.920 350.650 ;
        RECT 3320.260 350.370 3320.540 350.650 ;
        RECT 3324.460 350.370 3324.740 350.650 ;
        RECT 3325.080 350.370 3325.360 350.650 ;
        RECT 3325.700 350.370 3325.980 350.650 ;
        RECT 3326.320 350.370 3326.600 350.650 ;
        RECT 3326.940 350.370 3327.220 350.650 ;
        RECT 3327.560 350.370 3327.840 350.650 ;
        RECT 3328.180 350.370 3328.460 350.650 ;
        RECT 3328.800 350.370 3329.080 350.650 ;
        RECT 3329.420 350.370 3329.700 350.650 ;
        RECT 3330.040 350.370 3330.320 350.650 ;
        RECT 3330.660 350.370 3330.940 350.650 ;
        RECT 3331.280 350.370 3331.560 350.650 ;
        RECT 3331.900 350.370 3332.180 350.650 ;
        RECT 3332.520 350.370 3332.800 350.650 ;
        RECT 3333.140 350.370 3333.420 350.650 ;
        RECT 3333.760 350.370 3334.040 350.650 ;
        RECT 3336.310 350.370 3336.590 350.650 ;
        RECT 3336.930 350.370 3337.210 350.650 ;
        RECT 3337.550 350.370 3337.830 350.650 ;
        RECT 3338.170 350.370 3338.450 350.650 ;
        RECT 3338.790 350.370 3339.070 350.650 ;
        RECT 3339.410 350.370 3339.690 350.650 ;
        RECT 3340.030 350.370 3340.310 350.650 ;
        RECT 3340.650 350.370 3340.930 350.650 ;
        RECT 3341.270 350.370 3341.550 350.650 ;
        RECT 3341.890 350.370 3342.170 350.650 ;
        RECT 3342.510 350.370 3342.790 350.650 ;
        RECT 3343.130 350.370 3343.410 350.650 ;
        RECT 3343.750 350.370 3344.030 350.650 ;
        RECT 3344.370 350.370 3344.650 350.650 ;
        RECT 3344.990 350.370 3345.270 350.650 ;
        RECT 3345.610 350.370 3345.890 350.650 ;
        RECT 3349.330 350.370 3349.610 350.650 ;
        RECT 3349.950 350.370 3350.230 350.650 ;
        RECT 3350.570 350.370 3350.850 350.650 ;
        RECT 3351.190 350.370 3351.470 350.650 ;
        RECT 3351.810 350.370 3352.090 350.650 ;
        RECT 3352.430 350.370 3352.710 350.650 ;
        RECT 3353.050 350.370 3353.330 350.650 ;
        RECT 3353.670 350.370 3353.950 350.650 ;
        RECT 3354.290 350.370 3354.570 350.650 ;
        RECT 3354.910 350.370 3355.190 350.650 ;
        RECT 3355.530 350.370 3355.810 350.650 ;
        RECT 3356.150 350.370 3356.430 350.650 ;
        RECT 3356.770 350.370 3357.050 350.650 ;
        RECT 3357.390 350.370 3357.670 350.650 ;
        RECT 3358.010 350.370 3358.290 350.650 ;
      LAYER Metal3 ;
        RECT 1906.360 4749.000 1915.860 4750.000 ;
        RECT 1918.760 4749.000 1929.010 4750.000 ;
        RECT 1930.610 4749.000 1940.860 4750.000 ;
        RECT 1944.140 4749.000 1954.390 4750.000 ;
        RECT 1955.990 4749.000 1966.240 4750.000 ;
        RECT 1969.140 4749.000 1978.640 4750.000 ;
        RECT 3006.360 4749.000 3015.860 4750.000 ;
        RECT 3018.760 4749.000 3029.010 4750.000 ;
        RECT 3030.610 4749.000 3040.860 4750.000 ;
        RECT 3044.140 4749.000 3054.390 4750.000 ;
        RECT 3055.990 4749.000 3066.240 4750.000 ;
        RECT 3069.140 4749.000 3078.640 4750.000 ;
        RECT 350.000 4414.140 351.000 4423.640 ;
        RECT 350.000 4400.990 351.000 4411.240 ;
        RECT 3539.000 4409.140 3540.000 4418.640 ;
        RECT 350.000 4389.140 351.000 4399.390 ;
        RECT 3539.000 4395.990 3540.000 4406.240 ;
        RECT 350.000 4375.610 351.000 4385.860 ;
        RECT 3539.000 4384.140 3540.000 4394.390 ;
        RECT 350.000 4363.760 351.000 4374.010 ;
        RECT 3539.000 4370.610 3540.000 4380.860 ;
        RECT 350.000 4351.360 351.000 4360.860 ;
        RECT 3539.000 4358.760 3540.000 4369.010 ;
        RECT 3539.000 4346.360 3540.000 4355.860 ;
        RECT 350.000 4209.140 351.000 4218.640 ;
        RECT 350.000 4195.990 351.000 4206.240 ;
        RECT 350.000 4184.140 351.000 4194.390 ;
        RECT 350.000 4170.610 351.000 4180.860 ;
        RECT 350.000 4158.760 351.000 4169.010 ;
        RECT 350.000 4146.360 351.000 4155.860 ;
        RECT 350.000 4004.140 351.000 4013.640 ;
        RECT 350.000 3990.990 351.000 4001.240 ;
        RECT 350.000 3979.140 351.000 3989.390 ;
        RECT 3539.000 3979.140 3540.000 3988.640 ;
        RECT 350.000 3965.610 351.000 3975.860 ;
        RECT 3539.000 3965.990 3540.000 3976.240 ;
        RECT 350.000 3953.760 351.000 3964.010 ;
        RECT 3539.000 3954.140 3540.000 3964.390 ;
        RECT 350.000 3941.360 351.000 3950.860 ;
        RECT 3539.000 3940.610 3540.000 3950.860 ;
        RECT 3539.000 3928.760 3540.000 3939.010 ;
        RECT 3539.000 3916.360 3540.000 3925.860 ;
        RECT 3539.000 2474.140 3540.000 2483.640 ;
        RECT 3539.000 2460.990 3540.000 2471.240 ;
        RECT 3539.000 2449.140 3540.000 2459.390 ;
        RECT 3539.000 2435.610 3540.000 2445.860 ;
        RECT 3539.000 2423.760 3540.000 2434.010 ;
        RECT 3539.000 2411.360 3540.000 2420.860 ;
        RECT 350.000 2364.140 351.000 2373.640 ;
        RECT 350.000 2350.990 351.000 2361.240 ;
        RECT 350.000 2339.140 351.000 2349.390 ;
        RECT 350.000 2325.610 351.000 2335.860 ;
        RECT 350.000 2313.760 351.000 2324.010 ;
        RECT 350.000 2301.360 351.000 2310.860 ;
        RECT 3539.005 2259.140 3540.005 2268.640 ;
        RECT 3539.005 2245.990 3540.005 2256.240 ;
        RECT 3539.005 2234.140 3540.005 2244.390 ;
        RECT 3539.005 2220.610 3540.005 2230.860 ;
        RECT 3539.005 2208.760 3540.005 2219.010 ;
        RECT 3539.005 2196.360 3540.005 2205.860 ;
        RECT 350.000 2159.145 351.000 2168.645 ;
        RECT 350.000 2145.995 351.000 2156.245 ;
        RECT 350.000 2134.145 351.000 2144.395 ;
        RECT 350.000 2120.615 351.000 2130.865 ;
        RECT 350.000 2108.765 351.000 2119.015 ;
        RECT 350.000 2096.365 351.000 2105.865 ;
        RECT 3539.000 2044.140 3540.000 2053.640 ;
        RECT 3539.000 2030.990 3540.000 2041.240 ;
        RECT 3539.000 2019.140 3540.000 2029.390 ;
        RECT 3539.000 2005.610 3540.000 2015.860 ;
        RECT 3539.000 1993.760 3540.000 2004.010 ;
        RECT 3539.000 1981.360 3540.000 1990.860 ;
        RECT 350.000 724.140 351.000 733.640 ;
        RECT 350.000 710.990 351.000 721.240 ;
        RECT 350.000 699.140 351.000 709.390 ;
        RECT 350.000 685.610 351.000 695.860 ;
        RECT 350.000 673.760 351.000 684.010 ;
        RECT 350.000 661.360 351.000 670.860 ;
        RECT 350.000 519.140 351.000 528.640 ;
        RECT 350.000 505.990 351.000 516.240 ;
        RECT 350.000 494.140 351.000 504.390 ;
        RECT 350.000 480.610 351.000 490.860 ;
        RECT 350.000 468.760 351.000 479.010 ;
        RECT 350.000 456.360 351.000 465.860 ;
        RECT 536.360 350.000 545.860 351.000 ;
        RECT 548.760 350.000 559.010 351.000 ;
        RECT 560.610 350.000 570.860 351.000 ;
        RECT 574.140 350.000 584.390 351.000 ;
        RECT 585.990 350.000 596.240 351.000 ;
        RECT 599.140 350.000 608.640 351.000 ;
        RECT 1361.360 350.000 1370.860 351.000 ;
        RECT 1373.760 350.000 1384.010 351.000 ;
        RECT 1385.610 350.000 1395.860 351.000 ;
        RECT 1399.140 350.000 1409.390 351.000 ;
        RECT 1410.990 350.000 1421.240 351.000 ;
        RECT 1424.140 350.000 1433.640 351.000 ;
        RECT 3011.360 350.000 3020.860 351.000 ;
        RECT 3023.760 350.000 3034.010 351.000 ;
        RECT 3035.610 350.000 3045.860 351.000 ;
        RECT 3049.140 350.000 3059.390 351.000 ;
        RECT 3060.990 350.000 3071.240 351.000 ;
        RECT 3074.140 350.000 3083.640 351.000 ;
        RECT 3286.360 350.000 3295.860 351.000 ;
        RECT 3298.760 350.000 3309.010 351.000 ;
        RECT 3310.610 350.000 3320.860 351.000 ;
        RECT 3324.140 350.000 3334.390 351.000 ;
        RECT 3335.990 350.000 3346.240 351.000 ;
        RECT 3349.140 350.000 3358.640 351.000 ;
      LAYER VIA3 ;
        RECT 1906.710 4749.350 1906.990 4749.630 ;
        RECT 1907.330 4749.350 1907.610 4749.630 ;
        RECT 1907.950 4749.350 1908.230 4749.630 ;
        RECT 1908.570 4749.350 1908.850 4749.630 ;
        RECT 1909.190 4749.350 1909.470 4749.630 ;
        RECT 1909.810 4749.350 1910.090 4749.630 ;
        RECT 1910.430 4749.350 1910.710 4749.630 ;
        RECT 1911.050 4749.350 1911.330 4749.630 ;
        RECT 1911.670 4749.350 1911.950 4749.630 ;
        RECT 1912.290 4749.350 1912.570 4749.630 ;
        RECT 1912.910 4749.350 1913.190 4749.630 ;
        RECT 1913.530 4749.350 1913.810 4749.630 ;
        RECT 1914.150 4749.350 1914.430 4749.630 ;
        RECT 1914.770 4749.350 1915.050 4749.630 ;
        RECT 1915.390 4749.350 1915.670 4749.630 ;
        RECT 1919.110 4749.350 1919.390 4749.630 ;
        RECT 1919.730 4749.350 1920.010 4749.630 ;
        RECT 1920.350 4749.350 1920.630 4749.630 ;
        RECT 1920.970 4749.350 1921.250 4749.630 ;
        RECT 1921.590 4749.350 1921.870 4749.630 ;
        RECT 1922.210 4749.350 1922.490 4749.630 ;
        RECT 1922.830 4749.350 1923.110 4749.630 ;
        RECT 1923.450 4749.350 1923.730 4749.630 ;
        RECT 1924.070 4749.350 1924.350 4749.630 ;
        RECT 1924.690 4749.350 1924.970 4749.630 ;
        RECT 1925.310 4749.350 1925.590 4749.630 ;
        RECT 1925.930 4749.350 1926.210 4749.630 ;
        RECT 1926.550 4749.350 1926.830 4749.630 ;
        RECT 1927.170 4749.350 1927.450 4749.630 ;
        RECT 1927.790 4749.350 1928.070 4749.630 ;
        RECT 1928.410 4749.350 1928.690 4749.630 ;
        RECT 1930.960 4749.350 1931.240 4749.630 ;
        RECT 1931.580 4749.350 1931.860 4749.630 ;
        RECT 1932.200 4749.350 1932.480 4749.630 ;
        RECT 1932.820 4749.350 1933.100 4749.630 ;
        RECT 1933.440 4749.350 1933.720 4749.630 ;
        RECT 1934.060 4749.350 1934.340 4749.630 ;
        RECT 1934.680 4749.350 1934.960 4749.630 ;
        RECT 1935.300 4749.350 1935.580 4749.630 ;
        RECT 1935.920 4749.350 1936.200 4749.630 ;
        RECT 1936.540 4749.350 1936.820 4749.630 ;
        RECT 1937.160 4749.350 1937.440 4749.630 ;
        RECT 1937.780 4749.350 1938.060 4749.630 ;
        RECT 1938.400 4749.350 1938.680 4749.630 ;
        RECT 1939.020 4749.350 1939.300 4749.630 ;
        RECT 1939.640 4749.350 1939.920 4749.630 ;
        RECT 1940.260 4749.350 1940.540 4749.630 ;
        RECT 1944.460 4749.350 1944.740 4749.630 ;
        RECT 1945.080 4749.350 1945.360 4749.630 ;
        RECT 1945.700 4749.350 1945.980 4749.630 ;
        RECT 1946.320 4749.350 1946.600 4749.630 ;
        RECT 1946.940 4749.350 1947.220 4749.630 ;
        RECT 1947.560 4749.350 1947.840 4749.630 ;
        RECT 1948.180 4749.350 1948.460 4749.630 ;
        RECT 1948.800 4749.350 1949.080 4749.630 ;
        RECT 1949.420 4749.350 1949.700 4749.630 ;
        RECT 1950.040 4749.350 1950.320 4749.630 ;
        RECT 1950.660 4749.350 1950.940 4749.630 ;
        RECT 1951.280 4749.350 1951.560 4749.630 ;
        RECT 1951.900 4749.350 1952.180 4749.630 ;
        RECT 1952.520 4749.350 1952.800 4749.630 ;
        RECT 1953.140 4749.350 1953.420 4749.630 ;
        RECT 1953.760 4749.350 1954.040 4749.630 ;
        RECT 1956.310 4749.350 1956.590 4749.630 ;
        RECT 1956.930 4749.350 1957.210 4749.630 ;
        RECT 1957.550 4749.350 1957.830 4749.630 ;
        RECT 1958.170 4749.350 1958.450 4749.630 ;
        RECT 1958.790 4749.350 1959.070 4749.630 ;
        RECT 1959.410 4749.350 1959.690 4749.630 ;
        RECT 1960.030 4749.350 1960.310 4749.630 ;
        RECT 1960.650 4749.350 1960.930 4749.630 ;
        RECT 1961.270 4749.350 1961.550 4749.630 ;
        RECT 1961.890 4749.350 1962.170 4749.630 ;
        RECT 1962.510 4749.350 1962.790 4749.630 ;
        RECT 1963.130 4749.350 1963.410 4749.630 ;
        RECT 1963.750 4749.350 1964.030 4749.630 ;
        RECT 1964.370 4749.350 1964.650 4749.630 ;
        RECT 1964.990 4749.350 1965.270 4749.630 ;
        RECT 1965.610 4749.350 1965.890 4749.630 ;
        RECT 1969.330 4749.350 1969.610 4749.630 ;
        RECT 1969.950 4749.350 1970.230 4749.630 ;
        RECT 1970.570 4749.350 1970.850 4749.630 ;
        RECT 1971.190 4749.350 1971.470 4749.630 ;
        RECT 1971.810 4749.350 1972.090 4749.630 ;
        RECT 1972.430 4749.350 1972.710 4749.630 ;
        RECT 1973.050 4749.350 1973.330 4749.630 ;
        RECT 1973.670 4749.350 1973.950 4749.630 ;
        RECT 1974.290 4749.350 1974.570 4749.630 ;
        RECT 1974.910 4749.350 1975.190 4749.630 ;
        RECT 1975.530 4749.350 1975.810 4749.630 ;
        RECT 1976.150 4749.350 1976.430 4749.630 ;
        RECT 1976.770 4749.350 1977.050 4749.630 ;
        RECT 1977.390 4749.350 1977.670 4749.630 ;
        RECT 1978.010 4749.350 1978.290 4749.630 ;
        RECT 3006.710 4749.350 3006.990 4749.630 ;
        RECT 3007.330 4749.350 3007.610 4749.630 ;
        RECT 3007.950 4749.350 3008.230 4749.630 ;
        RECT 3008.570 4749.350 3008.850 4749.630 ;
        RECT 3009.190 4749.350 3009.470 4749.630 ;
        RECT 3009.810 4749.350 3010.090 4749.630 ;
        RECT 3010.430 4749.350 3010.710 4749.630 ;
        RECT 3011.050 4749.350 3011.330 4749.630 ;
        RECT 3011.670 4749.350 3011.950 4749.630 ;
        RECT 3012.290 4749.350 3012.570 4749.630 ;
        RECT 3012.910 4749.350 3013.190 4749.630 ;
        RECT 3013.530 4749.350 3013.810 4749.630 ;
        RECT 3014.150 4749.350 3014.430 4749.630 ;
        RECT 3014.770 4749.350 3015.050 4749.630 ;
        RECT 3015.390 4749.350 3015.670 4749.630 ;
        RECT 3019.110 4749.350 3019.390 4749.630 ;
        RECT 3019.730 4749.350 3020.010 4749.630 ;
        RECT 3020.350 4749.350 3020.630 4749.630 ;
        RECT 3020.970 4749.350 3021.250 4749.630 ;
        RECT 3021.590 4749.350 3021.870 4749.630 ;
        RECT 3022.210 4749.350 3022.490 4749.630 ;
        RECT 3022.830 4749.350 3023.110 4749.630 ;
        RECT 3023.450 4749.350 3023.730 4749.630 ;
        RECT 3024.070 4749.350 3024.350 4749.630 ;
        RECT 3024.690 4749.350 3024.970 4749.630 ;
        RECT 3025.310 4749.350 3025.590 4749.630 ;
        RECT 3025.930 4749.350 3026.210 4749.630 ;
        RECT 3026.550 4749.350 3026.830 4749.630 ;
        RECT 3027.170 4749.350 3027.450 4749.630 ;
        RECT 3027.790 4749.350 3028.070 4749.630 ;
        RECT 3028.410 4749.350 3028.690 4749.630 ;
        RECT 3030.960 4749.350 3031.240 4749.630 ;
        RECT 3031.580 4749.350 3031.860 4749.630 ;
        RECT 3032.200 4749.350 3032.480 4749.630 ;
        RECT 3032.820 4749.350 3033.100 4749.630 ;
        RECT 3033.440 4749.350 3033.720 4749.630 ;
        RECT 3034.060 4749.350 3034.340 4749.630 ;
        RECT 3034.680 4749.350 3034.960 4749.630 ;
        RECT 3035.300 4749.350 3035.580 4749.630 ;
        RECT 3035.920 4749.350 3036.200 4749.630 ;
        RECT 3036.540 4749.350 3036.820 4749.630 ;
        RECT 3037.160 4749.350 3037.440 4749.630 ;
        RECT 3037.780 4749.350 3038.060 4749.630 ;
        RECT 3038.400 4749.350 3038.680 4749.630 ;
        RECT 3039.020 4749.350 3039.300 4749.630 ;
        RECT 3039.640 4749.350 3039.920 4749.630 ;
        RECT 3040.260 4749.350 3040.540 4749.630 ;
        RECT 3044.460 4749.350 3044.740 4749.630 ;
        RECT 3045.080 4749.350 3045.360 4749.630 ;
        RECT 3045.700 4749.350 3045.980 4749.630 ;
        RECT 3046.320 4749.350 3046.600 4749.630 ;
        RECT 3046.940 4749.350 3047.220 4749.630 ;
        RECT 3047.560 4749.350 3047.840 4749.630 ;
        RECT 3048.180 4749.350 3048.460 4749.630 ;
        RECT 3048.800 4749.350 3049.080 4749.630 ;
        RECT 3049.420 4749.350 3049.700 4749.630 ;
        RECT 3050.040 4749.350 3050.320 4749.630 ;
        RECT 3050.660 4749.350 3050.940 4749.630 ;
        RECT 3051.280 4749.350 3051.560 4749.630 ;
        RECT 3051.900 4749.350 3052.180 4749.630 ;
        RECT 3052.520 4749.350 3052.800 4749.630 ;
        RECT 3053.140 4749.350 3053.420 4749.630 ;
        RECT 3053.760 4749.350 3054.040 4749.630 ;
        RECT 3056.310 4749.350 3056.590 4749.630 ;
        RECT 3056.930 4749.350 3057.210 4749.630 ;
        RECT 3057.550 4749.350 3057.830 4749.630 ;
        RECT 3058.170 4749.350 3058.450 4749.630 ;
        RECT 3058.790 4749.350 3059.070 4749.630 ;
        RECT 3059.410 4749.350 3059.690 4749.630 ;
        RECT 3060.030 4749.350 3060.310 4749.630 ;
        RECT 3060.650 4749.350 3060.930 4749.630 ;
        RECT 3061.270 4749.350 3061.550 4749.630 ;
        RECT 3061.890 4749.350 3062.170 4749.630 ;
        RECT 3062.510 4749.350 3062.790 4749.630 ;
        RECT 3063.130 4749.350 3063.410 4749.630 ;
        RECT 3063.750 4749.350 3064.030 4749.630 ;
        RECT 3064.370 4749.350 3064.650 4749.630 ;
        RECT 3064.990 4749.350 3065.270 4749.630 ;
        RECT 3065.610 4749.350 3065.890 4749.630 ;
        RECT 3069.330 4749.350 3069.610 4749.630 ;
        RECT 3069.950 4749.350 3070.230 4749.630 ;
        RECT 3070.570 4749.350 3070.850 4749.630 ;
        RECT 3071.190 4749.350 3071.470 4749.630 ;
        RECT 3071.810 4749.350 3072.090 4749.630 ;
        RECT 3072.430 4749.350 3072.710 4749.630 ;
        RECT 3073.050 4749.350 3073.330 4749.630 ;
        RECT 3073.670 4749.350 3073.950 4749.630 ;
        RECT 3074.290 4749.350 3074.570 4749.630 ;
        RECT 3074.910 4749.350 3075.190 4749.630 ;
        RECT 3075.530 4749.350 3075.810 4749.630 ;
        RECT 3076.150 4749.350 3076.430 4749.630 ;
        RECT 3076.770 4749.350 3077.050 4749.630 ;
        RECT 3077.390 4749.350 3077.670 4749.630 ;
        RECT 3078.010 4749.350 3078.290 4749.630 ;
        RECT 350.370 4423.010 350.650 4423.290 ;
        RECT 350.370 4422.390 350.650 4422.670 ;
        RECT 350.370 4421.770 350.650 4422.050 ;
        RECT 350.370 4421.150 350.650 4421.430 ;
        RECT 350.370 4420.530 350.650 4420.810 ;
        RECT 350.370 4419.910 350.650 4420.190 ;
        RECT 350.370 4419.290 350.650 4419.570 ;
        RECT 350.370 4418.670 350.650 4418.950 ;
        RECT 350.370 4418.050 350.650 4418.330 ;
        RECT 350.370 4417.430 350.650 4417.710 ;
        RECT 350.370 4416.810 350.650 4417.090 ;
        RECT 350.370 4416.190 350.650 4416.470 ;
        RECT 350.370 4415.570 350.650 4415.850 ;
        RECT 350.370 4414.950 350.650 4415.230 ;
        RECT 350.370 4414.330 350.650 4414.610 ;
        RECT 3539.350 4418.010 3539.630 4418.290 ;
        RECT 3539.350 4417.390 3539.630 4417.670 ;
        RECT 3539.350 4416.770 3539.630 4417.050 ;
        RECT 3539.350 4416.150 3539.630 4416.430 ;
        RECT 3539.350 4415.530 3539.630 4415.810 ;
        RECT 3539.350 4414.910 3539.630 4415.190 ;
        RECT 3539.350 4414.290 3539.630 4414.570 ;
        RECT 3539.350 4413.670 3539.630 4413.950 ;
        RECT 3539.350 4413.050 3539.630 4413.330 ;
        RECT 3539.350 4412.430 3539.630 4412.710 ;
        RECT 3539.350 4411.810 3539.630 4412.090 ;
        RECT 350.370 4410.640 350.650 4410.920 ;
        RECT 350.370 4410.020 350.650 4410.300 ;
        RECT 350.370 4409.400 350.650 4409.680 ;
        RECT 3539.350 4411.190 3539.630 4411.470 ;
        RECT 3539.350 4410.570 3539.630 4410.850 ;
        RECT 3539.350 4409.950 3539.630 4410.230 ;
        RECT 3539.350 4409.330 3539.630 4409.610 ;
        RECT 350.370 4408.780 350.650 4409.060 ;
        RECT 350.370 4408.160 350.650 4408.440 ;
        RECT 350.370 4407.540 350.650 4407.820 ;
        RECT 350.370 4406.920 350.650 4407.200 ;
        RECT 350.370 4406.300 350.650 4406.580 ;
        RECT 350.370 4405.680 350.650 4405.960 ;
        RECT 350.370 4405.060 350.650 4405.340 ;
        RECT 350.370 4404.440 350.650 4404.720 ;
        RECT 350.370 4403.820 350.650 4404.100 ;
        RECT 350.370 4403.200 350.650 4403.480 ;
        RECT 350.370 4402.580 350.650 4402.860 ;
        RECT 350.370 4401.960 350.650 4402.240 ;
        RECT 350.370 4401.340 350.650 4401.620 ;
        RECT 3539.350 4405.610 3539.630 4405.890 ;
        RECT 3539.350 4404.990 3539.630 4405.270 ;
        RECT 3539.350 4404.370 3539.630 4404.650 ;
        RECT 3539.350 4403.750 3539.630 4404.030 ;
        RECT 3539.350 4403.130 3539.630 4403.410 ;
        RECT 3539.350 4402.510 3539.630 4402.790 ;
        RECT 3539.350 4401.890 3539.630 4402.170 ;
        RECT 3539.350 4401.270 3539.630 4401.550 ;
        RECT 3539.350 4400.650 3539.630 4400.930 ;
        RECT 3539.350 4400.030 3539.630 4400.310 ;
        RECT 3539.350 4399.410 3539.630 4399.690 ;
        RECT 350.370 4398.790 350.650 4399.070 ;
        RECT 350.370 4398.170 350.650 4398.450 ;
        RECT 350.370 4397.550 350.650 4397.830 ;
        RECT 350.370 4396.930 350.650 4397.210 ;
        RECT 350.370 4396.310 350.650 4396.590 ;
        RECT 3539.350 4398.790 3539.630 4399.070 ;
        RECT 3539.350 4398.170 3539.630 4398.450 ;
        RECT 3539.350 4397.550 3539.630 4397.830 ;
        RECT 3539.350 4396.930 3539.630 4397.210 ;
        RECT 3539.350 4396.310 3539.630 4396.590 ;
        RECT 350.370 4395.690 350.650 4395.970 ;
        RECT 350.370 4395.070 350.650 4395.350 ;
        RECT 350.370 4394.450 350.650 4394.730 ;
        RECT 350.370 4393.830 350.650 4394.110 ;
        RECT 350.370 4393.210 350.650 4393.490 ;
        RECT 350.370 4392.590 350.650 4392.870 ;
        RECT 350.370 4391.970 350.650 4392.250 ;
        RECT 350.370 4391.350 350.650 4391.630 ;
        RECT 350.370 4390.730 350.650 4391.010 ;
        RECT 350.370 4390.110 350.650 4390.390 ;
        RECT 350.370 4389.490 350.650 4389.770 ;
        RECT 3539.350 4393.760 3539.630 4394.040 ;
        RECT 3539.350 4393.140 3539.630 4393.420 ;
        RECT 3539.350 4392.520 3539.630 4392.800 ;
        RECT 3539.350 4391.900 3539.630 4392.180 ;
        RECT 3539.350 4391.280 3539.630 4391.560 ;
        RECT 3539.350 4390.660 3539.630 4390.940 ;
        RECT 3539.350 4390.040 3539.630 4390.320 ;
        RECT 3539.350 4389.420 3539.630 4389.700 ;
        RECT 3539.350 4388.800 3539.630 4389.080 ;
        RECT 3539.350 4388.180 3539.630 4388.460 ;
        RECT 3539.350 4387.560 3539.630 4387.840 ;
        RECT 3539.350 4386.940 3539.630 4387.220 ;
        RECT 3539.350 4386.320 3539.630 4386.600 ;
        RECT 350.370 4385.260 350.650 4385.540 ;
        RECT 350.370 4384.640 350.650 4384.920 ;
        RECT 350.370 4384.020 350.650 4384.300 ;
        RECT 3539.350 4385.700 3539.630 4385.980 ;
        RECT 3539.350 4385.080 3539.630 4385.360 ;
        RECT 3539.350 4384.460 3539.630 4384.740 ;
        RECT 350.370 4383.400 350.650 4383.680 ;
        RECT 350.370 4382.780 350.650 4383.060 ;
        RECT 350.370 4382.160 350.650 4382.440 ;
        RECT 350.370 4381.540 350.650 4381.820 ;
        RECT 350.370 4380.920 350.650 4381.200 ;
        RECT 350.370 4380.300 350.650 4380.580 ;
        RECT 350.370 4379.680 350.650 4379.960 ;
        RECT 350.370 4379.060 350.650 4379.340 ;
        RECT 350.370 4378.440 350.650 4378.720 ;
        RECT 350.370 4377.820 350.650 4378.100 ;
        RECT 350.370 4377.200 350.650 4377.480 ;
        RECT 350.370 4376.580 350.650 4376.860 ;
        RECT 350.370 4375.960 350.650 4376.240 ;
        RECT 3539.350 4380.230 3539.630 4380.510 ;
        RECT 3539.350 4379.610 3539.630 4379.890 ;
        RECT 3539.350 4378.990 3539.630 4379.270 ;
        RECT 3539.350 4378.370 3539.630 4378.650 ;
        RECT 3539.350 4377.750 3539.630 4378.030 ;
        RECT 3539.350 4377.130 3539.630 4377.410 ;
        RECT 3539.350 4376.510 3539.630 4376.790 ;
        RECT 3539.350 4375.890 3539.630 4376.170 ;
        RECT 3539.350 4375.270 3539.630 4375.550 ;
        RECT 3539.350 4374.650 3539.630 4374.930 ;
        RECT 3539.350 4374.030 3539.630 4374.310 ;
        RECT 350.370 4373.410 350.650 4373.690 ;
        RECT 350.370 4372.790 350.650 4373.070 ;
        RECT 350.370 4372.170 350.650 4372.450 ;
        RECT 350.370 4371.550 350.650 4371.830 ;
        RECT 350.370 4370.930 350.650 4371.210 ;
        RECT 3539.350 4373.410 3539.630 4373.690 ;
        RECT 3539.350 4372.790 3539.630 4373.070 ;
        RECT 3539.350 4372.170 3539.630 4372.450 ;
        RECT 3539.350 4371.550 3539.630 4371.830 ;
        RECT 3539.350 4370.930 3539.630 4371.210 ;
        RECT 350.370 4370.310 350.650 4370.590 ;
        RECT 350.370 4369.690 350.650 4369.970 ;
        RECT 350.370 4369.070 350.650 4369.350 ;
        RECT 350.370 4368.450 350.650 4368.730 ;
        RECT 350.370 4367.830 350.650 4368.110 ;
        RECT 350.370 4367.210 350.650 4367.490 ;
        RECT 350.370 4366.590 350.650 4366.870 ;
        RECT 350.370 4365.970 350.650 4366.250 ;
        RECT 350.370 4365.350 350.650 4365.630 ;
        RECT 350.370 4364.730 350.650 4365.010 ;
        RECT 350.370 4364.110 350.650 4364.390 ;
        RECT 3539.350 4368.380 3539.630 4368.660 ;
        RECT 3539.350 4367.760 3539.630 4368.040 ;
        RECT 3539.350 4367.140 3539.630 4367.420 ;
        RECT 3539.350 4366.520 3539.630 4366.800 ;
        RECT 3539.350 4365.900 3539.630 4366.180 ;
        RECT 3539.350 4365.280 3539.630 4365.560 ;
        RECT 3539.350 4364.660 3539.630 4364.940 ;
        RECT 3539.350 4364.040 3539.630 4364.320 ;
        RECT 3539.350 4363.420 3539.630 4363.700 ;
        RECT 3539.350 4362.800 3539.630 4363.080 ;
        RECT 3539.350 4362.180 3539.630 4362.460 ;
        RECT 3539.350 4361.560 3539.630 4361.840 ;
        RECT 3539.350 4360.940 3539.630 4361.220 ;
        RECT 350.370 4360.390 350.650 4360.670 ;
        RECT 350.370 4359.770 350.650 4360.050 ;
        RECT 350.370 4359.150 350.650 4359.430 ;
        RECT 350.370 4358.530 350.650 4358.810 ;
        RECT 3539.350 4360.320 3539.630 4360.600 ;
        RECT 3539.350 4359.700 3539.630 4359.980 ;
        RECT 3539.350 4359.080 3539.630 4359.360 ;
        RECT 350.370 4357.910 350.650 4358.190 ;
        RECT 350.370 4357.290 350.650 4357.570 ;
        RECT 350.370 4356.670 350.650 4356.950 ;
        RECT 350.370 4356.050 350.650 4356.330 ;
        RECT 350.370 4355.430 350.650 4355.710 ;
        RECT 350.370 4354.810 350.650 4355.090 ;
        RECT 350.370 4354.190 350.650 4354.470 ;
        RECT 350.370 4353.570 350.650 4353.850 ;
        RECT 350.370 4352.950 350.650 4353.230 ;
        RECT 350.370 4352.330 350.650 4352.610 ;
        RECT 350.370 4351.710 350.650 4351.990 ;
        RECT 3539.350 4355.390 3539.630 4355.670 ;
        RECT 3539.350 4354.770 3539.630 4355.050 ;
        RECT 3539.350 4354.150 3539.630 4354.430 ;
        RECT 3539.350 4353.530 3539.630 4353.810 ;
        RECT 3539.350 4352.910 3539.630 4353.190 ;
        RECT 3539.350 4352.290 3539.630 4352.570 ;
        RECT 3539.350 4351.670 3539.630 4351.950 ;
        RECT 3539.350 4351.050 3539.630 4351.330 ;
        RECT 3539.350 4350.430 3539.630 4350.710 ;
        RECT 3539.350 4349.810 3539.630 4350.090 ;
        RECT 3539.350 4349.190 3539.630 4349.470 ;
        RECT 3539.350 4348.570 3539.630 4348.850 ;
        RECT 3539.350 4347.950 3539.630 4348.230 ;
        RECT 3539.350 4347.330 3539.630 4347.610 ;
        RECT 3539.350 4346.710 3539.630 4346.990 ;
        RECT 350.370 4218.010 350.650 4218.290 ;
        RECT 350.370 4217.390 350.650 4217.670 ;
        RECT 350.370 4216.770 350.650 4217.050 ;
        RECT 350.370 4216.150 350.650 4216.430 ;
        RECT 350.370 4215.530 350.650 4215.810 ;
        RECT 350.370 4214.910 350.650 4215.190 ;
        RECT 350.370 4214.290 350.650 4214.570 ;
        RECT 350.370 4213.670 350.650 4213.950 ;
        RECT 350.370 4213.050 350.650 4213.330 ;
        RECT 350.370 4212.430 350.650 4212.710 ;
        RECT 350.370 4211.810 350.650 4212.090 ;
        RECT 350.370 4211.190 350.650 4211.470 ;
        RECT 350.370 4210.570 350.650 4210.850 ;
        RECT 350.370 4209.950 350.650 4210.230 ;
        RECT 350.370 4209.330 350.650 4209.610 ;
        RECT 350.370 4205.640 350.650 4205.920 ;
        RECT 350.370 4205.020 350.650 4205.300 ;
        RECT 350.370 4204.400 350.650 4204.680 ;
        RECT 350.370 4203.780 350.650 4204.060 ;
        RECT 350.370 4203.160 350.650 4203.440 ;
        RECT 350.370 4202.540 350.650 4202.820 ;
        RECT 350.370 4201.920 350.650 4202.200 ;
        RECT 350.370 4201.300 350.650 4201.580 ;
        RECT 350.370 4200.680 350.650 4200.960 ;
        RECT 350.370 4200.060 350.650 4200.340 ;
        RECT 350.370 4199.440 350.650 4199.720 ;
        RECT 350.370 4198.820 350.650 4199.100 ;
        RECT 350.370 4198.200 350.650 4198.480 ;
        RECT 350.370 4197.580 350.650 4197.860 ;
        RECT 350.370 4196.960 350.650 4197.240 ;
        RECT 350.370 4196.340 350.650 4196.620 ;
        RECT 350.370 4193.790 350.650 4194.070 ;
        RECT 350.370 4193.170 350.650 4193.450 ;
        RECT 350.370 4192.550 350.650 4192.830 ;
        RECT 350.370 4191.930 350.650 4192.210 ;
        RECT 350.370 4191.310 350.650 4191.590 ;
        RECT 350.370 4190.690 350.650 4190.970 ;
        RECT 350.370 4190.070 350.650 4190.350 ;
        RECT 350.370 4189.450 350.650 4189.730 ;
        RECT 350.370 4188.830 350.650 4189.110 ;
        RECT 350.370 4188.210 350.650 4188.490 ;
        RECT 350.370 4187.590 350.650 4187.870 ;
        RECT 350.370 4186.970 350.650 4187.250 ;
        RECT 350.370 4186.350 350.650 4186.630 ;
        RECT 350.370 4185.730 350.650 4186.010 ;
        RECT 350.370 4185.110 350.650 4185.390 ;
        RECT 350.370 4184.490 350.650 4184.770 ;
        RECT 350.370 4180.260 350.650 4180.540 ;
        RECT 350.370 4179.640 350.650 4179.920 ;
        RECT 350.370 4179.020 350.650 4179.300 ;
        RECT 350.370 4178.400 350.650 4178.680 ;
        RECT 350.370 4177.780 350.650 4178.060 ;
        RECT 350.370 4177.160 350.650 4177.440 ;
        RECT 350.370 4176.540 350.650 4176.820 ;
        RECT 350.370 4175.920 350.650 4176.200 ;
        RECT 350.370 4175.300 350.650 4175.580 ;
        RECT 350.370 4174.680 350.650 4174.960 ;
        RECT 350.370 4174.060 350.650 4174.340 ;
        RECT 350.370 4173.440 350.650 4173.720 ;
        RECT 350.370 4172.820 350.650 4173.100 ;
        RECT 350.370 4172.200 350.650 4172.480 ;
        RECT 350.370 4171.580 350.650 4171.860 ;
        RECT 350.370 4170.960 350.650 4171.240 ;
        RECT 350.370 4168.410 350.650 4168.690 ;
        RECT 350.370 4167.790 350.650 4168.070 ;
        RECT 350.370 4167.170 350.650 4167.450 ;
        RECT 350.370 4166.550 350.650 4166.830 ;
        RECT 350.370 4165.930 350.650 4166.210 ;
        RECT 350.370 4165.310 350.650 4165.590 ;
        RECT 350.370 4164.690 350.650 4164.970 ;
        RECT 350.370 4164.070 350.650 4164.350 ;
        RECT 350.370 4163.450 350.650 4163.730 ;
        RECT 350.370 4162.830 350.650 4163.110 ;
        RECT 350.370 4162.210 350.650 4162.490 ;
        RECT 350.370 4161.590 350.650 4161.870 ;
        RECT 350.370 4160.970 350.650 4161.250 ;
        RECT 350.370 4160.350 350.650 4160.630 ;
        RECT 350.370 4159.730 350.650 4160.010 ;
        RECT 350.370 4159.110 350.650 4159.390 ;
        RECT 350.370 4155.390 350.650 4155.670 ;
        RECT 350.370 4154.770 350.650 4155.050 ;
        RECT 350.370 4154.150 350.650 4154.430 ;
        RECT 350.370 4153.530 350.650 4153.810 ;
        RECT 350.370 4152.910 350.650 4153.190 ;
        RECT 350.370 4152.290 350.650 4152.570 ;
        RECT 350.370 4151.670 350.650 4151.950 ;
        RECT 350.370 4151.050 350.650 4151.330 ;
        RECT 350.370 4150.430 350.650 4150.710 ;
        RECT 350.370 4149.810 350.650 4150.090 ;
        RECT 350.370 4149.190 350.650 4149.470 ;
        RECT 350.370 4148.570 350.650 4148.850 ;
        RECT 350.370 4147.950 350.650 4148.230 ;
        RECT 350.370 4147.330 350.650 4147.610 ;
        RECT 350.370 4146.710 350.650 4146.990 ;
        RECT 350.370 4013.010 350.650 4013.290 ;
        RECT 350.370 4012.390 350.650 4012.670 ;
        RECT 350.370 4011.770 350.650 4012.050 ;
        RECT 350.370 4011.150 350.650 4011.430 ;
        RECT 350.370 4010.530 350.650 4010.810 ;
        RECT 350.370 4009.910 350.650 4010.190 ;
        RECT 350.370 4009.290 350.650 4009.570 ;
        RECT 350.370 4008.670 350.650 4008.950 ;
        RECT 350.370 4008.050 350.650 4008.330 ;
        RECT 350.370 4007.430 350.650 4007.710 ;
        RECT 350.370 4006.810 350.650 4007.090 ;
        RECT 350.370 4006.190 350.650 4006.470 ;
        RECT 350.370 4005.570 350.650 4005.850 ;
        RECT 350.370 4004.950 350.650 4005.230 ;
        RECT 350.370 4004.330 350.650 4004.610 ;
        RECT 350.370 4000.640 350.650 4000.920 ;
        RECT 350.370 4000.020 350.650 4000.300 ;
        RECT 350.370 3999.400 350.650 3999.680 ;
        RECT 350.370 3998.780 350.650 3999.060 ;
        RECT 350.370 3998.160 350.650 3998.440 ;
        RECT 350.370 3997.540 350.650 3997.820 ;
        RECT 350.370 3996.920 350.650 3997.200 ;
        RECT 350.370 3996.300 350.650 3996.580 ;
        RECT 350.370 3995.680 350.650 3995.960 ;
        RECT 350.370 3995.060 350.650 3995.340 ;
        RECT 350.370 3994.440 350.650 3994.720 ;
        RECT 350.370 3993.820 350.650 3994.100 ;
        RECT 350.370 3993.200 350.650 3993.480 ;
        RECT 350.370 3992.580 350.650 3992.860 ;
        RECT 350.370 3991.960 350.650 3992.240 ;
        RECT 350.370 3991.340 350.650 3991.620 ;
        RECT 350.370 3988.790 350.650 3989.070 ;
        RECT 350.370 3988.170 350.650 3988.450 ;
        RECT 350.370 3987.550 350.650 3987.830 ;
        RECT 350.370 3986.930 350.650 3987.210 ;
        RECT 350.370 3986.310 350.650 3986.590 ;
        RECT 350.370 3985.690 350.650 3985.970 ;
        RECT 350.370 3985.070 350.650 3985.350 ;
        RECT 350.370 3984.450 350.650 3984.730 ;
        RECT 350.370 3983.830 350.650 3984.110 ;
        RECT 350.370 3983.210 350.650 3983.490 ;
        RECT 350.370 3982.590 350.650 3982.870 ;
        RECT 350.370 3981.970 350.650 3982.250 ;
        RECT 350.370 3981.350 350.650 3981.630 ;
        RECT 350.370 3980.730 350.650 3981.010 ;
        RECT 350.370 3980.110 350.650 3980.390 ;
        RECT 350.370 3979.490 350.650 3979.770 ;
        RECT 3539.350 3988.010 3539.630 3988.290 ;
        RECT 3539.350 3987.390 3539.630 3987.670 ;
        RECT 3539.350 3986.770 3539.630 3987.050 ;
        RECT 3539.350 3986.150 3539.630 3986.430 ;
        RECT 3539.350 3985.530 3539.630 3985.810 ;
        RECT 3539.350 3984.910 3539.630 3985.190 ;
        RECT 3539.350 3984.290 3539.630 3984.570 ;
        RECT 3539.350 3983.670 3539.630 3983.950 ;
        RECT 3539.350 3983.050 3539.630 3983.330 ;
        RECT 3539.350 3982.430 3539.630 3982.710 ;
        RECT 3539.350 3981.810 3539.630 3982.090 ;
        RECT 3539.350 3981.190 3539.630 3981.470 ;
        RECT 3539.350 3980.570 3539.630 3980.850 ;
        RECT 3539.350 3979.950 3539.630 3980.230 ;
        RECT 3539.350 3979.330 3539.630 3979.610 ;
        RECT 350.370 3975.260 350.650 3975.540 ;
        RECT 350.370 3974.640 350.650 3974.920 ;
        RECT 350.370 3974.020 350.650 3974.300 ;
        RECT 350.370 3973.400 350.650 3973.680 ;
        RECT 350.370 3972.780 350.650 3973.060 ;
        RECT 350.370 3972.160 350.650 3972.440 ;
        RECT 350.370 3971.540 350.650 3971.820 ;
        RECT 350.370 3970.920 350.650 3971.200 ;
        RECT 350.370 3970.300 350.650 3970.580 ;
        RECT 350.370 3969.680 350.650 3969.960 ;
        RECT 350.370 3969.060 350.650 3969.340 ;
        RECT 350.370 3968.440 350.650 3968.720 ;
        RECT 350.370 3967.820 350.650 3968.100 ;
        RECT 350.370 3967.200 350.650 3967.480 ;
        RECT 350.370 3966.580 350.650 3966.860 ;
        RECT 350.370 3965.960 350.650 3966.240 ;
        RECT 3539.350 3975.610 3539.630 3975.890 ;
        RECT 3539.350 3974.990 3539.630 3975.270 ;
        RECT 3539.350 3974.370 3539.630 3974.650 ;
        RECT 3539.350 3973.750 3539.630 3974.030 ;
        RECT 3539.350 3973.130 3539.630 3973.410 ;
        RECT 3539.350 3972.510 3539.630 3972.790 ;
        RECT 3539.350 3971.890 3539.630 3972.170 ;
        RECT 3539.350 3971.270 3539.630 3971.550 ;
        RECT 3539.350 3970.650 3539.630 3970.930 ;
        RECT 3539.350 3970.030 3539.630 3970.310 ;
        RECT 3539.350 3969.410 3539.630 3969.690 ;
        RECT 3539.350 3968.790 3539.630 3969.070 ;
        RECT 3539.350 3968.170 3539.630 3968.450 ;
        RECT 3539.350 3967.550 3539.630 3967.830 ;
        RECT 3539.350 3966.930 3539.630 3967.210 ;
        RECT 3539.350 3966.310 3539.630 3966.590 ;
        RECT 350.370 3963.410 350.650 3963.690 ;
        RECT 350.370 3962.790 350.650 3963.070 ;
        RECT 350.370 3962.170 350.650 3962.450 ;
        RECT 350.370 3961.550 350.650 3961.830 ;
        RECT 350.370 3960.930 350.650 3961.210 ;
        RECT 350.370 3960.310 350.650 3960.590 ;
        RECT 350.370 3959.690 350.650 3959.970 ;
        RECT 350.370 3959.070 350.650 3959.350 ;
        RECT 350.370 3958.450 350.650 3958.730 ;
        RECT 350.370 3957.830 350.650 3958.110 ;
        RECT 350.370 3957.210 350.650 3957.490 ;
        RECT 350.370 3956.590 350.650 3956.870 ;
        RECT 350.370 3955.970 350.650 3956.250 ;
        RECT 350.370 3955.350 350.650 3955.630 ;
        RECT 350.370 3954.730 350.650 3955.010 ;
        RECT 350.370 3954.110 350.650 3954.390 ;
        RECT 3539.350 3963.760 3539.630 3964.040 ;
        RECT 3539.350 3963.140 3539.630 3963.420 ;
        RECT 3539.350 3962.520 3539.630 3962.800 ;
        RECT 3539.350 3961.900 3539.630 3962.180 ;
        RECT 3539.350 3961.280 3539.630 3961.560 ;
        RECT 3539.350 3960.660 3539.630 3960.940 ;
        RECT 3539.350 3960.040 3539.630 3960.320 ;
        RECT 3539.350 3959.420 3539.630 3959.700 ;
        RECT 3539.350 3958.800 3539.630 3959.080 ;
        RECT 3539.350 3958.180 3539.630 3958.460 ;
        RECT 3539.350 3957.560 3539.630 3957.840 ;
        RECT 3539.350 3956.940 3539.630 3957.220 ;
        RECT 3539.350 3956.320 3539.630 3956.600 ;
        RECT 3539.350 3955.700 3539.630 3955.980 ;
        RECT 3539.350 3955.080 3539.630 3955.360 ;
        RECT 3539.350 3954.460 3539.630 3954.740 ;
        RECT 350.370 3950.390 350.650 3950.670 ;
        RECT 350.370 3949.770 350.650 3950.050 ;
        RECT 350.370 3949.150 350.650 3949.430 ;
        RECT 350.370 3948.530 350.650 3948.810 ;
        RECT 350.370 3947.910 350.650 3948.190 ;
        RECT 350.370 3947.290 350.650 3947.570 ;
        RECT 350.370 3946.670 350.650 3946.950 ;
        RECT 350.370 3946.050 350.650 3946.330 ;
        RECT 350.370 3945.430 350.650 3945.710 ;
        RECT 350.370 3944.810 350.650 3945.090 ;
        RECT 350.370 3944.190 350.650 3944.470 ;
        RECT 350.370 3943.570 350.650 3943.850 ;
        RECT 350.370 3942.950 350.650 3943.230 ;
        RECT 350.370 3942.330 350.650 3942.610 ;
        RECT 350.370 3941.710 350.650 3941.990 ;
        RECT 3539.350 3950.230 3539.630 3950.510 ;
        RECT 3539.350 3949.610 3539.630 3949.890 ;
        RECT 3539.350 3948.990 3539.630 3949.270 ;
        RECT 3539.350 3948.370 3539.630 3948.650 ;
        RECT 3539.350 3947.750 3539.630 3948.030 ;
        RECT 3539.350 3947.130 3539.630 3947.410 ;
        RECT 3539.350 3946.510 3539.630 3946.790 ;
        RECT 3539.350 3945.890 3539.630 3946.170 ;
        RECT 3539.350 3945.270 3539.630 3945.550 ;
        RECT 3539.350 3944.650 3539.630 3944.930 ;
        RECT 3539.350 3944.030 3539.630 3944.310 ;
        RECT 3539.350 3943.410 3539.630 3943.690 ;
        RECT 3539.350 3942.790 3539.630 3943.070 ;
        RECT 3539.350 3942.170 3539.630 3942.450 ;
        RECT 3539.350 3941.550 3539.630 3941.830 ;
        RECT 3539.350 3940.930 3539.630 3941.210 ;
        RECT 3539.350 3938.380 3539.630 3938.660 ;
        RECT 3539.350 3937.760 3539.630 3938.040 ;
        RECT 3539.350 3937.140 3539.630 3937.420 ;
        RECT 3539.350 3936.520 3539.630 3936.800 ;
        RECT 3539.350 3935.900 3539.630 3936.180 ;
        RECT 3539.350 3935.280 3539.630 3935.560 ;
        RECT 3539.350 3934.660 3539.630 3934.940 ;
        RECT 3539.350 3934.040 3539.630 3934.320 ;
        RECT 3539.350 3933.420 3539.630 3933.700 ;
        RECT 3539.350 3932.800 3539.630 3933.080 ;
        RECT 3539.350 3932.180 3539.630 3932.460 ;
        RECT 3539.350 3931.560 3539.630 3931.840 ;
        RECT 3539.350 3930.940 3539.630 3931.220 ;
        RECT 3539.350 3930.320 3539.630 3930.600 ;
        RECT 3539.350 3929.700 3539.630 3929.980 ;
        RECT 3539.350 3929.080 3539.630 3929.360 ;
        RECT 3539.350 3925.390 3539.630 3925.670 ;
        RECT 3539.350 3924.770 3539.630 3925.050 ;
        RECT 3539.350 3924.150 3539.630 3924.430 ;
        RECT 3539.350 3923.530 3539.630 3923.810 ;
        RECT 3539.350 3922.910 3539.630 3923.190 ;
        RECT 3539.350 3922.290 3539.630 3922.570 ;
        RECT 3539.350 3921.670 3539.630 3921.950 ;
        RECT 3539.350 3921.050 3539.630 3921.330 ;
        RECT 3539.350 3920.430 3539.630 3920.710 ;
        RECT 3539.350 3919.810 3539.630 3920.090 ;
        RECT 3539.350 3919.190 3539.630 3919.470 ;
        RECT 3539.350 3918.570 3539.630 3918.850 ;
        RECT 3539.350 3917.950 3539.630 3918.230 ;
        RECT 3539.350 3917.330 3539.630 3917.610 ;
        RECT 3539.350 3916.710 3539.630 3916.990 ;
        RECT 3539.350 2483.010 3539.630 2483.290 ;
        RECT 3539.350 2482.390 3539.630 2482.670 ;
        RECT 3539.350 2481.770 3539.630 2482.050 ;
        RECT 3539.350 2481.150 3539.630 2481.430 ;
        RECT 3539.350 2480.530 3539.630 2480.810 ;
        RECT 3539.350 2479.910 3539.630 2480.190 ;
        RECT 3539.350 2479.290 3539.630 2479.570 ;
        RECT 3539.350 2478.670 3539.630 2478.950 ;
        RECT 3539.350 2478.050 3539.630 2478.330 ;
        RECT 3539.350 2477.430 3539.630 2477.710 ;
        RECT 3539.350 2476.810 3539.630 2477.090 ;
        RECT 3539.350 2476.190 3539.630 2476.470 ;
        RECT 3539.350 2475.570 3539.630 2475.850 ;
        RECT 3539.350 2474.950 3539.630 2475.230 ;
        RECT 3539.350 2474.330 3539.630 2474.610 ;
        RECT 3539.350 2470.610 3539.630 2470.890 ;
        RECT 3539.350 2469.990 3539.630 2470.270 ;
        RECT 3539.350 2469.370 3539.630 2469.650 ;
        RECT 3539.350 2468.750 3539.630 2469.030 ;
        RECT 3539.350 2468.130 3539.630 2468.410 ;
        RECT 3539.350 2467.510 3539.630 2467.790 ;
        RECT 3539.350 2466.890 3539.630 2467.170 ;
        RECT 3539.350 2466.270 3539.630 2466.550 ;
        RECT 3539.350 2465.650 3539.630 2465.930 ;
        RECT 3539.350 2465.030 3539.630 2465.310 ;
        RECT 3539.350 2464.410 3539.630 2464.690 ;
        RECT 3539.350 2463.790 3539.630 2464.070 ;
        RECT 3539.350 2463.170 3539.630 2463.450 ;
        RECT 3539.350 2462.550 3539.630 2462.830 ;
        RECT 3539.350 2461.930 3539.630 2462.210 ;
        RECT 3539.350 2461.310 3539.630 2461.590 ;
        RECT 3539.350 2458.760 3539.630 2459.040 ;
        RECT 3539.350 2458.140 3539.630 2458.420 ;
        RECT 3539.350 2457.520 3539.630 2457.800 ;
        RECT 3539.350 2456.900 3539.630 2457.180 ;
        RECT 3539.350 2456.280 3539.630 2456.560 ;
        RECT 3539.350 2455.660 3539.630 2455.940 ;
        RECT 3539.350 2455.040 3539.630 2455.320 ;
        RECT 3539.350 2454.420 3539.630 2454.700 ;
        RECT 3539.350 2453.800 3539.630 2454.080 ;
        RECT 3539.350 2453.180 3539.630 2453.460 ;
        RECT 3539.350 2452.560 3539.630 2452.840 ;
        RECT 3539.350 2451.940 3539.630 2452.220 ;
        RECT 3539.350 2451.320 3539.630 2451.600 ;
        RECT 3539.350 2450.700 3539.630 2450.980 ;
        RECT 3539.350 2450.080 3539.630 2450.360 ;
        RECT 3539.350 2449.460 3539.630 2449.740 ;
        RECT 3539.350 2445.230 3539.630 2445.510 ;
        RECT 3539.350 2444.610 3539.630 2444.890 ;
        RECT 3539.350 2443.990 3539.630 2444.270 ;
        RECT 3539.350 2443.370 3539.630 2443.650 ;
        RECT 3539.350 2442.750 3539.630 2443.030 ;
        RECT 3539.350 2442.130 3539.630 2442.410 ;
        RECT 3539.350 2441.510 3539.630 2441.790 ;
        RECT 3539.350 2440.890 3539.630 2441.170 ;
        RECT 3539.350 2440.270 3539.630 2440.550 ;
        RECT 3539.350 2439.650 3539.630 2439.930 ;
        RECT 3539.350 2439.030 3539.630 2439.310 ;
        RECT 3539.350 2438.410 3539.630 2438.690 ;
        RECT 3539.350 2437.790 3539.630 2438.070 ;
        RECT 3539.350 2437.170 3539.630 2437.450 ;
        RECT 3539.350 2436.550 3539.630 2436.830 ;
        RECT 3539.350 2435.930 3539.630 2436.210 ;
        RECT 3539.350 2433.380 3539.630 2433.660 ;
        RECT 3539.350 2432.760 3539.630 2433.040 ;
        RECT 3539.350 2432.140 3539.630 2432.420 ;
        RECT 3539.350 2431.520 3539.630 2431.800 ;
        RECT 3539.350 2430.900 3539.630 2431.180 ;
        RECT 3539.350 2430.280 3539.630 2430.560 ;
        RECT 3539.350 2429.660 3539.630 2429.940 ;
        RECT 3539.350 2429.040 3539.630 2429.320 ;
        RECT 3539.350 2428.420 3539.630 2428.700 ;
        RECT 3539.350 2427.800 3539.630 2428.080 ;
        RECT 3539.350 2427.180 3539.630 2427.460 ;
        RECT 3539.350 2426.560 3539.630 2426.840 ;
        RECT 3539.350 2425.940 3539.630 2426.220 ;
        RECT 3539.350 2425.320 3539.630 2425.600 ;
        RECT 3539.350 2424.700 3539.630 2424.980 ;
        RECT 3539.350 2424.080 3539.630 2424.360 ;
        RECT 3539.350 2420.390 3539.630 2420.670 ;
        RECT 3539.350 2419.770 3539.630 2420.050 ;
        RECT 3539.350 2419.150 3539.630 2419.430 ;
        RECT 3539.350 2418.530 3539.630 2418.810 ;
        RECT 3539.350 2417.910 3539.630 2418.190 ;
        RECT 3539.350 2417.290 3539.630 2417.570 ;
        RECT 3539.350 2416.670 3539.630 2416.950 ;
        RECT 3539.350 2416.050 3539.630 2416.330 ;
        RECT 3539.350 2415.430 3539.630 2415.710 ;
        RECT 3539.350 2414.810 3539.630 2415.090 ;
        RECT 3539.350 2414.190 3539.630 2414.470 ;
        RECT 3539.350 2413.570 3539.630 2413.850 ;
        RECT 3539.350 2412.950 3539.630 2413.230 ;
        RECT 3539.350 2412.330 3539.630 2412.610 ;
        RECT 3539.350 2411.710 3539.630 2411.990 ;
        RECT 350.370 2373.010 350.650 2373.290 ;
        RECT 350.370 2372.390 350.650 2372.670 ;
        RECT 350.370 2371.770 350.650 2372.050 ;
        RECT 350.370 2371.150 350.650 2371.430 ;
        RECT 350.370 2370.530 350.650 2370.810 ;
        RECT 350.370 2369.910 350.650 2370.190 ;
        RECT 350.370 2369.290 350.650 2369.570 ;
        RECT 350.370 2368.670 350.650 2368.950 ;
        RECT 350.370 2368.050 350.650 2368.330 ;
        RECT 350.370 2367.430 350.650 2367.710 ;
        RECT 350.370 2366.810 350.650 2367.090 ;
        RECT 350.370 2366.190 350.650 2366.470 ;
        RECT 350.370 2365.570 350.650 2365.850 ;
        RECT 350.370 2364.950 350.650 2365.230 ;
        RECT 350.370 2364.330 350.650 2364.610 ;
        RECT 350.370 2360.640 350.650 2360.920 ;
        RECT 350.370 2360.020 350.650 2360.300 ;
        RECT 350.370 2359.400 350.650 2359.680 ;
        RECT 350.370 2358.780 350.650 2359.060 ;
        RECT 350.370 2358.160 350.650 2358.440 ;
        RECT 350.370 2357.540 350.650 2357.820 ;
        RECT 350.370 2356.920 350.650 2357.200 ;
        RECT 350.370 2356.300 350.650 2356.580 ;
        RECT 350.370 2355.680 350.650 2355.960 ;
        RECT 350.370 2355.060 350.650 2355.340 ;
        RECT 350.370 2354.440 350.650 2354.720 ;
        RECT 350.370 2353.820 350.650 2354.100 ;
        RECT 350.370 2353.200 350.650 2353.480 ;
        RECT 350.370 2352.580 350.650 2352.860 ;
        RECT 350.370 2351.960 350.650 2352.240 ;
        RECT 350.370 2351.340 350.650 2351.620 ;
        RECT 350.370 2348.790 350.650 2349.070 ;
        RECT 350.370 2348.170 350.650 2348.450 ;
        RECT 350.370 2347.550 350.650 2347.830 ;
        RECT 350.370 2346.930 350.650 2347.210 ;
        RECT 350.370 2346.310 350.650 2346.590 ;
        RECT 350.370 2345.690 350.650 2345.970 ;
        RECT 350.370 2345.070 350.650 2345.350 ;
        RECT 350.370 2344.450 350.650 2344.730 ;
        RECT 350.370 2343.830 350.650 2344.110 ;
        RECT 350.370 2343.210 350.650 2343.490 ;
        RECT 350.370 2342.590 350.650 2342.870 ;
        RECT 350.370 2341.970 350.650 2342.250 ;
        RECT 350.370 2341.350 350.650 2341.630 ;
        RECT 350.370 2340.730 350.650 2341.010 ;
        RECT 350.370 2340.110 350.650 2340.390 ;
        RECT 350.370 2339.490 350.650 2339.770 ;
        RECT 350.370 2335.260 350.650 2335.540 ;
        RECT 350.370 2334.640 350.650 2334.920 ;
        RECT 350.370 2334.020 350.650 2334.300 ;
        RECT 350.370 2333.400 350.650 2333.680 ;
        RECT 350.370 2332.780 350.650 2333.060 ;
        RECT 350.370 2332.160 350.650 2332.440 ;
        RECT 350.370 2331.540 350.650 2331.820 ;
        RECT 350.370 2330.920 350.650 2331.200 ;
        RECT 350.370 2330.300 350.650 2330.580 ;
        RECT 350.370 2329.680 350.650 2329.960 ;
        RECT 350.370 2329.060 350.650 2329.340 ;
        RECT 350.370 2328.440 350.650 2328.720 ;
        RECT 350.370 2327.820 350.650 2328.100 ;
        RECT 350.370 2327.200 350.650 2327.480 ;
        RECT 350.370 2326.580 350.650 2326.860 ;
        RECT 350.370 2325.960 350.650 2326.240 ;
        RECT 350.370 2323.410 350.650 2323.690 ;
        RECT 350.370 2322.790 350.650 2323.070 ;
        RECT 350.370 2322.170 350.650 2322.450 ;
        RECT 350.370 2321.550 350.650 2321.830 ;
        RECT 350.370 2320.930 350.650 2321.210 ;
        RECT 350.370 2320.310 350.650 2320.590 ;
        RECT 350.370 2319.690 350.650 2319.970 ;
        RECT 350.370 2319.070 350.650 2319.350 ;
        RECT 350.370 2318.450 350.650 2318.730 ;
        RECT 350.370 2317.830 350.650 2318.110 ;
        RECT 350.370 2317.210 350.650 2317.490 ;
        RECT 350.370 2316.590 350.650 2316.870 ;
        RECT 350.370 2315.970 350.650 2316.250 ;
        RECT 350.370 2315.350 350.650 2315.630 ;
        RECT 350.370 2314.730 350.650 2315.010 ;
        RECT 350.370 2314.110 350.650 2314.390 ;
        RECT 350.370 2310.390 350.650 2310.670 ;
        RECT 350.370 2309.770 350.650 2310.050 ;
        RECT 350.370 2309.150 350.650 2309.430 ;
        RECT 350.370 2308.530 350.650 2308.810 ;
        RECT 350.370 2307.910 350.650 2308.190 ;
        RECT 350.370 2307.290 350.650 2307.570 ;
        RECT 350.370 2306.670 350.650 2306.950 ;
        RECT 350.370 2306.050 350.650 2306.330 ;
        RECT 350.370 2305.430 350.650 2305.710 ;
        RECT 350.370 2304.810 350.650 2305.090 ;
        RECT 350.370 2304.190 350.650 2304.470 ;
        RECT 350.370 2303.570 350.650 2303.850 ;
        RECT 350.370 2302.950 350.650 2303.230 ;
        RECT 350.370 2302.330 350.650 2302.610 ;
        RECT 350.370 2301.710 350.650 2301.990 ;
        RECT 3539.350 2268.010 3539.630 2268.290 ;
        RECT 3539.350 2267.390 3539.630 2267.670 ;
        RECT 3539.350 2266.770 3539.630 2267.050 ;
        RECT 3539.350 2266.150 3539.630 2266.430 ;
        RECT 3539.350 2265.530 3539.630 2265.810 ;
        RECT 3539.350 2264.910 3539.630 2265.190 ;
        RECT 3539.350 2264.290 3539.630 2264.570 ;
        RECT 3539.350 2263.670 3539.630 2263.950 ;
        RECT 3539.350 2263.050 3539.630 2263.330 ;
        RECT 3539.350 2262.430 3539.630 2262.710 ;
        RECT 3539.350 2261.810 3539.630 2262.090 ;
        RECT 3539.350 2261.190 3539.630 2261.470 ;
        RECT 3539.350 2260.570 3539.630 2260.850 ;
        RECT 3539.350 2259.950 3539.630 2260.230 ;
        RECT 3539.350 2259.330 3539.630 2259.610 ;
        RECT 3539.350 2255.610 3539.630 2255.890 ;
        RECT 3539.350 2254.990 3539.630 2255.270 ;
        RECT 3539.350 2254.370 3539.630 2254.650 ;
        RECT 3539.350 2253.750 3539.630 2254.030 ;
        RECT 3539.350 2253.130 3539.630 2253.410 ;
        RECT 3539.350 2252.510 3539.630 2252.790 ;
        RECT 3539.350 2251.890 3539.630 2252.170 ;
        RECT 3539.350 2251.270 3539.630 2251.550 ;
        RECT 3539.350 2250.650 3539.630 2250.930 ;
        RECT 3539.350 2250.030 3539.630 2250.310 ;
        RECT 3539.350 2249.410 3539.630 2249.690 ;
        RECT 3539.350 2248.790 3539.630 2249.070 ;
        RECT 3539.350 2248.170 3539.630 2248.450 ;
        RECT 3539.350 2247.550 3539.630 2247.830 ;
        RECT 3539.350 2246.930 3539.630 2247.210 ;
        RECT 3539.350 2246.310 3539.630 2246.590 ;
        RECT 3539.350 2243.760 3539.630 2244.040 ;
        RECT 3539.350 2243.140 3539.630 2243.420 ;
        RECT 3539.350 2242.520 3539.630 2242.800 ;
        RECT 3539.350 2241.900 3539.630 2242.180 ;
        RECT 3539.350 2241.280 3539.630 2241.560 ;
        RECT 3539.350 2240.660 3539.630 2240.940 ;
        RECT 3539.350 2240.040 3539.630 2240.320 ;
        RECT 3539.350 2239.420 3539.630 2239.700 ;
        RECT 3539.350 2238.800 3539.630 2239.080 ;
        RECT 3539.350 2238.180 3539.630 2238.460 ;
        RECT 3539.350 2237.560 3539.630 2237.840 ;
        RECT 3539.350 2236.940 3539.630 2237.220 ;
        RECT 3539.350 2236.320 3539.630 2236.600 ;
        RECT 3539.350 2235.700 3539.630 2235.980 ;
        RECT 3539.350 2235.080 3539.630 2235.360 ;
        RECT 3539.350 2234.460 3539.630 2234.740 ;
        RECT 3539.350 2230.230 3539.630 2230.510 ;
        RECT 3539.350 2229.610 3539.630 2229.890 ;
        RECT 3539.350 2228.990 3539.630 2229.270 ;
        RECT 3539.350 2228.370 3539.630 2228.650 ;
        RECT 3539.350 2227.750 3539.630 2228.030 ;
        RECT 3539.350 2227.130 3539.630 2227.410 ;
        RECT 3539.350 2226.510 3539.630 2226.790 ;
        RECT 3539.350 2225.890 3539.630 2226.170 ;
        RECT 3539.350 2225.270 3539.630 2225.550 ;
        RECT 3539.350 2224.650 3539.630 2224.930 ;
        RECT 3539.350 2224.030 3539.630 2224.310 ;
        RECT 3539.350 2223.410 3539.630 2223.690 ;
        RECT 3539.350 2222.790 3539.630 2223.070 ;
        RECT 3539.350 2222.170 3539.630 2222.450 ;
        RECT 3539.350 2221.550 3539.630 2221.830 ;
        RECT 3539.350 2220.930 3539.630 2221.210 ;
        RECT 3539.350 2218.380 3539.630 2218.660 ;
        RECT 3539.350 2217.760 3539.630 2218.040 ;
        RECT 3539.350 2217.140 3539.630 2217.420 ;
        RECT 3539.350 2216.520 3539.630 2216.800 ;
        RECT 3539.350 2215.900 3539.630 2216.180 ;
        RECT 3539.350 2215.280 3539.630 2215.560 ;
        RECT 3539.350 2214.660 3539.630 2214.940 ;
        RECT 3539.350 2214.040 3539.630 2214.320 ;
        RECT 3539.350 2213.420 3539.630 2213.700 ;
        RECT 3539.350 2212.800 3539.630 2213.080 ;
        RECT 3539.350 2212.180 3539.630 2212.460 ;
        RECT 3539.350 2211.560 3539.630 2211.840 ;
        RECT 3539.350 2210.940 3539.630 2211.220 ;
        RECT 3539.350 2210.320 3539.630 2210.600 ;
        RECT 3539.350 2209.700 3539.630 2209.980 ;
        RECT 3539.350 2209.080 3539.630 2209.360 ;
        RECT 3539.350 2205.390 3539.630 2205.670 ;
        RECT 3539.350 2204.770 3539.630 2205.050 ;
        RECT 3539.350 2204.150 3539.630 2204.430 ;
        RECT 3539.350 2203.530 3539.630 2203.810 ;
        RECT 3539.350 2202.910 3539.630 2203.190 ;
        RECT 3539.350 2202.290 3539.630 2202.570 ;
        RECT 3539.350 2201.670 3539.630 2201.950 ;
        RECT 3539.350 2201.050 3539.630 2201.330 ;
        RECT 3539.350 2200.430 3539.630 2200.710 ;
        RECT 3539.350 2199.810 3539.630 2200.090 ;
        RECT 3539.350 2199.190 3539.630 2199.470 ;
        RECT 3539.350 2198.570 3539.630 2198.850 ;
        RECT 3539.350 2197.950 3539.630 2198.230 ;
        RECT 3539.350 2197.330 3539.630 2197.610 ;
        RECT 3539.350 2196.710 3539.630 2196.990 ;
        RECT 350.370 2168.010 350.650 2168.290 ;
        RECT 350.370 2167.390 350.650 2167.670 ;
        RECT 350.370 2166.770 350.650 2167.050 ;
        RECT 350.370 2166.150 350.650 2166.430 ;
        RECT 350.370 2165.530 350.650 2165.810 ;
        RECT 350.370 2164.910 350.650 2165.190 ;
        RECT 350.370 2164.290 350.650 2164.570 ;
        RECT 350.370 2163.670 350.650 2163.950 ;
        RECT 350.370 2163.050 350.650 2163.330 ;
        RECT 350.370 2162.430 350.650 2162.710 ;
        RECT 350.370 2161.810 350.650 2162.090 ;
        RECT 350.370 2161.190 350.650 2161.470 ;
        RECT 350.370 2160.570 350.650 2160.850 ;
        RECT 350.370 2159.950 350.650 2160.230 ;
        RECT 350.370 2159.330 350.650 2159.610 ;
        RECT 350.370 2155.640 350.650 2155.920 ;
        RECT 350.370 2155.020 350.650 2155.300 ;
        RECT 350.370 2154.400 350.650 2154.680 ;
        RECT 350.370 2153.780 350.650 2154.060 ;
        RECT 350.370 2153.160 350.650 2153.440 ;
        RECT 350.370 2152.540 350.650 2152.820 ;
        RECT 350.370 2151.920 350.650 2152.200 ;
        RECT 350.370 2151.300 350.650 2151.580 ;
        RECT 350.370 2150.680 350.650 2150.960 ;
        RECT 350.370 2150.060 350.650 2150.340 ;
        RECT 350.370 2149.440 350.650 2149.720 ;
        RECT 350.370 2148.820 350.650 2149.100 ;
        RECT 350.370 2148.200 350.650 2148.480 ;
        RECT 350.370 2147.580 350.650 2147.860 ;
        RECT 350.370 2146.960 350.650 2147.240 ;
        RECT 350.370 2146.340 350.650 2146.620 ;
        RECT 350.370 2143.790 350.650 2144.070 ;
        RECT 350.370 2143.170 350.650 2143.450 ;
        RECT 350.370 2142.550 350.650 2142.830 ;
        RECT 350.370 2141.930 350.650 2142.210 ;
        RECT 350.370 2141.310 350.650 2141.590 ;
        RECT 350.370 2140.690 350.650 2140.970 ;
        RECT 350.370 2140.070 350.650 2140.350 ;
        RECT 350.370 2139.450 350.650 2139.730 ;
        RECT 350.370 2138.830 350.650 2139.110 ;
        RECT 350.370 2138.210 350.650 2138.490 ;
        RECT 350.370 2137.590 350.650 2137.870 ;
        RECT 350.370 2136.970 350.650 2137.250 ;
        RECT 350.370 2136.350 350.650 2136.630 ;
        RECT 350.370 2135.730 350.650 2136.010 ;
        RECT 350.370 2135.110 350.650 2135.390 ;
        RECT 350.370 2134.490 350.650 2134.770 ;
        RECT 350.370 2130.260 350.650 2130.540 ;
        RECT 350.370 2129.640 350.650 2129.920 ;
        RECT 350.370 2129.020 350.650 2129.300 ;
        RECT 350.370 2128.400 350.650 2128.680 ;
        RECT 350.370 2127.780 350.650 2128.060 ;
        RECT 350.370 2127.160 350.650 2127.440 ;
        RECT 350.370 2126.540 350.650 2126.820 ;
        RECT 350.370 2125.920 350.650 2126.200 ;
        RECT 350.370 2125.300 350.650 2125.580 ;
        RECT 350.370 2124.680 350.650 2124.960 ;
        RECT 350.370 2124.060 350.650 2124.340 ;
        RECT 350.370 2123.440 350.650 2123.720 ;
        RECT 350.370 2122.820 350.650 2123.100 ;
        RECT 350.370 2122.200 350.650 2122.480 ;
        RECT 350.370 2121.580 350.650 2121.860 ;
        RECT 350.370 2120.960 350.650 2121.240 ;
        RECT 350.370 2118.410 350.650 2118.690 ;
        RECT 350.370 2117.790 350.650 2118.070 ;
        RECT 350.370 2117.170 350.650 2117.450 ;
        RECT 350.370 2116.550 350.650 2116.830 ;
        RECT 350.370 2115.930 350.650 2116.210 ;
        RECT 350.370 2115.310 350.650 2115.590 ;
        RECT 350.370 2114.690 350.650 2114.970 ;
        RECT 350.370 2114.070 350.650 2114.350 ;
        RECT 350.370 2113.450 350.650 2113.730 ;
        RECT 350.370 2112.830 350.650 2113.110 ;
        RECT 350.370 2112.210 350.650 2112.490 ;
        RECT 350.370 2111.590 350.650 2111.870 ;
        RECT 350.370 2110.970 350.650 2111.250 ;
        RECT 350.370 2110.350 350.650 2110.630 ;
        RECT 350.370 2109.730 350.650 2110.010 ;
        RECT 350.370 2109.110 350.650 2109.390 ;
        RECT 350.370 2105.390 350.650 2105.670 ;
        RECT 350.370 2104.770 350.650 2105.050 ;
        RECT 350.370 2104.150 350.650 2104.430 ;
        RECT 350.370 2103.530 350.650 2103.810 ;
        RECT 350.370 2102.910 350.650 2103.190 ;
        RECT 350.370 2102.290 350.650 2102.570 ;
        RECT 350.370 2101.670 350.650 2101.950 ;
        RECT 350.370 2101.050 350.650 2101.330 ;
        RECT 350.370 2100.430 350.650 2100.710 ;
        RECT 350.370 2099.810 350.650 2100.090 ;
        RECT 350.370 2099.190 350.650 2099.470 ;
        RECT 350.370 2098.570 350.650 2098.850 ;
        RECT 350.370 2097.950 350.650 2098.230 ;
        RECT 350.370 2097.330 350.650 2097.610 ;
        RECT 350.370 2096.710 350.650 2096.990 ;
        RECT 3539.350 2053.010 3539.630 2053.290 ;
        RECT 3539.350 2052.390 3539.630 2052.670 ;
        RECT 3539.350 2051.770 3539.630 2052.050 ;
        RECT 3539.350 2051.150 3539.630 2051.430 ;
        RECT 3539.350 2050.530 3539.630 2050.810 ;
        RECT 3539.350 2049.910 3539.630 2050.190 ;
        RECT 3539.350 2049.290 3539.630 2049.570 ;
        RECT 3539.350 2048.670 3539.630 2048.950 ;
        RECT 3539.350 2048.050 3539.630 2048.330 ;
        RECT 3539.350 2047.430 3539.630 2047.710 ;
        RECT 3539.350 2046.810 3539.630 2047.090 ;
        RECT 3539.350 2046.190 3539.630 2046.470 ;
        RECT 3539.350 2045.570 3539.630 2045.850 ;
        RECT 3539.350 2044.950 3539.630 2045.230 ;
        RECT 3539.350 2044.330 3539.630 2044.610 ;
        RECT 3539.350 2040.610 3539.630 2040.890 ;
        RECT 3539.350 2039.990 3539.630 2040.270 ;
        RECT 3539.350 2039.370 3539.630 2039.650 ;
        RECT 3539.350 2038.750 3539.630 2039.030 ;
        RECT 3539.350 2038.130 3539.630 2038.410 ;
        RECT 3539.350 2037.510 3539.630 2037.790 ;
        RECT 3539.350 2036.890 3539.630 2037.170 ;
        RECT 3539.350 2036.270 3539.630 2036.550 ;
        RECT 3539.350 2035.650 3539.630 2035.930 ;
        RECT 3539.350 2035.030 3539.630 2035.310 ;
        RECT 3539.350 2034.410 3539.630 2034.690 ;
        RECT 3539.350 2033.790 3539.630 2034.070 ;
        RECT 3539.350 2033.170 3539.630 2033.450 ;
        RECT 3539.350 2032.550 3539.630 2032.830 ;
        RECT 3539.350 2031.930 3539.630 2032.210 ;
        RECT 3539.350 2031.310 3539.630 2031.590 ;
        RECT 3539.350 2028.760 3539.630 2029.040 ;
        RECT 3539.350 2028.140 3539.630 2028.420 ;
        RECT 3539.350 2027.520 3539.630 2027.800 ;
        RECT 3539.350 2026.900 3539.630 2027.180 ;
        RECT 3539.350 2026.280 3539.630 2026.560 ;
        RECT 3539.350 2025.660 3539.630 2025.940 ;
        RECT 3539.350 2025.040 3539.630 2025.320 ;
        RECT 3539.350 2024.420 3539.630 2024.700 ;
        RECT 3539.350 2023.800 3539.630 2024.080 ;
        RECT 3539.350 2023.180 3539.630 2023.460 ;
        RECT 3539.350 2022.560 3539.630 2022.840 ;
        RECT 3539.350 2021.940 3539.630 2022.220 ;
        RECT 3539.350 2021.320 3539.630 2021.600 ;
        RECT 3539.350 2020.700 3539.630 2020.980 ;
        RECT 3539.350 2020.080 3539.630 2020.360 ;
        RECT 3539.350 2019.460 3539.630 2019.740 ;
        RECT 3539.350 2015.230 3539.630 2015.510 ;
        RECT 3539.350 2014.610 3539.630 2014.890 ;
        RECT 3539.350 2013.990 3539.630 2014.270 ;
        RECT 3539.350 2013.370 3539.630 2013.650 ;
        RECT 3539.350 2012.750 3539.630 2013.030 ;
        RECT 3539.350 2012.130 3539.630 2012.410 ;
        RECT 3539.350 2011.510 3539.630 2011.790 ;
        RECT 3539.350 2010.890 3539.630 2011.170 ;
        RECT 3539.350 2010.270 3539.630 2010.550 ;
        RECT 3539.350 2009.650 3539.630 2009.930 ;
        RECT 3539.350 2009.030 3539.630 2009.310 ;
        RECT 3539.350 2008.410 3539.630 2008.690 ;
        RECT 3539.350 2007.790 3539.630 2008.070 ;
        RECT 3539.350 2007.170 3539.630 2007.450 ;
        RECT 3539.350 2006.550 3539.630 2006.830 ;
        RECT 3539.350 2005.930 3539.630 2006.210 ;
        RECT 3539.350 2003.380 3539.630 2003.660 ;
        RECT 3539.350 2002.760 3539.630 2003.040 ;
        RECT 3539.350 2002.140 3539.630 2002.420 ;
        RECT 3539.350 2001.520 3539.630 2001.800 ;
        RECT 3539.350 2000.900 3539.630 2001.180 ;
        RECT 3539.350 2000.280 3539.630 2000.560 ;
        RECT 3539.350 1999.660 3539.630 1999.940 ;
        RECT 3539.350 1999.040 3539.630 1999.320 ;
        RECT 3539.350 1998.420 3539.630 1998.700 ;
        RECT 3539.350 1997.800 3539.630 1998.080 ;
        RECT 3539.350 1997.180 3539.630 1997.460 ;
        RECT 3539.350 1996.560 3539.630 1996.840 ;
        RECT 3539.350 1995.940 3539.630 1996.220 ;
        RECT 3539.350 1995.320 3539.630 1995.600 ;
        RECT 3539.350 1994.700 3539.630 1994.980 ;
        RECT 3539.350 1994.080 3539.630 1994.360 ;
        RECT 3539.350 1990.390 3539.630 1990.670 ;
        RECT 3539.350 1989.770 3539.630 1990.050 ;
        RECT 3539.350 1989.150 3539.630 1989.430 ;
        RECT 3539.350 1988.530 3539.630 1988.810 ;
        RECT 3539.350 1987.910 3539.630 1988.190 ;
        RECT 3539.350 1987.290 3539.630 1987.570 ;
        RECT 3539.350 1986.670 3539.630 1986.950 ;
        RECT 3539.350 1986.050 3539.630 1986.330 ;
        RECT 3539.350 1985.430 3539.630 1985.710 ;
        RECT 3539.350 1984.810 3539.630 1985.090 ;
        RECT 3539.350 1984.190 3539.630 1984.470 ;
        RECT 3539.350 1983.570 3539.630 1983.850 ;
        RECT 3539.350 1982.950 3539.630 1983.230 ;
        RECT 3539.350 1982.330 3539.630 1982.610 ;
        RECT 3539.350 1981.710 3539.630 1981.990 ;
        RECT 350.370 733.010 350.650 733.290 ;
        RECT 350.370 732.390 350.650 732.670 ;
        RECT 350.370 731.770 350.650 732.050 ;
        RECT 350.370 731.150 350.650 731.430 ;
        RECT 350.370 730.530 350.650 730.810 ;
        RECT 350.370 729.910 350.650 730.190 ;
        RECT 350.370 729.290 350.650 729.570 ;
        RECT 350.370 728.670 350.650 728.950 ;
        RECT 350.370 728.050 350.650 728.330 ;
        RECT 350.370 727.430 350.650 727.710 ;
        RECT 350.370 726.810 350.650 727.090 ;
        RECT 350.370 726.190 350.650 726.470 ;
        RECT 350.370 725.570 350.650 725.850 ;
        RECT 350.370 724.950 350.650 725.230 ;
        RECT 350.370 724.330 350.650 724.610 ;
        RECT 350.370 720.640 350.650 720.920 ;
        RECT 350.370 720.020 350.650 720.300 ;
        RECT 350.370 719.400 350.650 719.680 ;
        RECT 350.370 718.780 350.650 719.060 ;
        RECT 350.370 718.160 350.650 718.440 ;
        RECT 350.370 717.540 350.650 717.820 ;
        RECT 350.370 716.920 350.650 717.200 ;
        RECT 350.370 716.300 350.650 716.580 ;
        RECT 350.370 715.680 350.650 715.960 ;
        RECT 350.370 715.060 350.650 715.340 ;
        RECT 350.370 714.440 350.650 714.720 ;
        RECT 350.370 713.820 350.650 714.100 ;
        RECT 350.370 713.200 350.650 713.480 ;
        RECT 350.370 712.580 350.650 712.860 ;
        RECT 350.370 711.960 350.650 712.240 ;
        RECT 350.370 711.340 350.650 711.620 ;
        RECT 350.370 708.790 350.650 709.070 ;
        RECT 350.370 708.170 350.650 708.450 ;
        RECT 350.370 707.550 350.650 707.830 ;
        RECT 350.370 706.930 350.650 707.210 ;
        RECT 350.370 706.310 350.650 706.590 ;
        RECT 350.370 705.690 350.650 705.970 ;
        RECT 350.370 705.070 350.650 705.350 ;
        RECT 350.370 704.450 350.650 704.730 ;
        RECT 350.370 703.830 350.650 704.110 ;
        RECT 350.370 703.210 350.650 703.490 ;
        RECT 350.370 702.590 350.650 702.870 ;
        RECT 350.370 701.970 350.650 702.250 ;
        RECT 350.370 701.350 350.650 701.630 ;
        RECT 350.370 700.730 350.650 701.010 ;
        RECT 350.370 700.110 350.650 700.390 ;
        RECT 350.370 699.490 350.650 699.770 ;
        RECT 350.370 695.260 350.650 695.540 ;
        RECT 350.370 694.640 350.650 694.920 ;
        RECT 350.370 694.020 350.650 694.300 ;
        RECT 350.370 693.400 350.650 693.680 ;
        RECT 350.370 692.780 350.650 693.060 ;
        RECT 350.370 692.160 350.650 692.440 ;
        RECT 350.370 691.540 350.650 691.820 ;
        RECT 350.370 690.920 350.650 691.200 ;
        RECT 350.370 690.300 350.650 690.580 ;
        RECT 350.370 689.680 350.650 689.960 ;
        RECT 350.370 689.060 350.650 689.340 ;
        RECT 350.370 688.440 350.650 688.720 ;
        RECT 350.370 687.820 350.650 688.100 ;
        RECT 350.370 687.200 350.650 687.480 ;
        RECT 350.370 686.580 350.650 686.860 ;
        RECT 350.370 685.960 350.650 686.240 ;
        RECT 350.370 683.410 350.650 683.690 ;
        RECT 350.370 682.790 350.650 683.070 ;
        RECT 350.370 682.170 350.650 682.450 ;
        RECT 350.370 681.550 350.650 681.830 ;
        RECT 350.370 680.930 350.650 681.210 ;
        RECT 350.370 680.310 350.650 680.590 ;
        RECT 350.370 679.690 350.650 679.970 ;
        RECT 350.370 679.070 350.650 679.350 ;
        RECT 350.370 678.450 350.650 678.730 ;
        RECT 350.370 677.830 350.650 678.110 ;
        RECT 350.370 677.210 350.650 677.490 ;
        RECT 350.370 676.590 350.650 676.870 ;
        RECT 350.370 675.970 350.650 676.250 ;
        RECT 350.370 675.350 350.650 675.630 ;
        RECT 350.370 674.730 350.650 675.010 ;
        RECT 350.370 674.110 350.650 674.390 ;
        RECT 350.370 670.390 350.650 670.670 ;
        RECT 350.370 669.770 350.650 670.050 ;
        RECT 350.370 669.150 350.650 669.430 ;
        RECT 350.370 668.530 350.650 668.810 ;
        RECT 350.370 667.910 350.650 668.190 ;
        RECT 350.370 667.290 350.650 667.570 ;
        RECT 350.370 666.670 350.650 666.950 ;
        RECT 350.370 666.050 350.650 666.330 ;
        RECT 350.370 665.430 350.650 665.710 ;
        RECT 350.370 664.810 350.650 665.090 ;
        RECT 350.370 664.190 350.650 664.470 ;
        RECT 350.370 663.570 350.650 663.850 ;
        RECT 350.370 662.950 350.650 663.230 ;
        RECT 350.370 662.330 350.650 662.610 ;
        RECT 350.370 661.710 350.650 661.990 ;
        RECT 350.370 528.010 350.650 528.290 ;
        RECT 350.370 527.390 350.650 527.670 ;
        RECT 350.370 526.770 350.650 527.050 ;
        RECT 350.370 526.150 350.650 526.430 ;
        RECT 350.370 525.530 350.650 525.810 ;
        RECT 350.370 524.910 350.650 525.190 ;
        RECT 350.370 524.290 350.650 524.570 ;
        RECT 350.370 523.670 350.650 523.950 ;
        RECT 350.370 523.050 350.650 523.330 ;
        RECT 350.370 522.430 350.650 522.710 ;
        RECT 350.370 521.810 350.650 522.090 ;
        RECT 350.370 521.190 350.650 521.470 ;
        RECT 350.370 520.570 350.650 520.850 ;
        RECT 350.370 519.950 350.650 520.230 ;
        RECT 350.370 519.330 350.650 519.610 ;
        RECT 350.370 515.640 350.650 515.920 ;
        RECT 350.370 515.020 350.650 515.300 ;
        RECT 350.370 514.400 350.650 514.680 ;
        RECT 350.370 513.780 350.650 514.060 ;
        RECT 350.370 513.160 350.650 513.440 ;
        RECT 350.370 512.540 350.650 512.820 ;
        RECT 350.370 511.920 350.650 512.200 ;
        RECT 350.370 511.300 350.650 511.580 ;
        RECT 350.370 510.680 350.650 510.960 ;
        RECT 350.370 510.060 350.650 510.340 ;
        RECT 350.370 509.440 350.650 509.720 ;
        RECT 350.370 508.820 350.650 509.100 ;
        RECT 350.370 508.200 350.650 508.480 ;
        RECT 350.370 507.580 350.650 507.860 ;
        RECT 350.370 506.960 350.650 507.240 ;
        RECT 350.370 506.340 350.650 506.620 ;
        RECT 350.370 503.790 350.650 504.070 ;
        RECT 350.370 503.170 350.650 503.450 ;
        RECT 350.370 502.550 350.650 502.830 ;
        RECT 350.370 501.930 350.650 502.210 ;
        RECT 350.370 501.310 350.650 501.590 ;
        RECT 350.370 500.690 350.650 500.970 ;
        RECT 350.370 500.070 350.650 500.350 ;
        RECT 350.370 499.450 350.650 499.730 ;
        RECT 350.370 498.830 350.650 499.110 ;
        RECT 350.370 498.210 350.650 498.490 ;
        RECT 350.370 497.590 350.650 497.870 ;
        RECT 350.370 496.970 350.650 497.250 ;
        RECT 350.370 496.350 350.650 496.630 ;
        RECT 350.370 495.730 350.650 496.010 ;
        RECT 350.370 495.110 350.650 495.390 ;
        RECT 350.370 494.490 350.650 494.770 ;
        RECT 350.370 490.260 350.650 490.540 ;
        RECT 350.370 489.640 350.650 489.920 ;
        RECT 350.370 489.020 350.650 489.300 ;
        RECT 350.370 488.400 350.650 488.680 ;
        RECT 350.370 487.780 350.650 488.060 ;
        RECT 350.370 487.160 350.650 487.440 ;
        RECT 350.370 486.540 350.650 486.820 ;
        RECT 350.370 485.920 350.650 486.200 ;
        RECT 350.370 485.300 350.650 485.580 ;
        RECT 350.370 484.680 350.650 484.960 ;
        RECT 350.370 484.060 350.650 484.340 ;
        RECT 350.370 483.440 350.650 483.720 ;
        RECT 350.370 482.820 350.650 483.100 ;
        RECT 350.370 482.200 350.650 482.480 ;
        RECT 350.370 481.580 350.650 481.860 ;
        RECT 350.370 480.960 350.650 481.240 ;
        RECT 350.370 478.410 350.650 478.690 ;
        RECT 350.370 477.790 350.650 478.070 ;
        RECT 350.370 477.170 350.650 477.450 ;
        RECT 350.370 476.550 350.650 476.830 ;
        RECT 350.370 475.930 350.650 476.210 ;
        RECT 350.370 475.310 350.650 475.590 ;
        RECT 350.370 474.690 350.650 474.970 ;
        RECT 350.370 474.070 350.650 474.350 ;
        RECT 350.370 473.450 350.650 473.730 ;
        RECT 350.370 472.830 350.650 473.110 ;
        RECT 350.370 472.210 350.650 472.490 ;
        RECT 350.370 471.590 350.650 471.870 ;
        RECT 350.370 470.970 350.650 471.250 ;
        RECT 350.370 470.350 350.650 470.630 ;
        RECT 350.370 469.730 350.650 470.010 ;
        RECT 350.370 469.110 350.650 469.390 ;
        RECT 350.370 465.390 350.650 465.670 ;
        RECT 350.370 464.770 350.650 465.050 ;
        RECT 350.370 464.150 350.650 464.430 ;
        RECT 350.370 463.530 350.650 463.810 ;
        RECT 350.370 462.910 350.650 463.190 ;
        RECT 350.370 462.290 350.650 462.570 ;
        RECT 350.370 461.670 350.650 461.950 ;
        RECT 350.370 461.050 350.650 461.330 ;
        RECT 350.370 460.430 350.650 460.710 ;
        RECT 350.370 459.810 350.650 460.090 ;
        RECT 350.370 459.190 350.650 459.470 ;
        RECT 350.370 458.570 350.650 458.850 ;
        RECT 350.370 457.950 350.650 458.230 ;
        RECT 350.370 457.330 350.650 457.610 ;
        RECT 350.370 456.710 350.650 456.990 ;
        RECT 536.710 350.370 536.990 350.650 ;
        RECT 537.330 350.370 537.610 350.650 ;
        RECT 537.950 350.370 538.230 350.650 ;
        RECT 538.570 350.370 538.850 350.650 ;
        RECT 539.190 350.370 539.470 350.650 ;
        RECT 539.810 350.370 540.090 350.650 ;
        RECT 540.430 350.370 540.710 350.650 ;
        RECT 541.050 350.370 541.330 350.650 ;
        RECT 541.670 350.370 541.950 350.650 ;
        RECT 542.290 350.370 542.570 350.650 ;
        RECT 542.910 350.370 543.190 350.650 ;
        RECT 543.530 350.370 543.810 350.650 ;
        RECT 544.150 350.370 544.430 350.650 ;
        RECT 544.770 350.370 545.050 350.650 ;
        RECT 545.390 350.370 545.670 350.650 ;
        RECT 549.110 350.370 549.390 350.650 ;
        RECT 549.730 350.370 550.010 350.650 ;
        RECT 550.350 350.370 550.630 350.650 ;
        RECT 550.970 350.370 551.250 350.650 ;
        RECT 551.590 350.370 551.870 350.650 ;
        RECT 552.210 350.370 552.490 350.650 ;
        RECT 552.830 350.370 553.110 350.650 ;
        RECT 553.450 350.370 553.730 350.650 ;
        RECT 554.070 350.370 554.350 350.650 ;
        RECT 554.690 350.370 554.970 350.650 ;
        RECT 555.310 350.370 555.590 350.650 ;
        RECT 555.930 350.370 556.210 350.650 ;
        RECT 556.550 350.370 556.830 350.650 ;
        RECT 557.170 350.370 557.450 350.650 ;
        RECT 557.790 350.370 558.070 350.650 ;
        RECT 558.410 350.370 558.690 350.650 ;
        RECT 560.960 350.370 561.240 350.650 ;
        RECT 561.580 350.370 561.860 350.650 ;
        RECT 562.200 350.370 562.480 350.650 ;
        RECT 562.820 350.370 563.100 350.650 ;
        RECT 563.440 350.370 563.720 350.650 ;
        RECT 564.060 350.370 564.340 350.650 ;
        RECT 564.680 350.370 564.960 350.650 ;
        RECT 565.300 350.370 565.580 350.650 ;
        RECT 565.920 350.370 566.200 350.650 ;
        RECT 566.540 350.370 566.820 350.650 ;
        RECT 567.160 350.370 567.440 350.650 ;
        RECT 567.780 350.370 568.060 350.650 ;
        RECT 568.400 350.370 568.680 350.650 ;
        RECT 569.020 350.370 569.300 350.650 ;
        RECT 569.640 350.370 569.920 350.650 ;
        RECT 570.260 350.370 570.540 350.650 ;
        RECT 574.460 350.370 574.740 350.650 ;
        RECT 575.080 350.370 575.360 350.650 ;
        RECT 575.700 350.370 575.980 350.650 ;
        RECT 576.320 350.370 576.600 350.650 ;
        RECT 576.940 350.370 577.220 350.650 ;
        RECT 577.560 350.370 577.840 350.650 ;
        RECT 578.180 350.370 578.460 350.650 ;
        RECT 578.800 350.370 579.080 350.650 ;
        RECT 579.420 350.370 579.700 350.650 ;
        RECT 580.040 350.370 580.320 350.650 ;
        RECT 580.660 350.370 580.940 350.650 ;
        RECT 581.280 350.370 581.560 350.650 ;
        RECT 581.900 350.370 582.180 350.650 ;
        RECT 582.520 350.370 582.800 350.650 ;
        RECT 583.140 350.370 583.420 350.650 ;
        RECT 583.760 350.370 584.040 350.650 ;
        RECT 586.310 350.370 586.590 350.650 ;
        RECT 586.930 350.370 587.210 350.650 ;
        RECT 587.550 350.370 587.830 350.650 ;
        RECT 588.170 350.370 588.450 350.650 ;
        RECT 588.790 350.370 589.070 350.650 ;
        RECT 589.410 350.370 589.690 350.650 ;
        RECT 590.030 350.370 590.310 350.650 ;
        RECT 590.650 350.370 590.930 350.650 ;
        RECT 591.270 350.370 591.550 350.650 ;
        RECT 591.890 350.370 592.170 350.650 ;
        RECT 592.510 350.370 592.790 350.650 ;
        RECT 593.130 350.370 593.410 350.650 ;
        RECT 593.750 350.370 594.030 350.650 ;
        RECT 594.370 350.370 594.650 350.650 ;
        RECT 594.990 350.370 595.270 350.650 ;
        RECT 595.610 350.370 595.890 350.650 ;
        RECT 599.330 350.370 599.610 350.650 ;
        RECT 599.950 350.370 600.230 350.650 ;
        RECT 600.570 350.370 600.850 350.650 ;
        RECT 601.190 350.370 601.470 350.650 ;
        RECT 601.810 350.370 602.090 350.650 ;
        RECT 602.430 350.370 602.710 350.650 ;
        RECT 603.050 350.370 603.330 350.650 ;
        RECT 603.670 350.370 603.950 350.650 ;
        RECT 604.290 350.370 604.570 350.650 ;
        RECT 604.910 350.370 605.190 350.650 ;
        RECT 605.530 350.370 605.810 350.650 ;
        RECT 606.150 350.370 606.430 350.650 ;
        RECT 606.770 350.370 607.050 350.650 ;
        RECT 607.390 350.370 607.670 350.650 ;
        RECT 608.010 350.370 608.290 350.650 ;
        RECT 1361.710 350.370 1361.990 350.650 ;
        RECT 1362.330 350.370 1362.610 350.650 ;
        RECT 1362.950 350.370 1363.230 350.650 ;
        RECT 1363.570 350.370 1363.850 350.650 ;
        RECT 1364.190 350.370 1364.470 350.650 ;
        RECT 1364.810 350.370 1365.090 350.650 ;
        RECT 1365.430 350.370 1365.710 350.650 ;
        RECT 1366.050 350.370 1366.330 350.650 ;
        RECT 1366.670 350.370 1366.950 350.650 ;
        RECT 1367.290 350.370 1367.570 350.650 ;
        RECT 1367.910 350.370 1368.190 350.650 ;
        RECT 1368.530 350.370 1368.810 350.650 ;
        RECT 1369.150 350.370 1369.430 350.650 ;
        RECT 1369.770 350.370 1370.050 350.650 ;
        RECT 1370.390 350.370 1370.670 350.650 ;
        RECT 1374.110 350.370 1374.390 350.650 ;
        RECT 1374.730 350.370 1375.010 350.650 ;
        RECT 1375.350 350.370 1375.630 350.650 ;
        RECT 1375.970 350.370 1376.250 350.650 ;
        RECT 1376.590 350.370 1376.870 350.650 ;
        RECT 1377.210 350.370 1377.490 350.650 ;
        RECT 1377.830 350.370 1378.110 350.650 ;
        RECT 1378.450 350.370 1378.730 350.650 ;
        RECT 1379.070 350.370 1379.350 350.650 ;
        RECT 1379.690 350.370 1379.970 350.650 ;
        RECT 1380.310 350.370 1380.590 350.650 ;
        RECT 1380.930 350.370 1381.210 350.650 ;
        RECT 1381.550 350.370 1381.830 350.650 ;
        RECT 1382.170 350.370 1382.450 350.650 ;
        RECT 1382.790 350.370 1383.070 350.650 ;
        RECT 1383.410 350.370 1383.690 350.650 ;
        RECT 1385.960 350.370 1386.240 350.650 ;
        RECT 1386.580 350.370 1386.860 350.650 ;
        RECT 1387.200 350.370 1387.480 350.650 ;
        RECT 1387.820 350.370 1388.100 350.650 ;
        RECT 1388.440 350.370 1388.720 350.650 ;
        RECT 1389.060 350.370 1389.340 350.650 ;
        RECT 1389.680 350.370 1389.960 350.650 ;
        RECT 1390.300 350.370 1390.580 350.650 ;
        RECT 1390.920 350.370 1391.200 350.650 ;
        RECT 1391.540 350.370 1391.820 350.650 ;
        RECT 1392.160 350.370 1392.440 350.650 ;
        RECT 1392.780 350.370 1393.060 350.650 ;
        RECT 1393.400 350.370 1393.680 350.650 ;
        RECT 1394.020 350.370 1394.300 350.650 ;
        RECT 1394.640 350.370 1394.920 350.650 ;
        RECT 1395.260 350.370 1395.540 350.650 ;
        RECT 1399.460 350.370 1399.740 350.650 ;
        RECT 1400.080 350.370 1400.360 350.650 ;
        RECT 1400.700 350.370 1400.980 350.650 ;
        RECT 1401.320 350.370 1401.600 350.650 ;
        RECT 1401.940 350.370 1402.220 350.650 ;
        RECT 1402.560 350.370 1402.840 350.650 ;
        RECT 1403.180 350.370 1403.460 350.650 ;
        RECT 1403.800 350.370 1404.080 350.650 ;
        RECT 1404.420 350.370 1404.700 350.650 ;
        RECT 1405.040 350.370 1405.320 350.650 ;
        RECT 1405.660 350.370 1405.940 350.650 ;
        RECT 1406.280 350.370 1406.560 350.650 ;
        RECT 1406.900 350.370 1407.180 350.650 ;
        RECT 1407.520 350.370 1407.800 350.650 ;
        RECT 1408.140 350.370 1408.420 350.650 ;
        RECT 1408.760 350.370 1409.040 350.650 ;
        RECT 1411.310 350.370 1411.590 350.650 ;
        RECT 1411.930 350.370 1412.210 350.650 ;
        RECT 1412.550 350.370 1412.830 350.650 ;
        RECT 1413.170 350.370 1413.450 350.650 ;
        RECT 1413.790 350.370 1414.070 350.650 ;
        RECT 1414.410 350.370 1414.690 350.650 ;
        RECT 1415.030 350.370 1415.310 350.650 ;
        RECT 1415.650 350.370 1415.930 350.650 ;
        RECT 1416.270 350.370 1416.550 350.650 ;
        RECT 1416.890 350.370 1417.170 350.650 ;
        RECT 1417.510 350.370 1417.790 350.650 ;
        RECT 1418.130 350.370 1418.410 350.650 ;
        RECT 1418.750 350.370 1419.030 350.650 ;
        RECT 1419.370 350.370 1419.650 350.650 ;
        RECT 1419.990 350.370 1420.270 350.650 ;
        RECT 1420.610 350.370 1420.890 350.650 ;
        RECT 1424.330 350.370 1424.610 350.650 ;
        RECT 1424.950 350.370 1425.230 350.650 ;
        RECT 1425.570 350.370 1425.850 350.650 ;
        RECT 1426.190 350.370 1426.470 350.650 ;
        RECT 1426.810 350.370 1427.090 350.650 ;
        RECT 1427.430 350.370 1427.710 350.650 ;
        RECT 1428.050 350.370 1428.330 350.650 ;
        RECT 1428.670 350.370 1428.950 350.650 ;
        RECT 1429.290 350.370 1429.570 350.650 ;
        RECT 1429.910 350.370 1430.190 350.650 ;
        RECT 1430.530 350.370 1430.810 350.650 ;
        RECT 1431.150 350.370 1431.430 350.650 ;
        RECT 1431.770 350.370 1432.050 350.650 ;
        RECT 1432.390 350.370 1432.670 350.650 ;
        RECT 1433.010 350.370 1433.290 350.650 ;
        RECT 3011.710 350.370 3011.990 350.650 ;
        RECT 3012.330 350.370 3012.610 350.650 ;
        RECT 3012.950 350.370 3013.230 350.650 ;
        RECT 3013.570 350.370 3013.850 350.650 ;
        RECT 3014.190 350.370 3014.470 350.650 ;
        RECT 3014.810 350.370 3015.090 350.650 ;
        RECT 3015.430 350.370 3015.710 350.650 ;
        RECT 3016.050 350.370 3016.330 350.650 ;
        RECT 3016.670 350.370 3016.950 350.650 ;
        RECT 3017.290 350.370 3017.570 350.650 ;
        RECT 3017.910 350.370 3018.190 350.650 ;
        RECT 3018.530 350.370 3018.810 350.650 ;
        RECT 3019.150 350.370 3019.430 350.650 ;
        RECT 3019.770 350.370 3020.050 350.650 ;
        RECT 3020.390 350.370 3020.670 350.650 ;
        RECT 3024.110 350.370 3024.390 350.650 ;
        RECT 3024.730 350.370 3025.010 350.650 ;
        RECT 3025.350 350.370 3025.630 350.650 ;
        RECT 3025.970 350.370 3026.250 350.650 ;
        RECT 3026.590 350.370 3026.870 350.650 ;
        RECT 3027.210 350.370 3027.490 350.650 ;
        RECT 3027.830 350.370 3028.110 350.650 ;
        RECT 3028.450 350.370 3028.730 350.650 ;
        RECT 3029.070 350.370 3029.350 350.650 ;
        RECT 3029.690 350.370 3029.970 350.650 ;
        RECT 3030.310 350.370 3030.590 350.650 ;
        RECT 3030.930 350.370 3031.210 350.650 ;
        RECT 3031.550 350.370 3031.830 350.650 ;
        RECT 3032.170 350.370 3032.450 350.650 ;
        RECT 3032.790 350.370 3033.070 350.650 ;
        RECT 3033.410 350.370 3033.690 350.650 ;
        RECT 3035.960 350.370 3036.240 350.650 ;
        RECT 3036.580 350.370 3036.860 350.650 ;
        RECT 3037.200 350.370 3037.480 350.650 ;
        RECT 3037.820 350.370 3038.100 350.650 ;
        RECT 3038.440 350.370 3038.720 350.650 ;
        RECT 3039.060 350.370 3039.340 350.650 ;
        RECT 3039.680 350.370 3039.960 350.650 ;
        RECT 3040.300 350.370 3040.580 350.650 ;
        RECT 3040.920 350.370 3041.200 350.650 ;
        RECT 3041.540 350.370 3041.820 350.650 ;
        RECT 3042.160 350.370 3042.440 350.650 ;
        RECT 3042.780 350.370 3043.060 350.650 ;
        RECT 3043.400 350.370 3043.680 350.650 ;
        RECT 3044.020 350.370 3044.300 350.650 ;
        RECT 3044.640 350.370 3044.920 350.650 ;
        RECT 3045.260 350.370 3045.540 350.650 ;
        RECT 3049.460 350.370 3049.740 350.650 ;
        RECT 3050.080 350.370 3050.360 350.650 ;
        RECT 3050.700 350.370 3050.980 350.650 ;
        RECT 3051.320 350.370 3051.600 350.650 ;
        RECT 3051.940 350.370 3052.220 350.650 ;
        RECT 3052.560 350.370 3052.840 350.650 ;
        RECT 3053.180 350.370 3053.460 350.650 ;
        RECT 3053.800 350.370 3054.080 350.650 ;
        RECT 3054.420 350.370 3054.700 350.650 ;
        RECT 3055.040 350.370 3055.320 350.650 ;
        RECT 3055.660 350.370 3055.940 350.650 ;
        RECT 3056.280 350.370 3056.560 350.650 ;
        RECT 3056.900 350.370 3057.180 350.650 ;
        RECT 3057.520 350.370 3057.800 350.650 ;
        RECT 3058.140 350.370 3058.420 350.650 ;
        RECT 3058.760 350.370 3059.040 350.650 ;
        RECT 3061.310 350.370 3061.590 350.650 ;
        RECT 3061.930 350.370 3062.210 350.650 ;
        RECT 3062.550 350.370 3062.830 350.650 ;
        RECT 3063.170 350.370 3063.450 350.650 ;
        RECT 3063.790 350.370 3064.070 350.650 ;
        RECT 3064.410 350.370 3064.690 350.650 ;
        RECT 3065.030 350.370 3065.310 350.650 ;
        RECT 3065.650 350.370 3065.930 350.650 ;
        RECT 3066.270 350.370 3066.550 350.650 ;
        RECT 3066.890 350.370 3067.170 350.650 ;
        RECT 3067.510 350.370 3067.790 350.650 ;
        RECT 3068.130 350.370 3068.410 350.650 ;
        RECT 3068.750 350.370 3069.030 350.650 ;
        RECT 3069.370 350.370 3069.650 350.650 ;
        RECT 3069.990 350.370 3070.270 350.650 ;
        RECT 3070.610 350.370 3070.890 350.650 ;
        RECT 3074.330 350.370 3074.610 350.650 ;
        RECT 3074.950 350.370 3075.230 350.650 ;
        RECT 3075.570 350.370 3075.850 350.650 ;
        RECT 3076.190 350.370 3076.470 350.650 ;
        RECT 3076.810 350.370 3077.090 350.650 ;
        RECT 3077.430 350.370 3077.710 350.650 ;
        RECT 3078.050 350.370 3078.330 350.650 ;
        RECT 3078.670 350.370 3078.950 350.650 ;
        RECT 3079.290 350.370 3079.570 350.650 ;
        RECT 3079.910 350.370 3080.190 350.650 ;
        RECT 3080.530 350.370 3080.810 350.650 ;
        RECT 3081.150 350.370 3081.430 350.650 ;
        RECT 3081.770 350.370 3082.050 350.650 ;
        RECT 3082.390 350.370 3082.670 350.650 ;
        RECT 3083.010 350.370 3083.290 350.650 ;
        RECT 3286.710 350.370 3286.990 350.650 ;
        RECT 3287.330 350.370 3287.610 350.650 ;
        RECT 3287.950 350.370 3288.230 350.650 ;
        RECT 3288.570 350.370 3288.850 350.650 ;
        RECT 3289.190 350.370 3289.470 350.650 ;
        RECT 3289.810 350.370 3290.090 350.650 ;
        RECT 3290.430 350.370 3290.710 350.650 ;
        RECT 3291.050 350.370 3291.330 350.650 ;
        RECT 3291.670 350.370 3291.950 350.650 ;
        RECT 3292.290 350.370 3292.570 350.650 ;
        RECT 3292.910 350.370 3293.190 350.650 ;
        RECT 3293.530 350.370 3293.810 350.650 ;
        RECT 3294.150 350.370 3294.430 350.650 ;
        RECT 3294.770 350.370 3295.050 350.650 ;
        RECT 3295.390 350.370 3295.670 350.650 ;
        RECT 3299.110 350.370 3299.390 350.650 ;
        RECT 3299.730 350.370 3300.010 350.650 ;
        RECT 3300.350 350.370 3300.630 350.650 ;
        RECT 3300.970 350.370 3301.250 350.650 ;
        RECT 3301.590 350.370 3301.870 350.650 ;
        RECT 3302.210 350.370 3302.490 350.650 ;
        RECT 3302.830 350.370 3303.110 350.650 ;
        RECT 3303.450 350.370 3303.730 350.650 ;
        RECT 3304.070 350.370 3304.350 350.650 ;
        RECT 3304.690 350.370 3304.970 350.650 ;
        RECT 3305.310 350.370 3305.590 350.650 ;
        RECT 3305.930 350.370 3306.210 350.650 ;
        RECT 3306.550 350.370 3306.830 350.650 ;
        RECT 3307.170 350.370 3307.450 350.650 ;
        RECT 3307.790 350.370 3308.070 350.650 ;
        RECT 3308.410 350.370 3308.690 350.650 ;
        RECT 3310.960 350.370 3311.240 350.650 ;
        RECT 3311.580 350.370 3311.860 350.650 ;
        RECT 3312.200 350.370 3312.480 350.650 ;
        RECT 3312.820 350.370 3313.100 350.650 ;
        RECT 3313.440 350.370 3313.720 350.650 ;
        RECT 3314.060 350.370 3314.340 350.650 ;
        RECT 3314.680 350.370 3314.960 350.650 ;
        RECT 3315.300 350.370 3315.580 350.650 ;
        RECT 3315.920 350.370 3316.200 350.650 ;
        RECT 3316.540 350.370 3316.820 350.650 ;
        RECT 3317.160 350.370 3317.440 350.650 ;
        RECT 3317.780 350.370 3318.060 350.650 ;
        RECT 3318.400 350.370 3318.680 350.650 ;
        RECT 3319.020 350.370 3319.300 350.650 ;
        RECT 3319.640 350.370 3319.920 350.650 ;
        RECT 3320.260 350.370 3320.540 350.650 ;
        RECT 3324.460 350.370 3324.740 350.650 ;
        RECT 3325.080 350.370 3325.360 350.650 ;
        RECT 3325.700 350.370 3325.980 350.650 ;
        RECT 3326.320 350.370 3326.600 350.650 ;
        RECT 3326.940 350.370 3327.220 350.650 ;
        RECT 3327.560 350.370 3327.840 350.650 ;
        RECT 3328.180 350.370 3328.460 350.650 ;
        RECT 3328.800 350.370 3329.080 350.650 ;
        RECT 3329.420 350.370 3329.700 350.650 ;
        RECT 3330.040 350.370 3330.320 350.650 ;
        RECT 3330.660 350.370 3330.940 350.650 ;
        RECT 3331.280 350.370 3331.560 350.650 ;
        RECT 3331.900 350.370 3332.180 350.650 ;
        RECT 3332.520 350.370 3332.800 350.650 ;
        RECT 3333.140 350.370 3333.420 350.650 ;
        RECT 3333.760 350.370 3334.040 350.650 ;
        RECT 3336.310 350.370 3336.590 350.650 ;
        RECT 3336.930 350.370 3337.210 350.650 ;
        RECT 3337.550 350.370 3337.830 350.650 ;
        RECT 3338.170 350.370 3338.450 350.650 ;
        RECT 3338.790 350.370 3339.070 350.650 ;
        RECT 3339.410 350.370 3339.690 350.650 ;
        RECT 3340.030 350.370 3340.310 350.650 ;
        RECT 3340.650 350.370 3340.930 350.650 ;
        RECT 3341.270 350.370 3341.550 350.650 ;
        RECT 3341.890 350.370 3342.170 350.650 ;
        RECT 3342.510 350.370 3342.790 350.650 ;
        RECT 3343.130 350.370 3343.410 350.650 ;
        RECT 3343.750 350.370 3344.030 350.650 ;
        RECT 3344.370 350.370 3344.650 350.650 ;
        RECT 3344.990 350.370 3345.270 350.650 ;
        RECT 3345.610 350.370 3345.890 350.650 ;
        RECT 3349.330 350.370 3349.610 350.650 ;
        RECT 3349.950 350.370 3350.230 350.650 ;
        RECT 3350.570 350.370 3350.850 350.650 ;
        RECT 3351.190 350.370 3351.470 350.650 ;
        RECT 3351.810 350.370 3352.090 350.650 ;
        RECT 3352.430 350.370 3352.710 350.650 ;
        RECT 3353.050 350.370 3353.330 350.650 ;
        RECT 3353.670 350.370 3353.950 350.650 ;
        RECT 3354.290 350.370 3354.570 350.650 ;
        RECT 3354.910 350.370 3355.190 350.650 ;
        RECT 3355.530 350.370 3355.810 350.650 ;
        RECT 3356.150 350.370 3356.430 350.650 ;
        RECT 3356.770 350.370 3357.050 350.650 ;
        RECT 3357.390 350.370 3357.670 350.650 ;
        RECT 3358.010 350.370 3358.290 350.650 ;
      LAYER Metal4 ;
        RECT 350.000 4414.140 351.000 4423.640 ;
        RECT 350.000 4400.990 351.000 4411.240 ;
        RECT 350.000 4389.140 351.000 4399.390 ;
        RECT 350.000 4375.610 351.000 4385.860 ;
        RECT 350.000 4363.760 351.000 4374.010 ;
        RECT 350.000 4351.360 351.000 4360.860 ;
        RECT 350.000 4209.140 351.000 4218.640 ;
        RECT 350.000 4195.990 351.000 4206.240 ;
        RECT 350.000 4184.140 351.000 4194.390 ;
        RECT 350.000 4170.610 351.000 4180.860 ;
        RECT 350.000 4158.760 351.000 4169.010 ;
        RECT 350.000 4146.360 351.000 4155.860 ;
        RECT 350.000 4004.140 351.000 4013.640 ;
        RECT 350.000 3990.990 351.000 4001.240 ;
        RECT 350.000 3979.140 351.000 3989.390 ;
        RECT 350.000 3965.610 351.000 3975.860 ;
        RECT 350.000 3953.760 351.000 3964.010 ;
        RECT 350.000 3941.360 351.000 3950.860 ;
        RECT 350.000 2364.140 351.000 2373.640 ;
        RECT 350.000 2350.990 351.000 2361.240 ;
        RECT 350.000 2339.140 351.000 2349.390 ;
        RECT 350.000 2325.610 351.000 2335.860 ;
        RECT 350.000 2313.760 351.000 2324.010 ;
        RECT 350.000 2301.360 351.000 2310.860 ;
        RECT 350.000 2159.145 351.000 2168.645 ;
        RECT 350.000 2145.995 351.000 2156.245 ;
        RECT 350.000 2134.145 351.000 2144.395 ;
        RECT 350.000 2120.615 351.000 2130.865 ;
        RECT 350.000 2108.765 351.000 2119.015 ;
        RECT 350.000 2096.365 351.000 2105.865 ;
        RECT 350.000 724.140 351.000 733.640 ;
        RECT 350.000 710.990 351.000 721.240 ;
        RECT 350.000 699.140 351.000 709.390 ;
        RECT 350.000 685.610 351.000 695.860 ;
        RECT 350.000 673.760 351.000 684.010 ;
        RECT 350.000 661.360 351.000 670.860 ;
        RECT 350.000 519.140 351.000 528.640 ;
        RECT 350.000 505.990 351.000 516.240 ;
        RECT 350.000 494.140 351.000 504.390 ;
        RECT 350.000 480.610 351.000 490.860 ;
        RECT 350.000 468.760 351.000 479.010 ;
        RECT 350.000 456.360 351.000 465.860 ;
        RECT 388.390 388.390 393.390 4728.550 ;
        RECT 395.390 395.390 400.390 4730.550 ;
        RECT 701.695 4717.825 704.695 4719.425 ;
        RECT 976.695 4717.825 979.695 4719.425 ;
        RECT 1251.695 4717.825 1254.695 4719.425 ;
        RECT 1526.695 4717.825 1529.695 4719.425 ;
        RECT 1801.695 4717.825 1804.695 4719.425 ;
        RECT 440.030 4668.040 443.130 4711.610 ;
        RECT 530.030 4672.840 533.130 4704.610 ;
        RECT 552.120 4699.610 553.720 4717.520 ;
        RECT 587.120 4699.610 588.720 4717.520 ;
        RECT 622.120 4699.610 623.720 4717.520 ;
        RECT 701.695 4706.610 702.695 4715.425 ;
        RECT 703.695 4699.610 704.695 4717.825 ;
        RECT 710.030 4672.840 713.130 4704.610 ;
        RECT 800.030 4668.040 803.130 4711.610 ;
        RECT 827.120 4699.610 828.720 4717.520 ;
        RECT 862.120 4699.610 863.720 4717.520 ;
        RECT 890.030 4672.840 893.130 4704.610 ;
        RECT 897.120 4699.610 898.720 4717.520 ;
        RECT 976.695 4706.610 977.695 4715.425 ;
        RECT 978.695 4699.610 979.695 4717.825 ;
        RECT 1070.030 4672.840 1073.130 4704.610 ;
        RECT 1102.120 4699.610 1103.720 4717.520 ;
        RECT 1137.120 4699.610 1138.720 4717.520 ;
        RECT 1160.030 4668.040 1163.130 4711.610 ;
        RECT 1172.120 4699.610 1173.720 4717.520 ;
        RECT 1251.695 4706.610 1252.695 4715.425 ;
        RECT 1250.030 4672.840 1253.130 4704.610 ;
        RECT 1253.695 4699.610 1254.695 4717.825 ;
        RECT 1340.030 4668.040 1343.130 4711.610 ;
        RECT 1377.120 4699.610 1378.720 4717.520 ;
        RECT 1412.120 4699.610 1413.720 4717.520 ;
        RECT 1430.030 4672.840 1433.130 4704.610 ;
        RECT 1447.120 4699.610 1448.720 4717.520 ;
        RECT 1520.030 4668.040 1523.130 4711.610 ;
        RECT 1526.695 4706.610 1527.695 4715.425 ;
        RECT 1528.695 4699.610 1529.695 4717.825 ;
        RECT 1610.030 4672.840 1613.130 4704.610 ;
        RECT 1652.120 4699.610 1653.720 4717.520 ;
        RECT 1687.120 4699.610 1688.720 4717.520 ;
        RECT 1700.030 4668.040 1703.130 4711.610 ;
        RECT 1722.120 4699.610 1723.720 4717.520 ;
        RECT 1801.695 4706.610 1802.695 4715.425 ;
        RECT 1790.030 4672.840 1793.130 4704.610 ;
        RECT 1803.695 4699.610 1804.695 4717.825 ;
        RECT 1880.030 4668.040 1883.130 4711.610 ;
        RECT 1906.360 4699.610 1915.860 4750.000 ;
        RECT 1918.760 4699.610 1929.010 4750.000 ;
        RECT 1930.610 4699.610 1940.860 4750.000 ;
        RECT 1944.140 4699.610 1954.390 4750.000 ;
        RECT 1955.990 4699.610 1966.240 4750.000 ;
        RECT 1969.140 4699.610 1978.640 4750.000 ;
        RECT 2351.695 4717.825 2354.695 4719.425 ;
        RECT 2626.695 4717.825 2629.695 4719.425 ;
        RECT 2901.695 4717.825 2904.695 4719.425 ;
        RECT 1970.030 4672.840 1973.130 4699.610 ;
        RECT 2060.030 4668.040 2063.130 4711.610 ;
        RECT 2150.030 4672.840 2153.130 4704.610 ;
        RECT 2202.120 4699.610 2203.720 4717.520 ;
        RECT 2237.120 4699.610 2238.720 4717.520 ;
        RECT 2240.030 4668.040 2243.130 4711.610 ;
        RECT 2272.120 4699.610 2273.720 4717.520 ;
        RECT 2351.695 4706.610 2352.695 4715.425 ;
        RECT 2330.030 4672.840 2333.130 4704.610 ;
        RECT 2353.695 4699.610 2354.695 4717.825 ;
        RECT 2420.030 4668.040 2423.130 4711.610 ;
        RECT 2477.120 4699.610 2478.720 4717.520 ;
        RECT 2512.120 4704.610 2513.720 4717.520 ;
        RECT 2510.030 4699.610 2513.720 4704.610 ;
        RECT 2547.120 4699.610 2548.720 4717.520 ;
        RECT 2510.030 4672.840 2513.130 4699.610 ;
        RECT 2600.030 4668.040 2603.130 4711.610 ;
        RECT 2626.695 4706.610 2627.695 4715.425 ;
        RECT 2628.695 4699.610 2629.695 4717.825 ;
        RECT 2690.030 4672.840 2693.130 4704.610 ;
        RECT 2752.120 4699.610 2753.720 4717.520 ;
        RECT 2780.030 4668.040 2783.130 4711.610 ;
        RECT 2787.120 4699.610 2788.720 4717.520 ;
        RECT 2822.120 4699.610 2823.720 4717.520 ;
        RECT 2901.695 4706.610 2902.695 4715.425 ;
        RECT 2870.030 4672.840 2873.130 4704.610 ;
        RECT 2903.695 4699.610 2904.695 4717.825 ;
        RECT 2960.030 4668.040 2963.130 4711.610 ;
        RECT 3006.360 4699.610 3015.860 4750.000 ;
        RECT 3018.760 4699.610 3029.010 4750.000 ;
        RECT 3030.610 4699.610 3040.860 4750.000 ;
        RECT 3044.140 4699.610 3054.390 4750.000 ;
        RECT 3055.990 4699.610 3066.240 4750.000 ;
        RECT 3069.140 4699.610 3078.640 4750.000 ;
        RECT 3451.695 4717.825 3454.695 4719.425 ;
        RECT 3050.030 4672.840 3053.130 4699.610 ;
        RECT 3140.030 4668.040 3143.130 4711.610 ;
        RECT 3230.030 4672.840 3233.130 4704.610 ;
        RECT 3302.120 4699.610 3303.720 4717.520 ;
        RECT 3320.030 4668.040 3323.130 4711.610 ;
        RECT 3337.120 4699.610 3338.720 4717.520 ;
        RECT 3372.120 4699.610 3373.720 4717.520 ;
        RECT 3451.695 4706.610 3452.695 4715.425 ;
        RECT 3410.030 4672.840 3413.130 4704.610 ;
        RECT 3453.695 4699.610 3454.695 4717.825 ;
        RECT 440.030 1643.550 443.130 1672.600 ;
        RECT 530.030 1650.550 533.130 1667.800 ;
        RECT 620.030 1643.550 623.130 1672.600 ;
        RECT 710.030 1650.550 713.130 1667.800 ;
        RECT 572.775 1524.280 574.375 1571.420 ;
        RECT 580.750 1531.280 582.350 1571.420 ;
        RECT 588.725 1524.280 590.325 1571.420 ;
        RECT 596.700 1531.280 598.300 1571.420 ;
        RECT 604.675 1524.280 606.275 1571.420 ;
        RECT 612.650 1531.280 614.250 1571.420 ;
        RECT 620.625 1524.280 622.225 1571.420 ;
        RECT 785.440 1524.280 788.540 1648.550 ;
        RECT 790.540 1531.280 793.640 1655.550 ;
        RECT 800.030 1643.550 803.130 1672.600 ;
        RECT 890.030 1650.550 893.130 1667.800 ;
        RECT 980.030 1643.550 983.130 1672.600 ;
        RECT 1070.030 1650.550 1073.130 1667.800 ;
        RECT 1160.030 1643.550 1163.130 1672.600 ;
        RECT 1250.030 1650.550 1253.130 1667.800 ;
        RECT 1340.030 1643.550 1343.130 1672.600 ;
        RECT 1430.030 1650.550 1433.130 1667.800 ;
        RECT 1520.030 1643.550 1523.130 1672.600 ;
        RECT 1610.030 1650.550 1613.130 1667.800 ;
        RECT 1700.030 1643.550 1703.130 1672.600 ;
        RECT 1790.030 1650.550 1793.130 1667.800 ;
        RECT 1880.030 1643.550 1883.130 1672.600 ;
        RECT 1906.200 1531.280 1909.300 1655.550 ;
        RECT 1970.030 1650.550 1973.130 1667.800 ;
        RECT 1911.300 1524.280 1914.400 1648.550 ;
        RECT 2060.030 1643.550 2063.130 1672.600 ;
        RECT 2150.030 1650.550 2153.130 1667.800 ;
        RECT 2240.030 1643.550 2243.130 1672.600 ;
        RECT 2330.030 1650.550 2333.130 1667.800 ;
        RECT 2420.030 1643.550 2423.130 1672.600 ;
        RECT 2510.030 1650.550 2513.130 1667.800 ;
        RECT 2600.030 1643.550 2603.130 1672.600 ;
        RECT 2690.030 1650.550 2693.130 1667.800 ;
        RECT 2780.030 1643.550 2783.130 1672.600 ;
        RECT 2870.030 1650.550 2873.130 1667.800 ;
        RECT 2960.030 1643.550 2963.130 1672.600 ;
        RECT 3050.030 1650.550 3053.130 1667.800 ;
        RECT 3140.030 1643.550 3143.130 1672.600 ;
        RECT 3230.030 1650.550 3233.130 1667.800 ;
        RECT 3320.030 1643.550 3323.130 1672.600 ;
        RECT 3410.030 1650.550 3413.130 1667.800 ;
        RECT 1942.775 1524.280 1944.375 1571.420 ;
        RECT 1950.750 1531.280 1952.350 1571.420 ;
        RECT 1958.725 1524.280 1960.325 1571.420 ;
        RECT 1966.700 1531.280 1968.300 1571.420 ;
        RECT 1974.675 1524.280 1976.275 1571.420 ;
        RECT 1982.650 1531.280 1984.250 1571.420 ;
        RECT 1990.625 1524.280 1992.225 1571.420 ;
        RECT 2442.775 1524.280 2444.375 1571.420 ;
        RECT 2450.750 1531.280 2452.350 1571.420 ;
        RECT 2458.725 1524.280 2460.325 1571.420 ;
        RECT 2466.700 1531.280 2468.300 1571.420 ;
        RECT 2474.675 1524.280 2476.275 1571.420 ;
        RECT 2482.650 1531.280 2484.250 1571.420 ;
        RECT 2490.625 1524.280 2492.225 1571.420 ;
        RECT 471.120 1396.840 472.720 1410.210 ;
        RECT 496.120 1396.840 497.720 1417.210 ;
        RECT 521.120 1396.840 522.720 1410.210 ;
        RECT 546.120 1396.840 547.720 1417.210 ;
        RECT 571.120 1396.840 572.720 1410.210 ;
        RECT 596.120 1396.840 597.720 1417.210 ;
        RECT 621.120 1396.840 622.720 1410.210 ;
        RECT 646.120 1396.840 647.720 1417.210 ;
        RECT 671.120 1396.840 672.720 1410.210 ;
        RECT 696.120 1396.840 697.720 1417.210 ;
        RECT 721.120 1396.840 722.720 1410.210 ;
        RECT 746.120 1396.840 747.720 1417.210 ;
        RECT 771.120 1396.840 772.720 1410.210 ;
        RECT 796.120 1396.840 797.720 1417.210 ;
        RECT 821.120 1396.840 822.720 1410.210 ;
        RECT 846.120 1396.840 847.720 1417.210 ;
        RECT 871.120 1396.840 872.720 1410.210 ;
        RECT 896.120 1396.840 897.720 1417.210 ;
        RECT 921.120 1396.840 922.720 1410.210 ;
        RECT 946.120 1396.840 947.720 1417.210 ;
        RECT 971.120 1396.840 972.720 1410.210 ;
        RECT 996.120 1396.840 997.720 1417.210 ;
        RECT 1021.120 1396.840 1022.720 1410.210 ;
        RECT 1046.120 1396.840 1047.720 1417.210 ;
        RECT 1071.120 1396.840 1072.720 1410.210 ;
        RECT 1096.120 1396.840 1097.720 1417.210 ;
        RECT 1121.120 1396.840 1122.720 1410.210 ;
        RECT 1146.120 1396.840 1147.720 1417.210 ;
        RECT 1171.120 1396.840 1172.720 1410.210 ;
        RECT 1196.120 1396.840 1197.720 1417.210 ;
        RECT 1221.120 1396.840 1222.720 1410.210 ;
        RECT 1246.120 1396.840 1247.720 1417.210 ;
        RECT 1271.120 1396.840 1272.720 1410.210 ;
        RECT 1296.120 1396.840 1297.720 1417.210 ;
        RECT 1321.120 1396.840 1322.720 1410.210 ;
        RECT 1346.120 1396.840 1347.720 1417.210 ;
        RECT 1371.120 1396.840 1372.720 1410.210 ;
        RECT 1396.120 1396.840 1397.720 1417.210 ;
        RECT 1421.120 1396.840 1422.720 1410.210 ;
        RECT 1446.120 1396.840 1447.720 1417.210 ;
        RECT 1471.120 1396.840 1472.720 1410.210 ;
        RECT 1496.120 1396.840 1497.720 1417.210 ;
        RECT 1521.120 1396.840 1522.720 1410.210 ;
        RECT 1546.120 1396.840 1547.720 1417.210 ;
        RECT 1571.120 1396.840 1572.720 1410.210 ;
        RECT 1596.120 1396.840 1597.720 1417.210 ;
        RECT 1621.120 1396.840 1622.720 1410.210 ;
        RECT 1646.120 1396.840 1647.720 1417.210 ;
        RECT 1671.120 1396.840 1672.720 1410.210 ;
        RECT 1696.120 1396.840 1697.720 1417.210 ;
        RECT 1721.120 1396.840 1722.720 1410.210 ;
        RECT 1746.120 1396.840 1747.720 1417.210 ;
        RECT 1771.120 1396.840 1772.720 1410.210 ;
        RECT 1796.120 1396.840 1797.720 1417.210 ;
        RECT 1821.120 1396.840 1822.720 1410.210 ;
        RECT 1846.120 1396.840 1847.720 1417.210 ;
        RECT 1871.120 1396.840 1872.720 1410.210 ;
        RECT 1896.120 1396.840 1897.720 1417.210 ;
        RECT 1921.120 1396.840 1922.720 1410.210 ;
        RECT 1946.120 1396.840 1947.720 1417.210 ;
        RECT 1971.120 1396.840 1972.720 1410.210 ;
        RECT 1996.120 1396.840 1997.720 1417.210 ;
        RECT 2021.120 1396.840 2022.720 1410.210 ;
        RECT 2046.120 1396.840 2047.720 1417.210 ;
        RECT 2071.120 1396.840 2072.720 1410.210 ;
        RECT 2096.120 1396.840 2097.720 1417.210 ;
        RECT 2121.120 1396.840 2122.720 1410.210 ;
        RECT 2146.120 1396.840 2147.720 1417.210 ;
        RECT 2171.120 1396.840 2172.720 1410.210 ;
        RECT 2196.120 1396.840 2197.720 1417.210 ;
        RECT 2221.120 1396.840 2222.720 1410.210 ;
        RECT 2246.120 1396.840 2247.720 1417.210 ;
        RECT 2271.120 1396.840 2272.720 1410.210 ;
        RECT 2296.120 1396.840 2297.720 1417.210 ;
        RECT 2321.120 1396.840 2322.720 1410.210 ;
        RECT 2346.120 1396.840 2347.720 1417.210 ;
        RECT 2371.120 1396.840 2372.720 1410.210 ;
        RECT 2396.120 1396.840 2397.720 1417.210 ;
        RECT 2421.120 1396.840 2422.720 1410.210 ;
        RECT 2446.120 1396.840 2447.720 1417.210 ;
        RECT 2471.120 1396.840 2472.720 1410.210 ;
        RECT 2496.120 1396.840 2497.720 1417.210 ;
        RECT 2521.120 1396.840 2522.720 1410.210 ;
        RECT 2546.120 1396.840 2547.720 1417.210 ;
        RECT 2571.120 1396.840 2572.720 1410.210 ;
        RECT 2596.120 1396.840 2597.720 1417.210 ;
        RECT 2621.120 1396.840 2622.720 1410.210 ;
        RECT 2646.120 1396.840 2647.720 1417.210 ;
        RECT 2671.120 1396.840 2672.720 1410.210 ;
        RECT 2696.120 1396.840 2697.720 1417.210 ;
        RECT 2721.120 1396.840 2722.720 1410.210 ;
        RECT 2746.120 1396.840 2747.720 1417.210 ;
        RECT 2771.120 1396.840 2772.720 1410.210 ;
        RECT 471.120 388.390 472.720 408.760 ;
        RECT 496.120 395.390 497.720 408.760 ;
        RECT 521.120 388.390 522.720 408.760 ;
        RECT 536.360 350.000 545.860 400.390 ;
        RECT 548.760 350.000 559.010 400.390 ;
        RECT 560.610 350.000 570.860 400.390 ;
        RECT 574.140 350.000 584.390 400.390 ;
        RECT 585.990 350.000 596.240 400.390 ;
        RECT 599.140 350.000 608.640 400.390 ;
        RECT 621.120 388.390 622.720 408.760 ;
        RECT 646.120 395.390 647.720 408.760 ;
        RECT 671.120 388.390 672.720 408.760 ;
        RECT 696.120 395.390 697.720 408.760 ;
        RECT 721.120 388.390 722.720 408.760 ;
        RECT 746.120 395.390 747.720 408.760 ;
        RECT 771.120 388.390 772.720 408.760 ;
        RECT 796.120 395.390 797.720 408.760 ;
        RECT 821.120 388.390 822.720 408.760 ;
        RECT 846.120 395.390 847.720 408.760 ;
        RECT 871.120 388.390 872.720 408.760 ;
        RECT 896.120 395.390 897.720 408.760 ;
        RECT 921.120 388.390 922.720 408.760 ;
        RECT 946.120 395.390 947.720 408.760 ;
        RECT 971.120 388.390 972.720 408.760 ;
        RECT 996.120 395.390 997.720 408.760 ;
        RECT 1021.120 388.390 1022.720 408.760 ;
        RECT 1046.120 395.390 1047.720 408.760 ;
        RECT 1071.120 388.390 1072.720 408.760 ;
        RECT 1096.120 395.390 1097.720 408.760 ;
        RECT 1121.120 388.390 1122.720 408.760 ;
        RECT 1146.120 395.390 1147.720 408.760 ;
        RECT 1171.120 388.390 1172.720 408.760 ;
        RECT 1196.120 395.390 1197.720 408.760 ;
        RECT 1221.120 388.390 1222.720 408.760 ;
        RECT 1246.120 395.390 1247.720 408.760 ;
        RECT 1271.120 388.390 1272.720 408.760 ;
        RECT 1296.120 395.390 1297.720 408.760 ;
        RECT 1321.120 388.390 1322.720 408.760 ;
        RECT 1346.120 395.390 1347.720 408.760 ;
        RECT 1361.360 350.000 1370.860 400.390 ;
        RECT 1373.760 350.000 1384.010 400.390 ;
        RECT 1385.610 350.000 1395.860 400.390 ;
        RECT 1399.140 350.000 1409.390 400.390 ;
        RECT 1410.990 350.000 1421.240 400.390 ;
        RECT 1424.140 350.000 1433.640 400.390 ;
        RECT 1446.120 395.390 1447.720 408.760 ;
        RECT 1471.120 388.390 1472.720 408.760 ;
        RECT 1496.120 395.390 1497.720 408.760 ;
        RECT 1521.120 388.390 1522.720 408.760 ;
        RECT 1546.120 395.390 1547.720 408.760 ;
        RECT 1571.120 388.390 1572.720 408.760 ;
        RECT 1596.120 395.390 1597.720 408.760 ;
        RECT 1621.120 388.390 1622.720 408.760 ;
        RECT 1646.120 395.390 1647.720 408.760 ;
        RECT 1671.120 388.390 1672.720 408.760 ;
        RECT 1696.120 395.390 1697.720 408.760 ;
        RECT 1721.120 388.390 1722.720 408.760 ;
        RECT 1746.120 395.390 1747.720 408.760 ;
        RECT 1771.120 388.390 1772.720 408.760 ;
        RECT 1796.120 395.390 1797.720 408.760 ;
        RECT 1821.120 388.390 1822.720 408.760 ;
        RECT 1846.120 395.390 1847.720 408.760 ;
        RECT 1871.120 388.390 1872.720 408.760 ;
        RECT 1896.120 395.390 1897.720 408.760 ;
        RECT 1921.120 388.390 1922.720 408.760 ;
        RECT 1946.120 395.390 1947.720 408.760 ;
        RECT 1971.120 388.390 1972.720 408.760 ;
        RECT 1996.120 395.390 1997.720 408.760 ;
        RECT 2021.120 388.390 2022.720 408.760 ;
        RECT 2046.120 395.390 2047.720 408.760 ;
        RECT 2071.120 388.390 2072.720 408.760 ;
        RECT 2096.120 395.390 2097.720 408.760 ;
        RECT 2121.120 388.390 2122.720 408.760 ;
        RECT 2146.120 395.390 2147.720 408.760 ;
        RECT 2171.120 388.390 2172.720 408.760 ;
        RECT 2196.120 395.390 2197.720 408.760 ;
        RECT 2221.120 388.390 2222.720 408.760 ;
        RECT 2246.120 395.390 2247.720 408.760 ;
        RECT 2271.120 388.390 2272.720 408.760 ;
        RECT 2296.120 395.390 2297.720 408.760 ;
        RECT 2321.120 388.390 2322.720 408.760 ;
        RECT 2346.120 395.390 2347.720 408.760 ;
        RECT 2371.120 388.390 2372.720 408.760 ;
        RECT 2396.120 395.390 2397.720 408.760 ;
        RECT 2421.120 388.390 2422.720 408.760 ;
        RECT 2446.120 395.390 2447.720 408.760 ;
        RECT 2471.120 388.390 2472.720 408.760 ;
        RECT 2496.120 395.390 2497.720 408.760 ;
        RECT 2521.120 388.390 2522.720 408.760 ;
        RECT 2546.120 395.390 2547.720 408.760 ;
        RECT 2571.120 388.390 2572.720 408.760 ;
        RECT 2596.120 395.390 2597.720 408.760 ;
        RECT 2621.120 388.390 2622.720 408.760 ;
        RECT 2646.120 395.390 2647.720 408.760 ;
        RECT 2671.120 388.390 2672.720 408.760 ;
        RECT 2696.120 395.390 2697.720 408.760 ;
        RECT 2721.120 388.390 2722.720 408.760 ;
        RECT 2746.120 395.390 2747.720 408.760 ;
        RECT 2771.120 388.390 2772.720 408.760 ;
        RECT 2954.200 395.390 2959.200 1536.280 ;
        RECT 2961.200 388.390 2966.200 1529.280 ;
        RECT 3165.975 1524.280 3167.575 1571.420 ;
        RECT 3173.950 1531.280 3175.550 1571.420 ;
        RECT 3181.925 1524.280 3183.525 1571.420 ;
        RECT 3189.900 1531.280 3191.500 1571.420 ;
        RECT 3197.875 1524.280 3199.475 1571.420 ;
        RECT 3205.850 1531.280 3207.450 1571.420 ;
        RECT 3213.825 1524.280 3215.425 1571.420 ;
        RECT 3011.360 350.000 3020.860 400.390 ;
        RECT 3023.760 350.000 3034.010 400.390 ;
        RECT 3035.610 350.000 3045.860 400.390 ;
        RECT 3049.140 350.000 3059.390 400.390 ;
        RECT 3060.990 350.000 3071.240 400.390 ;
        RECT 3074.140 350.000 3083.640 400.390 ;
        RECT 3123.285 388.390 3124.885 423.750 ;
        RECT 3143.135 395.390 3144.735 423.750 ;
        RECT 3162.985 388.390 3164.585 423.750 ;
        RECT 3182.835 395.390 3184.435 423.750 ;
        RECT 3202.685 388.390 3204.285 423.750 ;
        RECT 3222.535 395.390 3224.135 423.750 ;
        RECT 3242.385 388.390 3243.985 423.750 ;
        RECT 3340.010 393.390 3344.010 497.895 ;
        RECT 3350.160 395.390 3354.160 497.895 ;
        RECT 3286.360 350.000 3295.860 393.390 ;
        RECT 3298.760 350.000 3309.010 393.390 ;
        RECT 3310.610 350.000 3320.860 393.390 ;
        RECT 3324.140 350.000 3334.390 393.390 ;
        RECT 3335.990 350.000 3346.240 393.390 ;
        RECT 3349.140 350.000 3358.640 393.390 ;
        RECT 3489.610 374.450 3494.610 4704.610 ;
        RECT 3496.610 376.450 3501.610 4711.610 ;
        RECT 3539.000 4409.140 3540.000 4418.640 ;
        RECT 3539.000 4395.990 3540.000 4406.240 ;
        RECT 3539.000 4384.140 3540.000 4394.390 ;
        RECT 3539.000 4370.610 3540.000 4380.860 ;
        RECT 3539.000 4358.760 3540.000 4369.010 ;
        RECT 3539.000 4346.360 3540.000 4355.860 ;
        RECT 3539.000 3979.140 3540.000 3988.640 ;
        RECT 3539.000 3965.990 3540.000 3976.240 ;
        RECT 3539.000 3954.140 3540.000 3964.390 ;
        RECT 3539.000 3940.610 3540.000 3950.860 ;
        RECT 3539.000 3928.760 3540.000 3939.010 ;
        RECT 3539.000 3916.360 3540.000 3925.860 ;
        RECT 3539.000 2474.140 3540.000 2483.640 ;
        RECT 3539.000 2460.990 3540.000 2471.240 ;
        RECT 3539.000 2449.140 3540.000 2459.390 ;
        RECT 3539.000 2435.610 3540.000 2445.860 ;
        RECT 3539.000 2423.760 3540.000 2434.010 ;
        RECT 3539.000 2411.360 3540.000 2420.860 ;
        RECT 3539.005 2259.140 3540.005 2268.640 ;
        RECT 3539.005 2245.990 3540.005 2256.240 ;
        RECT 3539.005 2234.140 3540.005 2244.390 ;
        RECT 3539.005 2220.610 3540.005 2230.860 ;
        RECT 3539.005 2208.760 3540.005 2219.010 ;
        RECT 3539.005 2196.360 3540.005 2205.860 ;
        RECT 3539.000 2044.140 3540.000 2053.640 ;
        RECT 3539.000 2030.990 3540.000 2041.240 ;
        RECT 3539.000 2019.140 3540.000 2029.390 ;
        RECT 3539.000 2005.610 3540.000 2015.860 ;
        RECT 3539.000 1993.760 3540.000 2004.010 ;
        RECT 3539.000 1981.360 3540.000 1990.860 ;
      LAYER VIA4 ;
        RECT 395.965 4729.920 396.245 4730.200 ;
        RECT 396.585 4729.920 396.865 4730.200 ;
        RECT 397.205 4729.920 397.485 4730.200 ;
        RECT 397.825 4729.920 398.105 4730.200 ;
        RECT 398.445 4729.920 398.725 4730.200 ;
        RECT 399.065 4729.920 399.345 4730.200 ;
        RECT 399.685 4729.920 399.965 4730.200 ;
        RECT 388.965 4727.920 389.245 4728.200 ;
        RECT 389.585 4727.920 389.865 4728.200 ;
        RECT 390.205 4727.920 390.485 4728.200 ;
        RECT 390.825 4727.920 391.105 4728.200 ;
        RECT 391.445 4727.920 391.725 4728.200 ;
        RECT 392.065 4727.920 392.345 4728.200 ;
        RECT 392.685 4727.920 392.965 4728.200 ;
        RECT 388.740 4710.980 389.020 4711.260 ;
        RECT 389.360 4710.980 389.640 4711.260 ;
        RECT 389.980 4710.980 390.260 4711.260 ;
        RECT 390.600 4710.980 390.880 4711.260 ;
        RECT 391.220 4710.980 391.500 4711.260 ;
        RECT 391.840 4710.980 392.120 4711.260 ;
        RECT 392.460 4710.980 392.740 4711.260 ;
        RECT 388.740 4710.360 389.020 4710.640 ;
        RECT 389.360 4710.360 389.640 4710.640 ;
        RECT 389.980 4710.360 390.260 4710.640 ;
        RECT 390.600 4710.360 390.880 4710.640 ;
        RECT 391.220 4710.360 391.500 4710.640 ;
        RECT 391.840 4710.360 392.120 4710.640 ;
        RECT 392.460 4710.360 392.740 4710.640 ;
        RECT 388.740 4709.740 389.020 4710.020 ;
        RECT 389.360 4709.740 389.640 4710.020 ;
        RECT 389.980 4709.740 390.260 4710.020 ;
        RECT 390.600 4709.740 390.880 4710.020 ;
        RECT 391.220 4709.740 391.500 4710.020 ;
        RECT 391.840 4709.740 392.120 4710.020 ;
        RECT 392.460 4709.740 392.740 4710.020 ;
        RECT 388.740 4709.120 389.020 4709.400 ;
        RECT 389.360 4709.120 389.640 4709.400 ;
        RECT 389.980 4709.120 390.260 4709.400 ;
        RECT 390.600 4709.120 390.880 4709.400 ;
        RECT 391.220 4709.120 391.500 4709.400 ;
        RECT 391.840 4709.120 392.120 4709.400 ;
        RECT 392.460 4709.120 392.740 4709.400 ;
        RECT 388.740 4708.500 389.020 4708.780 ;
        RECT 389.360 4708.500 389.640 4708.780 ;
        RECT 389.980 4708.500 390.260 4708.780 ;
        RECT 390.600 4708.500 390.880 4708.780 ;
        RECT 391.220 4708.500 391.500 4708.780 ;
        RECT 391.840 4708.500 392.120 4708.780 ;
        RECT 392.460 4708.500 392.740 4708.780 ;
        RECT 388.740 4707.880 389.020 4708.160 ;
        RECT 389.360 4707.880 389.640 4708.160 ;
        RECT 389.980 4707.880 390.260 4708.160 ;
        RECT 390.600 4707.880 390.880 4708.160 ;
        RECT 391.220 4707.880 391.500 4708.160 ;
        RECT 391.840 4707.880 392.120 4708.160 ;
        RECT 392.460 4707.880 392.740 4708.160 ;
        RECT 388.740 4707.260 389.020 4707.540 ;
        RECT 389.360 4707.260 389.640 4707.540 ;
        RECT 389.980 4707.260 390.260 4707.540 ;
        RECT 390.600 4707.260 390.880 4707.540 ;
        RECT 391.220 4707.260 391.500 4707.540 ;
        RECT 391.840 4707.260 392.120 4707.540 ;
        RECT 392.460 4707.260 392.740 4707.540 ;
        RECT 388.965 4630.590 389.245 4630.870 ;
        RECT 389.585 4630.590 389.865 4630.870 ;
        RECT 390.205 4630.590 390.485 4630.870 ;
        RECT 390.825 4630.590 391.105 4630.870 ;
        RECT 391.445 4630.590 391.725 4630.870 ;
        RECT 392.065 4630.590 392.345 4630.870 ;
        RECT 392.685 4630.590 392.965 4630.870 ;
        RECT 388.965 4629.970 389.245 4630.250 ;
        RECT 389.585 4629.970 389.865 4630.250 ;
        RECT 390.205 4629.970 390.485 4630.250 ;
        RECT 390.825 4629.970 391.105 4630.250 ;
        RECT 391.445 4629.970 391.725 4630.250 ;
        RECT 392.065 4629.970 392.345 4630.250 ;
        RECT 392.685 4629.970 392.965 4630.250 ;
        RECT 388.965 4595.590 389.245 4595.870 ;
        RECT 389.585 4595.590 389.865 4595.870 ;
        RECT 390.205 4595.590 390.485 4595.870 ;
        RECT 390.825 4595.590 391.105 4595.870 ;
        RECT 391.445 4595.590 391.725 4595.870 ;
        RECT 392.065 4595.590 392.345 4595.870 ;
        RECT 392.685 4595.590 392.965 4595.870 ;
        RECT 388.965 4594.970 389.245 4595.250 ;
        RECT 389.585 4594.970 389.865 4595.250 ;
        RECT 390.205 4594.970 390.485 4595.250 ;
        RECT 390.825 4594.970 391.105 4595.250 ;
        RECT 391.445 4594.970 391.725 4595.250 ;
        RECT 392.065 4594.970 392.345 4595.250 ;
        RECT 392.685 4594.970 392.965 4595.250 ;
        RECT 388.740 4572.670 389.020 4572.950 ;
        RECT 389.360 4572.670 389.640 4572.950 ;
        RECT 389.980 4572.670 390.260 4572.950 ;
        RECT 390.600 4572.670 390.880 4572.950 ;
        RECT 391.220 4572.670 391.500 4572.950 ;
        RECT 391.840 4572.670 392.120 4572.950 ;
        RECT 392.460 4572.670 392.740 4572.950 ;
        RECT 388.740 4572.050 389.020 4572.330 ;
        RECT 389.360 4572.050 389.640 4572.330 ;
        RECT 389.980 4572.050 390.260 4572.330 ;
        RECT 390.600 4572.050 390.880 4572.330 ;
        RECT 391.220 4572.050 391.500 4572.330 ;
        RECT 391.840 4572.050 392.120 4572.330 ;
        RECT 392.460 4572.050 392.740 4572.330 ;
        RECT 388.740 4571.430 389.020 4571.710 ;
        RECT 389.360 4571.430 389.640 4571.710 ;
        RECT 389.980 4571.430 390.260 4571.710 ;
        RECT 390.600 4571.430 390.880 4571.710 ;
        RECT 391.220 4571.430 391.500 4571.710 ;
        RECT 391.840 4571.430 392.120 4571.710 ;
        RECT 392.460 4571.430 392.740 4571.710 ;
        RECT 388.740 4570.810 389.020 4571.090 ;
        RECT 389.360 4570.810 389.640 4571.090 ;
        RECT 389.980 4570.810 390.260 4571.090 ;
        RECT 390.600 4570.810 390.880 4571.090 ;
        RECT 391.220 4570.810 391.500 4571.090 ;
        RECT 391.840 4570.810 392.120 4571.090 ;
        RECT 392.460 4570.810 392.740 4571.090 ;
        RECT 388.740 4570.190 389.020 4570.470 ;
        RECT 389.360 4570.190 389.640 4570.470 ;
        RECT 389.980 4570.190 390.260 4570.470 ;
        RECT 390.600 4570.190 390.880 4570.470 ;
        RECT 391.220 4570.190 391.500 4570.470 ;
        RECT 391.840 4570.190 392.120 4570.470 ;
        RECT 392.460 4570.190 392.740 4570.470 ;
        RECT 388.965 4560.590 389.245 4560.870 ;
        RECT 389.585 4560.590 389.865 4560.870 ;
        RECT 390.205 4560.590 390.485 4560.870 ;
        RECT 390.825 4560.590 391.105 4560.870 ;
        RECT 391.445 4560.590 391.725 4560.870 ;
        RECT 392.065 4560.590 392.345 4560.870 ;
        RECT 392.685 4560.590 392.965 4560.870 ;
        RECT 388.965 4559.970 389.245 4560.250 ;
        RECT 389.585 4559.970 389.865 4560.250 ;
        RECT 390.205 4559.970 390.485 4560.250 ;
        RECT 390.825 4559.970 391.105 4560.250 ;
        RECT 391.445 4559.970 391.725 4560.250 ;
        RECT 392.065 4559.970 392.345 4560.250 ;
        RECT 392.685 4559.970 392.965 4560.250 ;
        RECT 350.370 4423.010 350.650 4423.290 ;
        RECT 350.370 4422.390 350.650 4422.670 ;
        RECT 350.370 4421.770 350.650 4422.050 ;
        RECT 350.370 4421.150 350.650 4421.430 ;
        RECT 350.370 4420.530 350.650 4420.810 ;
        RECT 350.370 4419.910 350.650 4420.190 ;
        RECT 350.370 4419.290 350.650 4419.570 ;
        RECT 350.370 4418.670 350.650 4418.950 ;
        RECT 350.370 4418.050 350.650 4418.330 ;
        RECT 350.370 4417.430 350.650 4417.710 ;
        RECT 350.370 4416.810 350.650 4417.090 ;
        RECT 350.370 4416.190 350.650 4416.470 ;
        RECT 350.370 4415.570 350.650 4415.850 ;
        RECT 350.370 4414.950 350.650 4415.230 ;
        RECT 350.370 4414.330 350.650 4414.610 ;
        RECT 389.040 4423.070 389.320 4423.350 ;
        RECT 389.660 4423.070 389.940 4423.350 ;
        RECT 390.280 4423.070 390.560 4423.350 ;
        RECT 390.900 4423.070 391.180 4423.350 ;
        RECT 391.520 4423.070 391.800 4423.350 ;
        RECT 392.140 4423.070 392.420 4423.350 ;
        RECT 392.760 4423.070 393.040 4423.350 ;
        RECT 389.040 4422.450 389.320 4422.730 ;
        RECT 389.660 4422.450 389.940 4422.730 ;
        RECT 390.280 4422.450 390.560 4422.730 ;
        RECT 390.900 4422.450 391.180 4422.730 ;
        RECT 391.520 4422.450 391.800 4422.730 ;
        RECT 392.140 4422.450 392.420 4422.730 ;
        RECT 392.760 4422.450 393.040 4422.730 ;
        RECT 389.040 4421.830 389.320 4422.110 ;
        RECT 389.660 4421.830 389.940 4422.110 ;
        RECT 390.280 4421.830 390.560 4422.110 ;
        RECT 390.900 4421.830 391.180 4422.110 ;
        RECT 391.520 4421.830 391.800 4422.110 ;
        RECT 392.140 4421.830 392.420 4422.110 ;
        RECT 392.760 4421.830 393.040 4422.110 ;
        RECT 389.040 4421.210 389.320 4421.490 ;
        RECT 389.660 4421.210 389.940 4421.490 ;
        RECT 390.280 4421.210 390.560 4421.490 ;
        RECT 390.900 4421.210 391.180 4421.490 ;
        RECT 391.520 4421.210 391.800 4421.490 ;
        RECT 392.140 4421.210 392.420 4421.490 ;
        RECT 392.760 4421.210 393.040 4421.490 ;
        RECT 389.040 4420.590 389.320 4420.870 ;
        RECT 389.660 4420.590 389.940 4420.870 ;
        RECT 390.280 4420.590 390.560 4420.870 ;
        RECT 390.900 4420.590 391.180 4420.870 ;
        RECT 391.520 4420.590 391.800 4420.870 ;
        RECT 392.140 4420.590 392.420 4420.870 ;
        RECT 392.760 4420.590 393.040 4420.870 ;
        RECT 389.040 4419.970 389.320 4420.250 ;
        RECT 389.660 4419.970 389.940 4420.250 ;
        RECT 390.280 4419.970 390.560 4420.250 ;
        RECT 390.900 4419.970 391.180 4420.250 ;
        RECT 391.520 4419.970 391.800 4420.250 ;
        RECT 392.140 4419.970 392.420 4420.250 ;
        RECT 392.760 4419.970 393.040 4420.250 ;
        RECT 389.040 4419.350 389.320 4419.630 ;
        RECT 389.660 4419.350 389.940 4419.630 ;
        RECT 390.280 4419.350 390.560 4419.630 ;
        RECT 390.900 4419.350 391.180 4419.630 ;
        RECT 391.520 4419.350 391.800 4419.630 ;
        RECT 392.140 4419.350 392.420 4419.630 ;
        RECT 392.760 4419.350 393.040 4419.630 ;
        RECT 389.040 4418.730 389.320 4419.010 ;
        RECT 389.660 4418.730 389.940 4419.010 ;
        RECT 390.280 4418.730 390.560 4419.010 ;
        RECT 390.900 4418.730 391.180 4419.010 ;
        RECT 391.520 4418.730 391.800 4419.010 ;
        RECT 392.140 4418.730 392.420 4419.010 ;
        RECT 392.760 4418.730 393.040 4419.010 ;
        RECT 389.040 4418.110 389.320 4418.390 ;
        RECT 389.660 4418.110 389.940 4418.390 ;
        RECT 390.280 4418.110 390.560 4418.390 ;
        RECT 390.900 4418.110 391.180 4418.390 ;
        RECT 391.520 4418.110 391.800 4418.390 ;
        RECT 392.140 4418.110 392.420 4418.390 ;
        RECT 392.760 4418.110 393.040 4418.390 ;
        RECT 389.040 4417.490 389.320 4417.770 ;
        RECT 389.660 4417.490 389.940 4417.770 ;
        RECT 390.280 4417.490 390.560 4417.770 ;
        RECT 390.900 4417.490 391.180 4417.770 ;
        RECT 391.520 4417.490 391.800 4417.770 ;
        RECT 392.140 4417.490 392.420 4417.770 ;
        RECT 392.760 4417.490 393.040 4417.770 ;
        RECT 389.040 4416.870 389.320 4417.150 ;
        RECT 389.660 4416.870 389.940 4417.150 ;
        RECT 390.280 4416.870 390.560 4417.150 ;
        RECT 390.900 4416.870 391.180 4417.150 ;
        RECT 391.520 4416.870 391.800 4417.150 ;
        RECT 392.140 4416.870 392.420 4417.150 ;
        RECT 392.760 4416.870 393.040 4417.150 ;
        RECT 389.040 4416.250 389.320 4416.530 ;
        RECT 389.660 4416.250 389.940 4416.530 ;
        RECT 390.280 4416.250 390.560 4416.530 ;
        RECT 390.900 4416.250 391.180 4416.530 ;
        RECT 391.520 4416.250 391.800 4416.530 ;
        RECT 392.140 4416.250 392.420 4416.530 ;
        RECT 392.760 4416.250 393.040 4416.530 ;
        RECT 389.040 4415.630 389.320 4415.910 ;
        RECT 389.660 4415.630 389.940 4415.910 ;
        RECT 390.280 4415.630 390.560 4415.910 ;
        RECT 390.900 4415.630 391.180 4415.910 ;
        RECT 391.520 4415.630 391.800 4415.910 ;
        RECT 392.140 4415.630 392.420 4415.910 ;
        RECT 392.760 4415.630 393.040 4415.910 ;
        RECT 389.040 4415.010 389.320 4415.290 ;
        RECT 389.660 4415.010 389.940 4415.290 ;
        RECT 390.280 4415.010 390.560 4415.290 ;
        RECT 390.900 4415.010 391.180 4415.290 ;
        RECT 391.520 4415.010 391.800 4415.290 ;
        RECT 392.140 4415.010 392.420 4415.290 ;
        RECT 392.760 4415.010 393.040 4415.290 ;
        RECT 389.040 4414.390 389.320 4414.670 ;
        RECT 389.660 4414.390 389.940 4414.670 ;
        RECT 390.280 4414.390 390.560 4414.670 ;
        RECT 390.900 4414.390 391.180 4414.670 ;
        RECT 391.520 4414.390 391.800 4414.670 ;
        RECT 392.140 4414.390 392.420 4414.670 ;
        RECT 392.760 4414.390 393.040 4414.670 ;
        RECT 350.370 4410.640 350.650 4410.920 ;
        RECT 350.370 4410.020 350.650 4410.300 ;
        RECT 350.370 4409.400 350.650 4409.680 ;
        RECT 350.370 4408.780 350.650 4409.060 ;
        RECT 350.370 4408.160 350.650 4408.440 ;
        RECT 350.370 4407.540 350.650 4407.820 ;
        RECT 350.370 4406.920 350.650 4407.200 ;
        RECT 350.370 4406.300 350.650 4406.580 ;
        RECT 350.370 4405.680 350.650 4405.960 ;
        RECT 350.370 4405.060 350.650 4405.340 ;
        RECT 350.370 4404.440 350.650 4404.720 ;
        RECT 350.370 4403.820 350.650 4404.100 ;
        RECT 350.370 4403.200 350.650 4403.480 ;
        RECT 350.370 4402.580 350.650 4402.860 ;
        RECT 350.370 4401.960 350.650 4402.240 ;
        RECT 350.370 4401.340 350.650 4401.620 ;
        RECT 389.040 4410.670 389.320 4410.950 ;
        RECT 389.660 4410.670 389.940 4410.950 ;
        RECT 390.280 4410.670 390.560 4410.950 ;
        RECT 390.900 4410.670 391.180 4410.950 ;
        RECT 391.520 4410.670 391.800 4410.950 ;
        RECT 392.140 4410.670 392.420 4410.950 ;
        RECT 392.760 4410.670 393.040 4410.950 ;
        RECT 389.040 4410.050 389.320 4410.330 ;
        RECT 389.660 4410.050 389.940 4410.330 ;
        RECT 390.280 4410.050 390.560 4410.330 ;
        RECT 390.900 4410.050 391.180 4410.330 ;
        RECT 391.520 4410.050 391.800 4410.330 ;
        RECT 392.140 4410.050 392.420 4410.330 ;
        RECT 392.760 4410.050 393.040 4410.330 ;
        RECT 389.040 4409.430 389.320 4409.710 ;
        RECT 389.660 4409.430 389.940 4409.710 ;
        RECT 390.280 4409.430 390.560 4409.710 ;
        RECT 390.900 4409.430 391.180 4409.710 ;
        RECT 391.520 4409.430 391.800 4409.710 ;
        RECT 392.140 4409.430 392.420 4409.710 ;
        RECT 392.760 4409.430 393.040 4409.710 ;
        RECT 389.040 4408.810 389.320 4409.090 ;
        RECT 389.660 4408.810 389.940 4409.090 ;
        RECT 390.280 4408.810 390.560 4409.090 ;
        RECT 390.900 4408.810 391.180 4409.090 ;
        RECT 391.520 4408.810 391.800 4409.090 ;
        RECT 392.140 4408.810 392.420 4409.090 ;
        RECT 392.760 4408.810 393.040 4409.090 ;
        RECT 389.040 4408.190 389.320 4408.470 ;
        RECT 389.660 4408.190 389.940 4408.470 ;
        RECT 390.280 4408.190 390.560 4408.470 ;
        RECT 390.900 4408.190 391.180 4408.470 ;
        RECT 391.520 4408.190 391.800 4408.470 ;
        RECT 392.140 4408.190 392.420 4408.470 ;
        RECT 392.760 4408.190 393.040 4408.470 ;
        RECT 389.040 4407.570 389.320 4407.850 ;
        RECT 389.660 4407.570 389.940 4407.850 ;
        RECT 390.280 4407.570 390.560 4407.850 ;
        RECT 390.900 4407.570 391.180 4407.850 ;
        RECT 391.520 4407.570 391.800 4407.850 ;
        RECT 392.140 4407.570 392.420 4407.850 ;
        RECT 392.760 4407.570 393.040 4407.850 ;
        RECT 389.040 4406.950 389.320 4407.230 ;
        RECT 389.660 4406.950 389.940 4407.230 ;
        RECT 390.280 4406.950 390.560 4407.230 ;
        RECT 390.900 4406.950 391.180 4407.230 ;
        RECT 391.520 4406.950 391.800 4407.230 ;
        RECT 392.140 4406.950 392.420 4407.230 ;
        RECT 392.760 4406.950 393.040 4407.230 ;
        RECT 389.040 4406.330 389.320 4406.610 ;
        RECT 389.660 4406.330 389.940 4406.610 ;
        RECT 390.280 4406.330 390.560 4406.610 ;
        RECT 390.900 4406.330 391.180 4406.610 ;
        RECT 391.520 4406.330 391.800 4406.610 ;
        RECT 392.140 4406.330 392.420 4406.610 ;
        RECT 392.760 4406.330 393.040 4406.610 ;
        RECT 389.040 4405.710 389.320 4405.990 ;
        RECT 389.660 4405.710 389.940 4405.990 ;
        RECT 390.280 4405.710 390.560 4405.990 ;
        RECT 390.900 4405.710 391.180 4405.990 ;
        RECT 391.520 4405.710 391.800 4405.990 ;
        RECT 392.140 4405.710 392.420 4405.990 ;
        RECT 392.760 4405.710 393.040 4405.990 ;
        RECT 389.040 4405.090 389.320 4405.370 ;
        RECT 389.660 4405.090 389.940 4405.370 ;
        RECT 390.280 4405.090 390.560 4405.370 ;
        RECT 390.900 4405.090 391.180 4405.370 ;
        RECT 391.520 4405.090 391.800 4405.370 ;
        RECT 392.140 4405.090 392.420 4405.370 ;
        RECT 392.760 4405.090 393.040 4405.370 ;
        RECT 389.040 4404.470 389.320 4404.750 ;
        RECT 389.660 4404.470 389.940 4404.750 ;
        RECT 390.280 4404.470 390.560 4404.750 ;
        RECT 390.900 4404.470 391.180 4404.750 ;
        RECT 391.520 4404.470 391.800 4404.750 ;
        RECT 392.140 4404.470 392.420 4404.750 ;
        RECT 392.760 4404.470 393.040 4404.750 ;
        RECT 389.040 4403.850 389.320 4404.130 ;
        RECT 389.660 4403.850 389.940 4404.130 ;
        RECT 390.280 4403.850 390.560 4404.130 ;
        RECT 390.900 4403.850 391.180 4404.130 ;
        RECT 391.520 4403.850 391.800 4404.130 ;
        RECT 392.140 4403.850 392.420 4404.130 ;
        RECT 392.760 4403.850 393.040 4404.130 ;
        RECT 389.040 4403.230 389.320 4403.510 ;
        RECT 389.660 4403.230 389.940 4403.510 ;
        RECT 390.280 4403.230 390.560 4403.510 ;
        RECT 390.900 4403.230 391.180 4403.510 ;
        RECT 391.520 4403.230 391.800 4403.510 ;
        RECT 392.140 4403.230 392.420 4403.510 ;
        RECT 392.760 4403.230 393.040 4403.510 ;
        RECT 389.040 4402.610 389.320 4402.890 ;
        RECT 389.660 4402.610 389.940 4402.890 ;
        RECT 390.280 4402.610 390.560 4402.890 ;
        RECT 390.900 4402.610 391.180 4402.890 ;
        RECT 391.520 4402.610 391.800 4402.890 ;
        RECT 392.140 4402.610 392.420 4402.890 ;
        RECT 392.760 4402.610 393.040 4402.890 ;
        RECT 389.040 4401.990 389.320 4402.270 ;
        RECT 389.660 4401.990 389.940 4402.270 ;
        RECT 390.280 4401.990 390.560 4402.270 ;
        RECT 390.900 4401.990 391.180 4402.270 ;
        RECT 391.520 4401.990 391.800 4402.270 ;
        RECT 392.140 4401.990 392.420 4402.270 ;
        RECT 392.760 4401.990 393.040 4402.270 ;
        RECT 389.040 4401.370 389.320 4401.650 ;
        RECT 389.660 4401.370 389.940 4401.650 ;
        RECT 390.280 4401.370 390.560 4401.650 ;
        RECT 390.900 4401.370 391.180 4401.650 ;
        RECT 391.520 4401.370 391.800 4401.650 ;
        RECT 392.140 4401.370 392.420 4401.650 ;
        RECT 392.760 4401.370 393.040 4401.650 ;
        RECT 350.370 4398.790 350.650 4399.070 ;
        RECT 350.370 4398.170 350.650 4398.450 ;
        RECT 350.370 4397.550 350.650 4397.830 ;
        RECT 350.370 4396.930 350.650 4397.210 ;
        RECT 350.370 4396.310 350.650 4396.590 ;
        RECT 350.370 4395.690 350.650 4395.970 ;
        RECT 350.370 4395.070 350.650 4395.350 ;
        RECT 350.370 4394.450 350.650 4394.730 ;
        RECT 350.370 4393.830 350.650 4394.110 ;
        RECT 350.370 4393.210 350.650 4393.490 ;
        RECT 350.370 4392.590 350.650 4392.870 ;
        RECT 350.370 4391.970 350.650 4392.250 ;
        RECT 350.370 4391.350 350.650 4391.630 ;
        RECT 350.370 4390.730 350.650 4391.010 ;
        RECT 350.370 4390.110 350.650 4390.390 ;
        RECT 350.370 4389.490 350.650 4389.770 ;
        RECT 389.040 4398.820 389.320 4399.100 ;
        RECT 389.660 4398.820 389.940 4399.100 ;
        RECT 390.280 4398.820 390.560 4399.100 ;
        RECT 390.900 4398.820 391.180 4399.100 ;
        RECT 391.520 4398.820 391.800 4399.100 ;
        RECT 392.140 4398.820 392.420 4399.100 ;
        RECT 392.760 4398.820 393.040 4399.100 ;
        RECT 389.040 4398.200 389.320 4398.480 ;
        RECT 389.660 4398.200 389.940 4398.480 ;
        RECT 390.280 4398.200 390.560 4398.480 ;
        RECT 390.900 4398.200 391.180 4398.480 ;
        RECT 391.520 4398.200 391.800 4398.480 ;
        RECT 392.140 4398.200 392.420 4398.480 ;
        RECT 392.760 4398.200 393.040 4398.480 ;
        RECT 389.040 4397.580 389.320 4397.860 ;
        RECT 389.660 4397.580 389.940 4397.860 ;
        RECT 390.280 4397.580 390.560 4397.860 ;
        RECT 390.900 4397.580 391.180 4397.860 ;
        RECT 391.520 4397.580 391.800 4397.860 ;
        RECT 392.140 4397.580 392.420 4397.860 ;
        RECT 392.760 4397.580 393.040 4397.860 ;
        RECT 389.040 4396.960 389.320 4397.240 ;
        RECT 389.660 4396.960 389.940 4397.240 ;
        RECT 390.280 4396.960 390.560 4397.240 ;
        RECT 390.900 4396.960 391.180 4397.240 ;
        RECT 391.520 4396.960 391.800 4397.240 ;
        RECT 392.140 4396.960 392.420 4397.240 ;
        RECT 392.760 4396.960 393.040 4397.240 ;
        RECT 389.040 4396.340 389.320 4396.620 ;
        RECT 389.660 4396.340 389.940 4396.620 ;
        RECT 390.280 4396.340 390.560 4396.620 ;
        RECT 390.900 4396.340 391.180 4396.620 ;
        RECT 391.520 4396.340 391.800 4396.620 ;
        RECT 392.140 4396.340 392.420 4396.620 ;
        RECT 392.760 4396.340 393.040 4396.620 ;
        RECT 389.040 4395.720 389.320 4396.000 ;
        RECT 389.660 4395.720 389.940 4396.000 ;
        RECT 390.280 4395.720 390.560 4396.000 ;
        RECT 390.900 4395.720 391.180 4396.000 ;
        RECT 391.520 4395.720 391.800 4396.000 ;
        RECT 392.140 4395.720 392.420 4396.000 ;
        RECT 392.760 4395.720 393.040 4396.000 ;
        RECT 389.040 4395.100 389.320 4395.380 ;
        RECT 389.660 4395.100 389.940 4395.380 ;
        RECT 390.280 4395.100 390.560 4395.380 ;
        RECT 390.900 4395.100 391.180 4395.380 ;
        RECT 391.520 4395.100 391.800 4395.380 ;
        RECT 392.140 4395.100 392.420 4395.380 ;
        RECT 392.760 4395.100 393.040 4395.380 ;
        RECT 389.040 4394.480 389.320 4394.760 ;
        RECT 389.660 4394.480 389.940 4394.760 ;
        RECT 390.280 4394.480 390.560 4394.760 ;
        RECT 390.900 4394.480 391.180 4394.760 ;
        RECT 391.520 4394.480 391.800 4394.760 ;
        RECT 392.140 4394.480 392.420 4394.760 ;
        RECT 392.760 4394.480 393.040 4394.760 ;
        RECT 389.040 4393.860 389.320 4394.140 ;
        RECT 389.660 4393.860 389.940 4394.140 ;
        RECT 390.280 4393.860 390.560 4394.140 ;
        RECT 390.900 4393.860 391.180 4394.140 ;
        RECT 391.520 4393.860 391.800 4394.140 ;
        RECT 392.140 4393.860 392.420 4394.140 ;
        RECT 392.760 4393.860 393.040 4394.140 ;
        RECT 389.040 4393.240 389.320 4393.520 ;
        RECT 389.660 4393.240 389.940 4393.520 ;
        RECT 390.280 4393.240 390.560 4393.520 ;
        RECT 390.900 4393.240 391.180 4393.520 ;
        RECT 391.520 4393.240 391.800 4393.520 ;
        RECT 392.140 4393.240 392.420 4393.520 ;
        RECT 392.760 4393.240 393.040 4393.520 ;
        RECT 389.040 4392.620 389.320 4392.900 ;
        RECT 389.660 4392.620 389.940 4392.900 ;
        RECT 390.280 4392.620 390.560 4392.900 ;
        RECT 390.900 4392.620 391.180 4392.900 ;
        RECT 391.520 4392.620 391.800 4392.900 ;
        RECT 392.140 4392.620 392.420 4392.900 ;
        RECT 392.760 4392.620 393.040 4392.900 ;
        RECT 389.040 4392.000 389.320 4392.280 ;
        RECT 389.660 4392.000 389.940 4392.280 ;
        RECT 390.280 4392.000 390.560 4392.280 ;
        RECT 390.900 4392.000 391.180 4392.280 ;
        RECT 391.520 4392.000 391.800 4392.280 ;
        RECT 392.140 4392.000 392.420 4392.280 ;
        RECT 392.760 4392.000 393.040 4392.280 ;
        RECT 389.040 4391.380 389.320 4391.660 ;
        RECT 389.660 4391.380 389.940 4391.660 ;
        RECT 390.280 4391.380 390.560 4391.660 ;
        RECT 390.900 4391.380 391.180 4391.660 ;
        RECT 391.520 4391.380 391.800 4391.660 ;
        RECT 392.140 4391.380 392.420 4391.660 ;
        RECT 392.760 4391.380 393.040 4391.660 ;
        RECT 389.040 4390.760 389.320 4391.040 ;
        RECT 389.660 4390.760 389.940 4391.040 ;
        RECT 390.280 4390.760 390.560 4391.040 ;
        RECT 390.900 4390.760 391.180 4391.040 ;
        RECT 391.520 4390.760 391.800 4391.040 ;
        RECT 392.140 4390.760 392.420 4391.040 ;
        RECT 392.760 4390.760 393.040 4391.040 ;
        RECT 389.040 4390.140 389.320 4390.420 ;
        RECT 389.660 4390.140 389.940 4390.420 ;
        RECT 390.280 4390.140 390.560 4390.420 ;
        RECT 390.900 4390.140 391.180 4390.420 ;
        RECT 391.520 4390.140 391.800 4390.420 ;
        RECT 392.140 4390.140 392.420 4390.420 ;
        RECT 392.760 4390.140 393.040 4390.420 ;
        RECT 389.040 4389.520 389.320 4389.800 ;
        RECT 389.660 4389.520 389.940 4389.800 ;
        RECT 390.280 4389.520 390.560 4389.800 ;
        RECT 390.900 4389.520 391.180 4389.800 ;
        RECT 391.520 4389.520 391.800 4389.800 ;
        RECT 392.140 4389.520 392.420 4389.800 ;
        RECT 392.760 4389.520 393.040 4389.800 ;
        RECT 350.370 4385.260 350.650 4385.540 ;
        RECT 350.370 4384.640 350.650 4384.920 ;
        RECT 350.370 4384.020 350.650 4384.300 ;
        RECT 350.370 4383.400 350.650 4383.680 ;
        RECT 350.370 4382.780 350.650 4383.060 ;
        RECT 350.370 4382.160 350.650 4382.440 ;
        RECT 350.370 4381.540 350.650 4381.820 ;
        RECT 350.370 4380.920 350.650 4381.200 ;
        RECT 350.370 4380.300 350.650 4380.580 ;
        RECT 350.370 4379.680 350.650 4379.960 ;
        RECT 350.370 4379.060 350.650 4379.340 ;
        RECT 350.370 4378.440 350.650 4378.720 ;
        RECT 350.370 4377.820 350.650 4378.100 ;
        RECT 350.370 4377.200 350.650 4377.480 ;
        RECT 350.370 4376.580 350.650 4376.860 ;
        RECT 350.370 4375.960 350.650 4376.240 ;
        RECT 389.040 4385.290 389.320 4385.570 ;
        RECT 389.660 4385.290 389.940 4385.570 ;
        RECT 390.280 4385.290 390.560 4385.570 ;
        RECT 390.900 4385.290 391.180 4385.570 ;
        RECT 391.520 4385.290 391.800 4385.570 ;
        RECT 392.140 4385.290 392.420 4385.570 ;
        RECT 392.760 4385.290 393.040 4385.570 ;
        RECT 389.040 4384.670 389.320 4384.950 ;
        RECT 389.660 4384.670 389.940 4384.950 ;
        RECT 390.280 4384.670 390.560 4384.950 ;
        RECT 390.900 4384.670 391.180 4384.950 ;
        RECT 391.520 4384.670 391.800 4384.950 ;
        RECT 392.140 4384.670 392.420 4384.950 ;
        RECT 392.760 4384.670 393.040 4384.950 ;
        RECT 389.040 4384.050 389.320 4384.330 ;
        RECT 389.660 4384.050 389.940 4384.330 ;
        RECT 390.280 4384.050 390.560 4384.330 ;
        RECT 390.900 4384.050 391.180 4384.330 ;
        RECT 391.520 4384.050 391.800 4384.330 ;
        RECT 392.140 4384.050 392.420 4384.330 ;
        RECT 392.760 4384.050 393.040 4384.330 ;
        RECT 389.040 4383.430 389.320 4383.710 ;
        RECT 389.660 4383.430 389.940 4383.710 ;
        RECT 390.280 4383.430 390.560 4383.710 ;
        RECT 390.900 4383.430 391.180 4383.710 ;
        RECT 391.520 4383.430 391.800 4383.710 ;
        RECT 392.140 4383.430 392.420 4383.710 ;
        RECT 392.760 4383.430 393.040 4383.710 ;
        RECT 389.040 4382.810 389.320 4383.090 ;
        RECT 389.660 4382.810 389.940 4383.090 ;
        RECT 390.280 4382.810 390.560 4383.090 ;
        RECT 390.900 4382.810 391.180 4383.090 ;
        RECT 391.520 4382.810 391.800 4383.090 ;
        RECT 392.140 4382.810 392.420 4383.090 ;
        RECT 392.760 4382.810 393.040 4383.090 ;
        RECT 389.040 4382.190 389.320 4382.470 ;
        RECT 389.660 4382.190 389.940 4382.470 ;
        RECT 390.280 4382.190 390.560 4382.470 ;
        RECT 390.900 4382.190 391.180 4382.470 ;
        RECT 391.520 4382.190 391.800 4382.470 ;
        RECT 392.140 4382.190 392.420 4382.470 ;
        RECT 392.760 4382.190 393.040 4382.470 ;
        RECT 389.040 4381.570 389.320 4381.850 ;
        RECT 389.660 4381.570 389.940 4381.850 ;
        RECT 390.280 4381.570 390.560 4381.850 ;
        RECT 390.900 4381.570 391.180 4381.850 ;
        RECT 391.520 4381.570 391.800 4381.850 ;
        RECT 392.140 4381.570 392.420 4381.850 ;
        RECT 392.760 4381.570 393.040 4381.850 ;
        RECT 389.040 4380.950 389.320 4381.230 ;
        RECT 389.660 4380.950 389.940 4381.230 ;
        RECT 390.280 4380.950 390.560 4381.230 ;
        RECT 390.900 4380.950 391.180 4381.230 ;
        RECT 391.520 4380.950 391.800 4381.230 ;
        RECT 392.140 4380.950 392.420 4381.230 ;
        RECT 392.760 4380.950 393.040 4381.230 ;
        RECT 389.040 4380.330 389.320 4380.610 ;
        RECT 389.660 4380.330 389.940 4380.610 ;
        RECT 390.280 4380.330 390.560 4380.610 ;
        RECT 390.900 4380.330 391.180 4380.610 ;
        RECT 391.520 4380.330 391.800 4380.610 ;
        RECT 392.140 4380.330 392.420 4380.610 ;
        RECT 392.760 4380.330 393.040 4380.610 ;
        RECT 389.040 4379.710 389.320 4379.990 ;
        RECT 389.660 4379.710 389.940 4379.990 ;
        RECT 390.280 4379.710 390.560 4379.990 ;
        RECT 390.900 4379.710 391.180 4379.990 ;
        RECT 391.520 4379.710 391.800 4379.990 ;
        RECT 392.140 4379.710 392.420 4379.990 ;
        RECT 392.760 4379.710 393.040 4379.990 ;
        RECT 389.040 4379.090 389.320 4379.370 ;
        RECT 389.660 4379.090 389.940 4379.370 ;
        RECT 390.280 4379.090 390.560 4379.370 ;
        RECT 390.900 4379.090 391.180 4379.370 ;
        RECT 391.520 4379.090 391.800 4379.370 ;
        RECT 392.140 4379.090 392.420 4379.370 ;
        RECT 392.760 4379.090 393.040 4379.370 ;
        RECT 389.040 4378.470 389.320 4378.750 ;
        RECT 389.660 4378.470 389.940 4378.750 ;
        RECT 390.280 4378.470 390.560 4378.750 ;
        RECT 390.900 4378.470 391.180 4378.750 ;
        RECT 391.520 4378.470 391.800 4378.750 ;
        RECT 392.140 4378.470 392.420 4378.750 ;
        RECT 392.760 4378.470 393.040 4378.750 ;
        RECT 389.040 4377.850 389.320 4378.130 ;
        RECT 389.660 4377.850 389.940 4378.130 ;
        RECT 390.280 4377.850 390.560 4378.130 ;
        RECT 390.900 4377.850 391.180 4378.130 ;
        RECT 391.520 4377.850 391.800 4378.130 ;
        RECT 392.140 4377.850 392.420 4378.130 ;
        RECT 392.760 4377.850 393.040 4378.130 ;
        RECT 389.040 4377.230 389.320 4377.510 ;
        RECT 389.660 4377.230 389.940 4377.510 ;
        RECT 390.280 4377.230 390.560 4377.510 ;
        RECT 390.900 4377.230 391.180 4377.510 ;
        RECT 391.520 4377.230 391.800 4377.510 ;
        RECT 392.140 4377.230 392.420 4377.510 ;
        RECT 392.760 4377.230 393.040 4377.510 ;
        RECT 389.040 4376.610 389.320 4376.890 ;
        RECT 389.660 4376.610 389.940 4376.890 ;
        RECT 390.280 4376.610 390.560 4376.890 ;
        RECT 390.900 4376.610 391.180 4376.890 ;
        RECT 391.520 4376.610 391.800 4376.890 ;
        RECT 392.140 4376.610 392.420 4376.890 ;
        RECT 392.760 4376.610 393.040 4376.890 ;
        RECT 389.040 4375.990 389.320 4376.270 ;
        RECT 389.660 4375.990 389.940 4376.270 ;
        RECT 390.280 4375.990 390.560 4376.270 ;
        RECT 390.900 4375.990 391.180 4376.270 ;
        RECT 391.520 4375.990 391.800 4376.270 ;
        RECT 392.140 4375.990 392.420 4376.270 ;
        RECT 392.760 4375.990 393.040 4376.270 ;
        RECT 350.370 4373.410 350.650 4373.690 ;
        RECT 350.370 4372.790 350.650 4373.070 ;
        RECT 350.370 4372.170 350.650 4372.450 ;
        RECT 350.370 4371.550 350.650 4371.830 ;
        RECT 350.370 4370.930 350.650 4371.210 ;
        RECT 350.370 4370.310 350.650 4370.590 ;
        RECT 350.370 4369.690 350.650 4369.970 ;
        RECT 350.370 4369.070 350.650 4369.350 ;
        RECT 350.370 4368.450 350.650 4368.730 ;
        RECT 350.370 4367.830 350.650 4368.110 ;
        RECT 350.370 4367.210 350.650 4367.490 ;
        RECT 350.370 4366.590 350.650 4366.870 ;
        RECT 350.370 4365.970 350.650 4366.250 ;
        RECT 350.370 4365.350 350.650 4365.630 ;
        RECT 350.370 4364.730 350.650 4365.010 ;
        RECT 350.370 4364.110 350.650 4364.390 ;
        RECT 389.040 4373.440 389.320 4373.720 ;
        RECT 389.660 4373.440 389.940 4373.720 ;
        RECT 390.280 4373.440 390.560 4373.720 ;
        RECT 390.900 4373.440 391.180 4373.720 ;
        RECT 391.520 4373.440 391.800 4373.720 ;
        RECT 392.140 4373.440 392.420 4373.720 ;
        RECT 392.760 4373.440 393.040 4373.720 ;
        RECT 389.040 4372.820 389.320 4373.100 ;
        RECT 389.660 4372.820 389.940 4373.100 ;
        RECT 390.280 4372.820 390.560 4373.100 ;
        RECT 390.900 4372.820 391.180 4373.100 ;
        RECT 391.520 4372.820 391.800 4373.100 ;
        RECT 392.140 4372.820 392.420 4373.100 ;
        RECT 392.760 4372.820 393.040 4373.100 ;
        RECT 389.040 4372.200 389.320 4372.480 ;
        RECT 389.660 4372.200 389.940 4372.480 ;
        RECT 390.280 4372.200 390.560 4372.480 ;
        RECT 390.900 4372.200 391.180 4372.480 ;
        RECT 391.520 4372.200 391.800 4372.480 ;
        RECT 392.140 4372.200 392.420 4372.480 ;
        RECT 392.760 4372.200 393.040 4372.480 ;
        RECT 389.040 4371.580 389.320 4371.860 ;
        RECT 389.660 4371.580 389.940 4371.860 ;
        RECT 390.280 4371.580 390.560 4371.860 ;
        RECT 390.900 4371.580 391.180 4371.860 ;
        RECT 391.520 4371.580 391.800 4371.860 ;
        RECT 392.140 4371.580 392.420 4371.860 ;
        RECT 392.760 4371.580 393.040 4371.860 ;
        RECT 389.040 4370.960 389.320 4371.240 ;
        RECT 389.660 4370.960 389.940 4371.240 ;
        RECT 390.280 4370.960 390.560 4371.240 ;
        RECT 390.900 4370.960 391.180 4371.240 ;
        RECT 391.520 4370.960 391.800 4371.240 ;
        RECT 392.140 4370.960 392.420 4371.240 ;
        RECT 392.760 4370.960 393.040 4371.240 ;
        RECT 389.040 4370.340 389.320 4370.620 ;
        RECT 389.660 4370.340 389.940 4370.620 ;
        RECT 390.280 4370.340 390.560 4370.620 ;
        RECT 390.900 4370.340 391.180 4370.620 ;
        RECT 391.520 4370.340 391.800 4370.620 ;
        RECT 392.140 4370.340 392.420 4370.620 ;
        RECT 392.760 4370.340 393.040 4370.620 ;
        RECT 389.040 4369.720 389.320 4370.000 ;
        RECT 389.660 4369.720 389.940 4370.000 ;
        RECT 390.280 4369.720 390.560 4370.000 ;
        RECT 390.900 4369.720 391.180 4370.000 ;
        RECT 391.520 4369.720 391.800 4370.000 ;
        RECT 392.140 4369.720 392.420 4370.000 ;
        RECT 392.760 4369.720 393.040 4370.000 ;
        RECT 389.040 4369.100 389.320 4369.380 ;
        RECT 389.660 4369.100 389.940 4369.380 ;
        RECT 390.280 4369.100 390.560 4369.380 ;
        RECT 390.900 4369.100 391.180 4369.380 ;
        RECT 391.520 4369.100 391.800 4369.380 ;
        RECT 392.140 4369.100 392.420 4369.380 ;
        RECT 392.760 4369.100 393.040 4369.380 ;
        RECT 389.040 4368.480 389.320 4368.760 ;
        RECT 389.660 4368.480 389.940 4368.760 ;
        RECT 390.280 4368.480 390.560 4368.760 ;
        RECT 390.900 4368.480 391.180 4368.760 ;
        RECT 391.520 4368.480 391.800 4368.760 ;
        RECT 392.140 4368.480 392.420 4368.760 ;
        RECT 392.760 4368.480 393.040 4368.760 ;
        RECT 389.040 4367.860 389.320 4368.140 ;
        RECT 389.660 4367.860 389.940 4368.140 ;
        RECT 390.280 4367.860 390.560 4368.140 ;
        RECT 390.900 4367.860 391.180 4368.140 ;
        RECT 391.520 4367.860 391.800 4368.140 ;
        RECT 392.140 4367.860 392.420 4368.140 ;
        RECT 392.760 4367.860 393.040 4368.140 ;
        RECT 389.040 4367.240 389.320 4367.520 ;
        RECT 389.660 4367.240 389.940 4367.520 ;
        RECT 390.280 4367.240 390.560 4367.520 ;
        RECT 390.900 4367.240 391.180 4367.520 ;
        RECT 391.520 4367.240 391.800 4367.520 ;
        RECT 392.140 4367.240 392.420 4367.520 ;
        RECT 392.760 4367.240 393.040 4367.520 ;
        RECT 389.040 4366.620 389.320 4366.900 ;
        RECT 389.660 4366.620 389.940 4366.900 ;
        RECT 390.280 4366.620 390.560 4366.900 ;
        RECT 390.900 4366.620 391.180 4366.900 ;
        RECT 391.520 4366.620 391.800 4366.900 ;
        RECT 392.140 4366.620 392.420 4366.900 ;
        RECT 392.760 4366.620 393.040 4366.900 ;
        RECT 389.040 4366.000 389.320 4366.280 ;
        RECT 389.660 4366.000 389.940 4366.280 ;
        RECT 390.280 4366.000 390.560 4366.280 ;
        RECT 390.900 4366.000 391.180 4366.280 ;
        RECT 391.520 4366.000 391.800 4366.280 ;
        RECT 392.140 4366.000 392.420 4366.280 ;
        RECT 392.760 4366.000 393.040 4366.280 ;
        RECT 389.040 4365.380 389.320 4365.660 ;
        RECT 389.660 4365.380 389.940 4365.660 ;
        RECT 390.280 4365.380 390.560 4365.660 ;
        RECT 390.900 4365.380 391.180 4365.660 ;
        RECT 391.520 4365.380 391.800 4365.660 ;
        RECT 392.140 4365.380 392.420 4365.660 ;
        RECT 392.760 4365.380 393.040 4365.660 ;
        RECT 389.040 4364.760 389.320 4365.040 ;
        RECT 389.660 4364.760 389.940 4365.040 ;
        RECT 390.280 4364.760 390.560 4365.040 ;
        RECT 390.900 4364.760 391.180 4365.040 ;
        RECT 391.520 4364.760 391.800 4365.040 ;
        RECT 392.140 4364.760 392.420 4365.040 ;
        RECT 392.760 4364.760 393.040 4365.040 ;
        RECT 389.040 4364.140 389.320 4364.420 ;
        RECT 389.660 4364.140 389.940 4364.420 ;
        RECT 390.280 4364.140 390.560 4364.420 ;
        RECT 390.900 4364.140 391.180 4364.420 ;
        RECT 391.520 4364.140 391.800 4364.420 ;
        RECT 392.140 4364.140 392.420 4364.420 ;
        RECT 392.760 4364.140 393.040 4364.420 ;
        RECT 350.370 4360.390 350.650 4360.670 ;
        RECT 350.370 4359.770 350.650 4360.050 ;
        RECT 350.370 4359.150 350.650 4359.430 ;
        RECT 350.370 4358.530 350.650 4358.810 ;
        RECT 350.370 4357.910 350.650 4358.190 ;
        RECT 350.370 4357.290 350.650 4357.570 ;
        RECT 350.370 4356.670 350.650 4356.950 ;
        RECT 350.370 4356.050 350.650 4356.330 ;
        RECT 350.370 4355.430 350.650 4355.710 ;
        RECT 350.370 4354.810 350.650 4355.090 ;
        RECT 350.370 4354.190 350.650 4354.470 ;
        RECT 350.370 4353.570 350.650 4353.850 ;
        RECT 350.370 4352.950 350.650 4353.230 ;
        RECT 350.370 4352.330 350.650 4352.610 ;
        RECT 350.370 4351.710 350.650 4351.990 ;
        RECT 389.040 4360.420 389.320 4360.700 ;
        RECT 389.660 4360.420 389.940 4360.700 ;
        RECT 390.280 4360.420 390.560 4360.700 ;
        RECT 390.900 4360.420 391.180 4360.700 ;
        RECT 391.520 4360.420 391.800 4360.700 ;
        RECT 392.140 4360.420 392.420 4360.700 ;
        RECT 392.760 4360.420 393.040 4360.700 ;
        RECT 389.040 4359.800 389.320 4360.080 ;
        RECT 389.660 4359.800 389.940 4360.080 ;
        RECT 390.280 4359.800 390.560 4360.080 ;
        RECT 390.900 4359.800 391.180 4360.080 ;
        RECT 391.520 4359.800 391.800 4360.080 ;
        RECT 392.140 4359.800 392.420 4360.080 ;
        RECT 392.760 4359.800 393.040 4360.080 ;
        RECT 389.040 4359.180 389.320 4359.460 ;
        RECT 389.660 4359.180 389.940 4359.460 ;
        RECT 390.280 4359.180 390.560 4359.460 ;
        RECT 390.900 4359.180 391.180 4359.460 ;
        RECT 391.520 4359.180 391.800 4359.460 ;
        RECT 392.140 4359.180 392.420 4359.460 ;
        RECT 392.760 4359.180 393.040 4359.460 ;
        RECT 389.040 4358.560 389.320 4358.840 ;
        RECT 389.660 4358.560 389.940 4358.840 ;
        RECT 390.280 4358.560 390.560 4358.840 ;
        RECT 390.900 4358.560 391.180 4358.840 ;
        RECT 391.520 4358.560 391.800 4358.840 ;
        RECT 392.140 4358.560 392.420 4358.840 ;
        RECT 392.760 4358.560 393.040 4358.840 ;
        RECT 389.040 4357.940 389.320 4358.220 ;
        RECT 389.660 4357.940 389.940 4358.220 ;
        RECT 390.280 4357.940 390.560 4358.220 ;
        RECT 390.900 4357.940 391.180 4358.220 ;
        RECT 391.520 4357.940 391.800 4358.220 ;
        RECT 392.140 4357.940 392.420 4358.220 ;
        RECT 392.760 4357.940 393.040 4358.220 ;
        RECT 389.040 4357.320 389.320 4357.600 ;
        RECT 389.660 4357.320 389.940 4357.600 ;
        RECT 390.280 4357.320 390.560 4357.600 ;
        RECT 390.900 4357.320 391.180 4357.600 ;
        RECT 391.520 4357.320 391.800 4357.600 ;
        RECT 392.140 4357.320 392.420 4357.600 ;
        RECT 392.760 4357.320 393.040 4357.600 ;
        RECT 389.040 4356.700 389.320 4356.980 ;
        RECT 389.660 4356.700 389.940 4356.980 ;
        RECT 390.280 4356.700 390.560 4356.980 ;
        RECT 390.900 4356.700 391.180 4356.980 ;
        RECT 391.520 4356.700 391.800 4356.980 ;
        RECT 392.140 4356.700 392.420 4356.980 ;
        RECT 392.760 4356.700 393.040 4356.980 ;
        RECT 389.040 4356.080 389.320 4356.360 ;
        RECT 389.660 4356.080 389.940 4356.360 ;
        RECT 390.280 4356.080 390.560 4356.360 ;
        RECT 390.900 4356.080 391.180 4356.360 ;
        RECT 391.520 4356.080 391.800 4356.360 ;
        RECT 392.140 4356.080 392.420 4356.360 ;
        RECT 392.760 4356.080 393.040 4356.360 ;
        RECT 389.040 4355.460 389.320 4355.740 ;
        RECT 389.660 4355.460 389.940 4355.740 ;
        RECT 390.280 4355.460 390.560 4355.740 ;
        RECT 390.900 4355.460 391.180 4355.740 ;
        RECT 391.520 4355.460 391.800 4355.740 ;
        RECT 392.140 4355.460 392.420 4355.740 ;
        RECT 392.760 4355.460 393.040 4355.740 ;
        RECT 389.040 4354.840 389.320 4355.120 ;
        RECT 389.660 4354.840 389.940 4355.120 ;
        RECT 390.280 4354.840 390.560 4355.120 ;
        RECT 390.900 4354.840 391.180 4355.120 ;
        RECT 391.520 4354.840 391.800 4355.120 ;
        RECT 392.140 4354.840 392.420 4355.120 ;
        RECT 392.760 4354.840 393.040 4355.120 ;
        RECT 389.040 4354.220 389.320 4354.500 ;
        RECT 389.660 4354.220 389.940 4354.500 ;
        RECT 390.280 4354.220 390.560 4354.500 ;
        RECT 390.900 4354.220 391.180 4354.500 ;
        RECT 391.520 4354.220 391.800 4354.500 ;
        RECT 392.140 4354.220 392.420 4354.500 ;
        RECT 392.760 4354.220 393.040 4354.500 ;
        RECT 389.040 4353.600 389.320 4353.880 ;
        RECT 389.660 4353.600 389.940 4353.880 ;
        RECT 390.280 4353.600 390.560 4353.880 ;
        RECT 390.900 4353.600 391.180 4353.880 ;
        RECT 391.520 4353.600 391.800 4353.880 ;
        RECT 392.140 4353.600 392.420 4353.880 ;
        RECT 392.760 4353.600 393.040 4353.880 ;
        RECT 389.040 4352.980 389.320 4353.260 ;
        RECT 389.660 4352.980 389.940 4353.260 ;
        RECT 390.280 4352.980 390.560 4353.260 ;
        RECT 390.900 4352.980 391.180 4353.260 ;
        RECT 391.520 4352.980 391.800 4353.260 ;
        RECT 392.140 4352.980 392.420 4353.260 ;
        RECT 392.760 4352.980 393.040 4353.260 ;
        RECT 389.040 4352.360 389.320 4352.640 ;
        RECT 389.660 4352.360 389.940 4352.640 ;
        RECT 390.280 4352.360 390.560 4352.640 ;
        RECT 390.900 4352.360 391.180 4352.640 ;
        RECT 391.520 4352.360 391.800 4352.640 ;
        RECT 392.140 4352.360 392.420 4352.640 ;
        RECT 392.760 4352.360 393.040 4352.640 ;
        RECT 389.040 4351.740 389.320 4352.020 ;
        RECT 389.660 4351.740 389.940 4352.020 ;
        RECT 390.280 4351.740 390.560 4352.020 ;
        RECT 390.900 4351.740 391.180 4352.020 ;
        RECT 391.520 4351.740 391.800 4352.020 ;
        RECT 392.140 4351.740 392.420 4352.020 ;
        RECT 392.760 4351.740 393.040 4352.020 ;
        RECT 350.370 4218.010 350.650 4218.290 ;
        RECT 350.370 4217.390 350.650 4217.670 ;
        RECT 350.370 4216.770 350.650 4217.050 ;
        RECT 350.370 4216.150 350.650 4216.430 ;
        RECT 350.370 4215.530 350.650 4215.810 ;
        RECT 350.370 4214.910 350.650 4215.190 ;
        RECT 350.370 4214.290 350.650 4214.570 ;
        RECT 350.370 4213.670 350.650 4213.950 ;
        RECT 350.370 4213.050 350.650 4213.330 ;
        RECT 350.370 4212.430 350.650 4212.710 ;
        RECT 350.370 4211.810 350.650 4212.090 ;
        RECT 350.370 4211.190 350.650 4211.470 ;
        RECT 350.370 4210.570 350.650 4210.850 ;
        RECT 350.370 4209.950 350.650 4210.230 ;
        RECT 350.370 4209.330 350.650 4209.610 ;
        RECT 389.040 4218.070 389.320 4218.350 ;
        RECT 389.660 4218.070 389.940 4218.350 ;
        RECT 390.280 4218.070 390.560 4218.350 ;
        RECT 390.900 4218.070 391.180 4218.350 ;
        RECT 391.520 4218.070 391.800 4218.350 ;
        RECT 392.140 4218.070 392.420 4218.350 ;
        RECT 392.760 4218.070 393.040 4218.350 ;
        RECT 389.040 4217.450 389.320 4217.730 ;
        RECT 389.660 4217.450 389.940 4217.730 ;
        RECT 390.280 4217.450 390.560 4217.730 ;
        RECT 390.900 4217.450 391.180 4217.730 ;
        RECT 391.520 4217.450 391.800 4217.730 ;
        RECT 392.140 4217.450 392.420 4217.730 ;
        RECT 392.760 4217.450 393.040 4217.730 ;
        RECT 389.040 4216.830 389.320 4217.110 ;
        RECT 389.660 4216.830 389.940 4217.110 ;
        RECT 390.280 4216.830 390.560 4217.110 ;
        RECT 390.900 4216.830 391.180 4217.110 ;
        RECT 391.520 4216.830 391.800 4217.110 ;
        RECT 392.140 4216.830 392.420 4217.110 ;
        RECT 392.760 4216.830 393.040 4217.110 ;
        RECT 389.040 4216.210 389.320 4216.490 ;
        RECT 389.660 4216.210 389.940 4216.490 ;
        RECT 390.280 4216.210 390.560 4216.490 ;
        RECT 390.900 4216.210 391.180 4216.490 ;
        RECT 391.520 4216.210 391.800 4216.490 ;
        RECT 392.140 4216.210 392.420 4216.490 ;
        RECT 392.760 4216.210 393.040 4216.490 ;
        RECT 389.040 4215.590 389.320 4215.870 ;
        RECT 389.660 4215.590 389.940 4215.870 ;
        RECT 390.280 4215.590 390.560 4215.870 ;
        RECT 390.900 4215.590 391.180 4215.870 ;
        RECT 391.520 4215.590 391.800 4215.870 ;
        RECT 392.140 4215.590 392.420 4215.870 ;
        RECT 392.760 4215.590 393.040 4215.870 ;
        RECT 389.040 4214.970 389.320 4215.250 ;
        RECT 389.660 4214.970 389.940 4215.250 ;
        RECT 390.280 4214.970 390.560 4215.250 ;
        RECT 390.900 4214.970 391.180 4215.250 ;
        RECT 391.520 4214.970 391.800 4215.250 ;
        RECT 392.140 4214.970 392.420 4215.250 ;
        RECT 392.760 4214.970 393.040 4215.250 ;
        RECT 389.040 4214.350 389.320 4214.630 ;
        RECT 389.660 4214.350 389.940 4214.630 ;
        RECT 390.280 4214.350 390.560 4214.630 ;
        RECT 390.900 4214.350 391.180 4214.630 ;
        RECT 391.520 4214.350 391.800 4214.630 ;
        RECT 392.140 4214.350 392.420 4214.630 ;
        RECT 392.760 4214.350 393.040 4214.630 ;
        RECT 389.040 4213.730 389.320 4214.010 ;
        RECT 389.660 4213.730 389.940 4214.010 ;
        RECT 390.280 4213.730 390.560 4214.010 ;
        RECT 390.900 4213.730 391.180 4214.010 ;
        RECT 391.520 4213.730 391.800 4214.010 ;
        RECT 392.140 4213.730 392.420 4214.010 ;
        RECT 392.760 4213.730 393.040 4214.010 ;
        RECT 389.040 4213.110 389.320 4213.390 ;
        RECT 389.660 4213.110 389.940 4213.390 ;
        RECT 390.280 4213.110 390.560 4213.390 ;
        RECT 390.900 4213.110 391.180 4213.390 ;
        RECT 391.520 4213.110 391.800 4213.390 ;
        RECT 392.140 4213.110 392.420 4213.390 ;
        RECT 392.760 4213.110 393.040 4213.390 ;
        RECT 389.040 4212.490 389.320 4212.770 ;
        RECT 389.660 4212.490 389.940 4212.770 ;
        RECT 390.280 4212.490 390.560 4212.770 ;
        RECT 390.900 4212.490 391.180 4212.770 ;
        RECT 391.520 4212.490 391.800 4212.770 ;
        RECT 392.140 4212.490 392.420 4212.770 ;
        RECT 392.760 4212.490 393.040 4212.770 ;
        RECT 389.040 4211.870 389.320 4212.150 ;
        RECT 389.660 4211.870 389.940 4212.150 ;
        RECT 390.280 4211.870 390.560 4212.150 ;
        RECT 390.900 4211.870 391.180 4212.150 ;
        RECT 391.520 4211.870 391.800 4212.150 ;
        RECT 392.140 4211.870 392.420 4212.150 ;
        RECT 392.760 4211.870 393.040 4212.150 ;
        RECT 389.040 4211.250 389.320 4211.530 ;
        RECT 389.660 4211.250 389.940 4211.530 ;
        RECT 390.280 4211.250 390.560 4211.530 ;
        RECT 390.900 4211.250 391.180 4211.530 ;
        RECT 391.520 4211.250 391.800 4211.530 ;
        RECT 392.140 4211.250 392.420 4211.530 ;
        RECT 392.760 4211.250 393.040 4211.530 ;
        RECT 389.040 4210.630 389.320 4210.910 ;
        RECT 389.660 4210.630 389.940 4210.910 ;
        RECT 390.280 4210.630 390.560 4210.910 ;
        RECT 390.900 4210.630 391.180 4210.910 ;
        RECT 391.520 4210.630 391.800 4210.910 ;
        RECT 392.140 4210.630 392.420 4210.910 ;
        RECT 392.760 4210.630 393.040 4210.910 ;
        RECT 389.040 4210.010 389.320 4210.290 ;
        RECT 389.660 4210.010 389.940 4210.290 ;
        RECT 390.280 4210.010 390.560 4210.290 ;
        RECT 390.900 4210.010 391.180 4210.290 ;
        RECT 391.520 4210.010 391.800 4210.290 ;
        RECT 392.140 4210.010 392.420 4210.290 ;
        RECT 392.760 4210.010 393.040 4210.290 ;
        RECT 389.040 4209.390 389.320 4209.670 ;
        RECT 389.660 4209.390 389.940 4209.670 ;
        RECT 390.280 4209.390 390.560 4209.670 ;
        RECT 390.900 4209.390 391.180 4209.670 ;
        RECT 391.520 4209.390 391.800 4209.670 ;
        RECT 392.140 4209.390 392.420 4209.670 ;
        RECT 392.760 4209.390 393.040 4209.670 ;
        RECT 350.370 4205.640 350.650 4205.920 ;
        RECT 350.370 4205.020 350.650 4205.300 ;
        RECT 350.370 4204.400 350.650 4204.680 ;
        RECT 350.370 4203.780 350.650 4204.060 ;
        RECT 350.370 4203.160 350.650 4203.440 ;
        RECT 350.370 4202.540 350.650 4202.820 ;
        RECT 350.370 4201.920 350.650 4202.200 ;
        RECT 350.370 4201.300 350.650 4201.580 ;
        RECT 350.370 4200.680 350.650 4200.960 ;
        RECT 350.370 4200.060 350.650 4200.340 ;
        RECT 350.370 4199.440 350.650 4199.720 ;
        RECT 350.370 4198.820 350.650 4199.100 ;
        RECT 350.370 4198.200 350.650 4198.480 ;
        RECT 350.370 4197.580 350.650 4197.860 ;
        RECT 350.370 4196.960 350.650 4197.240 ;
        RECT 350.370 4196.340 350.650 4196.620 ;
        RECT 389.040 4205.670 389.320 4205.950 ;
        RECT 389.660 4205.670 389.940 4205.950 ;
        RECT 390.280 4205.670 390.560 4205.950 ;
        RECT 390.900 4205.670 391.180 4205.950 ;
        RECT 391.520 4205.670 391.800 4205.950 ;
        RECT 392.140 4205.670 392.420 4205.950 ;
        RECT 392.760 4205.670 393.040 4205.950 ;
        RECT 389.040 4205.050 389.320 4205.330 ;
        RECT 389.660 4205.050 389.940 4205.330 ;
        RECT 390.280 4205.050 390.560 4205.330 ;
        RECT 390.900 4205.050 391.180 4205.330 ;
        RECT 391.520 4205.050 391.800 4205.330 ;
        RECT 392.140 4205.050 392.420 4205.330 ;
        RECT 392.760 4205.050 393.040 4205.330 ;
        RECT 389.040 4204.430 389.320 4204.710 ;
        RECT 389.660 4204.430 389.940 4204.710 ;
        RECT 390.280 4204.430 390.560 4204.710 ;
        RECT 390.900 4204.430 391.180 4204.710 ;
        RECT 391.520 4204.430 391.800 4204.710 ;
        RECT 392.140 4204.430 392.420 4204.710 ;
        RECT 392.760 4204.430 393.040 4204.710 ;
        RECT 389.040 4203.810 389.320 4204.090 ;
        RECT 389.660 4203.810 389.940 4204.090 ;
        RECT 390.280 4203.810 390.560 4204.090 ;
        RECT 390.900 4203.810 391.180 4204.090 ;
        RECT 391.520 4203.810 391.800 4204.090 ;
        RECT 392.140 4203.810 392.420 4204.090 ;
        RECT 392.760 4203.810 393.040 4204.090 ;
        RECT 389.040 4203.190 389.320 4203.470 ;
        RECT 389.660 4203.190 389.940 4203.470 ;
        RECT 390.280 4203.190 390.560 4203.470 ;
        RECT 390.900 4203.190 391.180 4203.470 ;
        RECT 391.520 4203.190 391.800 4203.470 ;
        RECT 392.140 4203.190 392.420 4203.470 ;
        RECT 392.760 4203.190 393.040 4203.470 ;
        RECT 389.040 4202.570 389.320 4202.850 ;
        RECT 389.660 4202.570 389.940 4202.850 ;
        RECT 390.280 4202.570 390.560 4202.850 ;
        RECT 390.900 4202.570 391.180 4202.850 ;
        RECT 391.520 4202.570 391.800 4202.850 ;
        RECT 392.140 4202.570 392.420 4202.850 ;
        RECT 392.760 4202.570 393.040 4202.850 ;
        RECT 389.040 4201.950 389.320 4202.230 ;
        RECT 389.660 4201.950 389.940 4202.230 ;
        RECT 390.280 4201.950 390.560 4202.230 ;
        RECT 390.900 4201.950 391.180 4202.230 ;
        RECT 391.520 4201.950 391.800 4202.230 ;
        RECT 392.140 4201.950 392.420 4202.230 ;
        RECT 392.760 4201.950 393.040 4202.230 ;
        RECT 389.040 4201.330 389.320 4201.610 ;
        RECT 389.660 4201.330 389.940 4201.610 ;
        RECT 390.280 4201.330 390.560 4201.610 ;
        RECT 390.900 4201.330 391.180 4201.610 ;
        RECT 391.520 4201.330 391.800 4201.610 ;
        RECT 392.140 4201.330 392.420 4201.610 ;
        RECT 392.760 4201.330 393.040 4201.610 ;
        RECT 389.040 4200.710 389.320 4200.990 ;
        RECT 389.660 4200.710 389.940 4200.990 ;
        RECT 390.280 4200.710 390.560 4200.990 ;
        RECT 390.900 4200.710 391.180 4200.990 ;
        RECT 391.520 4200.710 391.800 4200.990 ;
        RECT 392.140 4200.710 392.420 4200.990 ;
        RECT 392.760 4200.710 393.040 4200.990 ;
        RECT 389.040 4200.090 389.320 4200.370 ;
        RECT 389.660 4200.090 389.940 4200.370 ;
        RECT 390.280 4200.090 390.560 4200.370 ;
        RECT 390.900 4200.090 391.180 4200.370 ;
        RECT 391.520 4200.090 391.800 4200.370 ;
        RECT 392.140 4200.090 392.420 4200.370 ;
        RECT 392.760 4200.090 393.040 4200.370 ;
        RECT 389.040 4199.470 389.320 4199.750 ;
        RECT 389.660 4199.470 389.940 4199.750 ;
        RECT 390.280 4199.470 390.560 4199.750 ;
        RECT 390.900 4199.470 391.180 4199.750 ;
        RECT 391.520 4199.470 391.800 4199.750 ;
        RECT 392.140 4199.470 392.420 4199.750 ;
        RECT 392.760 4199.470 393.040 4199.750 ;
        RECT 389.040 4198.850 389.320 4199.130 ;
        RECT 389.660 4198.850 389.940 4199.130 ;
        RECT 390.280 4198.850 390.560 4199.130 ;
        RECT 390.900 4198.850 391.180 4199.130 ;
        RECT 391.520 4198.850 391.800 4199.130 ;
        RECT 392.140 4198.850 392.420 4199.130 ;
        RECT 392.760 4198.850 393.040 4199.130 ;
        RECT 389.040 4198.230 389.320 4198.510 ;
        RECT 389.660 4198.230 389.940 4198.510 ;
        RECT 390.280 4198.230 390.560 4198.510 ;
        RECT 390.900 4198.230 391.180 4198.510 ;
        RECT 391.520 4198.230 391.800 4198.510 ;
        RECT 392.140 4198.230 392.420 4198.510 ;
        RECT 392.760 4198.230 393.040 4198.510 ;
        RECT 389.040 4197.610 389.320 4197.890 ;
        RECT 389.660 4197.610 389.940 4197.890 ;
        RECT 390.280 4197.610 390.560 4197.890 ;
        RECT 390.900 4197.610 391.180 4197.890 ;
        RECT 391.520 4197.610 391.800 4197.890 ;
        RECT 392.140 4197.610 392.420 4197.890 ;
        RECT 392.760 4197.610 393.040 4197.890 ;
        RECT 389.040 4196.990 389.320 4197.270 ;
        RECT 389.660 4196.990 389.940 4197.270 ;
        RECT 390.280 4196.990 390.560 4197.270 ;
        RECT 390.900 4196.990 391.180 4197.270 ;
        RECT 391.520 4196.990 391.800 4197.270 ;
        RECT 392.140 4196.990 392.420 4197.270 ;
        RECT 392.760 4196.990 393.040 4197.270 ;
        RECT 389.040 4196.370 389.320 4196.650 ;
        RECT 389.660 4196.370 389.940 4196.650 ;
        RECT 390.280 4196.370 390.560 4196.650 ;
        RECT 390.900 4196.370 391.180 4196.650 ;
        RECT 391.520 4196.370 391.800 4196.650 ;
        RECT 392.140 4196.370 392.420 4196.650 ;
        RECT 392.760 4196.370 393.040 4196.650 ;
        RECT 350.370 4193.790 350.650 4194.070 ;
        RECT 350.370 4193.170 350.650 4193.450 ;
        RECT 350.370 4192.550 350.650 4192.830 ;
        RECT 350.370 4191.930 350.650 4192.210 ;
        RECT 350.370 4191.310 350.650 4191.590 ;
        RECT 350.370 4190.690 350.650 4190.970 ;
        RECT 350.370 4190.070 350.650 4190.350 ;
        RECT 350.370 4189.450 350.650 4189.730 ;
        RECT 350.370 4188.830 350.650 4189.110 ;
        RECT 350.370 4188.210 350.650 4188.490 ;
        RECT 350.370 4187.590 350.650 4187.870 ;
        RECT 350.370 4186.970 350.650 4187.250 ;
        RECT 350.370 4186.350 350.650 4186.630 ;
        RECT 350.370 4185.730 350.650 4186.010 ;
        RECT 350.370 4185.110 350.650 4185.390 ;
        RECT 350.370 4184.490 350.650 4184.770 ;
        RECT 389.040 4193.820 389.320 4194.100 ;
        RECT 389.660 4193.820 389.940 4194.100 ;
        RECT 390.280 4193.820 390.560 4194.100 ;
        RECT 390.900 4193.820 391.180 4194.100 ;
        RECT 391.520 4193.820 391.800 4194.100 ;
        RECT 392.140 4193.820 392.420 4194.100 ;
        RECT 392.760 4193.820 393.040 4194.100 ;
        RECT 389.040 4193.200 389.320 4193.480 ;
        RECT 389.660 4193.200 389.940 4193.480 ;
        RECT 390.280 4193.200 390.560 4193.480 ;
        RECT 390.900 4193.200 391.180 4193.480 ;
        RECT 391.520 4193.200 391.800 4193.480 ;
        RECT 392.140 4193.200 392.420 4193.480 ;
        RECT 392.760 4193.200 393.040 4193.480 ;
        RECT 389.040 4192.580 389.320 4192.860 ;
        RECT 389.660 4192.580 389.940 4192.860 ;
        RECT 390.280 4192.580 390.560 4192.860 ;
        RECT 390.900 4192.580 391.180 4192.860 ;
        RECT 391.520 4192.580 391.800 4192.860 ;
        RECT 392.140 4192.580 392.420 4192.860 ;
        RECT 392.760 4192.580 393.040 4192.860 ;
        RECT 389.040 4191.960 389.320 4192.240 ;
        RECT 389.660 4191.960 389.940 4192.240 ;
        RECT 390.280 4191.960 390.560 4192.240 ;
        RECT 390.900 4191.960 391.180 4192.240 ;
        RECT 391.520 4191.960 391.800 4192.240 ;
        RECT 392.140 4191.960 392.420 4192.240 ;
        RECT 392.760 4191.960 393.040 4192.240 ;
        RECT 389.040 4191.340 389.320 4191.620 ;
        RECT 389.660 4191.340 389.940 4191.620 ;
        RECT 390.280 4191.340 390.560 4191.620 ;
        RECT 390.900 4191.340 391.180 4191.620 ;
        RECT 391.520 4191.340 391.800 4191.620 ;
        RECT 392.140 4191.340 392.420 4191.620 ;
        RECT 392.760 4191.340 393.040 4191.620 ;
        RECT 389.040 4190.720 389.320 4191.000 ;
        RECT 389.660 4190.720 389.940 4191.000 ;
        RECT 390.280 4190.720 390.560 4191.000 ;
        RECT 390.900 4190.720 391.180 4191.000 ;
        RECT 391.520 4190.720 391.800 4191.000 ;
        RECT 392.140 4190.720 392.420 4191.000 ;
        RECT 392.760 4190.720 393.040 4191.000 ;
        RECT 389.040 4190.100 389.320 4190.380 ;
        RECT 389.660 4190.100 389.940 4190.380 ;
        RECT 390.280 4190.100 390.560 4190.380 ;
        RECT 390.900 4190.100 391.180 4190.380 ;
        RECT 391.520 4190.100 391.800 4190.380 ;
        RECT 392.140 4190.100 392.420 4190.380 ;
        RECT 392.760 4190.100 393.040 4190.380 ;
        RECT 389.040 4189.480 389.320 4189.760 ;
        RECT 389.660 4189.480 389.940 4189.760 ;
        RECT 390.280 4189.480 390.560 4189.760 ;
        RECT 390.900 4189.480 391.180 4189.760 ;
        RECT 391.520 4189.480 391.800 4189.760 ;
        RECT 392.140 4189.480 392.420 4189.760 ;
        RECT 392.760 4189.480 393.040 4189.760 ;
        RECT 389.040 4188.860 389.320 4189.140 ;
        RECT 389.660 4188.860 389.940 4189.140 ;
        RECT 390.280 4188.860 390.560 4189.140 ;
        RECT 390.900 4188.860 391.180 4189.140 ;
        RECT 391.520 4188.860 391.800 4189.140 ;
        RECT 392.140 4188.860 392.420 4189.140 ;
        RECT 392.760 4188.860 393.040 4189.140 ;
        RECT 389.040 4188.240 389.320 4188.520 ;
        RECT 389.660 4188.240 389.940 4188.520 ;
        RECT 390.280 4188.240 390.560 4188.520 ;
        RECT 390.900 4188.240 391.180 4188.520 ;
        RECT 391.520 4188.240 391.800 4188.520 ;
        RECT 392.140 4188.240 392.420 4188.520 ;
        RECT 392.760 4188.240 393.040 4188.520 ;
        RECT 389.040 4187.620 389.320 4187.900 ;
        RECT 389.660 4187.620 389.940 4187.900 ;
        RECT 390.280 4187.620 390.560 4187.900 ;
        RECT 390.900 4187.620 391.180 4187.900 ;
        RECT 391.520 4187.620 391.800 4187.900 ;
        RECT 392.140 4187.620 392.420 4187.900 ;
        RECT 392.760 4187.620 393.040 4187.900 ;
        RECT 389.040 4187.000 389.320 4187.280 ;
        RECT 389.660 4187.000 389.940 4187.280 ;
        RECT 390.280 4187.000 390.560 4187.280 ;
        RECT 390.900 4187.000 391.180 4187.280 ;
        RECT 391.520 4187.000 391.800 4187.280 ;
        RECT 392.140 4187.000 392.420 4187.280 ;
        RECT 392.760 4187.000 393.040 4187.280 ;
        RECT 389.040 4186.380 389.320 4186.660 ;
        RECT 389.660 4186.380 389.940 4186.660 ;
        RECT 390.280 4186.380 390.560 4186.660 ;
        RECT 390.900 4186.380 391.180 4186.660 ;
        RECT 391.520 4186.380 391.800 4186.660 ;
        RECT 392.140 4186.380 392.420 4186.660 ;
        RECT 392.760 4186.380 393.040 4186.660 ;
        RECT 389.040 4185.760 389.320 4186.040 ;
        RECT 389.660 4185.760 389.940 4186.040 ;
        RECT 390.280 4185.760 390.560 4186.040 ;
        RECT 390.900 4185.760 391.180 4186.040 ;
        RECT 391.520 4185.760 391.800 4186.040 ;
        RECT 392.140 4185.760 392.420 4186.040 ;
        RECT 392.760 4185.760 393.040 4186.040 ;
        RECT 389.040 4185.140 389.320 4185.420 ;
        RECT 389.660 4185.140 389.940 4185.420 ;
        RECT 390.280 4185.140 390.560 4185.420 ;
        RECT 390.900 4185.140 391.180 4185.420 ;
        RECT 391.520 4185.140 391.800 4185.420 ;
        RECT 392.140 4185.140 392.420 4185.420 ;
        RECT 392.760 4185.140 393.040 4185.420 ;
        RECT 389.040 4184.520 389.320 4184.800 ;
        RECT 389.660 4184.520 389.940 4184.800 ;
        RECT 390.280 4184.520 390.560 4184.800 ;
        RECT 390.900 4184.520 391.180 4184.800 ;
        RECT 391.520 4184.520 391.800 4184.800 ;
        RECT 392.140 4184.520 392.420 4184.800 ;
        RECT 392.760 4184.520 393.040 4184.800 ;
        RECT 350.370 4180.260 350.650 4180.540 ;
        RECT 350.370 4179.640 350.650 4179.920 ;
        RECT 350.370 4179.020 350.650 4179.300 ;
        RECT 350.370 4178.400 350.650 4178.680 ;
        RECT 350.370 4177.780 350.650 4178.060 ;
        RECT 350.370 4177.160 350.650 4177.440 ;
        RECT 350.370 4176.540 350.650 4176.820 ;
        RECT 350.370 4175.920 350.650 4176.200 ;
        RECT 350.370 4175.300 350.650 4175.580 ;
        RECT 350.370 4174.680 350.650 4174.960 ;
        RECT 350.370 4174.060 350.650 4174.340 ;
        RECT 350.370 4173.440 350.650 4173.720 ;
        RECT 350.370 4172.820 350.650 4173.100 ;
        RECT 350.370 4172.200 350.650 4172.480 ;
        RECT 350.370 4171.580 350.650 4171.860 ;
        RECT 350.370 4170.960 350.650 4171.240 ;
        RECT 389.040 4180.290 389.320 4180.570 ;
        RECT 389.660 4180.290 389.940 4180.570 ;
        RECT 390.280 4180.290 390.560 4180.570 ;
        RECT 390.900 4180.290 391.180 4180.570 ;
        RECT 391.520 4180.290 391.800 4180.570 ;
        RECT 392.140 4180.290 392.420 4180.570 ;
        RECT 392.760 4180.290 393.040 4180.570 ;
        RECT 389.040 4179.670 389.320 4179.950 ;
        RECT 389.660 4179.670 389.940 4179.950 ;
        RECT 390.280 4179.670 390.560 4179.950 ;
        RECT 390.900 4179.670 391.180 4179.950 ;
        RECT 391.520 4179.670 391.800 4179.950 ;
        RECT 392.140 4179.670 392.420 4179.950 ;
        RECT 392.760 4179.670 393.040 4179.950 ;
        RECT 389.040 4179.050 389.320 4179.330 ;
        RECT 389.660 4179.050 389.940 4179.330 ;
        RECT 390.280 4179.050 390.560 4179.330 ;
        RECT 390.900 4179.050 391.180 4179.330 ;
        RECT 391.520 4179.050 391.800 4179.330 ;
        RECT 392.140 4179.050 392.420 4179.330 ;
        RECT 392.760 4179.050 393.040 4179.330 ;
        RECT 389.040 4178.430 389.320 4178.710 ;
        RECT 389.660 4178.430 389.940 4178.710 ;
        RECT 390.280 4178.430 390.560 4178.710 ;
        RECT 390.900 4178.430 391.180 4178.710 ;
        RECT 391.520 4178.430 391.800 4178.710 ;
        RECT 392.140 4178.430 392.420 4178.710 ;
        RECT 392.760 4178.430 393.040 4178.710 ;
        RECT 389.040 4177.810 389.320 4178.090 ;
        RECT 389.660 4177.810 389.940 4178.090 ;
        RECT 390.280 4177.810 390.560 4178.090 ;
        RECT 390.900 4177.810 391.180 4178.090 ;
        RECT 391.520 4177.810 391.800 4178.090 ;
        RECT 392.140 4177.810 392.420 4178.090 ;
        RECT 392.760 4177.810 393.040 4178.090 ;
        RECT 389.040 4177.190 389.320 4177.470 ;
        RECT 389.660 4177.190 389.940 4177.470 ;
        RECT 390.280 4177.190 390.560 4177.470 ;
        RECT 390.900 4177.190 391.180 4177.470 ;
        RECT 391.520 4177.190 391.800 4177.470 ;
        RECT 392.140 4177.190 392.420 4177.470 ;
        RECT 392.760 4177.190 393.040 4177.470 ;
        RECT 389.040 4176.570 389.320 4176.850 ;
        RECT 389.660 4176.570 389.940 4176.850 ;
        RECT 390.280 4176.570 390.560 4176.850 ;
        RECT 390.900 4176.570 391.180 4176.850 ;
        RECT 391.520 4176.570 391.800 4176.850 ;
        RECT 392.140 4176.570 392.420 4176.850 ;
        RECT 392.760 4176.570 393.040 4176.850 ;
        RECT 389.040 4175.950 389.320 4176.230 ;
        RECT 389.660 4175.950 389.940 4176.230 ;
        RECT 390.280 4175.950 390.560 4176.230 ;
        RECT 390.900 4175.950 391.180 4176.230 ;
        RECT 391.520 4175.950 391.800 4176.230 ;
        RECT 392.140 4175.950 392.420 4176.230 ;
        RECT 392.760 4175.950 393.040 4176.230 ;
        RECT 389.040 4175.330 389.320 4175.610 ;
        RECT 389.660 4175.330 389.940 4175.610 ;
        RECT 390.280 4175.330 390.560 4175.610 ;
        RECT 390.900 4175.330 391.180 4175.610 ;
        RECT 391.520 4175.330 391.800 4175.610 ;
        RECT 392.140 4175.330 392.420 4175.610 ;
        RECT 392.760 4175.330 393.040 4175.610 ;
        RECT 389.040 4174.710 389.320 4174.990 ;
        RECT 389.660 4174.710 389.940 4174.990 ;
        RECT 390.280 4174.710 390.560 4174.990 ;
        RECT 390.900 4174.710 391.180 4174.990 ;
        RECT 391.520 4174.710 391.800 4174.990 ;
        RECT 392.140 4174.710 392.420 4174.990 ;
        RECT 392.760 4174.710 393.040 4174.990 ;
        RECT 389.040 4174.090 389.320 4174.370 ;
        RECT 389.660 4174.090 389.940 4174.370 ;
        RECT 390.280 4174.090 390.560 4174.370 ;
        RECT 390.900 4174.090 391.180 4174.370 ;
        RECT 391.520 4174.090 391.800 4174.370 ;
        RECT 392.140 4174.090 392.420 4174.370 ;
        RECT 392.760 4174.090 393.040 4174.370 ;
        RECT 389.040 4173.470 389.320 4173.750 ;
        RECT 389.660 4173.470 389.940 4173.750 ;
        RECT 390.280 4173.470 390.560 4173.750 ;
        RECT 390.900 4173.470 391.180 4173.750 ;
        RECT 391.520 4173.470 391.800 4173.750 ;
        RECT 392.140 4173.470 392.420 4173.750 ;
        RECT 392.760 4173.470 393.040 4173.750 ;
        RECT 389.040 4172.850 389.320 4173.130 ;
        RECT 389.660 4172.850 389.940 4173.130 ;
        RECT 390.280 4172.850 390.560 4173.130 ;
        RECT 390.900 4172.850 391.180 4173.130 ;
        RECT 391.520 4172.850 391.800 4173.130 ;
        RECT 392.140 4172.850 392.420 4173.130 ;
        RECT 392.760 4172.850 393.040 4173.130 ;
        RECT 389.040 4172.230 389.320 4172.510 ;
        RECT 389.660 4172.230 389.940 4172.510 ;
        RECT 390.280 4172.230 390.560 4172.510 ;
        RECT 390.900 4172.230 391.180 4172.510 ;
        RECT 391.520 4172.230 391.800 4172.510 ;
        RECT 392.140 4172.230 392.420 4172.510 ;
        RECT 392.760 4172.230 393.040 4172.510 ;
        RECT 389.040 4171.610 389.320 4171.890 ;
        RECT 389.660 4171.610 389.940 4171.890 ;
        RECT 390.280 4171.610 390.560 4171.890 ;
        RECT 390.900 4171.610 391.180 4171.890 ;
        RECT 391.520 4171.610 391.800 4171.890 ;
        RECT 392.140 4171.610 392.420 4171.890 ;
        RECT 392.760 4171.610 393.040 4171.890 ;
        RECT 389.040 4170.990 389.320 4171.270 ;
        RECT 389.660 4170.990 389.940 4171.270 ;
        RECT 390.280 4170.990 390.560 4171.270 ;
        RECT 390.900 4170.990 391.180 4171.270 ;
        RECT 391.520 4170.990 391.800 4171.270 ;
        RECT 392.140 4170.990 392.420 4171.270 ;
        RECT 392.760 4170.990 393.040 4171.270 ;
        RECT 350.370 4168.410 350.650 4168.690 ;
        RECT 350.370 4167.790 350.650 4168.070 ;
        RECT 350.370 4167.170 350.650 4167.450 ;
        RECT 350.370 4166.550 350.650 4166.830 ;
        RECT 350.370 4165.930 350.650 4166.210 ;
        RECT 350.370 4165.310 350.650 4165.590 ;
        RECT 350.370 4164.690 350.650 4164.970 ;
        RECT 350.370 4164.070 350.650 4164.350 ;
        RECT 350.370 4163.450 350.650 4163.730 ;
        RECT 350.370 4162.830 350.650 4163.110 ;
        RECT 350.370 4162.210 350.650 4162.490 ;
        RECT 350.370 4161.590 350.650 4161.870 ;
        RECT 350.370 4160.970 350.650 4161.250 ;
        RECT 350.370 4160.350 350.650 4160.630 ;
        RECT 350.370 4159.730 350.650 4160.010 ;
        RECT 350.370 4159.110 350.650 4159.390 ;
        RECT 389.040 4168.440 389.320 4168.720 ;
        RECT 389.660 4168.440 389.940 4168.720 ;
        RECT 390.280 4168.440 390.560 4168.720 ;
        RECT 390.900 4168.440 391.180 4168.720 ;
        RECT 391.520 4168.440 391.800 4168.720 ;
        RECT 392.140 4168.440 392.420 4168.720 ;
        RECT 392.760 4168.440 393.040 4168.720 ;
        RECT 389.040 4167.820 389.320 4168.100 ;
        RECT 389.660 4167.820 389.940 4168.100 ;
        RECT 390.280 4167.820 390.560 4168.100 ;
        RECT 390.900 4167.820 391.180 4168.100 ;
        RECT 391.520 4167.820 391.800 4168.100 ;
        RECT 392.140 4167.820 392.420 4168.100 ;
        RECT 392.760 4167.820 393.040 4168.100 ;
        RECT 389.040 4167.200 389.320 4167.480 ;
        RECT 389.660 4167.200 389.940 4167.480 ;
        RECT 390.280 4167.200 390.560 4167.480 ;
        RECT 390.900 4167.200 391.180 4167.480 ;
        RECT 391.520 4167.200 391.800 4167.480 ;
        RECT 392.140 4167.200 392.420 4167.480 ;
        RECT 392.760 4167.200 393.040 4167.480 ;
        RECT 389.040 4166.580 389.320 4166.860 ;
        RECT 389.660 4166.580 389.940 4166.860 ;
        RECT 390.280 4166.580 390.560 4166.860 ;
        RECT 390.900 4166.580 391.180 4166.860 ;
        RECT 391.520 4166.580 391.800 4166.860 ;
        RECT 392.140 4166.580 392.420 4166.860 ;
        RECT 392.760 4166.580 393.040 4166.860 ;
        RECT 389.040 4165.960 389.320 4166.240 ;
        RECT 389.660 4165.960 389.940 4166.240 ;
        RECT 390.280 4165.960 390.560 4166.240 ;
        RECT 390.900 4165.960 391.180 4166.240 ;
        RECT 391.520 4165.960 391.800 4166.240 ;
        RECT 392.140 4165.960 392.420 4166.240 ;
        RECT 392.760 4165.960 393.040 4166.240 ;
        RECT 389.040 4165.340 389.320 4165.620 ;
        RECT 389.660 4165.340 389.940 4165.620 ;
        RECT 390.280 4165.340 390.560 4165.620 ;
        RECT 390.900 4165.340 391.180 4165.620 ;
        RECT 391.520 4165.340 391.800 4165.620 ;
        RECT 392.140 4165.340 392.420 4165.620 ;
        RECT 392.760 4165.340 393.040 4165.620 ;
        RECT 389.040 4164.720 389.320 4165.000 ;
        RECT 389.660 4164.720 389.940 4165.000 ;
        RECT 390.280 4164.720 390.560 4165.000 ;
        RECT 390.900 4164.720 391.180 4165.000 ;
        RECT 391.520 4164.720 391.800 4165.000 ;
        RECT 392.140 4164.720 392.420 4165.000 ;
        RECT 392.760 4164.720 393.040 4165.000 ;
        RECT 389.040 4164.100 389.320 4164.380 ;
        RECT 389.660 4164.100 389.940 4164.380 ;
        RECT 390.280 4164.100 390.560 4164.380 ;
        RECT 390.900 4164.100 391.180 4164.380 ;
        RECT 391.520 4164.100 391.800 4164.380 ;
        RECT 392.140 4164.100 392.420 4164.380 ;
        RECT 392.760 4164.100 393.040 4164.380 ;
        RECT 389.040 4163.480 389.320 4163.760 ;
        RECT 389.660 4163.480 389.940 4163.760 ;
        RECT 390.280 4163.480 390.560 4163.760 ;
        RECT 390.900 4163.480 391.180 4163.760 ;
        RECT 391.520 4163.480 391.800 4163.760 ;
        RECT 392.140 4163.480 392.420 4163.760 ;
        RECT 392.760 4163.480 393.040 4163.760 ;
        RECT 389.040 4162.860 389.320 4163.140 ;
        RECT 389.660 4162.860 389.940 4163.140 ;
        RECT 390.280 4162.860 390.560 4163.140 ;
        RECT 390.900 4162.860 391.180 4163.140 ;
        RECT 391.520 4162.860 391.800 4163.140 ;
        RECT 392.140 4162.860 392.420 4163.140 ;
        RECT 392.760 4162.860 393.040 4163.140 ;
        RECT 389.040 4162.240 389.320 4162.520 ;
        RECT 389.660 4162.240 389.940 4162.520 ;
        RECT 390.280 4162.240 390.560 4162.520 ;
        RECT 390.900 4162.240 391.180 4162.520 ;
        RECT 391.520 4162.240 391.800 4162.520 ;
        RECT 392.140 4162.240 392.420 4162.520 ;
        RECT 392.760 4162.240 393.040 4162.520 ;
        RECT 389.040 4161.620 389.320 4161.900 ;
        RECT 389.660 4161.620 389.940 4161.900 ;
        RECT 390.280 4161.620 390.560 4161.900 ;
        RECT 390.900 4161.620 391.180 4161.900 ;
        RECT 391.520 4161.620 391.800 4161.900 ;
        RECT 392.140 4161.620 392.420 4161.900 ;
        RECT 392.760 4161.620 393.040 4161.900 ;
        RECT 389.040 4161.000 389.320 4161.280 ;
        RECT 389.660 4161.000 389.940 4161.280 ;
        RECT 390.280 4161.000 390.560 4161.280 ;
        RECT 390.900 4161.000 391.180 4161.280 ;
        RECT 391.520 4161.000 391.800 4161.280 ;
        RECT 392.140 4161.000 392.420 4161.280 ;
        RECT 392.760 4161.000 393.040 4161.280 ;
        RECT 389.040 4160.380 389.320 4160.660 ;
        RECT 389.660 4160.380 389.940 4160.660 ;
        RECT 390.280 4160.380 390.560 4160.660 ;
        RECT 390.900 4160.380 391.180 4160.660 ;
        RECT 391.520 4160.380 391.800 4160.660 ;
        RECT 392.140 4160.380 392.420 4160.660 ;
        RECT 392.760 4160.380 393.040 4160.660 ;
        RECT 389.040 4159.760 389.320 4160.040 ;
        RECT 389.660 4159.760 389.940 4160.040 ;
        RECT 390.280 4159.760 390.560 4160.040 ;
        RECT 390.900 4159.760 391.180 4160.040 ;
        RECT 391.520 4159.760 391.800 4160.040 ;
        RECT 392.140 4159.760 392.420 4160.040 ;
        RECT 392.760 4159.760 393.040 4160.040 ;
        RECT 389.040 4159.140 389.320 4159.420 ;
        RECT 389.660 4159.140 389.940 4159.420 ;
        RECT 390.280 4159.140 390.560 4159.420 ;
        RECT 390.900 4159.140 391.180 4159.420 ;
        RECT 391.520 4159.140 391.800 4159.420 ;
        RECT 392.140 4159.140 392.420 4159.420 ;
        RECT 392.760 4159.140 393.040 4159.420 ;
        RECT 350.370 4155.390 350.650 4155.670 ;
        RECT 350.370 4154.770 350.650 4155.050 ;
        RECT 350.370 4154.150 350.650 4154.430 ;
        RECT 350.370 4153.530 350.650 4153.810 ;
        RECT 350.370 4152.910 350.650 4153.190 ;
        RECT 350.370 4152.290 350.650 4152.570 ;
        RECT 350.370 4151.670 350.650 4151.950 ;
        RECT 350.370 4151.050 350.650 4151.330 ;
        RECT 350.370 4150.430 350.650 4150.710 ;
        RECT 350.370 4149.810 350.650 4150.090 ;
        RECT 350.370 4149.190 350.650 4149.470 ;
        RECT 350.370 4148.570 350.650 4148.850 ;
        RECT 350.370 4147.950 350.650 4148.230 ;
        RECT 350.370 4147.330 350.650 4147.610 ;
        RECT 350.370 4146.710 350.650 4146.990 ;
        RECT 389.040 4155.420 389.320 4155.700 ;
        RECT 389.660 4155.420 389.940 4155.700 ;
        RECT 390.280 4155.420 390.560 4155.700 ;
        RECT 390.900 4155.420 391.180 4155.700 ;
        RECT 391.520 4155.420 391.800 4155.700 ;
        RECT 392.140 4155.420 392.420 4155.700 ;
        RECT 392.760 4155.420 393.040 4155.700 ;
        RECT 389.040 4154.800 389.320 4155.080 ;
        RECT 389.660 4154.800 389.940 4155.080 ;
        RECT 390.280 4154.800 390.560 4155.080 ;
        RECT 390.900 4154.800 391.180 4155.080 ;
        RECT 391.520 4154.800 391.800 4155.080 ;
        RECT 392.140 4154.800 392.420 4155.080 ;
        RECT 392.760 4154.800 393.040 4155.080 ;
        RECT 389.040 4154.180 389.320 4154.460 ;
        RECT 389.660 4154.180 389.940 4154.460 ;
        RECT 390.280 4154.180 390.560 4154.460 ;
        RECT 390.900 4154.180 391.180 4154.460 ;
        RECT 391.520 4154.180 391.800 4154.460 ;
        RECT 392.140 4154.180 392.420 4154.460 ;
        RECT 392.760 4154.180 393.040 4154.460 ;
        RECT 389.040 4153.560 389.320 4153.840 ;
        RECT 389.660 4153.560 389.940 4153.840 ;
        RECT 390.280 4153.560 390.560 4153.840 ;
        RECT 390.900 4153.560 391.180 4153.840 ;
        RECT 391.520 4153.560 391.800 4153.840 ;
        RECT 392.140 4153.560 392.420 4153.840 ;
        RECT 392.760 4153.560 393.040 4153.840 ;
        RECT 389.040 4152.940 389.320 4153.220 ;
        RECT 389.660 4152.940 389.940 4153.220 ;
        RECT 390.280 4152.940 390.560 4153.220 ;
        RECT 390.900 4152.940 391.180 4153.220 ;
        RECT 391.520 4152.940 391.800 4153.220 ;
        RECT 392.140 4152.940 392.420 4153.220 ;
        RECT 392.760 4152.940 393.040 4153.220 ;
        RECT 389.040 4152.320 389.320 4152.600 ;
        RECT 389.660 4152.320 389.940 4152.600 ;
        RECT 390.280 4152.320 390.560 4152.600 ;
        RECT 390.900 4152.320 391.180 4152.600 ;
        RECT 391.520 4152.320 391.800 4152.600 ;
        RECT 392.140 4152.320 392.420 4152.600 ;
        RECT 392.760 4152.320 393.040 4152.600 ;
        RECT 389.040 4151.700 389.320 4151.980 ;
        RECT 389.660 4151.700 389.940 4151.980 ;
        RECT 390.280 4151.700 390.560 4151.980 ;
        RECT 390.900 4151.700 391.180 4151.980 ;
        RECT 391.520 4151.700 391.800 4151.980 ;
        RECT 392.140 4151.700 392.420 4151.980 ;
        RECT 392.760 4151.700 393.040 4151.980 ;
        RECT 389.040 4151.080 389.320 4151.360 ;
        RECT 389.660 4151.080 389.940 4151.360 ;
        RECT 390.280 4151.080 390.560 4151.360 ;
        RECT 390.900 4151.080 391.180 4151.360 ;
        RECT 391.520 4151.080 391.800 4151.360 ;
        RECT 392.140 4151.080 392.420 4151.360 ;
        RECT 392.760 4151.080 393.040 4151.360 ;
        RECT 389.040 4150.460 389.320 4150.740 ;
        RECT 389.660 4150.460 389.940 4150.740 ;
        RECT 390.280 4150.460 390.560 4150.740 ;
        RECT 390.900 4150.460 391.180 4150.740 ;
        RECT 391.520 4150.460 391.800 4150.740 ;
        RECT 392.140 4150.460 392.420 4150.740 ;
        RECT 392.760 4150.460 393.040 4150.740 ;
        RECT 389.040 4149.840 389.320 4150.120 ;
        RECT 389.660 4149.840 389.940 4150.120 ;
        RECT 390.280 4149.840 390.560 4150.120 ;
        RECT 390.900 4149.840 391.180 4150.120 ;
        RECT 391.520 4149.840 391.800 4150.120 ;
        RECT 392.140 4149.840 392.420 4150.120 ;
        RECT 392.760 4149.840 393.040 4150.120 ;
        RECT 389.040 4149.220 389.320 4149.500 ;
        RECT 389.660 4149.220 389.940 4149.500 ;
        RECT 390.280 4149.220 390.560 4149.500 ;
        RECT 390.900 4149.220 391.180 4149.500 ;
        RECT 391.520 4149.220 391.800 4149.500 ;
        RECT 392.140 4149.220 392.420 4149.500 ;
        RECT 392.760 4149.220 393.040 4149.500 ;
        RECT 389.040 4148.600 389.320 4148.880 ;
        RECT 389.660 4148.600 389.940 4148.880 ;
        RECT 390.280 4148.600 390.560 4148.880 ;
        RECT 390.900 4148.600 391.180 4148.880 ;
        RECT 391.520 4148.600 391.800 4148.880 ;
        RECT 392.140 4148.600 392.420 4148.880 ;
        RECT 392.760 4148.600 393.040 4148.880 ;
        RECT 389.040 4147.980 389.320 4148.260 ;
        RECT 389.660 4147.980 389.940 4148.260 ;
        RECT 390.280 4147.980 390.560 4148.260 ;
        RECT 390.900 4147.980 391.180 4148.260 ;
        RECT 391.520 4147.980 391.800 4148.260 ;
        RECT 392.140 4147.980 392.420 4148.260 ;
        RECT 392.760 4147.980 393.040 4148.260 ;
        RECT 389.040 4147.360 389.320 4147.640 ;
        RECT 389.660 4147.360 389.940 4147.640 ;
        RECT 390.280 4147.360 390.560 4147.640 ;
        RECT 390.900 4147.360 391.180 4147.640 ;
        RECT 391.520 4147.360 391.800 4147.640 ;
        RECT 392.140 4147.360 392.420 4147.640 ;
        RECT 392.760 4147.360 393.040 4147.640 ;
        RECT 389.040 4146.740 389.320 4147.020 ;
        RECT 389.660 4146.740 389.940 4147.020 ;
        RECT 390.280 4146.740 390.560 4147.020 ;
        RECT 390.900 4146.740 391.180 4147.020 ;
        RECT 391.520 4146.740 391.800 4147.020 ;
        RECT 392.140 4146.740 392.420 4147.020 ;
        RECT 392.760 4146.740 393.040 4147.020 ;
        RECT 388.740 4032.670 389.020 4032.950 ;
        RECT 389.360 4032.670 389.640 4032.950 ;
        RECT 389.980 4032.670 390.260 4032.950 ;
        RECT 390.600 4032.670 390.880 4032.950 ;
        RECT 391.220 4032.670 391.500 4032.950 ;
        RECT 391.840 4032.670 392.120 4032.950 ;
        RECT 392.460 4032.670 392.740 4032.950 ;
        RECT 388.740 4032.050 389.020 4032.330 ;
        RECT 389.360 4032.050 389.640 4032.330 ;
        RECT 389.980 4032.050 390.260 4032.330 ;
        RECT 390.600 4032.050 390.880 4032.330 ;
        RECT 391.220 4032.050 391.500 4032.330 ;
        RECT 391.840 4032.050 392.120 4032.330 ;
        RECT 392.460 4032.050 392.740 4032.330 ;
        RECT 388.740 4031.430 389.020 4031.710 ;
        RECT 389.360 4031.430 389.640 4031.710 ;
        RECT 389.980 4031.430 390.260 4031.710 ;
        RECT 390.600 4031.430 390.880 4031.710 ;
        RECT 391.220 4031.430 391.500 4031.710 ;
        RECT 391.840 4031.430 392.120 4031.710 ;
        RECT 392.460 4031.430 392.740 4031.710 ;
        RECT 388.740 4030.810 389.020 4031.090 ;
        RECT 389.360 4030.810 389.640 4031.090 ;
        RECT 389.980 4030.810 390.260 4031.090 ;
        RECT 390.600 4030.810 390.880 4031.090 ;
        RECT 391.220 4030.810 391.500 4031.090 ;
        RECT 391.840 4030.810 392.120 4031.090 ;
        RECT 392.460 4030.810 392.740 4031.090 ;
        RECT 388.740 4030.190 389.020 4030.470 ;
        RECT 389.360 4030.190 389.640 4030.470 ;
        RECT 389.980 4030.190 390.260 4030.470 ;
        RECT 390.600 4030.190 390.880 4030.470 ;
        RECT 391.220 4030.190 391.500 4030.470 ;
        RECT 391.840 4030.190 392.120 4030.470 ;
        RECT 392.460 4030.190 392.740 4030.470 ;
        RECT 350.370 4013.010 350.650 4013.290 ;
        RECT 350.370 4012.390 350.650 4012.670 ;
        RECT 350.370 4011.770 350.650 4012.050 ;
        RECT 350.370 4011.150 350.650 4011.430 ;
        RECT 350.370 4010.530 350.650 4010.810 ;
        RECT 350.370 4009.910 350.650 4010.190 ;
        RECT 350.370 4009.290 350.650 4009.570 ;
        RECT 350.370 4008.670 350.650 4008.950 ;
        RECT 350.370 4008.050 350.650 4008.330 ;
        RECT 350.370 4007.430 350.650 4007.710 ;
        RECT 350.370 4006.810 350.650 4007.090 ;
        RECT 350.370 4006.190 350.650 4006.470 ;
        RECT 350.370 4005.570 350.650 4005.850 ;
        RECT 350.370 4004.950 350.650 4005.230 ;
        RECT 350.370 4004.330 350.650 4004.610 ;
        RECT 350.370 4000.640 350.650 4000.920 ;
        RECT 350.370 4000.020 350.650 4000.300 ;
        RECT 350.370 3999.400 350.650 3999.680 ;
        RECT 350.370 3998.780 350.650 3999.060 ;
        RECT 350.370 3998.160 350.650 3998.440 ;
        RECT 350.370 3997.540 350.650 3997.820 ;
        RECT 350.370 3996.920 350.650 3997.200 ;
        RECT 350.370 3996.300 350.650 3996.580 ;
        RECT 350.370 3995.680 350.650 3995.960 ;
        RECT 350.370 3995.060 350.650 3995.340 ;
        RECT 350.370 3994.440 350.650 3994.720 ;
        RECT 350.370 3993.820 350.650 3994.100 ;
        RECT 350.370 3993.200 350.650 3993.480 ;
        RECT 350.370 3992.580 350.650 3992.860 ;
        RECT 350.370 3991.960 350.650 3992.240 ;
        RECT 350.370 3991.340 350.650 3991.620 ;
        RECT 350.370 3988.790 350.650 3989.070 ;
        RECT 350.370 3988.170 350.650 3988.450 ;
        RECT 350.370 3987.550 350.650 3987.830 ;
        RECT 350.370 3986.930 350.650 3987.210 ;
        RECT 350.370 3986.310 350.650 3986.590 ;
        RECT 350.370 3985.690 350.650 3985.970 ;
        RECT 350.370 3985.070 350.650 3985.350 ;
        RECT 350.370 3984.450 350.650 3984.730 ;
        RECT 350.370 3983.830 350.650 3984.110 ;
        RECT 350.370 3983.210 350.650 3983.490 ;
        RECT 350.370 3982.590 350.650 3982.870 ;
        RECT 350.370 3981.970 350.650 3982.250 ;
        RECT 350.370 3981.350 350.650 3981.630 ;
        RECT 350.370 3980.730 350.650 3981.010 ;
        RECT 350.370 3980.110 350.650 3980.390 ;
        RECT 350.370 3979.490 350.650 3979.770 ;
        RECT 350.370 3975.260 350.650 3975.540 ;
        RECT 350.370 3974.640 350.650 3974.920 ;
        RECT 350.370 3974.020 350.650 3974.300 ;
        RECT 350.370 3973.400 350.650 3973.680 ;
        RECT 350.370 3972.780 350.650 3973.060 ;
        RECT 350.370 3972.160 350.650 3972.440 ;
        RECT 350.370 3971.540 350.650 3971.820 ;
        RECT 350.370 3970.920 350.650 3971.200 ;
        RECT 350.370 3970.300 350.650 3970.580 ;
        RECT 350.370 3969.680 350.650 3969.960 ;
        RECT 350.370 3969.060 350.650 3969.340 ;
        RECT 350.370 3968.440 350.650 3968.720 ;
        RECT 350.370 3967.820 350.650 3968.100 ;
        RECT 350.370 3967.200 350.650 3967.480 ;
        RECT 350.370 3966.580 350.650 3966.860 ;
        RECT 350.370 3965.960 350.650 3966.240 ;
        RECT 350.370 3963.410 350.650 3963.690 ;
        RECT 350.370 3962.790 350.650 3963.070 ;
        RECT 350.370 3962.170 350.650 3962.450 ;
        RECT 350.370 3961.550 350.650 3961.830 ;
        RECT 350.370 3960.930 350.650 3961.210 ;
        RECT 350.370 3960.310 350.650 3960.590 ;
        RECT 350.370 3959.690 350.650 3959.970 ;
        RECT 350.370 3959.070 350.650 3959.350 ;
        RECT 350.370 3958.450 350.650 3958.730 ;
        RECT 350.370 3957.830 350.650 3958.110 ;
        RECT 350.370 3957.210 350.650 3957.490 ;
        RECT 350.370 3956.590 350.650 3956.870 ;
        RECT 350.370 3955.970 350.650 3956.250 ;
        RECT 350.370 3955.350 350.650 3955.630 ;
        RECT 350.370 3954.730 350.650 3955.010 ;
        RECT 350.370 3954.110 350.650 3954.390 ;
        RECT 350.370 3950.390 350.650 3950.670 ;
        RECT 350.370 3949.770 350.650 3950.050 ;
        RECT 350.370 3949.150 350.650 3949.430 ;
        RECT 350.370 3948.530 350.650 3948.810 ;
        RECT 350.370 3947.910 350.650 3948.190 ;
        RECT 350.370 3947.290 350.650 3947.570 ;
        RECT 350.370 3946.670 350.650 3946.950 ;
        RECT 350.370 3946.050 350.650 3946.330 ;
        RECT 350.370 3945.430 350.650 3945.710 ;
        RECT 350.370 3944.810 350.650 3945.090 ;
        RECT 350.370 3944.190 350.650 3944.470 ;
        RECT 350.370 3943.570 350.650 3943.850 ;
        RECT 350.370 3942.950 350.650 3943.230 ;
        RECT 350.370 3942.330 350.650 3942.610 ;
        RECT 350.370 3941.710 350.650 3941.990 ;
        RECT 388.965 3907.920 389.245 3908.200 ;
        RECT 389.585 3907.920 389.865 3908.200 ;
        RECT 390.205 3907.920 390.485 3908.200 ;
        RECT 390.825 3907.920 391.105 3908.200 ;
        RECT 391.445 3907.920 391.725 3908.200 ;
        RECT 392.065 3907.920 392.345 3908.200 ;
        RECT 392.685 3907.920 392.965 3908.200 ;
        RECT 388.740 3852.670 389.020 3852.950 ;
        RECT 389.360 3852.670 389.640 3852.950 ;
        RECT 389.980 3852.670 390.260 3852.950 ;
        RECT 390.600 3852.670 390.880 3852.950 ;
        RECT 391.220 3852.670 391.500 3852.950 ;
        RECT 391.840 3852.670 392.120 3852.950 ;
        RECT 392.460 3852.670 392.740 3852.950 ;
        RECT 388.740 3852.050 389.020 3852.330 ;
        RECT 389.360 3852.050 389.640 3852.330 ;
        RECT 389.980 3852.050 390.260 3852.330 ;
        RECT 390.600 3852.050 390.880 3852.330 ;
        RECT 391.220 3852.050 391.500 3852.330 ;
        RECT 391.840 3852.050 392.120 3852.330 ;
        RECT 392.460 3852.050 392.740 3852.330 ;
        RECT 388.740 3851.430 389.020 3851.710 ;
        RECT 389.360 3851.430 389.640 3851.710 ;
        RECT 389.980 3851.430 390.260 3851.710 ;
        RECT 390.600 3851.430 390.880 3851.710 ;
        RECT 391.220 3851.430 391.500 3851.710 ;
        RECT 391.840 3851.430 392.120 3851.710 ;
        RECT 392.460 3851.430 392.740 3851.710 ;
        RECT 388.740 3850.810 389.020 3851.090 ;
        RECT 389.360 3850.810 389.640 3851.090 ;
        RECT 389.980 3850.810 390.260 3851.090 ;
        RECT 390.600 3850.810 390.880 3851.090 ;
        RECT 391.220 3850.810 391.500 3851.090 ;
        RECT 391.840 3850.810 392.120 3851.090 ;
        RECT 392.460 3850.810 392.740 3851.090 ;
        RECT 388.740 3850.190 389.020 3850.470 ;
        RECT 389.360 3850.190 389.640 3850.470 ;
        RECT 389.980 3850.190 390.260 3850.470 ;
        RECT 390.600 3850.190 390.880 3850.470 ;
        RECT 391.220 3850.190 391.500 3850.470 ;
        RECT 391.840 3850.190 392.120 3850.470 ;
        RECT 392.460 3850.190 392.740 3850.470 ;
        RECT 388.965 3810.590 389.245 3810.870 ;
        RECT 389.585 3810.590 389.865 3810.870 ;
        RECT 390.205 3810.590 390.485 3810.870 ;
        RECT 390.825 3810.590 391.105 3810.870 ;
        RECT 391.445 3810.590 391.725 3810.870 ;
        RECT 392.065 3810.590 392.345 3810.870 ;
        RECT 392.685 3810.590 392.965 3810.870 ;
        RECT 388.965 3809.970 389.245 3810.250 ;
        RECT 389.585 3809.970 389.865 3810.250 ;
        RECT 390.205 3809.970 390.485 3810.250 ;
        RECT 390.825 3809.970 391.105 3810.250 ;
        RECT 391.445 3809.970 391.725 3810.250 ;
        RECT 392.065 3809.970 392.345 3810.250 ;
        RECT 392.685 3809.970 392.965 3810.250 ;
        RECT 388.965 3775.590 389.245 3775.870 ;
        RECT 389.585 3775.590 389.865 3775.870 ;
        RECT 390.205 3775.590 390.485 3775.870 ;
        RECT 390.825 3775.590 391.105 3775.870 ;
        RECT 391.445 3775.590 391.725 3775.870 ;
        RECT 392.065 3775.590 392.345 3775.870 ;
        RECT 392.685 3775.590 392.965 3775.870 ;
        RECT 388.965 3774.970 389.245 3775.250 ;
        RECT 389.585 3774.970 389.865 3775.250 ;
        RECT 390.205 3774.970 390.485 3775.250 ;
        RECT 390.825 3774.970 391.105 3775.250 ;
        RECT 391.445 3774.970 391.725 3775.250 ;
        RECT 392.065 3774.970 392.345 3775.250 ;
        RECT 392.685 3774.970 392.965 3775.250 ;
        RECT 388.965 3740.590 389.245 3740.870 ;
        RECT 389.585 3740.590 389.865 3740.870 ;
        RECT 390.205 3740.590 390.485 3740.870 ;
        RECT 390.825 3740.590 391.105 3740.870 ;
        RECT 391.445 3740.590 391.725 3740.870 ;
        RECT 392.065 3740.590 392.345 3740.870 ;
        RECT 392.685 3740.590 392.965 3740.870 ;
        RECT 388.965 3739.970 389.245 3740.250 ;
        RECT 389.585 3739.970 389.865 3740.250 ;
        RECT 390.205 3739.970 390.485 3740.250 ;
        RECT 390.825 3739.970 391.105 3740.250 ;
        RECT 391.445 3739.970 391.725 3740.250 ;
        RECT 392.065 3739.970 392.345 3740.250 ;
        RECT 392.685 3739.970 392.965 3740.250 ;
        RECT 388.965 3702.920 389.245 3703.200 ;
        RECT 389.585 3702.920 389.865 3703.200 ;
        RECT 390.205 3702.920 390.485 3703.200 ;
        RECT 390.825 3702.920 391.105 3703.200 ;
        RECT 391.445 3702.920 391.725 3703.200 ;
        RECT 392.065 3702.920 392.345 3703.200 ;
        RECT 392.685 3702.920 392.965 3703.200 ;
        RECT 388.740 3672.670 389.020 3672.950 ;
        RECT 389.360 3672.670 389.640 3672.950 ;
        RECT 389.980 3672.670 390.260 3672.950 ;
        RECT 390.600 3672.670 390.880 3672.950 ;
        RECT 391.220 3672.670 391.500 3672.950 ;
        RECT 391.840 3672.670 392.120 3672.950 ;
        RECT 392.460 3672.670 392.740 3672.950 ;
        RECT 388.740 3672.050 389.020 3672.330 ;
        RECT 389.360 3672.050 389.640 3672.330 ;
        RECT 389.980 3672.050 390.260 3672.330 ;
        RECT 390.600 3672.050 390.880 3672.330 ;
        RECT 391.220 3672.050 391.500 3672.330 ;
        RECT 391.840 3672.050 392.120 3672.330 ;
        RECT 392.460 3672.050 392.740 3672.330 ;
        RECT 388.740 3671.430 389.020 3671.710 ;
        RECT 389.360 3671.430 389.640 3671.710 ;
        RECT 389.980 3671.430 390.260 3671.710 ;
        RECT 390.600 3671.430 390.880 3671.710 ;
        RECT 391.220 3671.430 391.500 3671.710 ;
        RECT 391.840 3671.430 392.120 3671.710 ;
        RECT 392.460 3671.430 392.740 3671.710 ;
        RECT 388.740 3670.810 389.020 3671.090 ;
        RECT 389.360 3670.810 389.640 3671.090 ;
        RECT 389.980 3670.810 390.260 3671.090 ;
        RECT 390.600 3670.810 390.880 3671.090 ;
        RECT 391.220 3670.810 391.500 3671.090 ;
        RECT 391.840 3670.810 392.120 3671.090 ;
        RECT 392.460 3670.810 392.740 3671.090 ;
        RECT 388.740 3670.190 389.020 3670.470 ;
        RECT 389.360 3670.190 389.640 3670.470 ;
        RECT 389.980 3670.190 390.260 3670.470 ;
        RECT 390.600 3670.190 390.880 3670.470 ;
        RECT 391.220 3670.190 391.500 3670.470 ;
        RECT 391.840 3670.190 392.120 3670.470 ;
        RECT 392.460 3670.190 392.740 3670.470 ;
        RECT 388.965 3605.590 389.245 3605.870 ;
        RECT 389.585 3605.590 389.865 3605.870 ;
        RECT 390.205 3605.590 390.485 3605.870 ;
        RECT 390.825 3605.590 391.105 3605.870 ;
        RECT 391.445 3605.590 391.725 3605.870 ;
        RECT 392.065 3605.590 392.345 3605.870 ;
        RECT 392.685 3605.590 392.965 3605.870 ;
        RECT 388.965 3604.970 389.245 3605.250 ;
        RECT 389.585 3604.970 389.865 3605.250 ;
        RECT 390.205 3604.970 390.485 3605.250 ;
        RECT 390.825 3604.970 391.105 3605.250 ;
        RECT 391.445 3604.970 391.725 3605.250 ;
        RECT 392.065 3604.970 392.345 3605.250 ;
        RECT 392.685 3604.970 392.965 3605.250 ;
        RECT 388.965 3570.590 389.245 3570.870 ;
        RECT 389.585 3570.590 389.865 3570.870 ;
        RECT 390.205 3570.590 390.485 3570.870 ;
        RECT 390.825 3570.590 391.105 3570.870 ;
        RECT 391.445 3570.590 391.725 3570.870 ;
        RECT 392.065 3570.590 392.345 3570.870 ;
        RECT 392.685 3570.590 392.965 3570.870 ;
        RECT 388.965 3569.970 389.245 3570.250 ;
        RECT 389.585 3569.970 389.865 3570.250 ;
        RECT 390.205 3569.970 390.485 3570.250 ;
        RECT 390.825 3569.970 391.105 3570.250 ;
        RECT 391.445 3569.970 391.725 3570.250 ;
        RECT 392.065 3569.970 392.345 3570.250 ;
        RECT 392.685 3569.970 392.965 3570.250 ;
        RECT 388.965 3535.590 389.245 3535.870 ;
        RECT 389.585 3535.590 389.865 3535.870 ;
        RECT 390.205 3535.590 390.485 3535.870 ;
        RECT 390.825 3535.590 391.105 3535.870 ;
        RECT 391.445 3535.590 391.725 3535.870 ;
        RECT 392.065 3535.590 392.345 3535.870 ;
        RECT 392.685 3535.590 392.965 3535.870 ;
        RECT 388.965 3534.970 389.245 3535.250 ;
        RECT 389.585 3534.970 389.865 3535.250 ;
        RECT 390.205 3534.970 390.485 3535.250 ;
        RECT 390.825 3534.970 391.105 3535.250 ;
        RECT 391.445 3534.970 391.725 3535.250 ;
        RECT 392.065 3534.970 392.345 3535.250 ;
        RECT 392.685 3534.970 392.965 3535.250 ;
        RECT 388.965 3497.920 389.245 3498.200 ;
        RECT 389.585 3497.920 389.865 3498.200 ;
        RECT 390.205 3497.920 390.485 3498.200 ;
        RECT 390.825 3497.920 391.105 3498.200 ;
        RECT 391.445 3497.920 391.725 3498.200 ;
        RECT 392.065 3497.920 392.345 3498.200 ;
        RECT 392.685 3497.920 392.965 3498.200 ;
        RECT 388.740 3492.670 389.020 3492.950 ;
        RECT 389.360 3492.670 389.640 3492.950 ;
        RECT 389.980 3492.670 390.260 3492.950 ;
        RECT 390.600 3492.670 390.880 3492.950 ;
        RECT 391.220 3492.670 391.500 3492.950 ;
        RECT 391.840 3492.670 392.120 3492.950 ;
        RECT 392.460 3492.670 392.740 3492.950 ;
        RECT 388.740 3492.050 389.020 3492.330 ;
        RECT 389.360 3492.050 389.640 3492.330 ;
        RECT 389.980 3492.050 390.260 3492.330 ;
        RECT 390.600 3492.050 390.880 3492.330 ;
        RECT 391.220 3492.050 391.500 3492.330 ;
        RECT 391.840 3492.050 392.120 3492.330 ;
        RECT 392.460 3492.050 392.740 3492.330 ;
        RECT 388.740 3491.430 389.020 3491.710 ;
        RECT 389.360 3491.430 389.640 3491.710 ;
        RECT 389.980 3491.430 390.260 3491.710 ;
        RECT 390.600 3491.430 390.880 3491.710 ;
        RECT 391.220 3491.430 391.500 3491.710 ;
        RECT 391.840 3491.430 392.120 3491.710 ;
        RECT 392.460 3491.430 392.740 3491.710 ;
        RECT 388.740 3490.810 389.020 3491.090 ;
        RECT 389.360 3490.810 389.640 3491.090 ;
        RECT 389.980 3490.810 390.260 3491.090 ;
        RECT 390.600 3490.810 390.880 3491.090 ;
        RECT 391.220 3490.810 391.500 3491.090 ;
        RECT 391.840 3490.810 392.120 3491.090 ;
        RECT 392.460 3490.810 392.740 3491.090 ;
        RECT 388.740 3490.190 389.020 3490.470 ;
        RECT 389.360 3490.190 389.640 3490.470 ;
        RECT 389.980 3490.190 390.260 3490.470 ;
        RECT 390.600 3490.190 390.880 3490.470 ;
        RECT 391.220 3490.190 391.500 3490.470 ;
        RECT 391.840 3490.190 392.120 3490.470 ;
        RECT 392.460 3490.190 392.740 3490.470 ;
        RECT 388.965 3400.590 389.245 3400.870 ;
        RECT 389.585 3400.590 389.865 3400.870 ;
        RECT 390.205 3400.590 390.485 3400.870 ;
        RECT 390.825 3400.590 391.105 3400.870 ;
        RECT 391.445 3400.590 391.725 3400.870 ;
        RECT 392.065 3400.590 392.345 3400.870 ;
        RECT 392.685 3400.590 392.965 3400.870 ;
        RECT 388.965 3399.970 389.245 3400.250 ;
        RECT 389.585 3399.970 389.865 3400.250 ;
        RECT 390.205 3399.970 390.485 3400.250 ;
        RECT 390.825 3399.970 391.105 3400.250 ;
        RECT 391.445 3399.970 391.725 3400.250 ;
        RECT 392.065 3399.970 392.345 3400.250 ;
        RECT 392.685 3399.970 392.965 3400.250 ;
        RECT 388.965 3365.590 389.245 3365.870 ;
        RECT 389.585 3365.590 389.865 3365.870 ;
        RECT 390.205 3365.590 390.485 3365.870 ;
        RECT 390.825 3365.590 391.105 3365.870 ;
        RECT 391.445 3365.590 391.725 3365.870 ;
        RECT 392.065 3365.590 392.345 3365.870 ;
        RECT 392.685 3365.590 392.965 3365.870 ;
        RECT 388.965 3364.970 389.245 3365.250 ;
        RECT 389.585 3364.970 389.865 3365.250 ;
        RECT 390.205 3364.970 390.485 3365.250 ;
        RECT 390.825 3364.970 391.105 3365.250 ;
        RECT 391.445 3364.970 391.725 3365.250 ;
        RECT 392.065 3364.970 392.345 3365.250 ;
        RECT 392.685 3364.970 392.965 3365.250 ;
        RECT 388.965 3330.590 389.245 3330.870 ;
        RECT 389.585 3330.590 389.865 3330.870 ;
        RECT 390.205 3330.590 390.485 3330.870 ;
        RECT 390.825 3330.590 391.105 3330.870 ;
        RECT 391.445 3330.590 391.725 3330.870 ;
        RECT 392.065 3330.590 392.345 3330.870 ;
        RECT 392.685 3330.590 392.965 3330.870 ;
        RECT 388.965 3329.970 389.245 3330.250 ;
        RECT 389.585 3329.970 389.865 3330.250 ;
        RECT 390.205 3329.970 390.485 3330.250 ;
        RECT 390.825 3329.970 391.105 3330.250 ;
        RECT 391.445 3329.970 391.725 3330.250 ;
        RECT 392.065 3329.970 392.345 3330.250 ;
        RECT 392.685 3329.970 392.965 3330.250 ;
        RECT 388.740 3312.670 389.020 3312.950 ;
        RECT 389.360 3312.670 389.640 3312.950 ;
        RECT 389.980 3312.670 390.260 3312.950 ;
        RECT 390.600 3312.670 390.880 3312.950 ;
        RECT 391.220 3312.670 391.500 3312.950 ;
        RECT 391.840 3312.670 392.120 3312.950 ;
        RECT 392.460 3312.670 392.740 3312.950 ;
        RECT 388.740 3312.050 389.020 3312.330 ;
        RECT 389.360 3312.050 389.640 3312.330 ;
        RECT 389.980 3312.050 390.260 3312.330 ;
        RECT 390.600 3312.050 390.880 3312.330 ;
        RECT 391.220 3312.050 391.500 3312.330 ;
        RECT 391.840 3312.050 392.120 3312.330 ;
        RECT 392.460 3312.050 392.740 3312.330 ;
        RECT 388.740 3311.430 389.020 3311.710 ;
        RECT 389.360 3311.430 389.640 3311.710 ;
        RECT 389.980 3311.430 390.260 3311.710 ;
        RECT 390.600 3311.430 390.880 3311.710 ;
        RECT 391.220 3311.430 391.500 3311.710 ;
        RECT 391.840 3311.430 392.120 3311.710 ;
        RECT 392.460 3311.430 392.740 3311.710 ;
        RECT 388.740 3310.810 389.020 3311.090 ;
        RECT 389.360 3310.810 389.640 3311.090 ;
        RECT 389.980 3310.810 390.260 3311.090 ;
        RECT 390.600 3310.810 390.880 3311.090 ;
        RECT 391.220 3310.810 391.500 3311.090 ;
        RECT 391.840 3310.810 392.120 3311.090 ;
        RECT 392.460 3310.810 392.740 3311.090 ;
        RECT 388.740 3310.190 389.020 3310.470 ;
        RECT 389.360 3310.190 389.640 3310.470 ;
        RECT 389.980 3310.190 390.260 3310.470 ;
        RECT 390.600 3310.190 390.880 3310.470 ;
        RECT 391.220 3310.190 391.500 3310.470 ;
        RECT 391.840 3310.190 392.120 3310.470 ;
        RECT 392.460 3310.190 392.740 3310.470 ;
        RECT 388.965 3292.920 389.245 3293.200 ;
        RECT 389.585 3292.920 389.865 3293.200 ;
        RECT 390.205 3292.920 390.485 3293.200 ;
        RECT 390.825 3292.920 391.105 3293.200 ;
        RECT 391.445 3292.920 391.725 3293.200 ;
        RECT 392.065 3292.920 392.345 3293.200 ;
        RECT 392.685 3292.920 392.965 3293.200 ;
        RECT 388.965 3195.590 389.245 3195.870 ;
        RECT 389.585 3195.590 389.865 3195.870 ;
        RECT 390.205 3195.590 390.485 3195.870 ;
        RECT 390.825 3195.590 391.105 3195.870 ;
        RECT 391.445 3195.590 391.725 3195.870 ;
        RECT 392.065 3195.590 392.345 3195.870 ;
        RECT 392.685 3195.590 392.965 3195.870 ;
        RECT 388.965 3194.970 389.245 3195.250 ;
        RECT 389.585 3194.970 389.865 3195.250 ;
        RECT 390.205 3194.970 390.485 3195.250 ;
        RECT 390.825 3194.970 391.105 3195.250 ;
        RECT 391.445 3194.970 391.725 3195.250 ;
        RECT 392.065 3194.970 392.345 3195.250 ;
        RECT 392.685 3194.970 392.965 3195.250 ;
        RECT 388.965 3160.590 389.245 3160.870 ;
        RECT 389.585 3160.590 389.865 3160.870 ;
        RECT 390.205 3160.590 390.485 3160.870 ;
        RECT 390.825 3160.590 391.105 3160.870 ;
        RECT 391.445 3160.590 391.725 3160.870 ;
        RECT 392.065 3160.590 392.345 3160.870 ;
        RECT 392.685 3160.590 392.965 3160.870 ;
        RECT 388.965 3159.970 389.245 3160.250 ;
        RECT 389.585 3159.970 389.865 3160.250 ;
        RECT 390.205 3159.970 390.485 3160.250 ;
        RECT 390.825 3159.970 391.105 3160.250 ;
        RECT 391.445 3159.970 391.725 3160.250 ;
        RECT 392.065 3159.970 392.345 3160.250 ;
        RECT 392.685 3159.970 392.965 3160.250 ;
        RECT 388.740 3132.670 389.020 3132.950 ;
        RECT 389.360 3132.670 389.640 3132.950 ;
        RECT 389.980 3132.670 390.260 3132.950 ;
        RECT 390.600 3132.670 390.880 3132.950 ;
        RECT 391.220 3132.670 391.500 3132.950 ;
        RECT 391.840 3132.670 392.120 3132.950 ;
        RECT 392.460 3132.670 392.740 3132.950 ;
        RECT 388.740 3132.050 389.020 3132.330 ;
        RECT 389.360 3132.050 389.640 3132.330 ;
        RECT 389.980 3132.050 390.260 3132.330 ;
        RECT 390.600 3132.050 390.880 3132.330 ;
        RECT 391.220 3132.050 391.500 3132.330 ;
        RECT 391.840 3132.050 392.120 3132.330 ;
        RECT 392.460 3132.050 392.740 3132.330 ;
        RECT 388.740 3131.430 389.020 3131.710 ;
        RECT 389.360 3131.430 389.640 3131.710 ;
        RECT 389.980 3131.430 390.260 3131.710 ;
        RECT 390.600 3131.430 390.880 3131.710 ;
        RECT 391.220 3131.430 391.500 3131.710 ;
        RECT 391.840 3131.430 392.120 3131.710 ;
        RECT 392.460 3131.430 392.740 3131.710 ;
        RECT 388.740 3130.810 389.020 3131.090 ;
        RECT 389.360 3130.810 389.640 3131.090 ;
        RECT 389.980 3130.810 390.260 3131.090 ;
        RECT 390.600 3130.810 390.880 3131.090 ;
        RECT 391.220 3130.810 391.500 3131.090 ;
        RECT 391.840 3130.810 392.120 3131.090 ;
        RECT 392.460 3130.810 392.740 3131.090 ;
        RECT 388.740 3130.190 389.020 3130.470 ;
        RECT 389.360 3130.190 389.640 3130.470 ;
        RECT 389.980 3130.190 390.260 3130.470 ;
        RECT 390.600 3130.190 390.880 3130.470 ;
        RECT 391.220 3130.190 391.500 3130.470 ;
        RECT 391.840 3130.190 392.120 3130.470 ;
        RECT 392.460 3130.190 392.740 3130.470 ;
        RECT 388.965 3125.590 389.245 3125.870 ;
        RECT 389.585 3125.590 389.865 3125.870 ;
        RECT 390.205 3125.590 390.485 3125.870 ;
        RECT 390.825 3125.590 391.105 3125.870 ;
        RECT 391.445 3125.590 391.725 3125.870 ;
        RECT 392.065 3125.590 392.345 3125.870 ;
        RECT 392.685 3125.590 392.965 3125.870 ;
        RECT 388.965 3124.970 389.245 3125.250 ;
        RECT 389.585 3124.970 389.865 3125.250 ;
        RECT 390.205 3124.970 390.485 3125.250 ;
        RECT 390.825 3124.970 391.105 3125.250 ;
        RECT 391.445 3124.970 391.725 3125.250 ;
        RECT 392.065 3124.970 392.345 3125.250 ;
        RECT 392.685 3124.970 392.965 3125.250 ;
        RECT 388.965 3087.920 389.245 3088.200 ;
        RECT 389.585 3087.920 389.865 3088.200 ;
        RECT 390.205 3087.920 390.485 3088.200 ;
        RECT 390.825 3087.920 391.105 3088.200 ;
        RECT 391.445 3087.920 391.725 3088.200 ;
        RECT 392.065 3087.920 392.345 3088.200 ;
        RECT 392.685 3087.920 392.965 3088.200 ;
        RECT 388.965 2990.590 389.245 2990.870 ;
        RECT 389.585 2990.590 389.865 2990.870 ;
        RECT 390.205 2990.590 390.485 2990.870 ;
        RECT 390.825 2990.590 391.105 2990.870 ;
        RECT 391.445 2990.590 391.725 2990.870 ;
        RECT 392.065 2990.590 392.345 2990.870 ;
        RECT 392.685 2990.590 392.965 2990.870 ;
        RECT 388.965 2989.970 389.245 2990.250 ;
        RECT 389.585 2989.970 389.865 2990.250 ;
        RECT 390.205 2989.970 390.485 2990.250 ;
        RECT 390.825 2989.970 391.105 2990.250 ;
        RECT 391.445 2989.970 391.725 2990.250 ;
        RECT 392.065 2989.970 392.345 2990.250 ;
        RECT 392.685 2989.970 392.965 2990.250 ;
        RECT 388.965 2955.590 389.245 2955.870 ;
        RECT 389.585 2955.590 389.865 2955.870 ;
        RECT 390.205 2955.590 390.485 2955.870 ;
        RECT 390.825 2955.590 391.105 2955.870 ;
        RECT 391.445 2955.590 391.725 2955.870 ;
        RECT 392.065 2955.590 392.345 2955.870 ;
        RECT 392.685 2955.590 392.965 2955.870 ;
        RECT 388.965 2954.970 389.245 2955.250 ;
        RECT 389.585 2954.970 389.865 2955.250 ;
        RECT 390.205 2954.970 390.485 2955.250 ;
        RECT 390.825 2954.970 391.105 2955.250 ;
        RECT 391.445 2954.970 391.725 2955.250 ;
        RECT 392.065 2954.970 392.345 2955.250 ;
        RECT 392.685 2954.970 392.965 2955.250 ;
        RECT 388.740 2952.670 389.020 2952.950 ;
        RECT 389.360 2952.670 389.640 2952.950 ;
        RECT 389.980 2952.670 390.260 2952.950 ;
        RECT 390.600 2952.670 390.880 2952.950 ;
        RECT 391.220 2952.670 391.500 2952.950 ;
        RECT 391.840 2952.670 392.120 2952.950 ;
        RECT 392.460 2952.670 392.740 2952.950 ;
        RECT 388.740 2952.050 389.020 2952.330 ;
        RECT 389.360 2952.050 389.640 2952.330 ;
        RECT 389.980 2952.050 390.260 2952.330 ;
        RECT 390.600 2952.050 390.880 2952.330 ;
        RECT 391.220 2952.050 391.500 2952.330 ;
        RECT 391.840 2952.050 392.120 2952.330 ;
        RECT 392.460 2952.050 392.740 2952.330 ;
        RECT 388.740 2951.430 389.020 2951.710 ;
        RECT 389.360 2951.430 389.640 2951.710 ;
        RECT 389.980 2951.430 390.260 2951.710 ;
        RECT 390.600 2951.430 390.880 2951.710 ;
        RECT 391.220 2951.430 391.500 2951.710 ;
        RECT 391.840 2951.430 392.120 2951.710 ;
        RECT 392.460 2951.430 392.740 2951.710 ;
        RECT 388.740 2950.810 389.020 2951.090 ;
        RECT 389.360 2950.810 389.640 2951.090 ;
        RECT 389.980 2950.810 390.260 2951.090 ;
        RECT 390.600 2950.810 390.880 2951.090 ;
        RECT 391.220 2950.810 391.500 2951.090 ;
        RECT 391.840 2950.810 392.120 2951.090 ;
        RECT 392.460 2950.810 392.740 2951.090 ;
        RECT 388.740 2950.190 389.020 2950.470 ;
        RECT 389.360 2950.190 389.640 2950.470 ;
        RECT 389.980 2950.190 390.260 2950.470 ;
        RECT 390.600 2950.190 390.880 2950.470 ;
        RECT 391.220 2950.190 391.500 2950.470 ;
        RECT 391.840 2950.190 392.120 2950.470 ;
        RECT 392.460 2950.190 392.740 2950.470 ;
        RECT 388.965 2920.590 389.245 2920.870 ;
        RECT 389.585 2920.590 389.865 2920.870 ;
        RECT 390.205 2920.590 390.485 2920.870 ;
        RECT 390.825 2920.590 391.105 2920.870 ;
        RECT 391.445 2920.590 391.725 2920.870 ;
        RECT 392.065 2920.590 392.345 2920.870 ;
        RECT 392.685 2920.590 392.965 2920.870 ;
        RECT 388.965 2919.970 389.245 2920.250 ;
        RECT 389.585 2919.970 389.865 2920.250 ;
        RECT 390.205 2919.970 390.485 2920.250 ;
        RECT 390.825 2919.970 391.105 2920.250 ;
        RECT 391.445 2919.970 391.725 2920.250 ;
        RECT 392.065 2919.970 392.345 2920.250 ;
        RECT 392.685 2919.970 392.965 2920.250 ;
        RECT 388.965 2882.920 389.245 2883.200 ;
        RECT 389.585 2882.920 389.865 2883.200 ;
        RECT 390.205 2882.920 390.485 2883.200 ;
        RECT 390.825 2882.920 391.105 2883.200 ;
        RECT 391.445 2882.920 391.725 2883.200 ;
        RECT 392.065 2882.920 392.345 2883.200 ;
        RECT 392.685 2882.920 392.965 2883.200 ;
        RECT 388.965 2785.590 389.245 2785.870 ;
        RECT 389.585 2785.590 389.865 2785.870 ;
        RECT 390.205 2785.590 390.485 2785.870 ;
        RECT 390.825 2785.590 391.105 2785.870 ;
        RECT 391.445 2785.590 391.725 2785.870 ;
        RECT 392.065 2785.590 392.345 2785.870 ;
        RECT 392.685 2785.590 392.965 2785.870 ;
        RECT 388.965 2784.970 389.245 2785.250 ;
        RECT 389.585 2784.970 389.865 2785.250 ;
        RECT 390.205 2784.970 390.485 2785.250 ;
        RECT 390.825 2784.970 391.105 2785.250 ;
        RECT 391.445 2784.970 391.725 2785.250 ;
        RECT 392.065 2784.970 392.345 2785.250 ;
        RECT 392.685 2784.970 392.965 2785.250 ;
        RECT 388.740 2772.670 389.020 2772.950 ;
        RECT 389.360 2772.670 389.640 2772.950 ;
        RECT 389.980 2772.670 390.260 2772.950 ;
        RECT 390.600 2772.670 390.880 2772.950 ;
        RECT 391.220 2772.670 391.500 2772.950 ;
        RECT 391.840 2772.670 392.120 2772.950 ;
        RECT 392.460 2772.670 392.740 2772.950 ;
        RECT 388.740 2772.050 389.020 2772.330 ;
        RECT 389.360 2772.050 389.640 2772.330 ;
        RECT 389.980 2772.050 390.260 2772.330 ;
        RECT 390.600 2772.050 390.880 2772.330 ;
        RECT 391.220 2772.050 391.500 2772.330 ;
        RECT 391.840 2772.050 392.120 2772.330 ;
        RECT 392.460 2772.050 392.740 2772.330 ;
        RECT 388.740 2771.430 389.020 2771.710 ;
        RECT 389.360 2771.430 389.640 2771.710 ;
        RECT 389.980 2771.430 390.260 2771.710 ;
        RECT 390.600 2771.430 390.880 2771.710 ;
        RECT 391.220 2771.430 391.500 2771.710 ;
        RECT 391.840 2771.430 392.120 2771.710 ;
        RECT 392.460 2771.430 392.740 2771.710 ;
        RECT 388.740 2770.810 389.020 2771.090 ;
        RECT 389.360 2770.810 389.640 2771.090 ;
        RECT 389.980 2770.810 390.260 2771.090 ;
        RECT 390.600 2770.810 390.880 2771.090 ;
        RECT 391.220 2770.810 391.500 2771.090 ;
        RECT 391.840 2770.810 392.120 2771.090 ;
        RECT 392.460 2770.810 392.740 2771.090 ;
        RECT 388.740 2770.190 389.020 2770.470 ;
        RECT 389.360 2770.190 389.640 2770.470 ;
        RECT 389.980 2770.190 390.260 2770.470 ;
        RECT 390.600 2770.190 390.880 2770.470 ;
        RECT 391.220 2770.190 391.500 2770.470 ;
        RECT 391.840 2770.190 392.120 2770.470 ;
        RECT 392.460 2770.190 392.740 2770.470 ;
        RECT 388.965 2750.590 389.245 2750.870 ;
        RECT 389.585 2750.590 389.865 2750.870 ;
        RECT 390.205 2750.590 390.485 2750.870 ;
        RECT 390.825 2750.590 391.105 2750.870 ;
        RECT 391.445 2750.590 391.725 2750.870 ;
        RECT 392.065 2750.590 392.345 2750.870 ;
        RECT 392.685 2750.590 392.965 2750.870 ;
        RECT 388.965 2749.970 389.245 2750.250 ;
        RECT 389.585 2749.970 389.865 2750.250 ;
        RECT 390.205 2749.970 390.485 2750.250 ;
        RECT 390.825 2749.970 391.105 2750.250 ;
        RECT 391.445 2749.970 391.725 2750.250 ;
        RECT 392.065 2749.970 392.345 2750.250 ;
        RECT 392.685 2749.970 392.965 2750.250 ;
        RECT 388.965 2715.590 389.245 2715.870 ;
        RECT 389.585 2715.590 389.865 2715.870 ;
        RECT 390.205 2715.590 390.485 2715.870 ;
        RECT 390.825 2715.590 391.105 2715.870 ;
        RECT 391.445 2715.590 391.725 2715.870 ;
        RECT 392.065 2715.590 392.345 2715.870 ;
        RECT 392.685 2715.590 392.965 2715.870 ;
        RECT 388.965 2714.970 389.245 2715.250 ;
        RECT 389.585 2714.970 389.865 2715.250 ;
        RECT 390.205 2714.970 390.485 2715.250 ;
        RECT 390.825 2714.970 391.105 2715.250 ;
        RECT 391.445 2714.970 391.725 2715.250 ;
        RECT 392.065 2714.970 392.345 2715.250 ;
        RECT 392.685 2714.970 392.965 2715.250 ;
        RECT 388.965 2677.920 389.245 2678.200 ;
        RECT 389.585 2677.920 389.865 2678.200 ;
        RECT 390.205 2677.920 390.485 2678.200 ;
        RECT 390.825 2677.920 391.105 2678.200 ;
        RECT 391.445 2677.920 391.725 2678.200 ;
        RECT 392.065 2677.920 392.345 2678.200 ;
        RECT 392.685 2677.920 392.965 2678.200 ;
        RECT 388.740 2592.670 389.020 2592.950 ;
        RECT 389.360 2592.670 389.640 2592.950 ;
        RECT 389.980 2592.670 390.260 2592.950 ;
        RECT 390.600 2592.670 390.880 2592.950 ;
        RECT 391.220 2592.670 391.500 2592.950 ;
        RECT 391.840 2592.670 392.120 2592.950 ;
        RECT 392.460 2592.670 392.740 2592.950 ;
        RECT 388.740 2592.050 389.020 2592.330 ;
        RECT 389.360 2592.050 389.640 2592.330 ;
        RECT 389.980 2592.050 390.260 2592.330 ;
        RECT 390.600 2592.050 390.880 2592.330 ;
        RECT 391.220 2592.050 391.500 2592.330 ;
        RECT 391.840 2592.050 392.120 2592.330 ;
        RECT 392.460 2592.050 392.740 2592.330 ;
        RECT 388.740 2591.430 389.020 2591.710 ;
        RECT 389.360 2591.430 389.640 2591.710 ;
        RECT 389.980 2591.430 390.260 2591.710 ;
        RECT 390.600 2591.430 390.880 2591.710 ;
        RECT 391.220 2591.430 391.500 2591.710 ;
        RECT 391.840 2591.430 392.120 2591.710 ;
        RECT 392.460 2591.430 392.740 2591.710 ;
        RECT 388.740 2590.810 389.020 2591.090 ;
        RECT 389.360 2590.810 389.640 2591.090 ;
        RECT 389.980 2590.810 390.260 2591.090 ;
        RECT 390.600 2590.810 390.880 2591.090 ;
        RECT 391.220 2590.810 391.500 2591.090 ;
        RECT 391.840 2590.810 392.120 2591.090 ;
        RECT 392.460 2590.810 392.740 2591.090 ;
        RECT 388.740 2590.190 389.020 2590.470 ;
        RECT 389.360 2590.190 389.640 2590.470 ;
        RECT 389.980 2590.190 390.260 2590.470 ;
        RECT 390.600 2590.190 390.880 2590.470 ;
        RECT 391.220 2590.190 391.500 2590.470 ;
        RECT 391.840 2590.190 392.120 2590.470 ;
        RECT 392.460 2590.190 392.740 2590.470 ;
        RECT 388.965 2580.590 389.245 2580.870 ;
        RECT 389.585 2580.590 389.865 2580.870 ;
        RECT 390.205 2580.590 390.485 2580.870 ;
        RECT 390.825 2580.590 391.105 2580.870 ;
        RECT 391.445 2580.590 391.725 2580.870 ;
        RECT 392.065 2580.590 392.345 2580.870 ;
        RECT 392.685 2580.590 392.965 2580.870 ;
        RECT 388.965 2579.970 389.245 2580.250 ;
        RECT 389.585 2579.970 389.865 2580.250 ;
        RECT 390.205 2579.970 390.485 2580.250 ;
        RECT 390.825 2579.970 391.105 2580.250 ;
        RECT 391.445 2579.970 391.725 2580.250 ;
        RECT 392.065 2579.970 392.345 2580.250 ;
        RECT 392.685 2579.970 392.965 2580.250 ;
        RECT 388.965 2545.590 389.245 2545.870 ;
        RECT 389.585 2545.590 389.865 2545.870 ;
        RECT 390.205 2545.590 390.485 2545.870 ;
        RECT 390.825 2545.590 391.105 2545.870 ;
        RECT 391.445 2545.590 391.725 2545.870 ;
        RECT 392.065 2545.590 392.345 2545.870 ;
        RECT 392.685 2545.590 392.965 2545.870 ;
        RECT 388.965 2544.970 389.245 2545.250 ;
        RECT 389.585 2544.970 389.865 2545.250 ;
        RECT 390.205 2544.970 390.485 2545.250 ;
        RECT 390.825 2544.970 391.105 2545.250 ;
        RECT 391.445 2544.970 391.725 2545.250 ;
        RECT 392.065 2544.970 392.345 2545.250 ;
        RECT 392.685 2544.970 392.965 2545.250 ;
        RECT 388.965 2510.590 389.245 2510.870 ;
        RECT 389.585 2510.590 389.865 2510.870 ;
        RECT 390.205 2510.590 390.485 2510.870 ;
        RECT 390.825 2510.590 391.105 2510.870 ;
        RECT 391.445 2510.590 391.725 2510.870 ;
        RECT 392.065 2510.590 392.345 2510.870 ;
        RECT 392.685 2510.590 392.965 2510.870 ;
        RECT 388.965 2509.970 389.245 2510.250 ;
        RECT 389.585 2509.970 389.865 2510.250 ;
        RECT 390.205 2509.970 390.485 2510.250 ;
        RECT 390.825 2509.970 391.105 2510.250 ;
        RECT 391.445 2509.970 391.725 2510.250 ;
        RECT 392.065 2509.970 392.345 2510.250 ;
        RECT 392.685 2509.970 392.965 2510.250 ;
        RECT 388.740 2412.670 389.020 2412.950 ;
        RECT 389.360 2412.670 389.640 2412.950 ;
        RECT 389.980 2412.670 390.260 2412.950 ;
        RECT 390.600 2412.670 390.880 2412.950 ;
        RECT 391.220 2412.670 391.500 2412.950 ;
        RECT 391.840 2412.670 392.120 2412.950 ;
        RECT 392.460 2412.670 392.740 2412.950 ;
        RECT 388.740 2412.050 389.020 2412.330 ;
        RECT 389.360 2412.050 389.640 2412.330 ;
        RECT 389.980 2412.050 390.260 2412.330 ;
        RECT 390.600 2412.050 390.880 2412.330 ;
        RECT 391.220 2412.050 391.500 2412.330 ;
        RECT 391.840 2412.050 392.120 2412.330 ;
        RECT 392.460 2412.050 392.740 2412.330 ;
        RECT 388.740 2411.430 389.020 2411.710 ;
        RECT 389.360 2411.430 389.640 2411.710 ;
        RECT 389.980 2411.430 390.260 2411.710 ;
        RECT 390.600 2411.430 390.880 2411.710 ;
        RECT 391.220 2411.430 391.500 2411.710 ;
        RECT 391.840 2411.430 392.120 2411.710 ;
        RECT 392.460 2411.430 392.740 2411.710 ;
        RECT 388.740 2410.810 389.020 2411.090 ;
        RECT 389.360 2410.810 389.640 2411.090 ;
        RECT 389.980 2410.810 390.260 2411.090 ;
        RECT 390.600 2410.810 390.880 2411.090 ;
        RECT 391.220 2410.810 391.500 2411.090 ;
        RECT 391.840 2410.810 392.120 2411.090 ;
        RECT 392.460 2410.810 392.740 2411.090 ;
        RECT 388.740 2410.190 389.020 2410.470 ;
        RECT 389.360 2410.190 389.640 2410.470 ;
        RECT 389.980 2410.190 390.260 2410.470 ;
        RECT 390.600 2410.190 390.880 2410.470 ;
        RECT 391.220 2410.190 391.500 2410.470 ;
        RECT 391.840 2410.190 392.120 2410.470 ;
        RECT 392.460 2410.190 392.740 2410.470 ;
        RECT 350.370 2373.010 350.650 2373.290 ;
        RECT 350.370 2372.390 350.650 2372.670 ;
        RECT 350.370 2371.770 350.650 2372.050 ;
        RECT 350.370 2371.150 350.650 2371.430 ;
        RECT 350.370 2370.530 350.650 2370.810 ;
        RECT 350.370 2369.910 350.650 2370.190 ;
        RECT 350.370 2369.290 350.650 2369.570 ;
        RECT 350.370 2368.670 350.650 2368.950 ;
        RECT 350.370 2368.050 350.650 2368.330 ;
        RECT 350.370 2367.430 350.650 2367.710 ;
        RECT 350.370 2366.810 350.650 2367.090 ;
        RECT 350.370 2366.190 350.650 2366.470 ;
        RECT 350.370 2365.570 350.650 2365.850 ;
        RECT 350.370 2364.950 350.650 2365.230 ;
        RECT 350.370 2364.330 350.650 2364.610 ;
        RECT 389.040 2373.070 389.320 2373.350 ;
        RECT 389.660 2373.070 389.940 2373.350 ;
        RECT 390.280 2373.070 390.560 2373.350 ;
        RECT 390.900 2373.070 391.180 2373.350 ;
        RECT 391.520 2373.070 391.800 2373.350 ;
        RECT 392.140 2373.070 392.420 2373.350 ;
        RECT 392.760 2373.070 393.040 2373.350 ;
        RECT 389.040 2372.450 389.320 2372.730 ;
        RECT 389.660 2372.450 389.940 2372.730 ;
        RECT 390.280 2372.450 390.560 2372.730 ;
        RECT 390.900 2372.450 391.180 2372.730 ;
        RECT 391.520 2372.450 391.800 2372.730 ;
        RECT 392.140 2372.450 392.420 2372.730 ;
        RECT 392.760 2372.450 393.040 2372.730 ;
        RECT 389.040 2371.830 389.320 2372.110 ;
        RECT 389.660 2371.830 389.940 2372.110 ;
        RECT 390.280 2371.830 390.560 2372.110 ;
        RECT 390.900 2371.830 391.180 2372.110 ;
        RECT 391.520 2371.830 391.800 2372.110 ;
        RECT 392.140 2371.830 392.420 2372.110 ;
        RECT 392.760 2371.830 393.040 2372.110 ;
        RECT 389.040 2371.210 389.320 2371.490 ;
        RECT 389.660 2371.210 389.940 2371.490 ;
        RECT 390.280 2371.210 390.560 2371.490 ;
        RECT 390.900 2371.210 391.180 2371.490 ;
        RECT 391.520 2371.210 391.800 2371.490 ;
        RECT 392.140 2371.210 392.420 2371.490 ;
        RECT 392.760 2371.210 393.040 2371.490 ;
        RECT 389.040 2370.590 389.320 2370.870 ;
        RECT 389.660 2370.590 389.940 2370.870 ;
        RECT 390.280 2370.590 390.560 2370.870 ;
        RECT 390.900 2370.590 391.180 2370.870 ;
        RECT 391.520 2370.590 391.800 2370.870 ;
        RECT 392.140 2370.590 392.420 2370.870 ;
        RECT 392.760 2370.590 393.040 2370.870 ;
        RECT 389.040 2369.970 389.320 2370.250 ;
        RECT 389.660 2369.970 389.940 2370.250 ;
        RECT 390.280 2369.970 390.560 2370.250 ;
        RECT 390.900 2369.970 391.180 2370.250 ;
        RECT 391.520 2369.970 391.800 2370.250 ;
        RECT 392.140 2369.970 392.420 2370.250 ;
        RECT 392.760 2369.970 393.040 2370.250 ;
        RECT 389.040 2369.350 389.320 2369.630 ;
        RECT 389.660 2369.350 389.940 2369.630 ;
        RECT 390.280 2369.350 390.560 2369.630 ;
        RECT 390.900 2369.350 391.180 2369.630 ;
        RECT 391.520 2369.350 391.800 2369.630 ;
        RECT 392.140 2369.350 392.420 2369.630 ;
        RECT 392.760 2369.350 393.040 2369.630 ;
        RECT 389.040 2368.730 389.320 2369.010 ;
        RECT 389.660 2368.730 389.940 2369.010 ;
        RECT 390.280 2368.730 390.560 2369.010 ;
        RECT 390.900 2368.730 391.180 2369.010 ;
        RECT 391.520 2368.730 391.800 2369.010 ;
        RECT 392.140 2368.730 392.420 2369.010 ;
        RECT 392.760 2368.730 393.040 2369.010 ;
        RECT 389.040 2368.110 389.320 2368.390 ;
        RECT 389.660 2368.110 389.940 2368.390 ;
        RECT 390.280 2368.110 390.560 2368.390 ;
        RECT 390.900 2368.110 391.180 2368.390 ;
        RECT 391.520 2368.110 391.800 2368.390 ;
        RECT 392.140 2368.110 392.420 2368.390 ;
        RECT 392.760 2368.110 393.040 2368.390 ;
        RECT 389.040 2367.490 389.320 2367.770 ;
        RECT 389.660 2367.490 389.940 2367.770 ;
        RECT 390.280 2367.490 390.560 2367.770 ;
        RECT 390.900 2367.490 391.180 2367.770 ;
        RECT 391.520 2367.490 391.800 2367.770 ;
        RECT 392.140 2367.490 392.420 2367.770 ;
        RECT 392.760 2367.490 393.040 2367.770 ;
        RECT 389.040 2366.870 389.320 2367.150 ;
        RECT 389.660 2366.870 389.940 2367.150 ;
        RECT 390.280 2366.870 390.560 2367.150 ;
        RECT 390.900 2366.870 391.180 2367.150 ;
        RECT 391.520 2366.870 391.800 2367.150 ;
        RECT 392.140 2366.870 392.420 2367.150 ;
        RECT 392.760 2366.870 393.040 2367.150 ;
        RECT 389.040 2366.250 389.320 2366.530 ;
        RECT 389.660 2366.250 389.940 2366.530 ;
        RECT 390.280 2366.250 390.560 2366.530 ;
        RECT 390.900 2366.250 391.180 2366.530 ;
        RECT 391.520 2366.250 391.800 2366.530 ;
        RECT 392.140 2366.250 392.420 2366.530 ;
        RECT 392.760 2366.250 393.040 2366.530 ;
        RECT 389.040 2365.630 389.320 2365.910 ;
        RECT 389.660 2365.630 389.940 2365.910 ;
        RECT 390.280 2365.630 390.560 2365.910 ;
        RECT 390.900 2365.630 391.180 2365.910 ;
        RECT 391.520 2365.630 391.800 2365.910 ;
        RECT 392.140 2365.630 392.420 2365.910 ;
        RECT 392.760 2365.630 393.040 2365.910 ;
        RECT 389.040 2365.010 389.320 2365.290 ;
        RECT 389.660 2365.010 389.940 2365.290 ;
        RECT 390.280 2365.010 390.560 2365.290 ;
        RECT 390.900 2365.010 391.180 2365.290 ;
        RECT 391.520 2365.010 391.800 2365.290 ;
        RECT 392.140 2365.010 392.420 2365.290 ;
        RECT 392.760 2365.010 393.040 2365.290 ;
        RECT 389.040 2364.390 389.320 2364.670 ;
        RECT 389.660 2364.390 389.940 2364.670 ;
        RECT 390.280 2364.390 390.560 2364.670 ;
        RECT 390.900 2364.390 391.180 2364.670 ;
        RECT 391.520 2364.390 391.800 2364.670 ;
        RECT 392.140 2364.390 392.420 2364.670 ;
        RECT 392.760 2364.390 393.040 2364.670 ;
        RECT 350.370 2360.640 350.650 2360.920 ;
        RECT 350.370 2360.020 350.650 2360.300 ;
        RECT 350.370 2359.400 350.650 2359.680 ;
        RECT 350.370 2358.780 350.650 2359.060 ;
        RECT 350.370 2358.160 350.650 2358.440 ;
        RECT 350.370 2357.540 350.650 2357.820 ;
        RECT 350.370 2356.920 350.650 2357.200 ;
        RECT 350.370 2356.300 350.650 2356.580 ;
        RECT 350.370 2355.680 350.650 2355.960 ;
        RECT 350.370 2355.060 350.650 2355.340 ;
        RECT 350.370 2354.440 350.650 2354.720 ;
        RECT 350.370 2353.820 350.650 2354.100 ;
        RECT 350.370 2353.200 350.650 2353.480 ;
        RECT 350.370 2352.580 350.650 2352.860 ;
        RECT 350.370 2351.960 350.650 2352.240 ;
        RECT 350.370 2351.340 350.650 2351.620 ;
        RECT 389.040 2360.670 389.320 2360.950 ;
        RECT 389.660 2360.670 389.940 2360.950 ;
        RECT 390.280 2360.670 390.560 2360.950 ;
        RECT 390.900 2360.670 391.180 2360.950 ;
        RECT 391.520 2360.670 391.800 2360.950 ;
        RECT 392.140 2360.670 392.420 2360.950 ;
        RECT 392.760 2360.670 393.040 2360.950 ;
        RECT 389.040 2360.050 389.320 2360.330 ;
        RECT 389.660 2360.050 389.940 2360.330 ;
        RECT 390.280 2360.050 390.560 2360.330 ;
        RECT 390.900 2360.050 391.180 2360.330 ;
        RECT 391.520 2360.050 391.800 2360.330 ;
        RECT 392.140 2360.050 392.420 2360.330 ;
        RECT 392.760 2360.050 393.040 2360.330 ;
        RECT 389.040 2359.430 389.320 2359.710 ;
        RECT 389.660 2359.430 389.940 2359.710 ;
        RECT 390.280 2359.430 390.560 2359.710 ;
        RECT 390.900 2359.430 391.180 2359.710 ;
        RECT 391.520 2359.430 391.800 2359.710 ;
        RECT 392.140 2359.430 392.420 2359.710 ;
        RECT 392.760 2359.430 393.040 2359.710 ;
        RECT 389.040 2358.810 389.320 2359.090 ;
        RECT 389.660 2358.810 389.940 2359.090 ;
        RECT 390.280 2358.810 390.560 2359.090 ;
        RECT 390.900 2358.810 391.180 2359.090 ;
        RECT 391.520 2358.810 391.800 2359.090 ;
        RECT 392.140 2358.810 392.420 2359.090 ;
        RECT 392.760 2358.810 393.040 2359.090 ;
        RECT 389.040 2358.190 389.320 2358.470 ;
        RECT 389.660 2358.190 389.940 2358.470 ;
        RECT 390.280 2358.190 390.560 2358.470 ;
        RECT 390.900 2358.190 391.180 2358.470 ;
        RECT 391.520 2358.190 391.800 2358.470 ;
        RECT 392.140 2358.190 392.420 2358.470 ;
        RECT 392.760 2358.190 393.040 2358.470 ;
        RECT 389.040 2357.570 389.320 2357.850 ;
        RECT 389.660 2357.570 389.940 2357.850 ;
        RECT 390.280 2357.570 390.560 2357.850 ;
        RECT 390.900 2357.570 391.180 2357.850 ;
        RECT 391.520 2357.570 391.800 2357.850 ;
        RECT 392.140 2357.570 392.420 2357.850 ;
        RECT 392.760 2357.570 393.040 2357.850 ;
        RECT 389.040 2356.950 389.320 2357.230 ;
        RECT 389.660 2356.950 389.940 2357.230 ;
        RECT 390.280 2356.950 390.560 2357.230 ;
        RECT 390.900 2356.950 391.180 2357.230 ;
        RECT 391.520 2356.950 391.800 2357.230 ;
        RECT 392.140 2356.950 392.420 2357.230 ;
        RECT 392.760 2356.950 393.040 2357.230 ;
        RECT 389.040 2356.330 389.320 2356.610 ;
        RECT 389.660 2356.330 389.940 2356.610 ;
        RECT 390.280 2356.330 390.560 2356.610 ;
        RECT 390.900 2356.330 391.180 2356.610 ;
        RECT 391.520 2356.330 391.800 2356.610 ;
        RECT 392.140 2356.330 392.420 2356.610 ;
        RECT 392.760 2356.330 393.040 2356.610 ;
        RECT 389.040 2355.710 389.320 2355.990 ;
        RECT 389.660 2355.710 389.940 2355.990 ;
        RECT 390.280 2355.710 390.560 2355.990 ;
        RECT 390.900 2355.710 391.180 2355.990 ;
        RECT 391.520 2355.710 391.800 2355.990 ;
        RECT 392.140 2355.710 392.420 2355.990 ;
        RECT 392.760 2355.710 393.040 2355.990 ;
        RECT 389.040 2355.090 389.320 2355.370 ;
        RECT 389.660 2355.090 389.940 2355.370 ;
        RECT 390.280 2355.090 390.560 2355.370 ;
        RECT 390.900 2355.090 391.180 2355.370 ;
        RECT 391.520 2355.090 391.800 2355.370 ;
        RECT 392.140 2355.090 392.420 2355.370 ;
        RECT 392.760 2355.090 393.040 2355.370 ;
        RECT 389.040 2354.470 389.320 2354.750 ;
        RECT 389.660 2354.470 389.940 2354.750 ;
        RECT 390.280 2354.470 390.560 2354.750 ;
        RECT 390.900 2354.470 391.180 2354.750 ;
        RECT 391.520 2354.470 391.800 2354.750 ;
        RECT 392.140 2354.470 392.420 2354.750 ;
        RECT 392.760 2354.470 393.040 2354.750 ;
        RECT 389.040 2353.850 389.320 2354.130 ;
        RECT 389.660 2353.850 389.940 2354.130 ;
        RECT 390.280 2353.850 390.560 2354.130 ;
        RECT 390.900 2353.850 391.180 2354.130 ;
        RECT 391.520 2353.850 391.800 2354.130 ;
        RECT 392.140 2353.850 392.420 2354.130 ;
        RECT 392.760 2353.850 393.040 2354.130 ;
        RECT 389.040 2353.230 389.320 2353.510 ;
        RECT 389.660 2353.230 389.940 2353.510 ;
        RECT 390.280 2353.230 390.560 2353.510 ;
        RECT 390.900 2353.230 391.180 2353.510 ;
        RECT 391.520 2353.230 391.800 2353.510 ;
        RECT 392.140 2353.230 392.420 2353.510 ;
        RECT 392.760 2353.230 393.040 2353.510 ;
        RECT 389.040 2352.610 389.320 2352.890 ;
        RECT 389.660 2352.610 389.940 2352.890 ;
        RECT 390.280 2352.610 390.560 2352.890 ;
        RECT 390.900 2352.610 391.180 2352.890 ;
        RECT 391.520 2352.610 391.800 2352.890 ;
        RECT 392.140 2352.610 392.420 2352.890 ;
        RECT 392.760 2352.610 393.040 2352.890 ;
        RECT 389.040 2351.990 389.320 2352.270 ;
        RECT 389.660 2351.990 389.940 2352.270 ;
        RECT 390.280 2351.990 390.560 2352.270 ;
        RECT 390.900 2351.990 391.180 2352.270 ;
        RECT 391.520 2351.990 391.800 2352.270 ;
        RECT 392.140 2351.990 392.420 2352.270 ;
        RECT 392.760 2351.990 393.040 2352.270 ;
        RECT 389.040 2351.370 389.320 2351.650 ;
        RECT 389.660 2351.370 389.940 2351.650 ;
        RECT 390.280 2351.370 390.560 2351.650 ;
        RECT 390.900 2351.370 391.180 2351.650 ;
        RECT 391.520 2351.370 391.800 2351.650 ;
        RECT 392.140 2351.370 392.420 2351.650 ;
        RECT 392.760 2351.370 393.040 2351.650 ;
        RECT 350.370 2348.790 350.650 2349.070 ;
        RECT 350.370 2348.170 350.650 2348.450 ;
        RECT 350.370 2347.550 350.650 2347.830 ;
        RECT 350.370 2346.930 350.650 2347.210 ;
        RECT 350.370 2346.310 350.650 2346.590 ;
        RECT 350.370 2345.690 350.650 2345.970 ;
        RECT 350.370 2345.070 350.650 2345.350 ;
        RECT 350.370 2344.450 350.650 2344.730 ;
        RECT 350.370 2343.830 350.650 2344.110 ;
        RECT 350.370 2343.210 350.650 2343.490 ;
        RECT 350.370 2342.590 350.650 2342.870 ;
        RECT 350.370 2341.970 350.650 2342.250 ;
        RECT 350.370 2341.350 350.650 2341.630 ;
        RECT 350.370 2340.730 350.650 2341.010 ;
        RECT 350.370 2340.110 350.650 2340.390 ;
        RECT 350.370 2339.490 350.650 2339.770 ;
        RECT 389.040 2348.820 389.320 2349.100 ;
        RECT 389.660 2348.820 389.940 2349.100 ;
        RECT 390.280 2348.820 390.560 2349.100 ;
        RECT 390.900 2348.820 391.180 2349.100 ;
        RECT 391.520 2348.820 391.800 2349.100 ;
        RECT 392.140 2348.820 392.420 2349.100 ;
        RECT 392.760 2348.820 393.040 2349.100 ;
        RECT 389.040 2348.200 389.320 2348.480 ;
        RECT 389.660 2348.200 389.940 2348.480 ;
        RECT 390.280 2348.200 390.560 2348.480 ;
        RECT 390.900 2348.200 391.180 2348.480 ;
        RECT 391.520 2348.200 391.800 2348.480 ;
        RECT 392.140 2348.200 392.420 2348.480 ;
        RECT 392.760 2348.200 393.040 2348.480 ;
        RECT 389.040 2347.580 389.320 2347.860 ;
        RECT 389.660 2347.580 389.940 2347.860 ;
        RECT 390.280 2347.580 390.560 2347.860 ;
        RECT 390.900 2347.580 391.180 2347.860 ;
        RECT 391.520 2347.580 391.800 2347.860 ;
        RECT 392.140 2347.580 392.420 2347.860 ;
        RECT 392.760 2347.580 393.040 2347.860 ;
        RECT 389.040 2346.960 389.320 2347.240 ;
        RECT 389.660 2346.960 389.940 2347.240 ;
        RECT 390.280 2346.960 390.560 2347.240 ;
        RECT 390.900 2346.960 391.180 2347.240 ;
        RECT 391.520 2346.960 391.800 2347.240 ;
        RECT 392.140 2346.960 392.420 2347.240 ;
        RECT 392.760 2346.960 393.040 2347.240 ;
        RECT 389.040 2346.340 389.320 2346.620 ;
        RECT 389.660 2346.340 389.940 2346.620 ;
        RECT 390.280 2346.340 390.560 2346.620 ;
        RECT 390.900 2346.340 391.180 2346.620 ;
        RECT 391.520 2346.340 391.800 2346.620 ;
        RECT 392.140 2346.340 392.420 2346.620 ;
        RECT 392.760 2346.340 393.040 2346.620 ;
        RECT 389.040 2345.720 389.320 2346.000 ;
        RECT 389.660 2345.720 389.940 2346.000 ;
        RECT 390.280 2345.720 390.560 2346.000 ;
        RECT 390.900 2345.720 391.180 2346.000 ;
        RECT 391.520 2345.720 391.800 2346.000 ;
        RECT 392.140 2345.720 392.420 2346.000 ;
        RECT 392.760 2345.720 393.040 2346.000 ;
        RECT 389.040 2345.100 389.320 2345.380 ;
        RECT 389.660 2345.100 389.940 2345.380 ;
        RECT 390.280 2345.100 390.560 2345.380 ;
        RECT 390.900 2345.100 391.180 2345.380 ;
        RECT 391.520 2345.100 391.800 2345.380 ;
        RECT 392.140 2345.100 392.420 2345.380 ;
        RECT 392.760 2345.100 393.040 2345.380 ;
        RECT 389.040 2344.480 389.320 2344.760 ;
        RECT 389.660 2344.480 389.940 2344.760 ;
        RECT 390.280 2344.480 390.560 2344.760 ;
        RECT 390.900 2344.480 391.180 2344.760 ;
        RECT 391.520 2344.480 391.800 2344.760 ;
        RECT 392.140 2344.480 392.420 2344.760 ;
        RECT 392.760 2344.480 393.040 2344.760 ;
        RECT 389.040 2343.860 389.320 2344.140 ;
        RECT 389.660 2343.860 389.940 2344.140 ;
        RECT 390.280 2343.860 390.560 2344.140 ;
        RECT 390.900 2343.860 391.180 2344.140 ;
        RECT 391.520 2343.860 391.800 2344.140 ;
        RECT 392.140 2343.860 392.420 2344.140 ;
        RECT 392.760 2343.860 393.040 2344.140 ;
        RECT 389.040 2343.240 389.320 2343.520 ;
        RECT 389.660 2343.240 389.940 2343.520 ;
        RECT 390.280 2343.240 390.560 2343.520 ;
        RECT 390.900 2343.240 391.180 2343.520 ;
        RECT 391.520 2343.240 391.800 2343.520 ;
        RECT 392.140 2343.240 392.420 2343.520 ;
        RECT 392.760 2343.240 393.040 2343.520 ;
        RECT 389.040 2342.620 389.320 2342.900 ;
        RECT 389.660 2342.620 389.940 2342.900 ;
        RECT 390.280 2342.620 390.560 2342.900 ;
        RECT 390.900 2342.620 391.180 2342.900 ;
        RECT 391.520 2342.620 391.800 2342.900 ;
        RECT 392.140 2342.620 392.420 2342.900 ;
        RECT 392.760 2342.620 393.040 2342.900 ;
        RECT 389.040 2342.000 389.320 2342.280 ;
        RECT 389.660 2342.000 389.940 2342.280 ;
        RECT 390.280 2342.000 390.560 2342.280 ;
        RECT 390.900 2342.000 391.180 2342.280 ;
        RECT 391.520 2342.000 391.800 2342.280 ;
        RECT 392.140 2342.000 392.420 2342.280 ;
        RECT 392.760 2342.000 393.040 2342.280 ;
        RECT 389.040 2341.380 389.320 2341.660 ;
        RECT 389.660 2341.380 389.940 2341.660 ;
        RECT 390.280 2341.380 390.560 2341.660 ;
        RECT 390.900 2341.380 391.180 2341.660 ;
        RECT 391.520 2341.380 391.800 2341.660 ;
        RECT 392.140 2341.380 392.420 2341.660 ;
        RECT 392.760 2341.380 393.040 2341.660 ;
        RECT 389.040 2340.760 389.320 2341.040 ;
        RECT 389.660 2340.760 389.940 2341.040 ;
        RECT 390.280 2340.760 390.560 2341.040 ;
        RECT 390.900 2340.760 391.180 2341.040 ;
        RECT 391.520 2340.760 391.800 2341.040 ;
        RECT 392.140 2340.760 392.420 2341.040 ;
        RECT 392.760 2340.760 393.040 2341.040 ;
        RECT 389.040 2340.140 389.320 2340.420 ;
        RECT 389.660 2340.140 389.940 2340.420 ;
        RECT 390.280 2340.140 390.560 2340.420 ;
        RECT 390.900 2340.140 391.180 2340.420 ;
        RECT 391.520 2340.140 391.800 2340.420 ;
        RECT 392.140 2340.140 392.420 2340.420 ;
        RECT 392.760 2340.140 393.040 2340.420 ;
        RECT 389.040 2339.520 389.320 2339.800 ;
        RECT 389.660 2339.520 389.940 2339.800 ;
        RECT 390.280 2339.520 390.560 2339.800 ;
        RECT 390.900 2339.520 391.180 2339.800 ;
        RECT 391.520 2339.520 391.800 2339.800 ;
        RECT 392.140 2339.520 392.420 2339.800 ;
        RECT 392.760 2339.520 393.040 2339.800 ;
        RECT 350.370 2335.260 350.650 2335.540 ;
        RECT 350.370 2334.640 350.650 2334.920 ;
        RECT 350.370 2334.020 350.650 2334.300 ;
        RECT 350.370 2333.400 350.650 2333.680 ;
        RECT 350.370 2332.780 350.650 2333.060 ;
        RECT 350.370 2332.160 350.650 2332.440 ;
        RECT 350.370 2331.540 350.650 2331.820 ;
        RECT 350.370 2330.920 350.650 2331.200 ;
        RECT 350.370 2330.300 350.650 2330.580 ;
        RECT 350.370 2329.680 350.650 2329.960 ;
        RECT 350.370 2329.060 350.650 2329.340 ;
        RECT 350.370 2328.440 350.650 2328.720 ;
        RECT 350.370 2327.820 350.650 2328.100 ;
        RECT 350.370 2327.200 350.650 2327.480 ;
        RECT 350.370 2326.580 350.650 2326.860 ;
        RECT 350.370 2325.960 350.650 2326.240 ;
        RECT 389.040 2335.290 389.320 2335.570 ;
        RECT 389.660 2335.290 389.940 2335.570 ;
        RECT 390.280 2335.290 390.560 2335.570 ;
        RECT 390.900 2335.290 391.180 2335.570 ;
        RECT 391.520 2335.290 391.800 2335.570 ;
        RECT 392.140 2335.290 392.420 2335.570 ;
        RECT 392.760 2335.290 393.040 2335.570 ;
        RECT 389.040 2334.670 389.320 2334.950 ;
        RECT 389.660 2334.670 389.940 2334.950 ;
        RECT 390.280 2334.670 390.560 2334.950 ;
        RECT 390.900 2334.670 391.180 2334.950 ;
        RECT 391.520 2334.670 391.800 2334.950 ;
        RECT 392.140 2334.670 392.420 2334.950 ;
        RECT 392.760 2334.670 393.040 2334.950 ;
        RECT 389.040 2334.050 389.320 2334.330 ;
        RECT 389.660 2334.050 389.940 2334.330 ;
        RECT 390.280 2334.050 390.560 2334.330 ;
        RECT 390.900 2334.050 391.180 2334.330 ;
        RECT 391.520 2334.050 391.800 2334.330 ;
        RECT 392.140 2334.050 392.420 2334.330 ;
        RECT 392.760 2334.050 393.040 2334.330 ;
        RECT 389.040 2333.430 389.320 2333.710 ;
        RECT 389.660 2333.430 389.940 2333.710 ;
        RECT 390.280 2333.430 390.560 2333.710 ;
        RECT 390.900 2333.430 391.180 2333.710 ;
        RECT 391.520 2333.430 391.800 2333.710 ;
        RECT 392.140 2333.430 392.420 2333.710 ;
        RECT 392.760 2333.430 393.040 2333.710 ;
        RECT 389.040 2332.810 389.320 2333.090 ;
        RECT 389.660 2332.810 389.940 2333.090 ;
        RECT 390.280 2332.810 390.560 2333.090 ;
        RECT 390.900 2332.810 391.180 2333.090 ;
        RECT 391.520 2332.810 391.800 2333.090 ;
        RECT 392.140 2332.810 392.420 2333.090 ;
        RECT 392.760 2332.810 393.040 2333.090 ;
        RECT 389.040 2332.190 389.320 2332.470 ;
        RECT 389.660 2332.190 389.940 2332.470 ;
        RECT 390.280 2332.190 390.560 2332.470 ;
        RECT 390.900 2332.190 391.180 2332.470 ;
        RECT 391.520 2332.190 391.800 2332.470 ;
        RECT 392.140 2332.190 392.420 2332.470 ;
        RECT 392.760 2332.190 393.040 2332.470 ;
        RECT 389.040 2331.570 389.320 2331.850 ;
        RECT 389.660 2331.570 389.940 2331.850 ;
        RECT 390.280 2331.570 390.560 2331.850 ;
        RECT 390.900 2331.570 391.180 2331.850 ;
        RECT 391.520 2331.570 391.800 2331.850 ;
        RECT 392.140 2331.570 392.420 2331.850 ;
        RECT 392.760 2331.570 393.040 2331.850 ;
        RECT 389.040 2330.950 389.320 2331.230 ;
        RECT 389.660 2330.950 389.940 2331.230 ;
        RECT 390.280 2330.950 390.560 2331.230 ;
        RECT 390.900 2330.950 391.180 2331.230 ;
        RECT 391.520 2330.950 391.800 2331.230 ;
        RECT 392.140 2330.950 392.420 2331.230 ;
        RECT 392.760 2330.950 393.040 2331.230 ;
        RECT 389.040 2330.330 389.320 2330.610 ;
        RECT 389.660 2330.330 389.940 2330.610 ;
        RECT 390.280 2330.330 390.560 2330.610 ;
        RECT 390.900 2330.330 391.180 2330.610 ;
        RECT 391.520 2330.330 391.800 2330.610 ;
        RECT 392.140 2330.330 392.420 2330.610 ;
        RECT 392.760 2330.330 393.040 2330.610 ;
        RECT 389.040 2329.710 389.320 2329.990 ;
        RECT 389.660 2329.710 389.940 2329.990 ;
        RECT 390.280 2329.710 390.560 2329.990 ;
        RECT 390.900 2329.710 391.180 2329.990 ;
        RECT 391.520 2329.710 391.800 2329.990 ;
        RECT 392.140 2329.710 392.420 2329.990 ;
        RECT 392.760 2329.710 393.040 2329.990 ;
        RECT 389.040 2329.090 389.320 2329.370 ;
        RECT 389.660 2329.090 389.940 2329.370 ;
        RECT 390.280 2329.090 390.560 2329.370 ;
        RECT 390.900 2329.090 391.180 2329.370 ;
        RECT 391.520 2329.090 391.800 2329.370 ;
        RECT 392.140 2329.090 392.420 2329.370 ;
        RECT 392.760 2329.090 393.040 2329.370 ;
        RECT 389.040 2328.470 389.320 2328.750 ;
        RECT 389.660 2328.470 389.940 2328.750 ;
        RECT 390.280 2328.470 390.560 2328.750 ;
        RECT 390.900 2328.470 391.180 2328.750 ;
        RECT 391.520 2328.470 391.800 2328.750 ;
        RECT 392.140 2328.470 392.420 2328.750 ;
        RECT 392.760 2328.470 393.040 2328.750 ;
        RECT 389.040 2327.850 389.320 2328.130 ;
        RECT 389.660 2327.850 389.940 2328.130 ;
        RECT 390.280 2327.850 390.560 2328.130 ;
        RECT 390.900 2327.850 391.180 2328.130 ;
        RECT 391.520 2327.850 391.800 2328.130 ;
        RECT 392.140 2327.850 392.420 2328.130 ;
        RECT 392.760 2327.850 393.040 2328.130 ;
        RECT 389.040 2327.230 389.320 2327.510 ;
        RECT 389.660 2327.230 389.940 2327.510 ;
        RECT 390.280 2327.230 390.560 2327.510 ;
        RECT 390.900 2327.230 391.180 2327.510 ;
        RECT 391.520 2327.230 391.800 2327.510 ;
        RECT 392.140 2327.230 392.420 2327.510 ;
        RECT 392.760 2327.230 393.040 2327.510 ;
        RECT 389.040 2326.610 389.320 2326.890 ;
        RECT 389.660 2326.610 389.940 2326.890 ;
        RECT 390.280 2326.610 390.560 2326.890 ;
        RECT 390.900 2326.610 391.180 2326.890 ;
        RECT 391.520 2326.610 391.800 2326.890 ;
        RECT 392.140 2326.610 392.420 2326.890 ;
        RECT 392.760 2326.610 393.040 2326.890 ;
        RECT 389.040 2325.990 389.320 2326.270 ;
        RECT 389.660 2325.990 389.940 2326.270 ;
        RECT 390.280 2325.990 390.560 2326.270 ;
        RECT 390.900 2325.990 391.180 2326.270 ;
        RECT 391.520 2325.990 391.800 2326.270 ;
        RECT 392.140 2325.990 392.420 2326.270 ;
        RECT 392.760 2325.990 393.040 2326.270 ;
        RECT 350.370 2323.410 350.650 2323.690 ;
        RECT 350.370 2322.790 350.650 2323.070 ;
        RECT 350.370 2322.170 350.650 2322.450 ;
        RECT 350.370 2321.550 350.650 2321.830 ;
        RECT 350.370 2320.930 350.650 2321.210 ;
        RECT 350.370 2320.310 350.650 2320.590 ;
        RECT 350.370 2319.690 350.650 2319.970 ;
        RECT 350.370 2319.070 350.650 2319.350 ;
        RECT 350.370 2318.450 350.650 2318.730 ;
        RECT 350.370 2317.830 350.650 2318.110 ;
        RECT 350.370 2317.210 350.650 2317.490 ;
        RECT 350.370 2316.590 350.650 2316.870 ;
        RECT 350.370 2315.970 350.650 2316.250 ;
        RECT 350.370 2315.350 350.650 2315.630 ;
        RECT 350.370 2314.730 350.650 2315.010 ;
        RECT 350.370 2314.110 350.650 2314.390 ;
        RECT 389.040 2323.440 389.320 2323.720 ;
        RECT 389.660 2323.440 389.940 2323.720 ;
        RECT 390.280 2323.440 390.560 2323.720 ;
        RECT 390.900 2323.440 391.180 2323.720 ;
        RECT 391.520 2323.440 391.800 2323.720 ;
        RECT 392.140 2323.440 392.420 2323.720 ;
        RECT 392.760 2323.440 393.040 2323.720 ;
        RECT 389.040 2322.820 389.320 2323.100 ;
        RECT 389.660 2322.820 389.940 2323.100 ;
        RECT 390.280 2322.820 390.560 2323.100 ;
        RECT 390.900 2322.820 391.180 2323.100 ;
        RECT 391.520 2322.820 391.800 2323.100 ;
        RECT 392.140 2322.820 392.420 2323.100 ;
        RECT 392.760 2322.820 393.040 2323.100 ;
        RECT 389.040 2322.200 389.320 2322.480 ;
        RECT 389.660 2322.200 389.940 2322.480 ;
        RECT 390.280 2322.200 390.560 2322.480 ;
        RECT 390.900 2322.200 391.180 2322.480 ;
        RECT 391.520 2322.200 391.800 2322.480 ;
        RECT 392.140 2322.200 392.420 2322.480 ;
        RECT 392.760 2322.200 393.040 2322.480 ;
        RECT 389.040 2321.580 389.320 2321.860 ;
        RECT 389.660 2321.580 389.940 2321.860 ;
        RECT 390.280 2321.580 390.560 2321.860 ;
        RECT 390.900 2321.580 391.180 2321.860 ;
        RECT 391.520 2321.580 391.800 2321.860 ;
        RECT 392.140 2321.580 392.420 2321.860 ;
        RECT 392.760 2321.580 393.040 2321.860 ;
        RECT 389.040 2320.960 389.320 2321.240 ;
        RECT 389.660 2320.960 389.940 2321.240 ;
        RECT 390.280 2320.960 390.560 2321.240 ;
        RECT 390.900 2320.960 391.180 2321.240 ;
        RECT 391.520 2320.960 391.800 2321.240 ;
        RECT 392.140 2320.960 392.420 2321.240 ;
        RECT 392.760 2320.960 393.040 2321.240 ;
        RECT 389.040 2320.340 389.320 2320.620 ;
        RECT 389.660 2320.340 389.940 2320.620 ;
        RECT 390.280 2320.340 390.560 2320.620 ;
        RECT 390.900 2320.340 391.180 2320.620 ;
        RECT 391.520 2320.340 391.800 2320.620 ;
        RECT 392.140 2320.340 392.420 2320.620 ;
        RECT 392.760 2320.340 393.040 2320.620 ;
        RECT 389.040 2319.720 389.320 2320.000 ;
        RECT 389.660 2319.720 389.940 2320.000 ;
        RECT 390.280 2319.720 390.560 2320.000 ;
        RECT 390.900 2319.720 391.180 2320.000 ;
        RECT 391.520 2319.720 391.800 2320.000 ;
        RECT 392.140 2319.720 392.420 2320.000 ;
        RECT 392.760 2319.720 393.040 2320.000 ;
        RECT 389.040 2319.100 389.320 2319.380 ;
        RECT 389.660 2319.100 389.940 2319.380 ;
        RECT 390.280 2319.100 390.560 2319.380 ;
        RECT 390.900 2319.100 391.180 2319.380 ;
        RECT 391.520 2319.100 391.800 2319.380 ;
        RECT 392.140 2319.100 392.420 2319.380 ;
        RECT 392.760 2319.100 393.040 2319.380 ;
        RECT 389.040 2318.480 389.320 2318.760 ;
        RECT 389.660 2318.480 389.940 2318.760 ;
        RECT 390.280 2318.480 390.560 2318.760 ;
        RECT 390.900 2318.480 391.180 2318.760 ;
        RECT 391.520 2318.480 391.800 2318.760 ;
        RECT 392.140 2318.480 392.420 2318.760 ;
        RECT 392.760 2318.480 393.040 2318.760 ;
        RECT 389.040 2317.860 389.320 2318.140 ;
        RECT 389.660 2317.860 389.940 2318.140 ;
        RECT 390.280 2317.860 390.560 2318.140 ;
        RECT 390.900 2317.860 391.180 2318.140 ;
        RECT 391.520 2317.860 391.800 2318.140 ;
        RECT 392.140 2317.860 392.420 2318.140 ;
        RECT 392.760 2317.860 393.040 2318.140 ;
        RECT 389.040 2317.240 389.320 2317.520 ;
        RECT 389.660 2317.240 389.940 2317.520 ;
        RECT 390.280 2317.240 390.560 2317.520 ;
        RECT 390.900 2317.240 391.180 2317.520 ;
        RECT 391.520 2317.240 391.800 2317.520 ;
        RECT 392.140 2317.240 392.420 2317.520 ;
        RECT 392.760 2317.240 393.040 2317.520 ;
        RECT 389.040 2316.620 389.320 2316.900 ;
        RECT 389.660 2316.620 389.940 2316.900 ;
        RECT 390.280 2316.620 390.560 2316.900 ;
        RECT 390.900 2316.620 391.180 2316.900 ;
        RECT 391.520 2316.620 391.800 2316.900 ;
        RECT 392.140 2316.620 392.420 2316.900 ;
        RECT 392.760 2316.620 393.040 2316.900 ;
        RECT 389.040 2316.000 389.320 2316.280 ;
        RECT 389.660 2316.000 389.940 2316.280 ;
        RECT 390.280 2316.000 390.560 2316.280 ;
        RECT 390.900 2316.000 391.180 2316.280 ;
        RECT 391.520 2316.000 391.800 2316.280 ;
        RECT 392.140 2316.000 392.420 2316.280 ;
        RECT 392.760 2316.000 393.040 2316.280 ;
        RECT 389.040 2315.380 389.320 2315.660 ;
        RECT 389.660 2315.380 389.940 2315.660 ;
        RECT 390.280 2315.380 390.560 2315.660 ;
        RECT 390.900 2315.380 391.180 2315.660 ;
        RECT 391.520 2315.380 391.800 2315.660 ;
        RECT 392.140 2315.380 392.420 2315.660 ;
        RECT 392.760 2315.380 393.040 2315.660 ;
        RECT 389.040 2314.760 389.320 2315.040 ;
        RECT 389.660 2314.760 389.940 2315.040 ;
        RECT 390.280 2314.760 390.560 2315.040 ;
        RECT 390.900 2314.760 391.180 2315.040 ;
        RECT 391.520 2314.760 391.800 2315.040 ;
        RECT 392.140 2314.760 392.420 2315.040 ;
        RECT 392.760 2314.760 393.040 2315.040 ;
        RECT 389.040 2314.140 389.320 2314.420 ;
        RECT 389.660 2314.140 389.940 2314.420 ;
        RECT 390.280 2314.140 390.560 2314.420 ;
        RECT 390.900 2314.140 391.180 2314.420 ;
        RECT 391.520 2314.140 391.800 2314.420 ;
        RECT 392.140 2314.140 392.420 2314.420 ;
        RECT 392.760 2314.140 393.040 2314.420 ;
        RECT 350.370 2310.390 350.650 2310.670 ;
        RECT 350.370 2309.770 350.650 2310.050 ;
        RECT 350.370 2309.150 350.650 2309.430 ;
        RECT 350.370 2308.530 350.650 2308.810 ;
        RECT 350.370 2307.910 350.650 2308.190 ;
        RECT 350.370 2307.290 350.650 2307.570 ;
        RECT 350.370 2306.670 350.650 2306.950 ;
        RECT 350.370 2306.050 350.650 2306.330 ;
        RECT 350.370 2305.430 350.650 2305.710 ;
        RECT 350.370 2304.810 350.650 2305.090 ;
        RECT 350.370 2304.190 350.650 2304.470 ;
        RECT 350.370 2303.570 350.650 2303.850 ;
        RECT 350.370 2302.950 350.650 2303.230 ;
        RECT 350.370 2302.330 350.650 2302.610 ;
        RECT 350.370 2301.710 350.650 2301.990 ;
        RECT 389.040 2310.420 389.320 2310.700 ;
        RECT 389.660 2310.420 389.940 2310.700 ;
        RECT 390.280 2310.420 390.560 2310.700 ;
        RECT 390.900 2310.420 391.180 2310.700 ;
        RECT 391.520 2310.420 391.800 2310.700 ;
        RECT 392.140 2310.420 392.420 2310.700 ;
        RECT 392.760 2310.420 393.040 2310.700 ;
        RECT 389.040 2309.800 389.320 2310.080 ;
        RECT 389.660 2309.800 389.940 2310.080 ;
        RECT 390.280 2309.800 390.560 2310.080 ;
        RECT 390.900 2309.800 391.180 2310.080 ;
        RECT 391.520 2309.800 391.800 2310.080 ;
        RECT 392.140 2309.800 392.420 2310.080 ;
        RECT 392.760 2309.800 393.040 2310.080 ;
        RECT 389.040 2309.180 389.320 2309.460 ;
        RECT 389.660 2309.180 389.940 2309.460 ;
        RECT 390.280 2309.180 390.560 2309.460 ;
        RECT 390.900 2309.180 391.180 2309.460 ;
        RECT 391.520 2309.180 391.800 2309.460 ;
        RECT 392.140 2309.180 392.420 2309.460 ;
        RECT 392.760 2309.180 393.040 2309.460 ;
        RECT 389.040 2308.560 389.320 2308.840 ;
        RECT 389.660 2308.560 389.940 2308.840 ;
        RECT 390.280 2308.560 390.560 2308.840 ;
        RECT 390.900 2308.560 391.180 2308.840 ;
        RECT 391.520 2308.560 391.800 2308.840 ;
        RECT 392.140 2308.560 392.420 2308.840 ;
        RECT 392.760 2308.560 393.040 2308.840 ;
        RECT 389.040 2307.940 389.320 2308.220 ;
        RECT 389.660 2307.940 389.940 2308.220 ;
        RECT 390.280 2307.940 390.560 2308.220 ;
        RECT 390.900 2307.940 391.180 2308.220 ;
        RECT 391.520 2307.940 391.800 2308.220 ;
        RECT 392.140 2307.940 392.420 2308.220 ;
        RECT 392.760 2307.940 393.040 2308.220 ;
        RECT 389.040 2307.320 389.320 2307.600 ;
        RECT 389.660 2307.320 389.940 2307.600 ;
        RECT 390.280 2307.320 390.560 2307.600 ;
        RECT 390.900 2307.320 391.180 2307.600 ;
        RECT 391.520 2307.320 391.800 2307.600 ;
        RECT 392.140 2307.320 392.420 2307.600 ;
        RECT 392.760 2307.320 393.040 2307.600 ;
        RECT 389.040 2306.700 389.320 2306.980 ;
        RECT 389.660 2306.700 389.940 2306.980 ;
        RECT 390.280 2306.700 390.560 2306.980 ;
        RECT 390.900 2306.700 391.180 2306.980 ;
        RECT 391.520 2306.700 391.800 2306.980 ;
        RECT 392.140 2306.700 392.420 2306.980 ;
        RECT 392.760 2306.700 393.040 2306.980 ;
        RECT 389.040 2306.080 389.320 2306.360 ;
        RECT 389.660 2306.080 389.940 2306.360 ;
        RECT 390.280 2306.080 390.560 2306.360 ;
        RECT 390.900 2306.080 391.180 2306.360 ;
        RECT 391.520 2306.080 391.800 2306.360 ;
        RECT 392.140 2306.080 392.420 2306.360 ;
        RECT 392.760 2306.080 393.040 2306.360 ;
        RECT 389.040 2305.460 389.320 2305.740 ;
        RECT 389.660 2305.460 389.940 2305.740 ;
        RECT 390.280 2305.460 390.560 2305.740 ;
        RECT 390.900 2305.460 391.180 2305.740 ;
        RECT 391.520 2305.460 391.800 2305.740 ;
        RECT 392.140 2305.460 392.420 2305.740 ;
        RECT 392.760 2305.460 393.040 2305.740 ;
        RECT 389.040 2304.840 389.320 2305.120 ;
        RECT 389.660 2304.840 389.940 2305.120 ;
        RECT 390.280 2304.840 390.560 2305.120 ;
        RECT 390.900 2304.840 391.180 2305.120 ;
        RECT 391.520 2304.840 391.800 2305.120 ;
        RECT 392.140 2304.840 392.420 2305.120 ;
        RECT 392.760 2304.840 393.040 2305.120 ;
        RECT 389.040 2304.220 389.320 2304.500 ;
        RECT 389.660 2304.220 389.940 2304.500 ;
        RECT 390.280 2304.220 390.560 2304.500 ;
        RECT 390.900 2304.220 391.180 2304.500 ;
        RECT 391.520 2304.220 391.800 2304.500 ;
        RECT 392.140 2304.220 392.420 2304.500 ;
        RECT 392.760 2304.220 393.040 2304.500 ;
        RECT 389.040 2303.600 389.320 2303.880 ;
        RECT 389.660 2303.600 389.940 2303.880 ;
        RECT 390.280 2303.600 390.560 2303.880 ;
        RECT 390.900 2303.600 391.180 2303.880 ;
        RECT 391.520 2303.600 391.800 2303.880 ;
        RECT 392.140 2303.600 392.420 2303.880 ;
        RECT 392.760 2303.600 393.040 2303.880 ;
        RECT 389.040 2302.980 389.320 2303.260 ;
        RECT 389.660 2302.980 389.940 2303.260 ;
        RECT 390.280 2302.980 390.560 2303.260 ;
        RECT 390.900 2302.980 391.180 2303.260 ;
        RECT 391.520 2302.980 391.800 2303.260 ;
        RECT 392.140 2302.980 392.420 2303.260 ;
        RECT 392.760 2302.980 393.040 2303.260 ;
        RECT 389.040 2302.360 389.320 2302.640 ;
        RECT 389.660 2302.360 389.940 2302.640 ;
        RECT 390.280 2302.360 390.560 2302.640 ;
        RECT 390.900 2302.360 391.180 2302.640 ;
        RECT 391.520 2302.360 391.800 2302.640 ;
        RECT 392.140 2302.360 392.420 2302.640 ;
        RECT 392.760 2302.360 393.040 2302.640 ;
        RECT 389.040 2301.740 389.320 2302.020 ;
        RECT 389.660 2301.740 389.940 2302.020 ;
        RECT 390.280 2301.740 390.560 2302.020 ;
        RECT 390.900 2301.740 391.180 2302.020 ;
        RECT 391.520 2301.740 391.800 2302.020 ;
        RECT 392.140 2301.740 392.420 2302.020 ;
        RECT 392.760 2301.740 393.040 2302.020 ;
        RECT 388.740 2232.670 389.020 2232.950 ;
        RECT 389.360 2232.670 389.640 2232.950 ;
        RECT 389.980 2232.670 390.260 2232.950 ;
        RECT 390.600 2232.670 390.880 2232.950 ;
        RECT 391.220 2232.670 391.500 2232.950 ;
        RECT 391.840 2232.670 392.120 2232.950 ;
        RECT 392.460 2232.670 392.740 2232.950 ;
        RECT 388.740 2232.050 389.020 2232.330 ;
        RECT 389.360 2232.050 389.640 2232.330 ;
        RECT 389.980 2232.050 390.260 2232.330 ;
        RECT 390.600 2232.050 390.880 2232.330 ;
        RECT 391.220 2232.050 391.500 2232.330 ;
        RECT 391.840 2232.050 392.120 2232.330 ;
        RECT 392.460 2232.050 392.740 2232.330 ;
        RECT 388.740 2231.430 389.020 2231.710 ;
        RECT 389.360 2231.430 389.640 2231.710 ;
        RECT 389.980 2231.430 390.260 2231.710 ;
        RECT 390.600 2231.430 390.880 2231.710 ;
        RECT 391.220 2231.430 391.500 2231.710 ;
        RECT 391.840 2231.430 392.120 2231.710 ;
        RECT 392.460 2231.430 392.740 2231.710 ;
        RECT 388.740 2230.810 389.020 2231.090 ;
        RECT 389.360 2230.810 389.640 2231.090 ;
        RECT 389.980 2230.810 390.260 2231.090 ;
        RECT 390.600 2230.810 390.880 2231.090 ;
        RECT 391.220 2230.810 391.500 2231.090 ;
        RECT 391.840 2230.810 392.120 2231.090 ;
        RECT 392.460 2230.810 392.740 2231.090 ;
        RECT 388.740 2230.190 389.020 2230.470 ;
        RECT 389.360 2230.190 389.640 2230.470 ;
        RECT 389.980 2230.190 390.260 2230.470 ;
        RECT 390.600 2230.190 390.880 2230.470 ;
        RECT 391.220 2230.190 391.500 2230.470 ;
        RECT 391.840 2230.190 392.120 2230.470 ;
        RECT 392.460 2230.190 392.740 2230.470 ;
        RECT 350.370 2168.010 350.650 2168.290 ;
        RECT 350.370 2167.390 350.650 2167.670 ;
        RECT 350.370 2166.770 350.650 2167.050 ;
        RECT 350.370 2166.150 350.650 2166.430 ;
        RECT 350.370 2165.530 350.650 2165.810 ;
        RECT 350.370 2164.910 350.650 2165.190 ;
        RECT 350.370 2164.290 350.650 2164.570 ;
        RECT 350.370 2163.670 350.650 2163.950 ;
        RECT 350.370 2163.050 350.650 2163.330 ;
        RECT 350.370 2162.430 350.650 2162.710 ;
        RECT 350.370 2161.810 350.650 2162.090 ;
        RECT 350.370 2161.190 350.650 2161.470 ;
        RECT 350.370 2160.570 350.650 2160.850 ;
        RECT 350.370 2159.950 350.650 2160.230 ;
        RECT 350.370 2159.330 350.650 2159.610 ;
        RECT 350.370 2155.640 350.650 2155.920 ;
        RECT 350.370 2155.020 350.650 2155.300 ;
        RECT 350.370 2154.400 350.650 2154.680 ;
        RECT 350.370 2153.780 350.650 2154.060 ;
        RECT 350.370 2153.160 350.650 2153.440 ;
        RECT 350.370 2152.540 350.650 2152.820 ;
        RECT 350.370 2151.920 350.650 2152.200 ;
        RECT 350.370 2151.300 350.650 2151.580 ;
        RECT 350.370 2150.680 350.650 2150.960 ;
        RECT 350.370 2150.060 350.650 2150.340 ;
        RECT 350.370 2149.440 350.650 2149.720 ;
        RECT 350.370 2148.820 350.650 2149.100 ;
        RECT 350.370 2148.200 350.650 2148.480 ;
        RECT 350.370 2147.580 350.650 2147.860 ;
        RECT 350.370 2146.960 350.650 2147.240 ;
        RECT 350.370 2146.340 350.650 2146.620 ;
        RECT 350.370 2143.790 350.650 2144.070 ;
        RECT 350.370 2143.170 350.650 2143.450 ;
        RECT 350.370 2142.550 350.650 2142.830 ;
        RECT 350.370 2141.930 350.650 2142.210 ;
        RECT 350.370 2141.310 350.650 2141.590 ;
        RECT 350.370 2140.690 350.650 2140.970 ;
        RECT 350.370 2140.070 350.650 2140.350 ;
        RECT 350.370 2139.450 350.650 2139.730 ;
        RECT 350.370 2138.830 350.650 2139.110 ;
        RECT 350.370 2138.210 350.650 2138.490 ;
        RECT 350.370 2137.590 350.650 2137.870 ;
        RECT 350.370 2136.970 350.650 2137.250 ;
        RECT 350.370 2136.350 350.650 2136.630 ;
        RECT 350.370 2135.730 350.650 2136.010 ;
        RECT 350.370 2135.110 350.650 2135.390 ;
        RECT 350.370 2134.490 350.650 2134.770 ;
        RECT 350.370 2130.260 350.650 2130.540 ;
        RECT 350.370 2129.640 350.650 2129.920 ;
        RECT 350.370 2129.020 350.650 2129.300 ;
        RECT 350.370 2128.400 350.650 2128.680 ;
        RECT 350.370 2127.780 350.650 2128.060 ;
        RECT 350.370 2127.160 350.650 2127.440 ;
        RECT 350.370 2126.540 350.650 2126.820 ;
        RECT 350.370 2125.920 350.650 2126.200 ;
        RECT 350.370 2125.300 350.650 2125.580 ;
        RECT 350.370 2124.680 350.650 2124.960 ;
        RECT 350.370 2124.060 350.650 2124.340 ;
        RECT 350.370 2123.440 350.650 2123.720 ;
        RECT 350.370 2122.820 350.650 2123.100 ;
        RECT 350.370 2122.200 350.650 2122.480 ;
        RECT 350.370 2121.580 350.650 2121.860 ;
        RECT 350.370 2120.960 350.650 2121.240 ;
        RECT 350.370 2118.410 350.650 2118.690 ;
        RECT 350.370 2117.790 350.650 2118.070 ;
        RECT 350.370 2117.170 350.650 2117.450 ;
        RECT 350.370 2116.550 350.650 2116.830 ;
        RECT 350.370 2115.930 350.650 2116.210 ;
        RECT 350.370 2115.310 350.650 2115.590 ;
        RECT 350.370 2114.690 350.650 2114.970 ;
        RECT 350.370 2114.070 350.650 2114.350 ;
        RECT 350.370 2113.450 350.650 2113.730 ;
        RECT 350.370 2112.830 350.650 2113.110 ;
        RECT 350.370 2112.210 350.650 2112.490 ;
        RECT 350.370 2111.590 350.650 2111.870 ;
        RECT 350.370 2110.970 350.650 2111.250 ;
        RECT 350.370 2110.350 350.650 2110.630 ;
        RECT 350.370 2109.730 350.650 2110.010 ;
        RECT 350.370 2109.110 350.650 2109.390 ;
        RECT 350.370 2105.390 350.650 2105.670 ;
        RECT 350.370 2104.770 350.650 2105.050 ;
        RECT 350.370 2104.150 350.650 2104.430 ;
        RECT 350.370 2103.530 350.650 2103.810 ;
        RECT 350.370 2102.910 350.650 2103.190 ;
        RECT 350.370 2102.290 350.650 2102.570 ;
        RECT 350.370 2101.670 350.650 2101.950 ;
        RECT 350.370 2101.050 350.650 2101.330 ;
        RECT 350.370 2100.430 350.650 2100.710 ;
        RECT 350.370 2099.810 350.650 2100.090 ;
        RECT 350.370 2099.190 350.650 2099.470 ;
        RECT 350.370 2098.570 350.650 2098.850 ;
        RECT 350.370 2097.950 350.650 2098.230 ;
        RECT 350.370 2097.330 350.650 2097.610 ;
        RECT 350.370 2096.710 350.650 2096.990 ;
        RECT 389.235 2062.885 389.515 2063.165 ;
        RECT 390.735 2062.885 391.015 2063.165 ;
        RECT 392.235 2062.885 392.515 2063.165 ;
        RECT 389.000 2051.865 389.280 2052.145 ;
        RECT 390.500 2051.865 390.780 2052.145 ;
        RECT 392.000 2051.865 392.280 2052.145 ;
        RECT 389.000 2050.865 389.280 2051.145 ;
        RECT 390.500 2050.865 390.780 2051.145 ;
        RECT 392.000 2050.865 392.280 2051.145 ;
        RECT 389.500 1965.230 389.780 1965.510 ;
        RECT 391.000 1965.230 391.280 1965.510 ;
        RECT 392.500 1965.230 392.780 1965.510 ;
        RECT 389.500 1930.230 389.780 1930.510 ;
        RECT 391.000 1930.230 391.280 1930.510 ;
        RECT 392.500 1930.230 392.780 1930.510 ;
        RECT 389.500 1895.230 389.780 1895.510 ;
        RECT 391.000 1895.230 391.280 1895.510 ;
        RECT 392.500 1895.230 392.780 1895.510 ;
        RECT 389.000 1871.865 389.280 1872.145 ;
        RECT 390.500 1871.865 390.780 1872.145 ;
        RECT 392.000 1871.865 392.280 1872.145 ;
        RECT 389.000 1870.865 389.280 1871.145 ;
        RECT 390.500 1870.865 390.780 1871.145 ;
        RECT 392.000 1870.865 392.280 1871.145 ;
        RECT 389.235 1857.885 389.515 1858.165 ;
        RECT 390.735 1857.885 391.015 1858.165 ;
        RECT 392.235 1857.885 392.515 1858.165 ;
        RECT 389.500 1760.230 389.780 1760.510 ;
        RECT 391.000 1760.230 391.280 1760.510 ;
        RECT 392.500 1760.230 392.780 1760.510 ;
        RECT 389.500 1725.230 389.780 1725.510 ;
        RECT 391.000 1725.230 391.280 1725.510 ;
        RECT 392.500 1725.230 392.780 1725.510 ;
        RECT 389.000 1691.865 389.280 1692.145 ;
        RECT 390.500 1691.865 390.780 1692.145 ;
        RECT 392.000 1691.865 392.280 1692.145 ;
        RECT 389.000 1690.865 389.280 1691.145 ;
        RECT 390.500 1690.865 390.780 1691.145 ;
        RECT 392.000 1690.865 392.280 1691.145 ;
        RECT 389.500 1690.230 389.780 1690.510 ;
        RECT 391.000 1690.230 391.280 1690.510 ;
        RECT 392.500 1690.230 392.780 1690.510 ;
        RECT 389.235 1652.885 389.515 1653.165 ;
        RECT 390.735 1652.885 391.015 1653.165 ;
        RECT 392.235 1652.885 392.515 1653.165 ;
        RECT 389.040 1647.920 389.320 1648.200 ;
        RECT 389.660 1647.920 389.940 1648.200 ;
        RECT 390.280 1647.920 390.560 1648.200 ;
        RECT 390.900 1647.920 391.180 1648.200 ;
        RECT 391.520 1647.920 391.800 1648.200 ;
        RECT 392.140 1647.920 392.420 1648.200 ;
        RECT 392.760 1647.920 393.040 1648.200 ;
        RECT 389.040 1647.300 389.320 1647.580 ;
        RECT 389.660 1647.300 389.940 1647.580 ;
        RECT 390.280 1647.300 390.560 1647.580 ;
        RECT 390.900 1647.300 391.180 1647.580 ;
        RECT 391.520 1647.300 391.800 1647.580 ;
        RECT 392.140 1647.300 392.420 1647.580 ;
        RECT 392.760 1647.300 393.040 1647.580 ;
        RECT 389.040 1646.680 389.320 1646.960 ;
        RECT 389.660 1646.680 389.940 1646.960 ;
        RECT 390.280 1646.680 390.560 1646.960 ;
        RECT 390.900 1646.680 391.180 1646.960 ;
        RECT 391.520 1646.680 391.800 1646.960 ;
        RECT 392.140 1646.680 392.420 1646.960 ;
        RECT 392.760 1646.680 393.040 1646.960 ;
        RECT 389.040 1646.060 389.320 1646.340 ;
        RECT 389.660 1646.060 389.940 1646.340 ;
        RECT 390.280 1646.060 390.560 1646.340 ;
        RECT 390.900 1646.060 391.180 1646.340 ;
        RECT 391.520 1646.060 391.800 1646.340 ;
        RECT 392.140 1646.060 392.420 1646.340 ;
        RECT 392.760 1646.060 393.040 1646.340 ;
        RECT 389.040 1645.440 389.320 1645.720 ;
        RECT 389.660 1645.440 389.940 1645.720 ;
        RECT 390.280 1645.440 390.560 1645.720 ;
        RECT 390.900 1645.440 391.180 1645.720 ;
        RECT 391.520 1645.440 391.800 1645.720 ;
        RECT 392.140 1645.440 392.420 1645.720 ;
        RECT 392.760 1645.440 393.040 1645.720 ;
        RECT 389.040 1644.820 389.320 1645.100 ;
        RECT 389.660 1644.820 389.940 1645.100 ;
        RECT 390.280 1644.820 390.560 1645.100 ;
        RECT 390.900 1644.820 391.180 1645.100 ;
        RECT 391.520 1644.820 391.800 1645.100 ;
        RECT 392.140 1644.820 392.420 1645.100 ;
        RECT 392.760 1644.820 393.040 1645.100 ;
        RECT 389.040 1644.200 389.320 1644.480 ;
        RECT 389.660 1644.200 389.940 1644.480 ;
        RECT 390.280 1644.200 390.560 1644.480 ;
        RECT 390.900 1644.200 391.180 1644.480 ;
        RECT 391.520 1644.200 391.800 1644.480 ;
        RECT 392.140 1644.200 392.420 1644.480 ;
        RECT 392.760 1644.200 393.040 1644.480 ;
        RECT 389.500 1555.230 389.780 1555.510 ;
        RECT 391.000 1555.230 391.280 1555.510 ;
        RECT 392.500 1555.230 392.780 1555.510 ;
        RECT 389.040 1528.650 389.320 1528.930 ;
        RECT 389.660 1528.650 389.940 1528.930 ;
        RECT 390.280 1528.650 390.560 1528.930 ;
        RECT 390.900 1528.650 391.180 1528.930 ;
        RECT 391.520 1528.650 391.800 1528.930 ;
        RECT 392.140 1528.650 392.420 1528.930 ;
        RECT 392.760 1528.650 393.040 1528.930 ;
        RECT 389.040 1528.030 389.320 1528.310 ;
        RECT 389.660 1528.030 389.940 1528.310 ;
        RECT 390.280 1528.030 390.560 1528.310 ;
        RECT 390.900 1528.030 391.180 1528.310 ;
        RECT 391.520 1528.030 391.800 1528.310 ;
        RECT 392.140 1528.030 392.420 1528.310 ;
        RECT 392.760 1528.030 393.040 1528.310 ;
        RECT 389.040 1527.410 389.320 1527.690 ;
        RECT 389.660 1527.410 389.940 1527.690 ;
        RECT 390.280 1527.410 390.560 1527.690 ;
        RECT 390.900 1527.410 391.180 1527.690 ;
        RECT 391.520 1527.410 391.800 1527.690 ;
        RECT 392.140 1527.410 392.420 1527.690 ;
        RECT 392.760 1527.410 393.040 1527.690 ;
        RECT 389.040 1526.790 389.320 1527.070 ;
        RECT 389.660 1526.790 389.940 1527.070 ;
        RECT 390.280 1526.790 390.560 1527.070 ;
        RECT 390.900 1526.790 391.180 1527.070 ;
        RECT 391.520 1526.790 391.800 1527.070 ;
        RECT 392.140 1526.790 392.420 1527.070 ;
        RECT 392.760 1526.790 393.040 1527.070 ;
        RECT 389.040 1526.170 389.320 1526.450 ;
        RECT 389.660 1526.170 389.940 1526.450 ;
        RECT 390.280 1526.170 390.560 1526.450 ;
        RECT 390.900 1526.170 391.180 1526.450 ;
        RECT 391.520 1526.170 391.800 1526.450 ;
        RECT 392.140 1526.170 392.420 1526.450 ;
        RECT 392.760 1526.170 393.040 1526.450 ;
        RECT 389.040 1525.550 389.320 1525.830 ;
        RECT 389.660 1525.550 389.940 1525.830 ;
        RECT 390.280 1525.550 390.560 1525.830 ;
        RECT 390.900 1525.550 391.180 1525.830 ;
        RECT 391.520 1525.550 391.800 1525.830 ;
        RECT 392.140 1525.550 392.420 1525.830 ;
        RECT 392.760 1525.550 393.040 1525.830 ;
        RECT 389.040 1524.930 389.320 1525.210 ;
        RECT 389.660 1524.930 389.940 1525.210 ;
        RECT 390.280 1524.930 390.560 1525.210 ;
        RECT 390.900 1524.930 391.180 1525.210 ;
        RECT 391.520 1524.930 391.800 1525.210 ;
        RECT 392.140 1524.930 392.420 1525.210 ;
        RECT 392.760 1524.930 393.040 1525.210 ;
        RECT 389.000 1520.330 389.280 1520.610 ;
        RECT 390.500 1520.330 390.780 1520.610 ;
        RECT 392.000 1520.330 392.280 1520.610 ;
        RECT 389.500 1485.230 389.780 1485.510 ;
        RECT 391.000 1485.230 391.280 1485.510 ;
        RECT 392.500 1485.230 392.780 1485.510 ;
        RECT 389.235 1447.885 389.515 1448.165 ;
        RECT 390.735 1447.885 391.015 1448.165 ;
        RECT 392.235 1447.885 392.515 1448.165 ;
        RECT 389.040 1409.580 389.320 1409.860 ;
        RECT 389.660 1409.580 389.940 1409.860 ;
        RECT 390.280 1409.580 390.560 1409.860 ;
        RECT 390.900 1409.580 391.180 1409.860 ;
        RECT 391.520 1409.580 391.800 1409.860 ;
        RECT 392.140 1409.580 392.420 1409.860 ;
        RECT 392.760 1409.580 393.040 1409.860 ;
        RECT 389.040 1408.960 389.320 1409.240 ;
        RECT 389.660 1408.960 389.940 1409.240 ;
        RECT 390.280 1408.960 390.560 1409.240 ;
        RECT 390.900 1408.960 391.180 1409.240 ;
        RECT 391.520 1408.960 391.800 1409.240 ;
        RECT 392.140 1408.960 392.420 1409.240 ;
        RECT 392.760 1408.960 393.040 1409.240 ;
        RECT 389.040 1408.340 389.320 1408.620 ;
        RECT 389.660 1408.340 389.940 1408.620 ;
        RECT 390.280 1408.340 390.560 1408.620 ;
        RECT 390.900 1408.340 391.180 1408.620 ;
        RECT 391.520 1408.340 391.800 1408.620 ;
        RECT 392.140 1408.340 392.420 1408.620 ;
        RECT 392.760 1408.340 393.040 1408.620 ;
        RECT 389.040 1407.720 389.320 1408.000 ;
        RECT 389.660 1407.720 389.940 1408.000 ;
        RECT 390.280 1407.720 390.560 1408.000 ;
        RECT 390.900 1407.720 391.180 1408.000 ;
        RECT 391.520 1407.720 391.800 1408.000 ;
        RECT 392.140 1407.720 392.420 1408.000 ;
        RECT 392.760 1407.720 393.040 1408.000 ;
        RECT 389.040 1407.100 389.320 1407.380 ;
        RECT 389.660 1407.100 389.940 1407.380 ;
        RECT 390.280 1407.100 390.560 1407.380 ;
        RECT 390.900 1407.100 391.180 1407.380 ;
        RECT 391.520 1407.100 391.800 1407.380 ;
        RECT 392.140 1407.100 392.420 1407.380 ;
        RECT 392.760 1407.100 393.040 1407.380 ;
        RECT 389.040 1406.480 389.320 1406.760 ;
        RECT 389.660 1406.480 389.940 1406.760 ;
        RECT 390.280 1406.480 390.560 1406.760 ;
        RECT 390.900 1406.480 391.180 1406.760 ;
        RECT 391.520 1406.480 391.800 1406.760 ;
        RECT 392.140 1406.480 392.420 1406.760 ;
        RECT 392.760 1406.480 393.040 1406.760 ;
        RECT 389.040 1405.860 389.320 1406.140 ;
        RECT 389.660 1405.860 389.940 1406.140 ;
        RECT 390.280 1405.860 390.560 1406.140 ;
        RECT 390.900 1405.860 391.180 1406.140 ;
        RECT 391.520 1405.860 391.800 1406.140 ;
        RECT 392.140 1405.860 392.420 1406.140 ;
        RECT 392.760 1405.860 393.040 1406.140 ;
        RECT 389.500 1350.230 389.780 1350.510 ;
        RECT 391.000 1350.230 391.280 1350.510 ;
        RECT 392.500 1350.230 392.780 1350.510 ;
        RECT 388.740 1341.580 389.020 1341.860 ;
        RECT 389.360 1341.580 389.640 1341.860 ;
        RECT 389.980 1341.580 390.260 1341.860 ;
        RECT 390.600 1341.580 390.880 1341.860 ;
        RECT 391.220 1341.580 391.500 1341.860 ;
        RECT 391.840 1341.580 392.120 1341.860 ;
        RECT 392.460 1341.580 392.740 1341.860 ;
        RECT 388.740 1340.960 389.020 1341.240 ;
        RECT 389.360 1340.960 389.640 1341.240 ;
        RECT 389.980 1340.960 390.260 1341.240 ;
        RECT 390.600 1340.960 390.880 1341.240 ;
        RECT 391.220 1340.960 391.500 1341.240 ;
        RECT 391.840 1340.960 392.120 1341.240 ;
        RECT 392.460 1340.960 392.740 1341.240 ;
        RECT 389.500 1315.230 389.780 1315.510 ;
        RECT 391.000 1315.230 391.280 1315.510 ;
        RECT 392.500 1315.230 392.780 1315.510 ;
        RECT 389.500 1280.230 389.780 1280.510 ;
        RECT 391.000 1280.230 391.280 1280.510 ;
        RECT 392.500 1280.230 392.780 1280.510 ;
        RECT 389.235 1242.885 389.515 1243.165 ;
        RECT 390.735 1242.885 391.015 1243.165 ;
        RECT 392.235 1242.885 392.515 1243.165 ;
        RECT 388.740 1211.580 389.020 1211.860 ;
        RECT 389.360 1211.580 389.640 1211.860 ;
        RECT 389.980 1211.580 390.260 1211.860 ;
        RECT 390.600 1211.580 390.880 1211.860 ;
        RECT 391.220 1211.580 391.500 1211.860 ;
        RECT 391.840 1211.580 392.120 1211.860 ;
        RECT 392.460 1211.580 392.740 1211.860 ;
        RECT 388.740 1210.960 389.020 1211.240 ;
        RECT 389.360 1210.960 389.640 1211.240 ;
        RECT 389.980 1210.960 390.260 1211.240 ;
        RECT 390.600 1210.960 390.880 1211.240 ;
        RECT 391.220 1210.960 391.500 1211.240 ;
        RECT 391.840 1210.960 392.120 1211.240 ;
        RECT 392.460 1210.960 392.740 1211.240 ;
        RECT 389.500 1145.230 389.780 1145.510 ;
        RECT 391.000 1145.230 391.280 1145.510 ;
        RECT 392.500 1145.230 392.780 1145.510 ;
        RECT 389.500 1110.230 389.780 1110.510 ;
        RECT 391.000 1110.230 391.280 1110.510 ;
        RECT 392.500 1110.230 392.780 1110.510 ;
        RECT 388.740 1081.580 389.020 1081.860 ;
        RECT 389.360 1081.580 389.640 1081.860 ;
        RECT 389.980 1081.580 390.260 1081.860 ;
        RECT 390.600 1081.580 390.880 1081.860 ;
        RECT 391.220 1081.580 391.500 1081.860 ;
        RECT 391.840 1081.580 392.120 1081.860 ;
        RECT 392.460 1081.580 392.740 1081.860 ;
        RECT 388.740 1080.960 389.020 1081.240 ;
        RECT 389.360 1080.960 389.640 1081.240 ;
        RECT 389.980 1080.960 390.260 1081.240 ;
        RECT 390.600 1080.960 390.880 1081.240 ;
        RECT 391.220 1080.960 391.500 1081.240 ;
        RECT 391.840 1080.960 392.120 1081.240 ;
        RECT 392.460 1080.960 392.740 1081.240 ;
        RECT 389.500 1075.230 389.780 1075.510 ;
        RECT 391.000 1075.230 391.280 1075.510 ;
        RECT 392.500 1075.230 392.780 1075.510 ;
        RECT 389.235 1037.885 389.515 1038.165 ;
        RECT 390.735 1037.885 391.015 1038.165 ;
        RECT 392.235 1037.885 392.515 1038.165 ;
        RECT 388.740 951.580 389.020 951.860 ;
        RECT 389.360 951.580 389.640 951.860 ;
        RECT 389.980 951.580 390.260 951.860 ;
        RECT 390.600 951.580 390.880 951.860 ;
        RECT 391.220 951.580 391.500 951.860 ;
        RECT 391.840 951.580 392.120 951.860 ;
        RECT 392.460 951.580 392.740 951.860 ;
        RECT 388.740 950.960 389.020 951.240 ;
        RECT 389.360 950.960 389.640 951.240 ;
        RECT 389.980 950.960 390.260 951.240 ;
        RECT 390.600 950.960 390.880 951.240 ;
        RECT 391.220 950.960 391.500 951.240 ;
        RECT 391.840 950.960 392.120 951.240 ;
        RECT 392.460 950.960 392.740 951.240 ;
        RECT 389.500 940.230 389.780 940.510 ;
        RECT 391.000 940.230 391.280 940.510 ;
        RECT 392.500 940.230 392.780 940.510 ;
        RECT 389.500 905.230 389.780 905.510 ;
        RECT 391.000 905.230 391.280 905.510 ;
        RECT 392.500 905.230 392.780 905.510 ;
        RECT 389.500 870.230 389.780 870.510 ;
        RECT 391.000 870.230 391.280 870.510 ;
        RECT 392.500 870.230 392.780 870.510 ;
        RECT 388.740 821.580 389.020 821.860 ;
        RECT 389.360 821.580 389.640 821.860 ;
        RECT 389.980 821.580 390.260 821.860 ;
        RECT 390.600 821.580 390.880 821.860 ;
        RECT 391.220 821.580 391.500 821.860 ;
        RECT 391.840 821.580 392.120 821.860 ;
        RECT 392.460 821.580 392.740 821.860 ;
        RECT 388.740 820.960 389.020 821.240 ;
        RECT 389.360 820.960 389.640 821.240 ;
        RECT 389.980 820.960 390.260 821.240 ;
        RECT 390.600 820.960 390.880 821.240 ;
        RECT 391.220 820.960 391.500 821.240 ;
        RECT 391.840 820.960 392.120 821.240 ;
        RECT 392.460 820.960 392.740 821.240 ;
        RECT 350.370 733.010 350.650 733.290 ;
        RECT 350.370 732.390 350.650 732.670 ;
        RECT 350.370 731.770 350.650 732.050 ;
        RECT 350.370 731.150 350.650 731.430 ;
        RECT 350.370 730.530 350.650 730.810 ;
        RECT 350.370 729.910 350.650 730.190 ;
        RECT 350.370 729.290 350.650 729.570 ;
        RECT 350.370 728.670 350.650 728.950 ;
        RECT 350.370 728.050 350.650 728.330 ;
        RECT 350.370 727.430 350.650 727.710 ;
        RECT 350.370 726.810 350.650 727.090 ;
        RECT 350.370 726.190 350.650 726.470 ;
        RECT 350.370 725.570 350.650 725.850 ;
        RECT 350.370 724.950 350.650 725.230 ;
        RECT 350.370 724.330 350.650 724.610 ;
        RECT 389.040 733.070 389.320 733.350 ;
        RECT 389.660 733.070 389.940 733.350 ;
        RECT 390.280 733.070 390.560 733.350 ;
        RECT 390.900 733.070 391.180 733.350 ;
        RECT 391.520 733.070 391.800 733.350 ;
        RECT 392.140 733.070 392.420 733.350 ;
        RECT 392.760 733.070 393.040 733.350 ;
        RECT 389.040 732.450 389.320 732.730 ;
        RECT 389.660 732.450 389.940 732.730 ;
        RECT 390.280 732.450 390.560 732.730 ;
        RECT 390.900 732.450 391.180 732.730 ;
        RECT 391.520 732.450 391.800 732.730 ;
        RECT 392.140 732.450 392.420 732.730 ;
        RECT 392.760 732.450 393.040 732.730 ;
        RECT 389.040 731.830 389.320 732.110 ;
        RECT 389.660 731.830 389.940 732.110 ;
        RECT 390.280 731.830 390.560 732.110 ;
        RECT 390.900 731.830 391.180 732.110 ;
        RECT 391.520 731.830 391.800 732.110 ;
        RECT 392.140 731.830 392.420 732.110 ;
        RECT 392.760 731.830 393.040 732.110 ;
        RECT 389.040 731.210 389.320 731.490 ;
        RECT 389.660 731.210 389.940 731.490 ;
        RECT 390.280 731.210 390.560 731.490 ;
        RECT 390.900 731.210 391.180 731.490 ;
        RECT 391.520 731.210 391.800 731.490 ;
        RECT 392.140 731.210 392.420 731.490 ;
        RECT 392.760 731.210 393.040 731.490 ;
        RECT 389.040 730.590 389.320 730.870 ;
        RECT 389.660 730.590 389.940 730.870 ;
        RECT 390.280 730.590 390.560 730.870 ;
        RECT 390.900 730.590 391.180 730.870 ;
        RECT 391.520 730.590 391.800 730.870 ;
        RECT 392.140 730.590 392.420 730.870 ;
        RECT 392.760 730.590 393.040 730.870 ;
        RECT 389.040 729.970 389.320 730.250 ;
        RECT 389.660 729.970 389.940 730.250 ;
        RECT 390.280 729.970 390.560 730.250 ;
        RECT 390.900 729.970 391.180 730.250 ;
        RECT 391.520 729.970 391.800 730.250 ;
        RECT 392.140 729.970 392.420 730.250 ;
        RECT 392.760 729.970 393.040 730.250 ;
        RECT 389.040 729.350 389.320 729.630 ;
        RECT 389.660 729.350 389.940 729.630 ;
        RECT 390.280 729.350 390.560 729.630 ;
        RECT 390.900 729.350 391.180 729.630 ;
        RECT 391.520 729.350 391.800 729.630 ;
        RECT 392.140 729.350 392.420 729.630 ;
        RECT 392.760 729.350 393.040 729.630 ;
        RECT 389.040 728.730 389.320 729.010 ;
        RECT 389.660 728.730 389.940 729.010 ;
        RECT 390.280 728.730 390.560 729.010 ;
        RECT 390.900 728.730 391.180 729.010 ;
        RECT 391.520 728.730 391.800 729.010 ;
        RECT 392.140 728.730 392.420 729.010 ;
        RECT 392.760 728.730 393.040 729.010 ;
        RECT 389.040 728.110 389.320 728.390 ;
        RECT 389.660 728.110 389.940 728.390 ;
        RECT 390.280 728.110 390.560 728.390 ;
        RECT 390.900 728.110 391.180 728.390 ;
        RECT 391.520 728.110 391.800 728.390 ;
        RECT 392.140 728.110 392.420 728.390 ;
        RECT 392.760 728.110 393.040 728.390 ;
        RECT 389.040 727.490 389.320 727.770 ;
        RECT 389.660 727.490 389.940 727.770 ;
        RECT 390.280 727.490 390.560 727.770 ;
        RECT 390.900 727.490 391.180 727.770 ;
        RECT 391.520 727.490 391.800 727.770 ;
        RECT 392.140 727.490 392.420 727.770 ;
        RECT 392.760 727.490 393.040 727.770 ;
        RECT 389.040 726.870 389.320 727.150 ;
        RECT 389.660 726.870 389.940 727.150 ;
        RECT 390.280 726.870 390.560 727.150 ;
        RECT 390.900 726.870 391.180 727.150 ;
        RECT 391.520 726.870 391.800 727.150 ;
        RECT 392.140 726.870 392.420 727.150 ;
        RECT 392.760 726.870 393.040 727.150 ;
        RECT 389.040 726.250 389.320 726.530 ;
        RECT 389.660 726.250 389.940 726.530 ;
        RECT 390.280 726.250 390.560 726.530 ;
        RECT 390.900 726.250 391.180 726.530 ;
        RECT 391.520 726.250 391.800 726.530 ;
        RECT 392.140 726.250 392.420 726.530 ;
        RECT 392.760 726.250 393.040 726.530 ;
        RECT 389.040 725.630 389.320 725.910 ;
        RECT 389.660 725.630 389.940 725.910 ;
        RECT 390.280 725.630 390.560 725.910 ;
        RECT 390.900 725.630 391.180 725.910 ;
        RECT 391.520 725.630 391.800 725.910 ;
        RECT 392.140 725.630 392.420 725.910 ;
        RECT 392.760 725.630 393.040 725.910 ;
        RECT 389.040 725.010 389.320 725.290 ;
        RECT 389.660 725.010 389.940 725.290 ;
        RECT 390.280 725.010 390.560 725.290 ;
        RECT 390.900 725.010 391.180 725.290 ;
        RECT 391.520 725.010 391.800 725.290 ;
        RECT 392.140 725.010 392.420 725.290 ;
        RECT 392.760 725.010 393.040 725.290 ;
        RECT 389.040 724.390 389.320 724.670 ;
        RECT 389.660 724.390 389.940 724.670 ;
        RECT 390.280 724.390 390.560 724.670 ;
        RECT 390.900 724.390 391.180 724.670 ;
        RECT 391.520 724.390 391.800 724.670 ;
        RECT 392.140 724.390 392.420 724.670 ;
        RECT 392.760 724.390 393.040 724.670 ;
        RECT 350.370 720.640 350.650 720.920 ;
        RECT 350.370 720.020 350.650 720.300 ;
        RECT 350.370 719.400 350.650 719.680 ;
        RECT 350.370 718.780 350.650 719.060 ;
        RECT 350.370 718.160 350.650 718.440 ;
        RECT 350.370 717.540 350.650 717.820 ;
        RECT 350.370 716.920 350.650 717.200 ;
        RECT 350.370 716.300 350.650 716.580 ;
        RECT 350.370 715.680 350.650 715.960 ;
        RECT 350.370 715.060 350.650 715.340 ;
        RECT 350.370 714.440 350.650 714.720 ;
        RECT 350.370 713.820 350.650 714.100 ;
        RECT 350.370 713.200 350.650 713.480 ;
        RECT 350.370 712.580 350.650 712.860 ;
        RECT 350.370 711.960 350.650 712.240 ;
        RECT 350.370 711.340 350.650 711.620 ;
        RECT 389.040 720.670 389.320 720.950 ;
        RECT 389.660 720.670 389.940 720.950 ;
        RECT 390.280 720.670 390.560 720.950 ;
        RECT 390.900 720.670 391.180 720.950 ;
        RECT 391.520 720.670 391.800 720.950 ;
        RECT 392.140 720.670 392.420 720.950 ;
        RECT 392.760 720.670 393.040 720.950 ;
        RECT 389.040 720.050 389.320 720.330 ;
        RECT 389.660 720.050 389.940 720.330 ;
        RECT 390.280 720.050 390.560 720.330 ;
        RECT 390.900 720.050 391.180 720.330 ;
        RECT 391.520 720.050 391.800 720.330 ;
        RECT 392.140 720.050 392.420 720.330 ;
        RECT 392.760 720.050 393.040 720.330 ;
        RECT 389.040 719.430 389.320 719.710 ;
        RECT 389.660 719.430 389.940 719.710 ;
        RECT 390.280 719.430 390.560 719.710 ;
        RECT 390.900 719.430 391.180 719.710 ;
        RECT 391.520 719.430 391.800 719.710 ;
        RECT 392.140 719.430 392.420 719.710 ;
        RECT 392.760 719.430 393.040 719.710 ;
        RECT 389.040 718.810 389.320 719.090 ;
        RECT 389.660 718.810 389.940 719.090 ;
        RECT 390.280 718.810 390.560 719.090 ;
        RECT 390.900 718.810 391.180 719.090 ;
        RECT 391.520 718.810 391.800 719.090 ;
        RECT 392.140 718.810 392.420 719.090 ;
        RECT 392.760 718.810 393.040 719.090 ;
        RECT 389.040 718.190 389.320 718.470 ;
        RECT 389.660 718.190 389.940 718.470 ;
        RECT 390.280 718.190 390.560 718.470 ;
        RECT 390.900 718.190 391.180 718.470 ;
        RECT 391.520 718.190 391.800 718.470 ;
        RECT 392.140 718.190 392.420 718.470 ;
        RECT 392.760 718.190 393.040 718.470 ;
        RECT 389.040 717.570 389.320 717.850 ;
        RECT 389.660 717.570 389.940 717.850 ;
        RECT 390.280 717.570 390.560 717.850 ;
        RECT 390.900 717.570 391.180 717.850 ;
        RECT 391.520 717.570 391.800 717.850 ;
        RECT 392.140 717.570 392.420 717.850 ;
        RECT 392.760 717.570 393.040 717.850 ;
        RECT 389.040 716.950 389.320 717.230 ;
        RECT 389.660 716.950 389.940 717.230 ;
        RECT 390.280 716.950 390.560 717.230 ;
        RECT 390.900 716.950 391.180 717.230 ;
        RECT 391.520 716.950 391.800 717.230 ;
        RECT 392.140 716.950 392.420 717.230 ;
        RECT 392.760 716.950 393.040 717.230 ;
        RECT 389.040 716.330 389.320 716.610 ;
        RECT 389.660 716.330 389.940 716.610 ;
        RECT 390.280 716.330 390.560 716.610 ;
        RECT 390.900 716.330 391.180 716.610 ;
        RECT 391.520 716.330 391.800 716.610 ;
        RECT 392.140 716.330 392.420 716.610 ;
        RECT 392.760 716.330 393.040 716.610 ;
        RECT 389.040 715.710 389.320 715.990 ;
        RECT 389.660 715.710 389.940 715.990 ;
        RECT 390.280 715.710 390.560 715.990 ;
        RECT 390.900 715.710 391.180 715.990 ;
        RECT 391.520 715.710 391.800 715.990 ;
        RECT 392.140 715.710 392.420 715.990 ;
        RECT 392.760 715.710 393.040 715.990 ;
        RECT 389.040 715.090 389.320 715.370 ;
        RECT 389.660 715.090 389.940 715.370 ;
        RECT 390.280 715.090 390.560 715.370 ;
        RECT 390.900 715.090 391.180 715.370 ;
        RECT 391.520 715.090 391.800 715.370 ;
        RECT 392.140 715.090 392.420 715.370 ;
        RECT 392.760 715.090 393.040 715.370 ;
        RECT 389.040 714.470 389.320 714.750 ;
        RECT 389.660 714.470 389.940 714.750 ;
        RECT 390.280 714.470 390.560 714.750 ;
        RECT 390.900 714.470 391.180 714.750 ;
        RECT 391.520 714.470 391.800 714.750 ;
        RECT 392.140 714.470 392.420 714.750 ;
        RECT 392.760 714.470 393.040 714.750 ;
        RECT 389.040 713.850 389.320 714.130 ;
        RECT 389.660 713.850 389.940 714.130 ;
        RECT 390.280 713.850 390.560 714.130 ;
        RECT 390.900 713.850 391.180 714.130 ;
        RECT 391.520 713.850 391.800 714.130 ;
        RECT 392.140 713.850 392.420 714.130 ;
        RECT 392.760 713.850 393.040 714.130 ;
        RECT 389.040 713.230 389.320 713.510 ;
        RECT 389.660 713.230 389.940 713.510 ;
        RECT 390.280 713.230 390.560 713.510 ;
        RECT 390.900 713.230 391.180 713.510 ;
        RECT 391.520 713.230 391.800 713.510 ;
        RECT 392.140 713.230 392.420 713.510 ;
        RECT 392.760 713.230 393.040 713.510 ;
        RECT 389.040 712.610 389.320 712.890 ;
        RECT 389.660 712.610 389.940 712.890 ;
        RECT 390.280 712.610 390.560 712.890 ;
        RECT 390.900 712.610 391.180 712.890 ;
        RECT 391.520 712.610 391.800 712.890 ;
        RECT 392.140 712.610 392.420 712.890 ;
        RECT 392.760 712.610 393.040 712.890 ;
        RECT 389.040 711.990 389.320 712.270 ;
        RECT 389.660 711.990 389.940 712.270 ;
        RECT 390.280 711.990 390.560 712.270 ;
        RECT 390.900 711.990 391.180 712.270 ;
        RECT 391.520 711.990 391.800 712.270 ;
        RECT 392.140 711.990 392.420 712.270 ;
        RECT 392.760 711.990 393.040 712.270 ;
        RECT 389.040 711.370 389.320 711.650 ;
        RECT 389.660 711.370 389.940 711.650 ;
        RECT 390.280 711.370 390.560 711.650 ;
        RECT 390.900 711.370 391.180 711.650 ;
        RECT 391.520 711.370 391.800 711.650 ;
        RECT 392.140 711.370 392.420 711.650 ;
        RECT 392.760 711.370 393.040 711.650 ;
        RECT 350.370 708.790 350.650 709.070 ;
        RECT 350.370 708.170 350.650 708.450 ;
        RECT 350.370 707.550 350.650 707.830 ;
        RECT 350.370 706.930 350.650 707.210 ;
        RECT 350.370 706.310 350.650 706.590 ;
        RECT 350.370 705.690 350.650 705.970 ;
        RECT 350.370 705.070 350.650 705.350 ;
        RECT 350.370 704.450 350.650 704.730 ;
        RECT 350.370 703.830 350.650 704.110 ;
        RECT 350.370 703.210 350.650 703.490 ;
        RECT 350.370 702.590 350.650 702.870 ;
        RECT 350.370 701.970 350.650 702.250 ;
        RECT 350.370 701.350 350.650 701.630 ;
        RECT 350.370 700.730 350.650 701.010 ;
        RECT 350.370 700.110 350.650 700.390 ;
        RECT 350.370 699.490 350.650 699.770 ;
        RECT 389.040 708.820 389.320 709.100 ;
        RECT 389.660 708.820 389.940 709.100 ;
        RECT 390.280 708.820 390.560 709.100 ;
        RECT 390.900 708.820 391.180 709.100 ;
        RECT 391.520 708.820 391.800 709.100 ;
        RECT 392.140 708.820 392.420 709.100 ;
        RECT 392.760 708.820 393.040 709.100 ;
        RECT 389.040 708.200 389.320 708.480 ;
        RECT 389.660 708.200 389.940 708.480 ;
        RECT 390.280 708.200 390.560 708.480 ;
        RECT 390.900 708.200 391.180 708.480 ;
        RECT 391.520 708.200 391.800 708.480 ;
        RECT 392.140 708.200 392.420 708.480 ;
        RECT 392.760 708.200 393.040 708.480 ;
        RECT 389.040 707.580 389.320 707.860 ;
        RECT 389.660 707.580 389.940 707.860 ;
        RECT 390.280 707.580 390.560 707.860 ;
        RECT 390.900 707.580 391.180 707.860 ;
        RECT 391.520 707.580 391.800 707.860 ;
        RECT 392.140 707.580 392.420 707.860 ;
        RECT 392.760 707.580 393.040 707.860 ;
        RECT 389.040 706.960 389.320 707.240 ;
        RECT 389.660 706.960 389.940 707.240 ;
        RECT 390.280 706.960 390.560 707.240 ;
        RECT 390.900 706.960 391.180 707.240 ;
        RECT 391.520 706.960 391.800 707.240 ;
        RECT 392.140 706.960 392.420 707.240 ;
        RECT 392.760 706.960 393.040 707.240 ;
        RECT 389.040 706.340 389.320 706.620 ;
        RECT 389.660 706.340 389.940 706.620 ;
        RECT 390.280 706.340 390.560 706.620 ;
        RECT 390.900 706.340 391.180 706.620 ;
        RECT 391.520 706.340 391.800 706.620 ;
        RECT 392.140 706.340 392.420 706.620 ;
        RECT 392.760 706.340 393.040 706.620 ;
        RECT 389.040 705.720 389.320 706.000 ;
        RECT 389.660 705.720 389.940 706.000 ;
        RECT 390.280 705.720 390.560 706.000 ;
        RECT 390.900 705.720 391.180 706.000 ;
        RECT 391.520 705.720 391.800 706.000 ;
        RECT 392.140 705.720 392.420 706.000 ;
        RECT 392.760 705.720 393.040 706.000 ;
        RECT 389.040 705.100 389.320 705.380 ;
        RECT 389.660 705.100 389.940 705.380 ;
        RECT 390.280 705.100 390.560 705.380 ;
        RECT 390.900 705.100 391.180 705.380 ;
        RECT 391.520 705.100 391.800 705.380 ;
        RECT 392.140 705.100 392.420 705.380 ;
        RECT 392.760 705.100 393.040 705.380 ;
        RECT 389.040 704.480 389.320 704.760 ;
        RECT 389.660 704.480 389.940 704.760 ;
        RECT 390.280 704.480 390.560 704.760 ;
        RECT 390.900 704.480 391.180 704.760 ;
        RECT 391.520 704.480 391.800 704.760 ;
        RECT 392.140 704.480 392.420 704.760 ;
        RECT 392.760 704.480 393.040 704.760 ;
        RECT 389.040 703.860 389.320 704.140 ;
        RECT 389.660 703.860 389.940 704.140 ;
        RECT 390.280 703.860 390.560 704.140 ;
        RECT 390.900 703.860 391.180 704.140 ;
        RECT 391.520 703.860 391.800 704.140 ;
        RECT 392.140 703.860 392.420 704.140 ;
        RECT 392.760 703.860 393.040 704.140 ;
        RECT 389.040 703.240 389.320 703.520 ;
        RECT 389.660 703.240 389.940 703.520 ;
        RECT 390.280 703.240 390.560 703.520 ;
        RECT 390.900 703.240 391.180 703.520 ;
        RECT 391.520 703.240 391.800 703.520 ;
        RECT 392.140 703.240 392.420 703.520 ;
        RECT 392.760 703.240 393.040 703.520 ;
        RECT 389.040 702.620 389.320 702.900 ;
        RECT 389.660 702.620 389.940 702.900 ;
        RECT 390.280 702.620 390.560 702.900 ;
        RECT 390.900 702.620 391.180 702.900 ;
        RECT 391.520 702.620 391.800 702.900 ;
        RECT 392.140 702.620 392.420 702.900 ;
        RECT 392.760 702.620 393.040 702.900 ;
        RECT 389.040 702.000 389.320 702.280 ;
        RECT 389.660 702.000 389.940 702.280 ;
        RECT 390.280 702.000 390.560 702.280 ;
        RECT 390.900 702.000 391.180 702.280 ;
        RECT 391.520 702.000 391.800 702.280 ;
        RECT 392.140 702.000 392.420 702.280 ;
        RECT 392.760 702.000 393.040 702.280 ;
        RECT 389.040 701.380 389.320 701.660 ;
        RECT 389.660 701.380 389.940 701.660 ;
        RECT 390.280 701.380 390.560 701.660 ;
        RECT 390.900 701.380 391.180 701.660 ;
        RECT 391.520 701.380 391.800 701.660 ;
        RECT 392.140 701.380 392.420 701.660 ;
        RECT 392.760 701.380 393.040 701.660 ;
        RECT 389.040 700.760 389.320 701.040 ;
        RECT 389.660 700.760 389.940 701.040 ;
        RECT 390.280 700.760 390.560 701.040 ;
        RECT 390.900 700.760 391.180 701.040 ;
        RECT 391.520 700.760 391.800 701.040 ;
        RECT 392.140 700.760 392.420 701.040 ;
        RECT 392.760 700.760 393.040 701.040 ;
        RECT 389.040 700.140 389.320 700.420 ;
        RECT 389.660 700.140 389.940 700.420 ;
        RECT 390.280 700.140 390.560 700.420 ;
        RECT 390.900 700.140 391.180 700.420 ;
        RECT 391.520 700.140 391.800 700.420 ;
        RECT 392.140 700.140 392.420 700.420 ;
        RECT 392.760 700.140 393.040 700.420 ;
        RECT 389.040 699.520 389.320 699.800 ;
        RECT 389.660 699.520 389.940 699.800 ;
        RECT 390.280 699.520 390.560 699.800 ;
        RECT 390.900 699.520 391.180 699.800 ;
        RECT 391.520 699.520 391.800 699.800 ;
        RECT 392.140 699.520 392.420 699.800 ;
        RECT 392.760 699.520 393.040 699.800 ;
        RECT 350.370 695.260 350.650 695.540 ;
        RECT 350.370 694.640 350.650 694.920 ;
        RECT 350.370 694.020 350.650 694.300 ;
        RECT 350.370 693.400 350.650 693.680 ;
        RECT 350.370 692.780 350.650 693.060 ;
        RECT 350.370 692.160 350.650 692.440 ;
        RECT 350.370 691.540 350.650 691.820 ;
        RECT 350.370 690.920 350.650 691.200 ;
        RECT 350.370 690.300 350.650 690.580 ;
        RECT 350.370 689.680 350.650 689.960 ;
        RECT 350.370 689.060 350.650 689.340 ;
        RECT 350.370 688.440 350.650 688.720 ;
        RECT 350.370 687.820 350.650 688.100 ;
        RECT 350.370 687.200 350.650 687.480 ;
        RECT 350.370 686.580 350.650 686.860 ;
        RECT 350.370 685.960 350.650 686.240 ;
        RECT 389.040 695.290 389.320 695.570 ;
        RECT 389.660 695.290 389.940 695.570 ;
        RECT 390.280 695.290 390.560 695.570 ;
        RECT 390.900 695.290 391.180 695.570 ;
        RECT 391.520 695.290 391.800 695.570 ;
        RECT 392.140 695.290 392.420 695.570 ;
        RECT 392.760 695.290 393.040 695.570 ;
        RECT 389.040 694.670 389.320 694.950 ;
        RECT 389.660 694.670 389.940 694.950 ;
        RECT 390.280 694.670 390.560 694.950 ;
        RECT 390.900 694.670 391.180 694.950 ;
        RECT 391.520 694.670 391.800 694.950 ;
        RECT 392.140 694.670 392.420 694.950 ;
        RECT 392.760 694.670 393.040 694.950 ;
        RECT 389.040 694.050 389.320 694.330 ;
        RECT 389.660 694.050 389.940 694.330 ;
        RECT 390.280 694.050 390.560 694.330 ;
        RECT 390.900 694.050 391.180 694.330 ;
        RECT 391.520 694.050 391.800 694.330 ;
        RECT 392.140 694.050 392.420 694.330 ;
        RECT 392.760 694.050 393.040 694.330 ;
        RECT 389.040 693.430 389.320 693.710 ;
        RECT 389.660 693.430 389.940 693.710 ;
        RECT 390.280 693.430 390.560 693.710 ;
        RECT 390.900 693.430 391.180 693.710 ;
        RECT 391.520 693.430 391.800 693.710 ;
        RECT 392.140 693.430 392.420 693.710 ;
        RECT 392.760 693.430 393.040 693.710 ;
        RECT 389.040 692.810 389.320 693.090 ;
        RECT 389.660 692.810 389.940 693.090 ;
        RECT 390.280 692.810 390.560 693.090 ;
        RECT 390.900 692.810 391.180 693.090 ;
        RECT 391.520 692.810 391.800 693.090 ;
        RECT 392.140 692.810 392.420 693.090 ;
        RECT 392.760 692.810 393.040 693.090 ;
        RECT 389.040 692.190 389.320 692.470 ;
        RECT 389.660 692.190 389.940 692.470 ;
        RECT 390.280 692.190 390.560 692.470 ;
        RECT 390.900 692.190 391.180 692.470 ;
        RECT 391.520 692.190 391.800 692.470 ;
        RECT 392.140 692.190 392.420 692.470 ;
        RECT 392.760 692.190 393.040 692.470 ;
        RECT 389.040 691.570 389.320 691.850 ;
        RECT 389.660 691.570 389.940 691.850 ;
        RECT 390.280 691.570 390.560 691.850 ;
        RECT 390.900 691.570 391.180 691.850 ;
        RECT 391.520 691.570 391.800 691.850 ;
        RECT 392.140 691.570 392.420 691.850 ;
        RECT 392.760 691.570 393.040 691.850 ;
        RECT 389.040 690.950 389.320 691.230 ;
        RECT 389.660 690.950 389.940 691.230 ;
        RECT 390.280 690.950 390.560 691.230 ;
        RECT 390.900 690.950 391.180 691.230 ;
        RECT 391.520 690.950 391.800 691.230 ;
        RECT 392.140 690.950 392.420 691.230 ;
        RECT 392.760 690.950 393.040 691.230 ;
        RECT 389.040 690.330 389.320 690.610 ;
        RECT 389.660 690.330 389.940 690.610 ;
        RECT 390.280 690.330 390.560 690.610 ;
        RECT 390.900 690.330 391.180 690.610 ;
        RECT 391.520 690.330 391.800 690.610 ;
        RECT 392.140 690.330 392.420 690.610 ;
        RECT 392.760 690.330 393.040 690.610 ;
        RECT 389.040 689.710 389.320 689.990 ;
        RECT 389.660 689.710 389.940 689.990 ;
        RECT 390.280 689.710 390.560 689.990 ;
        RECT 390.900 689.710 391.180 689.990 ;
        RECT 391.520 689.710 391.800 689.990 ;
        RECT 392.140 689.710 392.420 689.990 ;
        RECT 392.760 689.710 393.040 689.990 ;
        RECT 389.040 689.090 389.320 689.370 ;
        RECT 389.660 689.090 389.940 689.370 ;
        RECT 390.280 689.090 390.560 689.370 ;
        RECT 390.900 689.090 391.180 689.370 ;
        RECT 391.520 689.090 391.800 689.370 ;
        RECT 392.140 689.090 392.420 689.370 ;
        RECT 392.760 689.090 393.040 689.370 ;
        RECT 389.040 688.470 389.320 688.750 ;
        RECT 389.660 688.470 389.940 688.750 ;
        RECT 390.280 688.470 390.560 688.750 ;
        RECT 390.900 688.470 391.180 688.750 ;
        RECT 391.520 688.470 391.800 688.750 ;
        RECT 392.140 688.470 392.420 688.750 ;
        RECT 392.760 688.470 393.040 688.750 ;
        RECT 389.040 687.850 389.320 688.130 ;
        RECT 389.660 687.850 389.940 688.130 ;
        RECT 390.280 687.850 390.560 688.130 ;
        RECT 390.900 687.850 391.180 688.130 ;
        RECT 391.520 687.850 391.800 688.130 ;
        RECT 392.140 687.850 392.420 688.130 ;
        RECT 392.760 687.850 393.040 688.130 ;
        RECT 389.040 687.230 389.320 687.510 ;
        RECT 389.660 687.230 389.940 687.510 ;
        RECT 390.280 687.230 390.560 687.510 ;
        RECT 390.900 687.230 391.180 687.510 ;
        RECT 391.520 687.230 391.800 687.510 ;
        RECT 392.140 687.230 392.420 687.510 ;
        RECT 392.760 687.230 393.040 687.510 ;
        RECT 389.040 686.610 389.320 686.890 ;
        RECT 389.660 686.610 389.940 686.890 ;
        RECT 390.280 686.610 390.560 686.890 ;
        RECT 390.900 686.610 391.180 686.890 ;
        RECT 391.520 686.610 391.800 686.890 ;
        RECT 392.140 686.610 392.420 686.890 ;
        RECT 392.760 686.610 393.040 686.890 ;
        RECT 389.040 685.990 389.320 686.270 ;
        RECT 389.660 685.990 389.940 686.270 ;
        RECT 390.280 685.990 390.560 686.270 ;
        RECT 390.900 685.990 391.180 686.270 ;
        RECT 391.520 685.990 391.800 686.270 ;
        RECT 392.140 685.990 392.420 686.270 ;
        RECT 392.760 685.990 393.040 686.270 ;
        RECT 350.370 683.410 350.650 683.690 ;
        RECT 350.370 682.790 350.650 683.070 ;
        RECT 350.370 682.170 350.650 682.450 ;
        RECT 350.370 681.550 350.650 681.830 ;
        RECT 350.370 680.930 350.650 681.210 ;
        RECT 350.370 680.310 350.650 680.590 ;
        RECT 350.370 679.690 350.650 679.970 ;
        RECT 350.370 679.070 350.650 679.350 ;
        RECT 350.370 678.450 350.650 678.730 ;
        RECT 350.370 677.830 350.650 678.110 ;
        RECT 350.370 677.210 350.650 677.490 ;
        RECT 350.370 676.590 350.650 676.870 ;
        RECT 350.370 675.970 350.650 676.250 ;
        RECT 350.370 675.350 350.650 675.630 ;
        RECT 350.370 674.730 350.650 675.010 ;
        RECT 350.370 674.110 350.650 674.390 ;
        RECT 389.040 683.440 389.320 683.720 ;
        RECT 389.660 683.440 389.940 683.720 ;
        RECT 390.280 683.440 390.560 683.720 ;
        RECT 390.900 683.440 391.180 683.720 ;
        RECT 391.520 683.440 391.800 683.720 ;
        RECT 392.140 683.440 392.420 683.720 ;
        RECT 392.760 683.440 393.040 683.720 ;
        RECT 389.040 682.820 389.320 683.100 ;
        RECT 389.660 682.820 389.940 683.100 ;
        RECT 390.280 682.820 390.560 683.100 ;
        RECT 390.900 682.820 391.180 683.100 ;
        RECT 391.520 682.820 391.800 683.100 ;
        RECT 392.140 682.820 392.420 683.100 ;
        RECT 392.760 682.820 393.040 683.100 ;
        RECT 389.040 682.200 389.320 682.480 ;
        RECT 389.660 682.200 389.940 682.480 ;
        RECT 390.280 682.200 390.560 682.480 ;
        RECT 390.900 682.200 391.180 682.480 ;
        RECT 391.520 682.200 391.800 682.480 ;
        RECT 392.140 682.200 392.420 682.480 ;
        RECT 392.760 682.200 393.040 682.480 ;
        RECT 389.040 681.580 389.320 681.860 ;
        RECT 389.660 681.580 389.940 681.860 ;
        RECT 390.280 681.580 390.560 681.860 ;
        RECT 390.900 681.580 391.180 681.860 ;
        RECT 391.520 681.580 391.800 681.860 ;
        RECT 392.140 681.580 392.420 681.860 ;
        RECT 392.760 681.580 393.040 681.860 ;
        RECT 389.040 680.960 389.320 681.240 ;
        RECT 389.660 680.960 389.940 681.240 ;
        RECT 390.280 680.960 390.560 681.240 ;
        RECT 390.900 680.960 391.180 681.240 ;
        RECT 391.520 680.960 391.800 681.240 ;
        RECT 392.140 680.960 392.420 681.240 ;
        RECT 392.760 680.960 393.040 681.240 ;
        RECT 389.040 680.340 389.320 680.620 ;
        RECT 389.660 680.340 389.940 680.620 ;
        RECT 390.280 680.340 390.560 680.620 ;
        RECT 390.900 680.340 391.180 680.620 ;
        RECT 391.520 680.340 391.800 680.620 ;
        RECT 392.140 680.340 392.420 680.620 ;
        RECT 392.760 680.340 393.040 680.620 ;
        RECT 389.040 679.720 389.320 680.000 ;
        RECT 389.660 679.720 389.940 680.000 ;
        RECT 390.280 679.720 390.560 680.000 ;
        RECT 390.900 679.720 391.180 680.000 ;
        RECT 391.520 679.720 391.800 680.000 ;
        RECT 392.140 679.720 392.420 680.000 ;
        RECT 392.760 679.720 393.040 680.000 ;
        RECT 389.040 679.100 389.320 679.380 ;
        RECT 389.660 679.100 389.940 679.380 ;
        RECT 390.280 679.100 390.560 679.380 ;
        RECT 390.900 679.100 391.180 679.380 ;
        RECT 391.520 679.100 391.800 679.380 ;
        RECT 392.140 679.100 392.420 679.380 ;
        RECT 392.760 679.100 393.040 679.380 ;
        RECT 389.040 678.480 389.320 678.760 ;
        RECT 389.660 678.480 389.940 678.760 ;
        RECT 390.280 678.480 390.560 678.760 ;
        RECT 390.900 678.480 391.180 678.760 ;
        RECT 391.520 678.480 391.800 678.760 ;
        RECT 392.140 678.480 392.420 678.760 ;
        RECT 392.760 678.480 393.040 678.760 ;
        RECT 389.040 677.860 389.320 678.140 ;
        RECT 389.660 677.860 389.940 678.140 ;
        RECT 390.280 677.860 390.560 678.140 ;
        RECT 390.900 677.860 391.180 678.140 ;
        RECT 391.520 677.860 391.800 678.140 ;
        RECT 392.140 677.860 392.420 678.140 ;
        RECT 392.760 677.860 393.040 678.140 ;
        RECT 389.040 677.240 389.320 677.520 ;
        RECT 389.660 677.240 389.940 677.520 ;
        RECT 390.280 677.240 390.560 677.520 ;
        RECT 390.900 677.240 391.180 677.520 ;
        RECT 391.520 677.240 391.800 677.520 ;
        RECT 392.140 677.240 392.420 677.520 ;
        RECT 392.760 677.240 393.040 677.520 ;
        RECT 389.040 676.620 389.320 676.900 ;
        RECT 389.660 676.620 389.940 676.900 ;
        RECT 390.280 676.620 390.560 676.900 ;
        RECT 390.900 676.620 391.180 676.900 ;
        RECT 391.520 676.620 391.800 676.900 ;
        RECT 392.140 676.620 392.420 676.900 ;
        RECT 392.760 676.620 393.040 676.900 ;
        RECT 389.040 676.000 389.320 676.280 ;
        RECT 389.660 676.000 389.940 676.280 ;
        RECT 390.280 676.000 390.560 676.280 ;
        RECT 390.900 676.000 391.180 676.280 ;
        RECT 391.520 676.000 391.800 676.280 ;
        RECT 392.140 676.000 392.420 676.280 ;
        RECT 392.760 676.000 393.040 676.280 ;
        RECT 389.040 675.380 389.320 675.660 ;
        RECT 389.660 675.380 389.940 675.660 ;
        RECT 390.280 675.380 390.560 675.660 ;
        RECT 390.900 675.380 391.180 675.660 ;
        RECT 391.520 675.380 391.800 675.660 ;
        RECT 392.140 675.380 392.420 675.660 ;
        RECT 392.760 675.380 393.040 675.660 ;
        RECT 389.040 674.760 389.320 675.040 ;
        RECT 389.660 674.760 389.940 675.040 ;
        RECT 390.280 674.760 390.560 675.040 ;
        RECT 390.900 674.760 391.180 675.040 ;
        RECT 391.520 674.760 391.800 675.040 ;
        RECT 392.140 674.760 392.420 675.040 ;
        RECT 392.760 674.760 393.040 675.040 ;
        RECT 389.040 674.140 389.320 674.420 ;
        RECT 389.660 674.140 389.940 674.420 ;
        RECT 390.280 674.140 390.560 674.420 ;
        RECT 390.900 674.140 391.180 674.420 ;
        RECT 391.520 674.140 391.800 674.420 ;
        RECT 392.140 674.140 392.420 674.420 ;
        RECT 392.760 674.140 393.040 674.420 ;
        RECT 350.370 670.390 350.650 670.670 ;
        RECT 350.370 669.770 350.650 670.050 ;
        RECT 350.370 669.150 350.650 669.430 ;
        RECT 350.370 668.530 350.650 668.810 ;
        RECT 350.370 667.910 350.650 668.190 ;
        RECT 350.370 667.290 350.650 667.570 ;
        RECT 350.370 666.670 350.650 666.950 ;
        RECT 350.370 666.050 350.650 666.330 ;
        RECT 350.370 665.430 350.650 665.710 ;
        RECT 350.370 664.810 350.650 665.090 ;
        RECT 350.370 664.190 350.650 664.470 ;
        RECT 350.370 663.570 350.650 663.850 ;
        RECT 350.370 662.950 350.650 663.230 ;
        RECT 350.370 662.330 350.650 662.610 ;
        RECT 350.370 661.710 350.650 661.990 ;
        RECT 389.040 670.420 389.320 670.700 ;
        RECT 389.660 670.420 389.940 670.700 ;
        RECT 390.280 670.420 390.560 670.700 ;
        RECT 390.900 670.420 391.180 670.700 ;
        RECT 391.520 670.420 391.800 670.700 ;
        RECT 392.140 670.420 392.420 670.700 ;
        RECT 392.760 670.420 393.040 670.700 ;
        RECT 389.040 669.800 389.320 670.080 ;
        RECT 389.660 669.800 389.940 670.080 ;
        RECT 390.280 669.800 390.560 670.080 ;
        RECT 390.900 669.800 391.180 670.080 ;
        RECT 391.520 669.800 391.800 670.080 ;
        RECT 392.140 669.800 392.420 670.080 ;
        RECT 392.760 669.800 393.040 670.080 ;
        RECT 389.040 669.180 389.320 669.460 ;
        RECT 389.660 669.180 389.940 669.460 ;
        RECT 390.280 669.180 390.560 669.460 ;
        RECT 390.900 669.180 391.180 669.460 ;
        RECT 391.520 669.180 391.800 669.460 ;
        RECT 392.140 669.180 392.420 669.460 ;
        RECT 392.760 669.180 393.040 669.460 ;
        RECT 389.040 668.560 389.320 668.840 ;
        RECT 389.660 668.560 389.940 668.840 ;
        RECT 390.280 668.560 390.560 668.840 ;
        RECT 390.900 668.560 391.180 668.840 ;
        RECT 391.520 668.560 391.800 668.840 ;
        RECT 392.140 668.560 392.420 668.840 ;
        RECT 392.760 668.560 393.040 668.840 ;
        RECT 389.040 667.940 389.320 668.220 ;
        RECT 389.660 667.940 389.940 668.220 ;
        RECT 390.280 667.940 390.560 668.220 ;
        RECT 390.900 667.940 391.180 668.220 ;
        RECT 391.520 667.940 391.800 668.220 ;
        RECT 392.140 667.940 392.420 668.220 ;
        RECT 392.760 667.940 393.040 668.220 ;
        RECT 389.040 667.320 389.320 667.600 ;
        RECT 389.660 667.320 389.940 667.600 ;
        RECT 390.280 667.320 390.560 667.600 ;
        RECT 390.900 667.320 391.180 667.600 ;
        RECT 391.520 667.320 391.800 667.600 ;
        RECT 392.140 667.320 392.420 667.600 ;
        RECT 392.760 667.320 393.040 667.600 ;
        RECT 389.040 666.700 389.320 666.980 ;
        RECT 389.660 666.700 389.940 666.980 ;
        RECT 390.280 666.700 390.560 666.980 ;
        RECT 390.900 666.700 391.180 666.980 ;
        RECT 391.520 666.700 391.800 666.980 ;
        RECT 392.140 666.700 392.420 666.980 ;
        RECT 392.760 666.700 393.040 666.980 ;
        RECT 389.040 666.080 389.320 666.360 ;
        RECT 389.660 666.080 389.940 666.360 ;
        RECT 390.280 666.080 390.560 666.360 ;
        RECT 390.900 666.080 391.180 666.360 ;
        RECT 391.520 666.080 391.800 666.360 ;
        RECT 392.140 666.080 392.420 666.360 ;
        RECT 392.760 666.080 393.040 666.360 ;
        RECT 389.040 665.460 389.320 665.740 ;
        RECT 389.660 665.460 389.940 665.740 ;
        RECT 390.280 665.460 390.560 665.740 ;
        RECT 390.900 665.460 391.180 665.740 ;
        RECT 391.520 665.460 391.800 665.740 ;
        RECT 392.140 665.460 392.420 665.740 ;
        RECT 392.760 665.460 393.040 665.740 ;
        RECT 389.040 664.840 389.320 665.120 ;
        RECT 389.660 664.840 389.940 665.120 ;
        RECT 390.280 664.840 390.560 665.120 ;
        RECT 390.900 664.840 391.180 665.120 ;
        RECT 391.520 664.840 391.800 665.120 ;
        RECT 392.140 664.840 392.420 665.120 ;
        RECT 392.760 664.840 393.040 665.120 ;
        RECT 389.040 664.220 389.320 664.500 ;
        RECT 389.660 664.220 389.940 664.500 ;
        RECT 390.280 664.220 390.560 664.500 ;
        RECT 390.900 664.220 391.180 664.500 ;
        RECT 391.520 664.220 391.800 664.500 ;
        RECT 392.140 664.220 392.420 664.500 ;
        RECT 392.760 664.220 393.040 664.500 ;
        RECT 389.040 663.600 389.320 663.880 ;
        RECT 389.660 663.600 389.940 663.880 ;
        RECT 390.280 663.600 390.560 663.880 ;
        RECT 390.900 663.600 391.180 663.880 ;
        RECT 391.520 663.600 391.800 663.880 ;
        RECT 392.140 663.600 392.420 663.880 ;
        RECT 392.760 663.600 393.040 663.880 ;
        RECT 389.040 662.980 389.320 663.260 ;
        RECT 389.660 662.980 389.940 663.260 ;
        RECT 390.280 662.980 390.560 663.260 ;
        RECT 390.900 662.980 391.180 663.260 ;
        RECT 391.520 662.980 391.800 663.260 ;
        RECT 392.140 662.980 392.420 663.260 ;
        RECT 392.760 662.980 393.040 663.260 ;
        RECT 389.040 662.360 389.320 662.640 ;
        RECT 389.660 662.360 389.940 662.640 ;
        RECT 390.280 662.360 390.560 662.640 ;
        RECT 390.900 662.360 391.180 662.640 ;
        RECT 391.520 662.360 391.800 662.640 ;
        RECT 392.140 662.360 392.420 662.640 ;
        RECT 392.760 662.360 393.040 662.640 ;
        RECT 389.040 661.740 389.320 662.020 ;
        RECT 389.660 661.740 389.940 662.020 ;
        RECT 390.280 661.740 390.560 662.020 ;
        RECT 390.900 661.740 391.180 662.020 ;
        RECT 391.520 661.740 391.800 662.020 ;
        RECT 392.140 661.740 392.420 662.020 ;
        RECT 392.760 661.740 393.040 662.020 ;
        RECT 388.740 561.580 389.020 561.860 ;
        RECT 389.360 561.580 389.640 561.860 ;
        RECT 389.980 561.580 390.260 561.860 ;
        RECT 390.600 561.580 390.880 561.860 ;
        RECT 391.220 561.580 391.500 561.860 ;
        RECT 391.840 561.580 392.120 561.860 ;
        RECT 392.460 561.580 392.740 561.860 ;
        RECT 388.740 560.960 389.020 561.240 ;
        RECT 389.360 560.960 389.640 561.240 ;
        RECT 389.980 560.960 390.260 561.240 ;
        RECT 390.600 560.960 390.880 561.240 ;
        RECT 391.220 560.960 391.500 561.240 ;
        RECT 391.840 560.960 392.120 561.240 ;
        RECT 392.460 560.960 392.740 561.240 ;
        RECT 350.370 528.010 350.650 528.290 ;
        RECT 350.370 527.390 350.650 527.670 ;
        RECT 350.370 526.770 350.650 527.050 ;
        RECT 350.370 526.150 350.650 526.430 ;
        RECT 350.370 525.530 350.650 525.810 ;
        RECT 350.370 524.910 350.650 525.190 ;
        RECT 350.370 524.290 350.650 524.570 ;
        RECT 350.370 523.670 350.650 523.950 ;
        RECT 350.370 523.050 350.650 523.330 ;
        RECT 350.370 522.430 350.650 522.710 ;
        RECT 350.370 521.810 350.650 522.090 ;
        RECT 350.370 521.190 350.650 521.470 ;
        RECT 350.370 520.570 350.650 520.850 ;
        RECT 350.370 519.950 350.650 520.230 ;
        RECT 350.370 519.330 350.650 519.610 ;
        RECT 389.040 528.070 389.320 528.350 ;
        RECT 389.660 528.070 389.940 528.350 ;
        RECT 390.280 528.070 390.560 528.350 ;
        RECT 390.900 528.070 391.180 528.350 ;
        RECT 391.520 528.070 391.800 528.350 ;
        RECT 392.140 528.070 392.420 528.350 ;
        RECT 392.760 528.070 393.040 528.350 ;
        RECT 389.040 527.450 389.320 527.730 ;
        RECT 389.660 527.450 389.940 527.730 ;
        RECT 390.280 527.450 390.560 527.730 ;
        RECT 390.900 527.450 391.180 527.730 ;
        RECT 391.520 527.450 391.800 527.730 ;
        RECT 392.140 527.450 392.420 527.730 ;
        RECT 392.760 527.450 393.040 527.730 ;
        RECT 389.040 526.830 389.320 527.110 ;
        RECT 389.660 526.830 389.940 527.110 ;
        RECT 390.280 526.830 390.560 527.110 ;
        RECT 390.900 526.830 391.180 527.110 ;
        RECT 391.520 526.830 391.800 527.110 ;
        RECT 392.140 526.830 392.420 527.110 ;
        RECT 392.760 526.830 393.040 527.110 ;
        RECT 389.040 526.210 389.320 526.490 ;
        RECT 389.660 526.210 389.940 526.490 ;
        RECT 390.280 526.210 390.560 526.490 ;
        RECT 390.900 526.210 391.180 526.490 ;
        RECT 391.520 526.210 391.800 526.490 ;
        RECT 392.140 526.210 392.420 526.490 ;
        RECT 392.760 526.210 393.040 526.490 ;
        RECT 389.040 525.590 389.320 525.870 ;
        RECT 389.660 525.590 389.940 525.870 ;
        RECT 390.280 525.590 390.560 525.870 ;
        RECT 390.900 525.590 391.180 525.870 ;
        RECT 391.520 525.590 391.800 525.870 ;
        RECT 392.140 525.590 392.420 525.870 ;
        RECT 392.760 525.590 393.040 525.870 ;
        RECT 389.040 524.970 389.320 525.250 ;
        RECT 389.660 524.970 389.940 525.250 ;
        RECT 390.280 524.970 390.560 525.250 ;
        RECT 390.900 524.970 391.180 525.250 ;
        RECT 391.520 524.970 391.800 525.250 ;
        RECT 392.140 524.970 392.420 525.250 ;
        RECT 392.760 524.970 393.040 525.250 ;
        RECT 389.040 524.350 389.320 524.630 ;
        RECT 389.660 524.350 389.940 524.630 ;
        RECT 390.280 524.350 390.560 524.630 ;
        RECT 390.900 524.350 391.180 524.630 ;
        RECT 391.520 524.350 391.800 524.630 ;
        RECT 392.140 524.350 392.420 524.630 ;
        RECT 392.760 524.350 393.040 524.630 ;
        RECT 389.040 523.730 389.320 524.010 ;
        RECT 389.660 523.730 389.940 524.010 ;
        RECT 390.280 523.730 390.560 524.010 ;
        RECT 390.900 523.730 391.180 524.010 ;
        RECT 391.520 523.730 391.800 524.010 ;
        RECT 392.140 523.730 392.420 524.010 ;
        RECT 392.760 523.730 393.040 524.010 ;
        RECT 389.040 523.110 389.320 523.390 ;
        RECT 389.660 523.110 389.940 523.390 ;
        RECT 390.280 523.110 390.560 523.390 ;
        RECT 390.900 523.110 391.180 523.390 ;
        RECT 391.520 523.110 391.800 523.390 ;
        RECT 392.140 523.110 392.420 523.390 ;
        RECT 392.760 523.110 393.040 523.390 ;
        RECT 389.040 522.490 389.320 522.770 ;
        RECT 389.660 522.490 389.940 522.770 ;
        RECT 390.280 522.490 390.560 522.770 ;
        RECT 390.900 522.490 391.180 522.770 ;
        RECT 391.520 522.490 391.800 522.770 ;
        RECT 392.140 522.490 392.420 522.770 ;
        RECT 392.760 522.490 393.040 522.770 ;
        RECT 389.040 521.870 389.320 522.150 ;
        RECT 389.660 521.870 389.940 522.150 ;
        RECT 390.280 521.870 390.560 522.150 ;
        RECT 390.900 521.870 391.180 522.150 ;
        RECT 391.520 521.870 391.800 522.150 ;
        RECT 392.140 521.870 392.420 522.150 ;
        RECT 392.760 521.870 393.040 522.150 ;
        RECT 389.040 521.250 389.320 521.530 ;
        RECT 389.660 521.250 389.940 521.530 ;
        RECT 390.280 521.250 390.560 521.530 ;
        RECT 390.900 521.250 391.180 521.530 ;
        RECT 391.520 521.250 391.800 521.530 ;
        RECT 392.140 521.250 392.420 521.530 ;
        RECT 392.760 521.250 393.040 521.530 ;
        RECT 389.040 520.630 389.320 520.910 ;
        RECT 389.660 520.630 389.940 520.910 ;
        RECT 390.280 520.630 390.560 520.910 ;
        RECT 390.900 520.630 391.180 520.910 ;
        RECT 391.520 520.630 391.800 520.910 ;
        RECT 392.140 520.630 392.420 520.910 ;
        RECT 392.760 520.630 393.040 520.910 ;
        RECT 389.040 520.010 389.320 520.290 ;
        RECT 389.660 520.010 389.940 520.290 ;
        RECT 390.280 520.010 390.560 520.290 ;
        RECT 390.900 520.010 391.180 520.290 ;
        RECT 391.520 520.010 391.800 520.290 ;
        RECT 392.140 520.010 392.420 520.290 ;
        RECT 392.760 520.010 393.040 520.290 ;
        RECT 389.040 519.390 389.320 519.670 ;
        RECT 389.660 519.390 389.940 519.670 ;
        RECT 390.280 519.390 390.560 519.670 ;
        RECT 390.900 519.390 391.180 519.670 ;
        RECT 391.520 519.390 391.800 519.670 ;
        RECT 392.140 519.390 392.420 519.670 ;
        RECT 392.760 519.390 393.040 519.670 ;
        RECT 350.370 515.640 350.650 515.920 ;
        RECT 350.370 515.020 350.650 515.300 ;
        RECT 350.370 514.400 350.650 514.680 ;
        RECT 350.370 513.780 350.650 514.060 ;
        RECT 350.370 513.160 350.650 513.440 ;
        RECT 350.370 512.540 350.650 512.820 ;
        RECT 350.370 511.920 350.650 512.200 ;
        RECT 350.370 511.300 350.650 511.580 ;
        RECT 350.370 510.680 350.650 510.960 ;
        RECT 350.370 510.060 350.650 510.340 ;
        RECT 350.370 509.440 350.650 509.720 ;
        RECT 350.370 508.820 350.650 509.100 ;
        RECT 350.370 508.200 350.650 508.480 ;
        RECT 350.370 507.580 350.650 507.860 ;
        RECT 350.370 506.960 350.650 507.240 ;
        RECT 350.370 506.340 350.650 506.620 ;
        RECT 389.040 515.670 389.320 515.950 ;
        RECT 389.660 515.670 389.940 515.950 ;
        RECT 390.280 515.670 390.560 515.950 ;
        RECT 390.900 515.670 391.180 515.950 ;
        RECT 391.520 515.670 391.800 515.950 ;
        RECT 392.140 515.670 392.420 515.950 ;
        RECT 392.760 515.670 393.040 515.950 ;
        RECT 389.040 515.050 389.320 515.330 ;
        RECT 389.660 515.050 389.940 515.330 ;
        RECT 390.280 515.050 390.560 515.330 ;
        RECT 390.900 515.050 391.180 515.330 ;
        RECT 391.520 515.050 391.800 515.330 ;
        RECT 392.140 515.050 392.420 515.330 ;
        RECT 392.760 515.050 393.040 515.330 ;
        RECT 389.040 514.430 389.320 514.710 ;
        RECT 389.660 514.430 389.940 514.710 ;
        RECT 390.280 514.430 390.560 514.710 ;
        RECT 390.900 514.430 391.180 514.710 ;
        RECT 391.520 514.430 391.800 514.710 ;
        RECT 392.140 514.430 392.420 514.710 ;
        RECT 392.760 514.430 393.040 514.710 ;
        RECT 389.040 513.810 389.320 514.090 ;
        RECT 389.660 513.810 389.940 514.090 ;
        RECT 390.280 513.810 390.560 514.090 ;
        RECT 390.900 513.810 391.180 514.090 ;
        RECT 391.520 513.810 391.800 514.090 ;
        RECT 392.140 513.810 392.420 514.090 ;
        RECT 392.760 513.810 393.040 514.090 ;
        RECT 389.040 513.190 389.320 513.470 ;
        RECT 389.660 513.190 389.940 513.470 ;
        RECT 390.280 513.190 390.560 513.470 ;
        RECT 390.900 513.190 391.180 513.470 ;
        RECT 391.520 513.190 391.800 513.470 ;
        RECT 392.140 513.190 392.420 513.470 ;
        RECT 392.760 513.190 393.040 513.470 ;
        RECT 389.040 512.570 389.320 512.850 ;
        RECT 389.660 512.570 389.940 512.850 ;
        RECT 390.280 512.570 390.560 512.850 ;
        RECT 390.900 512.570 391.180 512.850 ;
        RECT 391.520 512.570 391.800 512.850 ;
        RECT 392.140 512.570 392.420 512.850 ;
        RECT 392.760 512.570 393.040 512.850 ;
        RECT 389.040 511.950 389.320 512.230 ;
        RECT 389.660 511.950 389.940 512.230 ;
        RECT 390.280 511.950 390.560 512.230 ;
        RECT 390.900 511.950 391.180 512.230 ;
        RECT 391.520 511.950 391.800 512.230 ;
        RECT 392.140 511.950 392.420 512.230 ;
        RECT 392.760 511.950 393.040 512.230 ;
        RECT 389.040 511.330 389.320 511.610 ;
        RECT 389.660 511.330 389.940 511.610 ;
        RECT 390.280 511.330 390.560 511.610 ;
        RECT 390.900 511.330 391.180 511.610 ;
        RECT 391.520 511.330 391.800 511.610 ;
        RECT 392.140 511.330 392.420 511.610 ;
        RECT 392.760 511.330 393.040 511.610 ;
        RECT 389.040 510.710 389.320 510.990 ;
        RECT 389.660 510.710 389.940 510.990 ;
        RECT 390.280 510.710 390.560 510.990 ;
        RECT 390.900 510.710 391.180 510.990 ;
        RECT 391.520 510.710 391.800 510.990 ;
        RECT 392.140 510.710 392.420 510.990 ;
        RECT 392.760 510.710 393.040 510.990 ;
        RECT 389.040 510.090 389.320 510.370 ;
        RECT 389.660 510.090 389.940 510.370 ;
        RECT 390.280 510.090 390.560 510.370 ;
        RECT 390.900 510.090 391.180 510.370 ;
        RECT 391.520 510.090 391.800 510.370 ;
        RECT 392.140 510.090 392.420 510.370 ;
        RECT 392.760 510.090 393.040 510.370 ;
        RECT 389.040 509.470 389.320 509.750 ;
        RECT 389.660 509.470 389.940 509.750 ;
        RECT 390.280 509.470 390.560 509.750 ;
        RECT 390.900 509.470 391.180 509.750 ;
        RECT 391.520 509.470 391.800 509.750 ;
        RECT 392.140 509.470 392.420 509.750 ;
        RECT 392.760 509.470 393.040 509.750 ;
        RECT 389.040 508.850 389.320 509.130 ;
        RECT 389.660 508.850 389.940 509.130 ;
        RECT 390.280 508.850 390.560 509.130 ;
        RECT 390.900 508.850 391.180 509.130 ;
        RECT 391.520 508.850 391.800 509.130 ;
        RECT 392.140 508.850 392.420 509.130 ;
        RECT 392.760 508.850 393.040 509.130 ;
        RECT 389.040 508.230 389.320 508.510 ;
        RECT 389.660 508.230 389.940 508.510 ;
        RECT 390.280 508.230 390.560 508.510 ;
        RECT 390.900 508.230 391.180 508.510 ;
        RECT 391.520 508.230 391.800 508.510 ;
        RECT 392.140 508.230 392.420 508.510 ;
        RECT 392.760 508.230 393.040 508.510 ;
        RECT 389.040 507.610 389.320 507.890 ;
        RECT 389.660 507.610 389.940 507.890 ;
        RECT 390.280 507.610 390.560 507.890 ;
        RECT 390.900 507.610 391.180 507.890 ;
        RECT 391.520 507.610 391.800 507.890 ;
        RECT 392.140 507.610 392.420 507.890 ;
        RECT 392.760 507.610 393.040 507.890 ;
        RECT 389.040 506.990 389.320 507.270 ;
        RECT 389.660 506.990 389.940 507.270 ;
        RECT 390.280 506.990 390.560 507.270 ;
        RECT 390.900 506.990 391.180 507.270 ;
        RECT 391.520 506.990 391.800 507.270 ;
        RECT 392.140 506.990 392.420 507.270 ;
        RECT 392.760 506.990 393.040 507.270 ;
        RECT 389.040 506.370 389.320 506.650 ;
        RECT 389.660 506.370 389.940 506.650 ;
        RECT 390.280 506.370 390.560 506.650 ;
        RECT 390.900 506.370 391.180 506.650 ;
        RECT 391.520 506.370 391.800 506.650 ;
        RECT 392.140 506.370 392.420 506.650 ;
        RECT 392.760 506.370 393.040 506.650 ;
        RECT 350.370 503.790 350.650 504.070 ;
        RECT 350.370 503.170 350.650 503.450 ;
        RECT 350.370 502.550 350.650 502.830 ;
        RECT 350.370 501.930 350.650 502.210 ;
        RECT 350.370 501.310 350.650 501.590 ;
        RECT 350.370 500.690 350.650 500.970 ;
        RECT 350.370 500.070 350.650 500.350 ;
        RECT 350.370 499.450 350.650 499.730 ;
        RECT 350.370 498.830 350.650 499.110 ;
        RECT 350.370 498.210 350.650 498.490 ;
        RECT 350.370 497.590 350.650 497.870 ;
        RECT 350.370 496.970 350.650 497.250 ;
        RECT 350.370 496.350 350.650 496.630 ;
        RECT 350.370 495.730 350.650 496.010 ;
        RECT 350.370 495.110 350.650 495.390 ;
        RECT 350.370 494.490 350.650 494.770 ;
        RECT 389.040 503.820 389.320 504.100 ;
        RECT 389.660 503.820 389.940 504.100 ;
        RECT 390.280 503.820 390.560 504.100 ;
        RECT 390.900 503.820 391.180 504.100 ;
        RECT 391.520 503.820 391.800 504.100 ;
        RECT 392.140 503.820 392.420 504.100 ;
        RECT 392.760 503.820 393.040 504.100 ;
        RECT 389.040 503.200 389.320 503.480 ;
        RECT 389.660 503.200 389.940 503.480 ;
        RECT 390.280 503.200 390.560 503.480 ;
        RECT 390.900 503.200 391.180 503.480 ;
        RECT 391.520 503.200 391.800 503.480 ;
        RECT 392.140 503.200 392.420 503.480 ;
        RECT 392.760 503.200 393.040 503.480 ;
        RECT 389.040 502.580 389.320 502.860 ;
        RECT 389.660 502.580 389.940 502.860 ;
        RECT 390.280 502.580 390.560 502.860 ;
        RECT 390.900 502.580 391.180 502.860 ;
        RECT 391.520 502.580 391.800 502.860 ;
        RECT 392.140 502.580 392.420 502.860 ;
        RECT 392.760 502.580 393.040 502.860 ;
        RECT 389.040 501.960 389.320 502.240 ;
        RECT 389.660 501.960 389.940 502.240 ;
        RECT 390.280 501.960 390.560 502.240 ;
        RECT 390.900 501.960 391.180 502.240 ;
        RECT 391.520 501.960 391.800 502.240 ;
        RECT 392.140 501.960 392.420 502.240 ;
        RECT 392.760 501.960 393.040 502.240 ;
        RECT 389.040 501.340 389.320 501.620 ;
        RECT 389.660 501.340 389.940 501.620 ;
        RECT 390.280 501.340 390.560 501.620 ;
        RECT 390.900 501.340 391.180 501.620 ;
        RECT 391.520 501.340 391.800 501.620 ;
        RECT 392.140 501.340 392.420 501.620 ;
        RECT 392.760 501.340 393.040 501.620 ;
        RECT 389.040 500.720 389.320 501.000 ;
        RECT 389.660 500.720 389.940 501.000 ;
        RECT 390.280 500.720 390.560 501.000 ;
        RECT 390.900 500.720 391.180 501.000 ;
        RECT 391.520 500.720 391.800 501.000 ;
        RECT 392.140 500.720 392.420 501.000 ;
        RECT 392.760 500.720 393.040 501.000 ;
        RECT 389.040 500.100 389.320 500.380 ;
        RECT 389.660 500.100 389.940 500.380 ;
        RECT 390.280 500.100 390.560 500.380 ;
        RECT 390.900 500.100 391.180 500.380 ;
        RECT 391.520 500.100 391.800 500.380 ;
        RECT 392.140 500.100 392.420 500.380 ;
        RECT 392.760 500.100 393.040 500.380 ;
        RECT 389.040 499.480 389.320 499.760 ;
        RECT 389.660 499.480 389.940 499.760 ;
        RECT 390.280 499.480 390.560 499.760 ;
        RECT 390.900 499.480 391.180 499.760 ;
        RECT 391.520 499.480 391.800 499.760 ;
        RECT 392.140 499.480 392.420 499.760 ;
        RECT 392.760 499.480 393.040 499.760 ;
        RECT 389.040 498.860 389.320 499.140 ;
        RECT 389.660 498.860 389.940 499.140 ;
        RECT 390.280 498.860 390.560 499.140 ;
        RECT 390.900 498.860 391.180 499.140 ;
        RECT 391.520 498.860 391.800 499.140 ;
        RECT 392.140 498.860 392.420 499.140 ;
        RECT 392.760 498.860 393.040 499.140 ;
        RECT 389.040 498.240 389.320 498.520 ;
        RECT 389.660 498.240 389.940 498.520 ;
        RECT 390.280 498.240 390.560 498.520 ;
        RECT 390.900 498.240 391.180 498.520 ;
        RECT 391.520 498.240 391.800 498.520 ;
        RECT 392.140 498.240 392.420 498.520 ;
        RECT 392.760 498.240 393.040 498.520 ;
        RECT 389.040 497.620 389.320 497.900 ;
        RECT 389.660 497.620 389.940 497.900 ;
        RECT 390.280 497.620 390.560 497.900 ;
        RECT 390.900 497.620 391.180 497.900 ;
        RECT 391.520 497.620 391.800 497.900 ;
        RECT 392.140 497.620 392.420 497.900 ;
        RECT 392.760 497.620 393.040 497.900 ;
        RECT 389.040 497.000 389.320 497.280 ;
        RECT 389.660 497.000 389.940 497.280 ;
        RECT 390.280 497.000 390.560 497.280 ;
        RECT 390.900 497.000 391.180 497.280 ;
        RECT 391.520 497.000 391.800 497.280 ;
        RECT 392.140 497.000 392.420 497.280 ;
        RECT 392.760 497.000 393.040 497.280 ;
        RECT 389.040 496.380 389.320 496.660 ;
        RECT 389.660 496.380 389.940 496.660 ;
        RECT 390.280 496.380 390.560 496.660 ;
        RECT 390.900 496.380 391.180 496.660 ;
        RECT 391.520 496.380 391.800 496.660 ;
        RECT 392.140 496.380 392.420 496.660 ;
        RECT 392.760 496.380 393.040 496.660 ;
        RECT 389.040 495.760 389.320 496.040 ;
        RECT 389.660 495.760 389.940 496.040 ;
        RECT 390.280 495.760 390.560 496.040 ;
        RECT 390.900 495.760 391.180 496.040 ;
        RECT 391.520 495.760 391.800 496.040 ;
        RECT 392.140 495.760 392.420 496.040 ;
        RECT 392.760 495.760 393.040 496.040 ;
        RECT 389.040 495.140 389.320 495.420 ;
        RECT 389.660 495.140 389.940 495.420 ;
        RECT 390.280 495.140 390.560 495.420 ;
        RECT 390.900 495.140 391.180 495.420 ;
        RECT 391.520 495.140 391.800 495.420 ;
        RECT 392.140 495.140 392.420 495.420 ;
        RECT 392.760 495.140 393.040 495.420 ;
        RECT 389.040 494.520 389.320 494.800 ;
        RECT 389.660 494.520 389.940 494.800 ;
        RECT 390.280 494.520 390.560 494.800 ;
        RECT 390.900 494.520 391.180 494.800 ;
        RECT 391.520 494.520 391.800 494.800 ;
        RECT 392.140 494.520 392.420 494.800 ;
        RECT 392.760 494.520 393.040 494.800 ;
        RECT 350.370 490.260 350.650 490.540 ;
        RECT 350.370 489.640 350.650 489.920 ;
        RECT 350.370 489.020 350.650 489.300 ;
        RECT 350.370 488.400 350.650 488.680 ;
        RECT 350.370 487.780 350.650 488.060 ;
        RECT 350.370 487.160 350.650 487.440 ;
        RECT 350.370 486.540 350.650 486.820 ;
        RECT 350.370 485.920 350.650 486.200 ;
        RECT 350.370 485.300 350.650 485.580 ;
        RECT 350.370 484.680 350.650 484.960 ;
        RECT 350.370 484.060 350.650 484.340 ;
        RECT 350.370 483.440 350.650 483.720 ;
        RECT 350.370 482.820 350.650 483.100 ;
        RECT 350.370 482.200 350.650 482.480 ;
        RECT 350.370 481.580 350.650 481.860 ;
        RECT 350.370 480.960 350.650 481.240 ;
        RECT 389.040 490.290 389.320 490.570 ;
        RECT 389.660 490.290 389.940 490.570 ;
        RECT 390.280 490.290 390.560 490.570 ;
        RECT 390.900 490.290 391.180 490.570 ;
        RECT 391.520 490.290 391.800 490.570 ;
        RECT 392.140 490.290 392.420 490.570 ;
        RECT 392.760 490.290 393.040 490.570 ;
        RECT 389.040 489.670 389.320 489.950 ;
        RECT 389.660 489.670 389.940 489.950 ;
        RECT 390.280 489.670 390.560 489.950 ;
        RECT 390.900 489.670 391.180 489.950 ;
        RECT 391.520 489.670 391.800 489.950 ;
        RECT 392.140 489.670 392.420 489.950 ;
        RECT 392.760 489.670 393.040 489.950 ;
        RECT 389.040 489.050 389.320 489.330 ;
        RECT 389.660 489.050 389.940 489.330 ;
        RECT 390.280 489.050 390.560 489.330 ;
        RECT 390.900 489.050 391.180 489.330 ;
        RECT 391.520 489.050 391.800 489.330 ;
        RECT 392.140 489.050 392.420 489.330 ;
        RECT 392.760 489.050 393.040 489.330 ;
        RECT 389.040 488.430 389.320 488.710 ;
        RECT 389.660 488.430 389.940 488.710 ;
        RECT 390.280 488.430 390.560 488.710 ;
        RECT 390.900 488.430 391.180 488.710 ;
        RECT 391.520 488.430 391.800 488.710 ;
        RECT 392.140 488.430 392.420 488.710 ;
        RECT 392.760 488.430 393.040 488.710 ;
        RECT 389.040 487.810 389.320 488.090 ;
        RECT 389.660 487.810 389.940 488.090 ;
        RECT 390.280 487.810 390.560 488.090 ;
        RECT 390.900 487.810 391.180 488.090 ;
        RECT 391.520 487.810 391.800 488.090 ;
        RECT 392.140 487.810 392.420 488.090 ;
        RECT 392.760 487.810 393.040 488.090 ;
        RECT 389.040 487.190 389.320 487.470 ;
        RECT 389.660 487.190 389.940 487.470 ;
        RECT 390.280 487.190 390.560 487.470 ;
        RECT 390.900 487.190 391.180 487.470 ;
        RECT 391.520 487.190 391.800 487.470 ;
        RECT 392.140 487.190 392.420 487.470 ;
        RECT 392.760 487.190 393.040 487.470 ;
        RECT 389.040 486.570 389.320 486.850 ;
        RECT 389.660 486.570 389.940 486.850 ;
        RECT 390.280 486.570 390.560 486.850 ;
        RECT 390.900 486.570 391.180 486.850 ;
        RECT 391.520 486.570 391.800 486.850 ;
        RECT 392.140 486.570 392.420 486.850 ;
        RECT 392.760 486.570 393.040 486.850 ;
        RECT 389.040 485.950 389.320 486.230 ;
        RECT 389.660 485.950 389.940 486.230 ;
        RECT 390.280 485.950 390.560 486.230 ;
        RECT 390.900 485.950 391.180 486.230 ;
        RECT 391.520 485.950 391.800 486.230 ;
        RECT 392.140 485.950 392.420 486.230 ;
        RECT 392.760 485.950 393.040 486.230 ;
        RECT 389.040 485.330 389.320 485.610 ;
        RECT 389.660 485.330 389.940 485.610 ;
        RECT 390.280 485.330 390.560 485.610 ;
        RECT 390.900 485.330 391.180 485.610 ;
        RECT 391.520 485.330 391.800 485.610 ;
        RECT 392.140 485.330 392.420 485.610 ;
        RECT 392.760 485.330 393.040 485.610 ;
        RECT 389.040 484.710 389.320 484.990 ;
        RECT 389.660 484.710 389.940 484.990 ;
        RECT 390.280 484.710 390.560 484.990 ;
        RECT 390.900 484.710 391.180 484.990 ;
        RECT 391.520 484.710 391.800 484.990 ;
        RECT 392.140 484.710 392.420 484.990 ;
        RECT 392.760 484.710 393.040 484.990 ;
        RECT 389.040 484.090 389.320 484.370 ;
        RECT 389.660 484.090 389.940 484.370 ;
        RECT 390.280 484.090 390.560 484.370 ;
        RECT 390.900 484.090 391.180 484.370 ;
        RECT 391.520 484.090 391.800 484.370 ;
        RECT 392.140 484.090 392.420 484.370 ;
        RECT 392.760 484.090 393.040 484.370 ;
        RECT 389.040 483.470 389.320 483.750 ;
        RECT 389.660 483.470 389.940 483.750 ;
        RECT 390.280 483.470 390.560 483.750 ;
        RECT 390.900 483.470 391.180 483.750 ;
        RECT 391.520 483.470 391.800 483.750 ;
        RECT 392.140 483.470 392.420 483.750 ;
        RECT 392.760 483.470 393.040 483.750 ;
        RECT 389.040 482.850 389.320 483.130 ;
        RECT 389.660 482.850 389.940 483.130 ;
        RECT 390.280 482.850 390.560 483.130 ;
        RECT 390.900 482.850 391.180 483.130 ;
        RECT 391.520 482.850 391.800 483.130 ;
        RECT 392.140 482.850 392.420 483.130 ;
        RECT 392.760 482.850 393.040 483.130 ;
        RECT 389.040 482.230 389.320 482.510 ;
        RECT 389.660 482.230 389.940 482.510 ;
        RECT 390.280 482.230 390.560 482.510 ;
        RECT 390.900 482.230 391.180 482.510 ;
        RECT 391.520 482.230 391.800 482.510 ;
        RECT 392.140 482.230 392.420 482.510 ;
        RECT 392.760 482.230 393.040 482.510 ;
        RECT 389.040 481.610 389.320 481.890 ;
        RECT 389.660 481.610 389.940 481.890 ;
        RECT 390.280 481.610 390.560 481.890 ;
        RECT 390.900 481.610 391.180 481.890 ;
        RECT 391.520 481.610 391.800 481.890 ;
        RECT 392.140 481.610 392.420 481.890 ;
        RECT 392.760 481.610 393.040 481.890 ;
        RECT 389.040 480.990 389.320 481.270 ;
        RECT 389.660 480.990 389.940 481.270 ;
        RECT 390.280 480.990 390.560 481.270 ;
        RECT 390.900 480.990 391.180 481.270 ;
        RECT 391.520 480.990 391.800 481.270 ;
        RECT 392.140 480.990 392.420 481.270 ;
        RECT 392.760 480.990 393.040 481.270 ;
        RECT 350.370 478.410 350.650 478.690 ;
        RECT 350.370 477.790 350.650 478.070 ;
        RECT 350.370 477.170 350.650 477.450 ;
        RECT 350.370 476.550 350.650 476.830 ;
        RECT 350.370 475.930 350.650 476.210 ;
        RECT 350.370 475.310 350.650 475.590 ;
        RECT 350.370 474.690 350.650 474.970 ;
        RECT 350.370 474.070 350.650 474.350 ;
        RECT 350.370 473.450 350.650 473.730 ;
        RECT 350.370 472.830 350.650 473.110 ;
        RECT 350.370 472.210 350.650 472.490 ;
        RECT 350.370 471.590 350.650 471.870 ;
        RECT 350.370 470.970 350.650 471.250 ;
        RECT 350.370 470.350 350.650 470.630 ;
        RECT 350.370 469.730 350.650 470.010 ;
        RECT 350.370 469.110 350.650 469.390 ;
        RECT 389.040 478.440 389.320 478.720 ;
        RECT 389.660 478.440 389.940 478.720 ;
        RECT 390.280 478.440 390.560 478.720 ;
        RECT 390.900 478.440 391.180 478.720 ;
        RECT 391.520 478.440 391.800 478.720 ;
        RECT 392.140 478.440 392.420 478.720 ;
        RECT 392.760 478.440 393.040 478.720 ;
        RECT 389.040 477.820 389.320 478.100 ;
        RECT 389.660 477.820 389.940 478.100 ;
        RECT 390.280 477.820 390.560 478.100 ;
        RECT 390.900 477.820 391.180 478.100 ;
        RECT 391.520 477.820 391.800 478.100 ;
        RECT 392.140 477.820 392.420 478.100 ;
        RECT 392.760 477.820 393.040 478.100 ;
        RECT 389.040 477.200 389.320 477.480 ;
        RECT 389.660 477.200 389.940 477.480 ;
        RECT 390.280 477.200 390.560 477.480 ;
        RECT 390.900 477.200 391.180 477.480 ;
        RECT 391.520 477.200 391.800 477.480 ;
        RECT 392.140 477.200 392.420 477.480 ;
        RECT 392.760 477.200 393.040 477.480 ;
        RECT 389.040 476.580 389.320 476.860 ;
        RECT 389.660 476.580 389.940 476.860 ;
        RECT 390.280 476.580 390.560 476.860 ;
        RECT 390.900 476.580 391.180 476.860 ;
        RECT 391.520 476.580 391.800 476.860 ;
        RECT 392.140 476.580 392.420 476.860 ;
        RECT 392.760 476.580 393.040 476.860 ;
        RECT 389.040 475.960 389.320 476.240 ;
        RECT 389.660 475.960 389.940 476.240 ;
        RECT 390.280 475.960 390.560 476.240 ;
        RECT 390.900 475.960 391.180 476.240 ;
        RECT 391.520 475.960 391.800 476.240 ;
        RECT 392.140 475.960 392.420 476.240 ;
        RECT 392.760 475.960 393.040 476.240 ;
        RECT 389.040 475.340 389.320 475.620 ;
        RECT 389.660 475.340 389.940 475.620 ;
        RECT 390.280 475.340 390.560 475.620 ;
        RECT 390.900 475.340 391.180 475.620 ;
        RECT 391.520 475.340 391.800 475.620 ;
        RECT 392.140 475.340 392.420 475.620 ;
        RECT 392.760 475.340 393.040 475.620 ;
        RECT 389.040 474.720 389.320 475.000 ;
        RECT 389.660 474.720 389.940 475.000 ;
        RECT 390.280 474.720 390.560 475.000 ;
        RECT 390.900 474.720 391.180 475.000 ;
        RECT 391.520 474.720 391.800 475.000 ;
        RECT 392.140 474.720 392.420 475.000 ;
        RECT 392.760 474.720 393.040 475.000 ;
        RECT 389.040 474.100 389.320 474.380 ;
        RECT 389.660 474.100 389.940 474.380 ;
        RECT 390.280 474.100 390.560 474.380 ;
        RECT 390.900 474.100 391.180 474.380 ;
        RECT 391.520 474.100 391.800 474.380 ;
        RECT 392.140 474.100 392.420 474.380 ;
        RECT 392.760 474.100 393.040 474.380 ;
        RECT 389.040 473.480 389.320 473.760 ;
        RECT 389.660 473.480 389.940 473.760 ;
        RECT 390.280 473.480 390.560 473.760 ;
        RECT 390.900 473.480 391.180 473.760 ;
        RECT 391.520 473.480 391.800 473.760 ;
        RECT 392.140 473.480 392.420 473.760 ;
        RECT 392.760 473.480 393.040 473.760 ;
        RECT 389.040 472.860 389.320 473.140 ;
        RECT 389.660 472.860 389.940 473.140 ;
        RECT 390.280 472.860 390.560 473.140 ;
        RECT 390.900 472.860 391.180 473.140 ;
        RECT 391.520 472.860 391.800 473.140 ;
        RECT 392.140 472.860 392.420 473.140 ;
        RECT 392.760 472.860 393.040 473.140 ;
        RECT 389.040 472.240 389.320 472.520 ;
        RECT 389.660 472.240 389.940 472.520 ;
        RECT 390.280 472.240 390.560 472.520 ;
        RECT 390.900 472.240 391.180 472.520 ;
        RECT 391.520 472.240 391.800 472.520 ;
        RECT 392.140 472.240 392.420 472.520 ;
        RECT 392.760 472.240 393.040 472.520 ;
        RECT 389.040 471.620 389.320 471.900 ;
        RECT 389.660 471.620 389.940 471.900 ;
        RECT 390.280 471.620 390.560 471.900 ;
        RECT 390.900 471.620 391.180 471.900 ;
        RECT 391.520 471.620 391.800 471.900 ;
        RECT 392.140 471.620 392.420 471.900 ;
        RECT 392.760 471.620 393.040 471.900 ;
        RECT 389.040 471.000 389.320 471.280 ;
        RECT 389.660 471.000 389.940 471.280 ;
        RECT 390.280 471.000 390.560 471.280 ;
        RECT 390.900 471.000 391.180 471.280 ;
        RECT 391.520 471.000 391.800 471.280 ;
        RECT 392.140 471.000 392.420 471.280 ;
        RECT 392.760 471.000 393.040 471.280 ;
        RECT 389.040 470.380 389.320 470.660 ;
        RECT 389.660 470.380 389.940 470.660 ;
        RECT 390.280 470.380 390.560 470.660 ;
        RECT 390.900 470.380 391.180 470.660 ;
        RECT 391.520 470.380 391.800 470.660 ;
        RECT 392.140 470.380 392.420 470.660 ;
        RECT 392.760 470.380 393.040 470.660 ;
        RECT 389.040 469.760 389.320 470.040 ;
        RECT 389.660 469.760 389.940 470.040 ;
        RECT 390.280 469.760 390.560 470.040 ;
        RECT 390.900 469.760 391.180 470.040 ;
        RECT 391.520 469.760 391.800 470.040 ;
        RECT 392.140 469.760 392.420 470.040 ;
        RECT 392.760 469.760 393.040 470.040 ;
        RECT 389.040 469.140 389.320 469.420 ;
        RECT 389.660 469.140 389.940 469.420 ;
        RECT 390.280 469.140 390.560 469.420 ;
        RECT 390.900 469.140 391.180 469.420 ;
        RECT 391.520 469.140 391.800 469.420 ;
        RECT 392.140 469.140 392.420 469.420 ;
        RECT 392.760 469.140 393.040 469.420 ;
        RECT 350.370 465.390 350.650 465.670 ;
        RECT 350.370 464.770 350.650 465.050 ;
        RECT 350.370 464.150 350.650 464.430 ;
        RECT 350.370 463.530 350.650 463.810 ;
        RECT 350.370 462.910 350.650 463.190 ;
        RECT 350.370 462.290 350.650 462.570 ;
        RECT 350.370 461.670 350.650 461.950 ;
        RECT 350.370 461.050 350.650 461.330 ;
        RECT 350.370 460.430 350.650 460.710 ;
        RECT 350.370 459.810 350.650 460.090 ;
        RECT 350.370 459.190 350.650 459.470 ;
        RECT 350.370 458.570 350.650 458.850 ;
        RECT 350.370 457.950 350.650 458.230 ;
        RECT 350.370 457.330 350.650 457.610 ;
        RECT 350.370 456.710 350.650 456.990 ;
        RECT 389.040 465.420 389.320 465.700 ;
        RECT 389.660 465.420 389.940 465.700 ;
        RECT 390.280 465.420 390.560 465.700 ;
        RECT 390.900 465.420 391.180 465.700 ;
        RECT 391.520 465.420 391.800 465.700 ;
        RECT 392.140 465.420 392.420 465.700 ;
        RECT 392.760 465.420 393.040 465.700 ;
        RECT 389.040 464.800 389.320 465.080 ;
        RECT 389.660 464.800 389.940 465.080 ;
        RECT 390.280 464.800 390.560 465.080 ;
        RECT 390.900 464.800 391.180 465.080 ;
        RECT 391.520 464.800 391.800 465.080 ;
        RECT 392.140 464.800 392.420 465.080 ;
        RECT 392.760 464.800 393.040 465.080 ;
        RECT 389.040 464.180 389.320 464.460 ;
        RECT 389.660 464.180 389.940 464.460 ;
        RECT 390.280 464.180 390.560 464.460 ;
        RECT 390.900 464.180 391.180 464.460 ;
        RECT 391.520 464.180 391.800 464.460 ;
        RECT 392.140 464.180 392.420 464.460 ;
        RECT 392.760 464.180 393.040 464.460 ;
        RECT 389.040 463.560 389.320 463.840 ;
        RECT 389.660 463.560 389.940 463.840 ;
        RECT 390.280 463.560 390.560 463.840 ;
        RECT 390.900 463.560 391.180 463.840 ;
        RECT 391.520 463.560 391.800 463.840 ;
        RECT 392.140 463.560 392.420 463.840 ;
        RECT 392.760 463.560 393.040 463.840 ;
        RECT 389.040 462.940 389.320 463.220 ;
        RECT 389.660 462.940 389.940 463.220 ;
        RECT 390.280 462.940 390.560 463.220 ;
        RECT 390.900 462.940 391.180 463.220 ;
        RECT 391.520 462.940 391.800 463.220 ;
        RECT 392.140 462.940 392.420 463.220 ;
        RECT 392.760 462.940 393.040 463.220 ;
        RECT 389.040 462.320 389.320 462.600 ;
        RECT 389.660 462.320 389.940 462.600 ;
        RECT 390.280 462.320 390.560 462.600 ;
        RECT 390.900 462.320 391.180 462.600 ;
        RECT 391.520 462.320 391.800 462.600 ;
        RECT 392.140 462.320 392.420 462.600 ;
        RECT 392.760 462.320 393.040 462.600 ;
        RECT 389.040 461.700 389.320 461.980 ;
        RECT 389.660 461.700 389.940 461.980 ;
        RECT 390.280 461.700 390.560 461.980 ;
        RECT 390.900 461.700 391.180 461.980 ;
        RECT 391.520 461.700 391.800 461.980 ;
        RECT 392.140 461.700 392.420 461.980 ;
        RECT 392.760 461.700 393.040 461.980 ;
        RECT 389.040 461.080 389.320 461.360 ;
        RECT 389.660 461.080 389.940 461.360 ;
        RECT 390.280 461.080 390.560 461.360 ;
        RECT 390.900 461.080 391.180 461.360 ;
        RECT 391.520 461.080 391.800 461.360 ;
        RECT 392.140 461.080 392.420 461.360 ;
        RECT 392.760 461.080 393.040 461.360 ;
        RECT 389.040 460.460 389.320 460.740 ;
        RECT 389.660 460.460 389.940 460.740 ;
        RECT 390.280 460.460 390.560 460.740 ;
        RECT 390.900 460.460 391.180 460.740 ;
        RECT 391.520 460.460 391.800 460.740 ;
        RECT 392.140 460.460 392.420 460.740 ;
        RECT 392.760 460.460 393.040 460.740 ;
        RECT 389.040 459.840 389.320 460.120 ;
        RECT 389.660 459.840 389.940 460.120 ;
        RECT 390.280 459.840 390.560 460.120 ;
        RECT 390.900 459.840 391.180 460.120 ;
        RECT 391.520 459.840 391.800 460.120 ;
        RECT 392.140 459.840 392.420 460.120 ;
        RECT 392.760 459.840 393.040 460.120 ;
        RECT 389.040 459.220 389.320 459.500 ;
        RECT 389.660 459.220 389.940 459.500 ;
        RECT 390.280 459.220 390.560 459.500 ;
        RECT 390.900 459.220 391.180 459.500 ;
        RECT 391.520 459.220 391.800 459.500 ;
        RECT 392.140 459.220 392.420 459.500 ;
        RECT 392.760 459.220 393.040 459.500 ;
        RECT 389.040 458.600 389.320 458.880 ;
        RECT 389.660 458.600 389.940 458.880 ;
        RECT 390.280 458.600 390.560 458.880 ;
        RECT 390.900 458.600 391.180 458.880 ;
        RECT 391.520 458.600 391.800 458.880 ;
        RECT 392.140 458.600 392.420 458.880 ;
        RECT 392.760 458.600 393.040 458.880 ;
        RECT 389.040 457.980 389.320 458.260 ;
        RECT 389.660 457.980 389.940 458.260 ;
        RECT 390.280 457.980 390.560 458.260 ;
        RECT 390.900 457.980 391.180 458.260 ;
        RECT 391.520 457.980 391.800 458.260 ;
        RECT 392.140 457.980 392.420 458.260 ;
        RECT 392.760 457.980 393.040 458.260 ;
        RECT 389.040 457.360 389.320 457.640 ;
        RECT 389.660 457.360 389.940 457.640 ;
        RECT 390.280 457.360 390.560 457.640 ;
        RECT 390.900 457.360 391.180 457.640 ;
        RECT 391.520 457.360 391.800 457.640 ;
        RECT 392.140 457.360 392.420 457.640 ;
        RECT 392.760 457.360 393.040 457.640 ;
        RECT 389.040 456.740 389.320 457.020 ;
        RECT 389.660 456.740 389.940 457.020 ;
        RECT 390.280 456.740 390.560 457.020 ;
        RECT 390.900 456.740 391.180 457.020 ;
        RECT 391.520 456.740 391.800 457.020 ;
        RECT 392.140 456.740 392.420 457.020 ;
        RECT 392.760 456.740 393.040 457.020 ;
        RECT 388.740 431.580 389.020 431.860 ;
        RECT 389.360 431.580 389.640 431.860 ;
        RECT 389.980 431.580 390.260 431.860 ;
        RECT 390.600 431.580 390.880 431.860 ;
        RECT 391.220 431.580 391.500 431.860 ;
        RECT 391.840 431.580 392.120 431.860 ;
        RECT 392.460 431.580 392.740 431.860 ;
        RECT 388.740 430.960 389.020 431.240 ;
        RECT 389.360 430.960 389.640 431.240 ;
        RECT 389.980 430.960 390.260 431.240 ;
        RECT 390.600 430.960 390.880 431.240 ;
        RECT 391.220 430.960 391.500 431.240 ;
        RECT 391.840 430.960 392.120 431.240 ;
        RECT 392.460 430.960 392.740 431.240 ;
        RECT 552.740 4716.895 553.020 4717.175 ;
        RECT 395.740 4703.980 396.020 4704.260 ;
        RECT 396.360 4703.980 396.640 4704.260 ;
        RECT 396.980 4703.980 397.260 4704.260 ;
        RECT 397.600 4703.980 397.880 4704.260 ;
        RECT 398.220 4703.980 398.500 4704.260 ;
        RECT 398.840 4703.980 399.120 4704.260 ;
        RECT 399.460 4703.980 399.740 4704.260 ;
        RECT 395.740 4703.360 396.020 4703.640 ;
        RECT 396.360 4703.360 396.640 4703.640 ;
        RECT 396.980 4703.360 397.260 4703.640 ;
        RECT 397.600 4703.360 397.880 4703.640 ;
        RECT 398.220 4703.360 398.500 4703.640 ;
        RECT 398.840 4703.360 399.120 4703.640 ;
        RECT 399.460 4703.360 399.740 4703.640 ;
        RECT 395.740 4702.740 396.020 4703.020 ;
        RECT 396.360 4702.740 396.640 4703.020 ;
        RECT 396.980 4702.740 397.260 4703.020 ;
        RECT 397.600 4702.740 397.880 4703.020 ;
        RECT 398.220 4702.740 398.500 4703.020 ;
        RECT 398.840 4702.740 399.120 4703.020 ;
        RECT 399.460 4702.740 399.740 4703.020 ;
        RECT 395.740 4702.120 396.020 4702.400 ;
        RECT 396.360 4702.120 396.640 4702.400 ;
        RECT 396.980 4702.120 397.260 4702.400 ;
        RECT 397.600 4702.120 397.880 4702.400 ;
        RECT 398.220 4702.120 398.500 4702.400 ;
        RECT 398.840 4702.120 399.120 4702.400 ;
        RECT 399.460 4702.120 399.740 4702.400 ;
        RECT 395.740 4701.500 396.020 4701.780 ;
        RECT 396.360 4701.500 396.640 4701.780 ;
        RECT 396.980 4701.500 397.260 4701.780 ;
        RECT 397.600 4701.500 397.880 4701.780 ;
        RECT 398.220 4701.500 398.500 4701.780 ;
        RECT 398.840 4701.500 399.120 4701.780 ;
        RECT 399.460 4701.500 399.740 4701.780 ;
        RECT 395.740 4700.880 396.020 4701.160 ;
        RECT 396.360 4700.880 396.640 4701.160 ;
        RECT 396.980 4700.880 397.260 4701.160 ;
        RECT 397.600 4700.880 397.880 4701.160 ;
        RECT 398.220 4700.880 398.500 4701.160 ;
        RECT 398.840 4700.880 399.120 4701.160 ;
        RECT 399.460 4700.880 399.740 4701.160 ;
        RECT 395.740 4700.260 396.020 4700.540 ;
        RECT 396.360 4700.260 396.640 4700.540 ;
        RECT 396.980 4700.260 397.260 4700.540 ;
        RECT 397.600 4700.260 397.880 4700.540 ;
        RECT 398.220 4700.260 398.500 4700.540 ;
        RECT 398.840 4700.260 399.120 4700.540 ;
        RECT 399.460 4700.260 399.740 4700.540 ;
        RECT 441.035 4710.720 441.315 4711.000 ;
        RECT 442.035 4710.720 442.315 4711.000 ;
        RECT 441.035 4709.220 441.315 4709.500 ;
        RECT 442.035 4709.220 442.315 4709.500 ;
        RECT 441.035 4707.720 441.315 4708.000 ;
        RECT 442.035 4707.720 442.315 4708.000 ;
        RECT 531.035 4703.720 531.315 4704.000 ;
        RECT 532.035 4703.720 532.315 4704.000 ;
        RECT 531.035 4702.220 531.315 4702.500 ;
        RECT 532.035 4702.220 532.315 4702.500 ;
        RECT 531.035 4700.720 531.315 4701.000 ;
        RECT 532.035 4700.720 532.315 4701.000 ;
        RECT 552.730 4703.270 553.010 4703.550 ;
        RECT 552.730 4701.770 553.010 4702.050 ;
        RECT 552.730 4700.270 553.010 4700.550 ;
        RECT 587.740 4716.895 588.020 4717.175 ;
        RECT 587.730 4703.270 588.010 4703.550 ;
        RECT 587.730 4701.770 588.010 4702.050 ;
        RECT 587.730 4700.270 588.010 4700.550 ;
        RECT 622.740 4716.895 623.020 4717.175 ;
        RECT 702.030 4710.485 702.310 4710.765 ;
        RECT 702.030 4708.985 702.310 4709.265 ;
        RECT 702.030 4707.485 702.310 4707.765 ;
        RECT 622.730 4703.270 623.010 4703.550 ;
        RECT 622.730 4701.770 623.010 4702.050 ;
        RECT 622.730 4700.270 623.010 4700.550 ;
        RECT 827.740 4716.895 828.020 4717.175 ;
        RECT 801.035 4710.720 801.315 4711.000 ;
        RECT 802.035 4710.720 802.315 4711.000 ;
        RECT 801.035 4709.220 801.315 4709.500 ;
        RECT 802.035 4709.220 802.315 4709.500 ;
        RECT 801.035 4707.720 801.315 4708.000 ;
        RECT 802.035 4707.720 802.315 4708.000 ;
        RECT 704.105 4703.300 704.385 4703.580 ;
        RECT 704.105 4701.800 704.385 4702.080 ;
        RECT 704.105 4700.300 704.385 4700.580 ;
        RECT 711.035 4703.720 711.315 4704.000 ;
        RECT 712.035 4703.720 712.315 4704.000 ;
        RECT 711.035 4702.220 711.315 4702.500 ;
        RECT 712.035 4702.220 712.315 4702.500 ;
        RECT 711.035 4700.720 711.315 4701.000 ;
        RECT 712.035 4700.720 712.315 4701.000 ;
        RECT 827.730 4703.270 828.010 4703.550 ;
        RECT 827.730 4701.770 828.010 4702.050 ;
        RECT 827.730 4700.270 828.010 4700.550 ;
        RECT 862.740 4716.895 863.020 4717.175 ;
        RECT 897.740 4716.895 898.020 4717.175 ;
        RECT 862.730 4703.270 863.010 4703.550 ;
        RECT 862.730 4701.770 863.010 4702.050 ;
        RECT 862.730 4700.270 863.010 4700.550 ;
        RECT 891.035 4703.720 891.315 4704.000 ;
        RECT 892.035 4703.720 892.315 4704.000 ;
        RECT 891.035 4702.220 891.315 4702.500 ;
        RECT 892.035 4702.220 892.315 4702.500 ;
        RECT 891.035 4700.720 891.315 4701.000 ;
        RECT 892.035 4700.720 892.315 4701.000 ;
        RECT 977.030 4710.485 977.310 4710.765 ;
        RECT 977.030 4708.985 977.310 4709.265 ;
        RECT 977.030 4707.485 977.310 4707.765 ;
        RECT 897.730 4703.270 898.010 4703.550 ;
        RECT 897.730 4701.770 898.010 4702.050 ;
        RECT 897.730 4700.270 898.010 4700.550 ;
        RECT 1102.740 4716.895 1103.020 4717.175 ;
        RECT 979.105 4703.300 979.385 4703.580 ;
        RECT 979.105 4701.800 979.385 4702.080 ;
        RECT 979.105 4700.300 979.385 4700.580 ;
        RECT 1071.035 4703.720 1071.315 4704.000 ;
        RECT 1072.035 4703.720 1072.315 4704.000 ;
        RECT 1071.035 4702.220 1071.315 4702.500 ;
        RECT 1072.035 4702.220 1072.315 4702.500 ;
        RECT 1071.035 4700.720 1071.315 4701.000 ;
        RECT 1072.035 4700.720 1072.315 4701.000 ;
        RECT 1102.730 4703.270 1103.010 4703.550 ;
        RECT 1102.730 4701.770 1103.010 4702.050 ;
        RECT 1102.730 4700.270 1103.010 4700.550 ;
        RECT 1137.740 4716.895 1138.020 4717.175 ;
        RECT 1172.740 4716.895 1173.020 4717.175 ;
        RECT 1137.730 4703.270 1138.010 4703.550 ;
        RECT 1137.730 4701.770 1138.010 4702.050 ;
        RECT 1137.730 4700.270 1138.010 4700.550 ;
        RECT 1161.035 4710.720 1161.315 4711.000 ;
        RECT 1162.035 4710.720 1162.315 4711.000 ;
        RECT 1161.035 4709.220 1161.315 4709.500 ;
        RECT 1162.035 4709.220 1162.315 4709.500 ;
        RECT 1161.035 4707.720 1161.315 4708.000 ;
        RECT 1162.035 4707.720 1162.315 4708.000 ;
        RECT 1252.030 4710.485 1252.310 4710.765 ;
        RECT 1252.030 4708.985 1252.310 4709.265 ;
        RECT 1252.030 4707.485 1252.310 4707.765 ;
        RECT 1172.730 4703.270 1173.010 4703.550 ;
        RECT 1172.730 4701.770 1173.010 4702.050 ;
        RECT 1172.730 4700.270 1173.010 4700.550 ;
        RECT 1251.035 4703.720 1251.315 4704.000 ;
        RECT 1252.035 4703.720 1252.315 4704.000 ;
        RECT 1251.035 4702.220 1251.315 4702.500 ;
        RECT 1252.035 4702.220 1252.315 4702.500 ;
        RECT 1251.035 4700.720 1251.315 4701.000 ;
        RECT 1252.035 4700.720 1252.315 4701.000 ;
        RECT 1377.740 4716.895 1378.020 4717.175 ;
        RECT 1254.105 4703.300 1254.385 4703.580 ;
        RECT 1254.105 4701.800 1254.385 4702.080 ;
        RECT 1254.105 4700.300 1254.385 4700.580 ;
        RECT 1341.035 4710.720 1341.315 4711.000 ;
        RECT 1342.035 4710.720 1342.315 4711.000 ;
        RECT 1341.035 4709.220 1341.315 4709.500 ;
        RECT 1342.035 4709.220 1342.315 4709.500 ;
        RECT 1341.035 4707.720 1341.315 4708.000 ;
        RECT 1342.035 4707.720 1342.315 4708.000 ;
        RECT 1377.730 4703.270 1378.010 4703.550 ;
        RECT 1377.730 4701.770 1378.010 4702.050 ;
        RECT 1377.730 4700.270 1378.010 4700.550 ;
        RECT 1412.740 4716.895 1413.020 4717.175 ;
        RECT 1447.740 4716.895 1448.020 4717.175 ;
        RECT 1412.730 4703.270 1413.010 4703.550 ;
        RECT 1412.730 4701.770 1413.010 4702.050 ;
        RECT 1412.730 4700.270 1413.010 4700.550 ;
        RECT 1431.035 4703.720 1431.315 4704.000 ;
        RECT 1432.035 4703.720 1432.315 4704.000 ;
        RECT 1431.035 4702.220 1431.315 4702.500 ;
        RECT 1432.035 4702.220 1432.315 4702.500 ;
        RECT 1431.035 4700.720 1431.315 4701.000 ;
        RECT 1432.035 4700.720 1432.315 4701.000 ;
        RECT 1447.730 4703.270 1448.010 4703.550 ;
        RECT 1447.730 4701.770 1448.010 4702.050 ;
        RECT 1447.730 4700.270 1448.010 4700.550 ;
        RECT 1521.035 4710.720 1521.315 4711.000 ;
        RECT 1522.035 4710.720 1522.315 4711.000 ;
        RECT 1521.035 4709.220 1521.315 4709.500 ;
        RECT 1522.035 4709.220 1522.315 4709.500 ;
        RECT 1521.035 4707.720 1521.315 4708.000 ;
        RECT 1522.035 4707.720 1522.315 4708.000 ;
        RECT 1527.030 4710.485 1527.310 4710.765 ;
        RECT 1527.030 4708.985 1527.310 4709.265 ;
        RECT 1527.030 4707.485 1527.310 4707.765 ;
        RECT 1652.740 4716.895 1653.020 4717.175 ;
        RECT 1529.105 4703.300 1529.385 4703.580 ;
        RECT 1529.105 4701.800 1529.385 4702.080 ;
        RECT 1529.105 4700.300 1529.385 4700.580 ;
        RECT 1611.035 4703.720 1611.315 4704.000 ;
        RECT 1612.035 4703.720 1612.315 4704.000 ;
        RECT 1611.035 4702.220 1611.315 4702.500 ;
        RECT 1612.035 4702.220 1612.315 4702.500 ;
        RECT 1611.035 4700.720 1611.315 4701.000 ;
        RECT 1612.035 4700.720 1612.315 4701.000 ;
        RECT 1652.730 4703.270 1653.010 4703.550 ;
        RECT 1652.730 4701.770 1653.010 4702.050 ;
        RECT 1652.730 4700.270 1653.010 4700.550 ;
        RECT 1687.740 4716.895 1688.020 4717.175 ;
        RECT 1722.740 4716.895 1723.020 4717.175 ;
        RECT 1687.730 4703.270 1688.010 4703.550 ;
        RECT 1687.730 4701.770 1688.010 4702.050 ;
        RECT 1687.730 4700.270 1688.010 4700.550 ;
        RECT 1701.035 4710.720 1701.315 4711.000 ;
        RECT 1702.035 4710.720 1702.315 4711.000 ;
        RECT 1701.035 4709.220 1701.315 4709.500 ;
        RECT 1702.035 4709.220 1702.315 4709.500 ;
        RECT 1701.035 4707.720 1701.315 4708.000 ;
        RECT 1702.035 4707.720 1702.315 4708.000 ;
        RECT 1802.030 4710.485 1802.310 4710.765 ;
        RECT 1802.030 4708.985 1802.310 4709.265 ;
        RECT 1802.030 4707.485 1802.310 4707.765 ;
        RECT 1722.730 4703.270 1723.010 4703.550 ;
        RECT 1722.730 4701.770 1723.010 4702.050 ;
        RECT 1722.730 4700.270 1723.010 4700.550 ;
        RECT 1791.035 4703.720 1791.315 4704.000 ;
        RECT 1792.035 4703.720 1792.315 4704.000 ;
        RECT 1791.035 4702.220 1791.315 4702.500 ;
        RECT 1792.035 4702.220 1792.315 4702.500 ;
        RECT 1791.035 4700.720 1791.315 4701.000 ;
        RECT 1792.035 4700.720 1792.315 4701.000 ;
        RECT 1804.105 4703.300 1804.385 4703.580 ;
        RECT 1804.105 4701.800 1804.385 4702.080 ;
        RECT 1804.105 4700.300 1804.385 4700.580 ;
        RECT 1881.035 4710.720 1881.315 4711.000 ;
        RECT 1882.035 4710.720 1882.315 4711.000 ;
        RECT 1881.035 4709.220 1881.315 4709.500 ;
        RECT 1882.035 4709.220 1882.315 4709.500 ;
        RECT 1881.035 4707.720 1881.315 4708.000 ;
        RECT 1882.035 4707.720 1882.315 4708.000 ;
        RECT 1906.740 4703.680 1907.020 4703.960 ;
        RECT 1907.360 4703.680 1907.640 4703.960 ;
        RECT 1907.980 4703.680 1908.260 4703.960 ;
        RECT 1908.600 4703.680 1908.880 4703.960 ;
        RECT 1909.220 4703.680 1909.500 4703.960 ;
        RECT 1909.840 4703.680 1910.120 4703.960 ;
        RECT 1910.460 4703.680 1910.740 4703.960 ;
        RECT 1911.080 4703.680 1911.360 4703.960 ;
        RECT 1911.700 4703.680 1911.980 4703.960 ;
        RECT 1912.320 4703.680 1912.600 4703.960 ;
        RECT 1912.940 4703.680 1913.220 4703.960 ;
        RECT 1913.560 4703.680 1913.840 4703.960 ;
        RECT 1914.180 4703.680 1914.460 4703.960 ;
        RECT 1914.800 4703.680 1915.080 4703.960 ;
        RECT 1915.420 4703.680 1915.700 4703.960 ;
        RECT 1906.740 4703.060 1907.020 4703.340 ;
        RECT 1907.360 4703.060 1907.640 4703.340 ;
        RECT 1907.980 4703.060 1908.260 4703.340 ;
        RECT 1908.600 4703.060 1908.880 4703.340 ;
        RECT 1909.220 4703.060 1909.500 4703.340 ;
        RECT 1909.840 4703.060 1910.120 4703.340 ;
        RECT 1910.460 4703.060 1910.740 4703.340 ;
        RECT 1911.080 4703.060 1911.360 4703.340 ;
        RECT 1911.700 4703.060 1911.980 4703.340 ;
        RECT 1912.320 4703.060 1912.600 4703.340 ;
        RECT 1912.940 4703.060 1913.220 4703.340 ;
        RECT 1913.560 4703.060 1913.840 4703.340 ;
        RECT 1914.180 4703.060 1914.460 4703.340 ;
        RECT 1914.800 4703.060 1915.080 4703.340 ;
        RECT 1915.420 4703.060 1915.700 4703.340 ;
        RECT 1906.740 4702.440 1907.020 4702.720 ;
        RECT 1907.360 4702.440 1907.640 4702.720 ;
        RECT 1907.980 4702.440 1908.260 4702.720 ;
        RECT 1908.600 4702.440 1908.880 4702.720 ;
        RECT 1909.220 4702.440 1909.500 4702.720 ;
        RECT 1909.840 4702.440 1910.120 4702.720 ;
        RECT 1910.460 4702.440 1910.740 4702.720 ;
        RECT 1911.080 4702.440 1911.360 4702.720 ;
        RECT 1911.700 4702.440 1911.980 4702.720 ;
        RECT 1912.320 4702.440 1912.600 4702.720 ;
        RECT 1912.940 4702.440 1913.220 4702.720 ;
        RECT 1913.560 4702.440 1913.840 4702.720 ;
        RECT 1914.180 4702.440 1914.460 4702.720 ;
        RECT 1914.800 4702.440 1915.080 4702.720 ;
        RECT 1915.420 4702.440 1915.700 4702.720 ;
        RECT 1906.740 4701.820 1907.020 4702.100 ;
        RECT 1907.360 4701.820 1907.640 4702.100 ;
        RECT 1907.980 4701.820 1908.260 4702.100 ;
        RECT 1908.600 4701.820 1908.880 4702.100 ;
        RECT 1909.220 4701.820 1909.500 4702.100 ;
        RECT 1909.840 4701.820 1910.120 4702.100 ;
        RECT 1910.460 4701.820 1910.740 4702.100 ;
        RECT 1911.080 4701.820 1911.360 4702.100 ;
        RECT 1911.700 4701.820 1911.980 4702.100 ;
        RECT 1912.320 4701.820 1912.600 4702.100 ;
        RECT 1912.940 4701.820 1913.220 4702.100 ;
        RECT 1913.560 4701.820 1913.840 4702.100 ;
        RECT 1914.180 4701.820 1914.460 4702.100 ;
        RECT 1914.800 4701.820 1915.080 4702.100 ;
        RECT 1915.420 4701.820 1915.700 4702.100 ;
        RECT 1906.740 4701.200 1907.020 4701.480 ;
        RECT 1907.360 4701.200 1907.640 4701.480 ;
        RECT 1907.980 4701.200 1908.260 4701.480 ;
        RECT 1908.600 4701.200 1908.880 4701.480 ;
        RECT 1909.220 4701.200 1909.500 4701.480 ;
        RECT 1909.840 4701.200 1910.120 4701.480 ;
        RECT 1910.460 4701.200 1910.740 4701.480 ;
        RECT 1911.080 4701.200 1911.360 4701.480 ;
        RECT 1911.700 4701.200 1911.980 4701.480 ;
        RECT 1912.320 4701.200 1912.600 4701.480 ;
        RECT 1912.940 4701.200 1913.220 4701.480 ;
        RECT 1913.560 4701.200 1913.840 4701.480 ;
        RECT 1914.180 4701.200 1914.460 4701.480 ;
        RECT 1914.800 4701.200 1915.080 4701.480 ;
        RECT 1915.420 4701.200 1915.700 4701.480 ;
        RECT 1906.740 4700.580 1907.020 4700.860 ;
        RECT 1907.360 4700.580 1907.640 4700.860 ;
        RECT 1907.980 4700.580 1908.260 4700.860 ;
        RECT 1908.600 4700.580 1908.880 4700.860 ;
        RECT 1909.220 4700.580 1909.500 4700.860 ;
        RECT 1909.840 4700.580 1910.120 4700.860 ;
        RECT 1910.460 4700.580 1910.740 4700.860 ;
        RECT 1911.080 4700.580 1911.360 4700.860 ;
        RECT 1911.700 4700.580 1911.980 4700.860 ;
        RECT 1912.320 4700.580 1912.600 4700.860 ;
        RECT 1912.940 4700.580 1913.220 4700.860 ;
        RECT 1913.560 4700.580 1913.840 4700.860 ;
        RECT 1914.180 4700.580 1914.460 4700.860 ;
        RECT 1914.800 4700.580 1915.080 4700.860 ;
        RECT 1915.420 4700.580 1915.700 4700.860 ;
        RECT 1906.740 4699.960 1907.020 4700.240 ;
        RECT 1907.360 4699.960 1907.640 4700.240 ;
        RECT 1907.980 4699.960 1908.260 4700.240 ;
        RECT 1908.600 4699.960 1908.880 4700.240 ;
        RECT 1909.220 4699.960 1909.500 4700.240 ;
        RECT 1909.840 4699.960 1910.120 4700.240 ;
        RECT 1910.460 4699.960 1910.740 4700.240 ;
        RECT 1911.080 4699.960 1911.360 4700.240 ;
        RECT 1911.700 4699.960 1911.980 4700.240 ;
        RECT 1912.320 4699.960 1912.600 4700.240 ;
        RECT 1912.940 4699.960 1913.220 4700.240 ;
        RECT 1913.560 4699.960 1913.840 4700.240 ;
        RECT 1914.180 4699.960 1914.460 4700.240 ;
        RECT 1914.800 4699.960 1915.080 4700.240 ;
        RECT 1915.420 4699.960 1915.700 4700.240 ;
        RECT 1919.140 4703.680 1919.420 4703.960 ;
        RECT 1919.760 4703.680 1920.040 4703.960 ;
        RECT 1920.380 4703.680 1920.660 4703.960 ;
        RECT 1921.000 4703.680 1921.280 4703.960 ;
        RECT 1921.620 4703.680 1921.900 4703.960 ;
        RECT 1922.240 4703.680 1922.520 4703.960 ;
        RECT 1922.860 4703.680 1923.140 4703.960 ;
        RECT 1923.480 4703.680 1923.760 4703.960 ;
        RECT 1924.100 4703.680 1924.380 4703.960 ;
        RECT 1924.720 4703.680 1925.000 4703.960 ;
        RECT 1925.340 4703.680 1925.620 4703.960 ;
        RECT 1925.960 4703.680 1926.240 4703.960 ;
        RECT 1926.580 4703.680 1926.860 4703.960 ;
        RECT 1927.200 4703.680 1927.480 4703.960 ;
        RECT 1927.820 4703.680 1928.100 4703.960 ;
        RECT 1928.440 4703.680 1928.720 4703.960 ;
        RECT 1919.140 4703.060 1919.420 4703.340 ;
        RECT 1919.760 4703.060 1920.040 4703.340 ;
        RECT 1920.380 4703.060 1920.660 4703.340 ;
        RECT 1921.000 4703.060 1921.280 4703.340 ;
        RECT 1921.620 4703.060 1921.900 4703.340 ;
        RECT 1922.240 4703.060 1922.520 4703.340 ;
        RECT 1922.860 4703.060 1923.140 4703.340 ;
        RECT 1923.480 4703.060 1923.760 4703.340 ;
        RECT 1924.100 4703.060 1924.380 4703.340 ;
        RECT 1924.720 4703.060 1925.000 4703.340 ;
        RECT 1925.340 4703.060 1925.620 4703.340 ;
        RECT 1925.960 4703.060 1926.240 4703.340 ;
        RECT 1926.580 4703.060 1926.860 4703.340 ;
        RECT 1927.200 4703.060 1927.480 4703.340 ;
        RECT 1927.820 4703.060 1928.100 4703.340 ;
        RECT 1928.440 4703.060 1928.720 4703.340 ;
        RECT 1919.140 4702.440 1919.420 4702.720 ;
        RECT 1919.760 4702.440 1920.040 4702.720 ;
        RECT 1920.380 4702.440 1920.660 4702.720 ;
        RECT 1921.000 4702.440 1921.280 4702.720 ;
        RECT 1921.620 4702.440 1921.900 4702.720 ;
        RECT 1922.240 4702.440 1922.520 4702.720 ;
        RECT 1922.860 4702.440 1923.140 4702.720 ;
        RECT 1923.480 4702.440 1923.760 4702.720 ;
        RECT 1924.100 4702.440 1924.380 4702.720 ;
        RECT 1924.720 4702.440 1925.000 4702.720 ;
        RECT 1925.340 4702.440 1925.620 4702.720 ;
        RECT 1925.960 4702.440 1926.240 4702.720 ;
        RECT 1926.580 4702.440 1926.860 4702.720 ;
        RECT 1927.200 4702.440 1927.480 4702.720 ;
        RECT 1927.820 4702.440 1928.100 4702.720 ;
        RECT 1928.440 4702.440 1928.720 4702.720 ;
        RECT 1919.140 4701.820 1919.420 4702.100 ;
        RECT 1919.760 4701.820 1920.040 4702.100 ;
        RECT 1920.380 4701.820 1920.660 4702.100 ;
        RECT 1921.000 4701.820 1921.280 4702.100 ;
        RECT 1921.620 4701.820 1921.900 4702.100 ;
        RECT 1922.240 4701.820 1922.520 4702.100 ;
        RECT 1922.860 4701.820 1923.140 4702.100 ;
        RECT 1923.480 4701.820 1923.760 4702.100 ;
        RECT 1924.100 4701.820 1924.380 4702.100 ;
        RECT 1924.720 4701.820 1925.000 4702.100 ;
        RECT 1925.340 4701.820 1925.620 4702.100 ;
        RECT 1925.960 4701.820 1926.240 4702.100 ;
        RECT 1926.580 4701.820 1926.860 4702.100 ;
        RECT 1927.200 4701.820 1927.480 4702.100 ;
        RECT 1927.820 4701.820 1928.100 4702.100 ;
        RECT 1928.440 4701.820 1928.720 4702.100 ;
        RECT 1919.140 4701.200 1919.420 4701.480 ;
        RECT 1919.760 4701.200 1920.040 4701.480 ;
        RECT 1920.380 4701.200 1920.660 4701.480 ;
        RECT 1921.000 4701.200 1921.280 4701.480 ;
        RECT 1921.620 4701.200 1921.900 4701.480 ;
        RECT 1922.240 4701.200 1922.520 4701.480 ;
        RECT 1922.860 4701.200 1923.140 4701.480 ;
        RECT 1923.480 4701.200 1923.760 4701.480 ;
        RECT 1924.100 4701.200 1924.380 4701.480 ;
        RECT 1924.720 4701.200 1925.000 4701.480 ;
        RECT 1925.340 4701.200 1925.620 4701.480 ;
        RECT 1925.960 4701.200 1926.240 4701.480 ;
        RECT 1926.580 4701.200 1926.860 4701.480 ;
        RECT 1927.200 4701.200 1927.480 4701.480 ;
        RECT 1927.820 4701.200 1928.100 4701.480 ;
        RECT 1928.440 4701.200 1928.720 4701.480 ;
        RECT 1919.140 4700.580 1919.420 4700.860 ;
        RECT 1919.760 4700.580 1920.040 4700.860 ;
        RECT 1920.380 4700.580 1920.660 4700.860 ;
        RECT 1921.000 4700.580 1921.280 4700.860 ;
        RECT 1921.620 4700.580 1921.900 4700.860 ;
        RECT 1922.240 4700.580 1922.520 4700.860 ;
        RECT 1922.860 4700.580 1923.140 4700.860 ;
        RECT 1923.480 4700.580 1923.760 4700.860 ;
        RECT 1924.100 4700.580 1924.380 4700.860 ;
        RECT 1924.720 4700.580 1925.000 4700.860 ;
        RECT 1925.340 4700.580 1925.620 4700.860 ;
        RECT 1925.960 4700.580 1926.240 4700.860 ;
        RECT 1926.580 4700.580 1926.860 4700.860 ;
        RECT 1927.200 4700.580 1927.480 4700.860 ;
        RECT 1927.820 4700.580 1928.100 4700.860 ;
        RECT 1928.440 4700.580 1928.720 4700.860 ;
        RECT 1919.140 4699.960 1919.420 4700.240 ;
        RECT 1919.760 4699.960 1920.040 4700.240 ;
        RECT 1920.380 4699.960 1920.660 4700.240 ;
        RECT 1921.000 4699.960 1921.280 4700.240 ;
        RECT 1921.620 4699.960 1921.900 4700.240 ;
        RECT 1922.240 4699.960 1922.520 4700.240 ;
        RECT 1922.860 4699.960 1923.140 4700.240 ;
        RECT 1923.480 4699.960 1923.760 4700.240 ;
        RECT 1924.100 4699.960 1924.380 4700.240 ;
        RECT 1924.720 4699.960 1925.000 4700.240 ;
        RECT 1925.340 4699.960 1925.620 4700.240 ;
        RECT 1925.960 4699.960 1926.240 4700.240 ;
        RECT 1926.580 4699.960 1926.860 4700.240 ;
        RECT 1927.200 4699.960 1927.480 4700.240 ;
        RECT 1927.820 4699.960 1928.100 4700.240 ;
        RECT 1928.440 4699.960 1928.720 4700.240 ;
        RECT 1930.990 4703.680 1931.270 4703.960 ;
        RECT 1931.610 4703.680 1931.890 4703.960 ;
        RECT 1932.230 4703.680 1932.510 4703.960 ;
        RECT 1932.850 4703.680 1933.130 4703.960 ;
        RECT 1933.470 4703.680 1933.750 4703.960 ;
        RECT 1934.090 4703.680 1934.370 4703.960 ;
        RECT 1934.710 4703.680 1934.990 4703.960 ;
        RECT 1935.330 4703.680 1935.610 4703.960 ;
        RECT 1935.950 4703.680 1936.230 4703.960 ;
        RECT 1936.570 4703.680 1936.850 4703.960 ;
        RECT 1937.190 4703.680 1937.470 4703.960 ;
        RECT 1937.810 4703.680 1938.090 4703.960 ;
        RECT 1938.430 4703.680 1938.710 4703.960 ;
        RECT 1939.050 4703.680 1939.330 4703.960 ;
        RECT 1939.670 4703.680 1939.950 4703.960 ;
        RECT 1940.290 4703.680 1940.570 4703.960 ;
        RECT 1930.990 4703.060 1931.270 4703.340 ;
        RECT 1931.610 4703.060 1931.890 4703.340 ;
        RECT 1932.230 4703.060 1932.510 4703.340 ;
        RECT 1932.850 4703.060 1933.130 4703.340 ;
        RECT 1933.470 4703.060 1933.750 4703.340 ;
        RECT 1934.090 4703.060 1934.370 4703.340 ;
        RECT 1934.710 4703.060 1934.990 4703.340 ;
        RECT 1935.330 4703.060 1935.610 4703.340 ;
        RECT 1935.950 4703.060 1936.230 4703.340 ;
        RECT 1936.570 4703.060 1936.850 4703.340 ;
        RECT 1937.190 4703.060 1937.470 4703.340 ;
        RECT 1937.810 4703.060 1938.090 4703.340 ;
        RECT 1938.430 4703.060 1938.710 4703.340 ;
        RECT 1939.050 4703.060 1939.330 4703.340 ;
        RECT 1939.670 4703.060 1939.950 4703.340 ;
        RECT 1940.290 4703.060 1940.570 4703.340 ;
        RECT 1930.990 4702.440 1931.270 4702.720 ;
        RECT 1931.610 4702.440 1931.890 4702.720 ;
        RECT 1932.230 4702.440 1932.510 4702.720 ;
        RECT 1932.850 4702.440 1933.130 4702.720 ;
        RECT 1933.470 4702.440 1933.750 4702.720 ;
        RECT 1934.090 4702.440 1934.370 4702.720 ;
        RECT 1934.710 4702.440 1934.990 4702.720 ;
        RECT 1935.330 4702.440 1935.610 4702.720 ;
        RECT 1935.950 4702.440 1936.230 4702.720 ;
        RECT 1936.570 4702.440 1936.850 4702.720 ;
        RECT 1937.190 4702.440 1937.470 4702.720 ;
        RECT 1937.810 4702.440 1938.090 4702.720 ;
        RECT 1938.430 4702.440 1938.710 4702.720 ;
        RECT 1939.050 4702.440 1939.330 4702.720 ;
        RECT 1939.670 4702.440 1939.950 4702.720 ;
        RECT 1940.290 4702.440 1940.570 4702.720 ;
        RECT 1930.990 4701.820 1931.270 4702.100 ;
        RECT 1931.610 4701.820 1931.890 4702.100 ;
        RECT 1932.230 4701.820 1932.510 4702.100 ;
        RECT 1932.850 4701.820 1933.130 4702.100 ;
        RECT 1933.470 4701.820 1933.750 4702.100 ;
        RECT 1934.090 4701.820 1934.370 4702.100 ;
        RECT 1934.710 4701.820 1934.990 4702.100 ;
        RECT 1935.330 4701.820 1935.610 4702.100 ;
        RECT 1935.950 4701.820 1936.230 4702.100 ;
        RECT 1936.570 4701.820 1936.850 4702.100 ;
        RECT 1937.190 4701.820 1937.470 4702.100 ;
        RECT 1937.810 4701.820 1938.090 4702.100 ;
        RECT 1938.430 4701.820 1938.710 4702.100 ;
        RECT 1939.050 4701.820 1939.330 4702.100 ;
        RECT 1939.670 4701.820 1939.950 4702.100 ;
        RECT 1940.290 4701.820 1940.570 4702.100 ;
        RECT 1930.990 4701.200 1931.270 4701.480 ;
        RECT 1931.610 4701.200 1931.890 4701.480 ;
        RECT 1932.230 4701.200 1932.510 4701.480 ;
        RECT 1932.850 4701.200 1933.130 4701.480 ;
        RECT 1933.470 4701.200 1933.750 4701.480 ;
        RECT 1934.090 4701.200 1934.370 4701.480 ;
        RECT 1934.710 4701.200 1934.990 4701.480 ;
        RECT 1935.330 4701.200 1935.610 4701.480 ;
        RECT 1935.950 4701.200 1936.230 4701.480 ;
        RECT 1936.570 4701.200 1936.850 4701.480 ;
        RECT 1937.190 4701.200 1937.470 4701.480 ;
        RECT 1937.810 4701.200 1938.090 4701.480 ;
        RECT 1938.430 4701.200 1938.710 4701.480 ;
        RECT 1939.050 4701.200 1939.330 4701.480 ;
        RECT 1939.670 4701.200 1939.950 4701.480 ;
        RECT 1940.290 4701.200 1940.570 4701.480 ;
        RECT 1930.990 4700.580 1931.270 4700.860 ;
        RECT 1931.610 4700.580 1931.890 4700.860 ;
        RECT 1932.230 4700.580 1932.510 4700.860 ;
        RECT 1932.850 4700.580 1933.130 4700.860 ;
        RECT 1933.470 4700.580 1933.750 4700.860 ;
        RECT 1934.090 4700.580 1934.370 4700.860 ;
        RECT 1934.710 4700.580 1934.990 4700.860 ;
        RECT 1935.330 4700.580 1935.610 4700.860 ;
        RECT 1935.950 4700.580 1936.230 4700.860 ;
        RECT 1936.570 4700.580 1936.850 4700.860 ;
        RECT 1937.190 4700.580 1937.470 4700.860 ;
        RECT 1937.810 4700.580 1938.090 4700.860 ;
        RECT 1938.430 4700.580 1938.710 4700.860 ;
        RECT 1939.050 4700.580 1939.330 4700.860 ;
        RECT 1939.670 4700.580 1939.950 4700.860 ;
        RECT 1940.290 4700.580 1940.570 4700.860 ;
        RECT 1930.990 4699.960 1931.270 4700.240 ;
        RECT 1931.610 4699.960 1931.890 4700.240 ;
        RECT 1932.230 4699.960 1932.510 4700.240 ;
        RECT 1932.850 4699.960 1933.130 4700.240 ;
        RECT 1933.470 4699.960 1933.750 4700.240 ;
        RECT 1934.090 4699.960 1934.370 4700.240 ;
        RECT 1934.710 4699.960 1934.990 4700.240 ;
        RECT 1935.330 4699.960 1935.610 4700.240 ;
        RECT 1935.950 4699.960 1936.230 4700.240 ;
        RECT 1936.570 4699.960 1936.850 4700.240 ;
        RECT 1937.190 4699.960 1937.470 4700.240 ;
        RECT 1937.810 4699.960 1938.090 4700.240 ;
        RECT 1938.430 4699.960 1938.710 4700.240 ;
        RECT 1939.050 4699.960 1939.330 4700.240 ;
        RECT 1939.670 4699.960 1939.950 4700.240 ;
        RECT 1940.290 4699.960 1940.570 4700.240 ;
        RECT 1944.520 4703.680 1944.800 4703.960 ;
        RECT 1945.140 4703.680 1945.420 4703.960 ;
        RECT 1945.760 4703.680 1946.040 4703.960 ;
        RECT 1946.380 4703.680 1946.660 4703.960 ;
        RECT 1947.000 4703.680 1947.280 4703.960 ;
        RECT 1947.620 4703.680 1947.900 4703.960 ;
        RECT 1948.240 4703.680 1948.520 4703.960 ;
        RECT 1948.860 4703.680 1949.140 4703.960 ;
        RECT 1949.480 4703.680 1949.760 4703.960 ;
        RECT 1950.100 4703.680 1950.380 4703.960 ;
        RECT 1950.720 4703.680 1951.000 4703.960 ;
        RECT 1951.340 4703.680 1951.620 4703.960 ;
        RECT 1951.960 4703.680 1952.240 4703.960 ;
        RECT 1952.580 4703.680 1952.860 4703.960 ;
        RECT 1953.200 4703.680 1953.480 4703.960 ;
        RECT 1953.820 4703.680 1954.100 4703.960 ;
        RECT 1944.520 4703.060 1944.800 4703.340 ;
        RECT 1945.140 4703.060 1945.420 4703.340 ;
        RECT 1945.760 4703.060 1946.040 4703.340 ;
        RECT 1946.380 4703.060 1946.660 4703.340 ;
        RECT 1947.000 4703.060 1947.280 4703.340 ;
        RECT 1947.620 4703.060 1947.900 4703.340 ;
        RECT 1948.240 4703.060 1948.520 4703.340 ;
        RECT 1948.860 4703.060 1949.140 4703.340 ;
        RECT 1949.480 4703.060 1949.760 4703.340 ;
        RECT 1950.100 4703.060 1950.380 4703.340 ;
        RECT 1950.720 4703.060 1951.000 4703.340 ;
        RECT 1951.340 4703.060 1951.620 4703.340 ;
        RECT 1951.960 4703.060 1952.240 4703.340 ;
        RECT 1952.580 4703.060 1952.860 4703.340 ;
        RECT 1953.200 4703.060 1953.480 4703.340 ;
        RECT 1953.820 4703.060 1954.100 4703.340 ;
        RECT 1944.520 4702.440 1944.800 4702.720 ;
        RECT 1945.140 4702.440 1945.420 4702.720 ;
        RECT 1945.760 4702.440 1946.040 4702.720 ;
        RECT 1946.380 4702.440 1946.660 4702.720 ;
        RECT 1947.000 4702.440 1947.280 4702.720 ;
        RECT 1947.620 4702.440 1947.900 4702.720 ;
        RECT 1948.240 4702.440 1948.520 4702.720 ;
        RECT 1948.860 4702.440 1949.140 4702.720 ;
        RECT 1949.480 4702.440 1949.760 4702.720 ;
        RECT 1950.100 4702.440 1950.380 4702.720 ;
        RECT 1950.720 4702.440 1951.000 4702.720 ;
        RECT 1951.340 4702.440 1951.620 4702.720 ;
        RECT 1951.960 4702.440 1952.240 4702.720 ;
        RECT 1952.580 4702.440 1952.860 4702.720 ;
        RECT 1953.200 4702.440 1953.480 4702.720 ;
        RECT 1953.820 4702.440 1954.100 4702.720 ;
        RECT 1944.520 4701.820 1944.800 4702.100 ;
        RECT 1945.140 4701.820 1945.420 4702.100 ;
        RECT 1945.760 4701.820 1946.040 4702.100 ;
        RECT 1946.380 4701.820 1946.660 4702.100 ;
        RECT 1947.000 4701.820 1947.280 4702.100 ;
        RECT 1947.620 4701.820 1947.900 4702.100 ;
        RECT 1948.240 4701.820 1948.520 4702.100 ;
        RECT 1948.860 4701.820 1949.140 4702.100 ;
        RECT 1949.480 4701.820 1949.760 4702.100 ;
        RECT 1950.100 4701.820 1950.380 4702.100 ;
        RECT 1950.720 4701.820 1951.000 4702.100 ;
        RECT 1951.340 4701.820 1951.620 4702.100 ;
        RECT 1951.960 4701.820 1952.240 4702.100 ;
        RECT 1952.580 4701.820 1952.860 4702.100 ;
        RECT 1953.200 4701.820 1953.480 4702.100 ;
        RECT 1953.820 4701.820 1954.100 4702.100 ;
        RECT 1944.520 4701.200 1944.800 4701.480 ;
        RECT 1945.140 4701.200 1945.420 4701.480 ;
        RECT 1945.760 4701.200 1946.040 4701.480 ;
        RECT 1946.380 4701.200 1946.660 4701.480 ;
        RECT 1947.000 4701.200 1947.280 4701.480 ;
        RECT 1947.620 4701.200 1947.900 4701.480 ;
        RECT 1948.240 4701.200 1948.520 4701.480 ;
        RECT 1948.860 4701.200 1949.140 4701.480 ;
        RECT 1949.480 4701.200 1949.760 4701.480 ;
        RECT 1950.100 4701.200 1950.380 4701.480 ;
        RECT 1950.720 4701.200 1951.000 4701.480 ;
        RECT 1951.340 4701.200 1951.620 4701.480 ;
        RECT 1951.960 4701.200 1952.240 4701.480 ;
        RECT 1952.580 4701.200 1952.860 4701.480 ;
        RECT 1953.200 4701.200 1953.480 4701.480 ;
        RECT 1953.820 4701.200 1954.100 4701.480 ;
        RECT 1944.520 4700.580 1944.800 4700.860 ;
        RECT 1945.140 4700.580 1945.420 4700.860 ;
        RECT 1945.760 4700.580 1946.040 4700.860 ;
        RECT 1946.380 4700.580 1946.660 4700.860 ;
        RECT 1947.000 4700.580 1947.280 4700.860 ;
        RECT 1947.620 4700.580 1947.900 4700.860 ;
        RECT 1948.240 4700.580 1948.520 4700.860 ;
        RECT 1948.860 4700.580 1949.140 4700.860 ;
        RECT 1949.480 4700.580 1949.760 4700.860 ;
        RECT 1950.100 4700.580 1950.380 4700.860 ;
        RECT 1950.720 4700.580 1951.000 4700.860 ;
        RECT 1951.340 4700.580 1951.620 4700.860 ;
        RECT 1951.960 4700.580 1952.240 4700.860 ;
        RECT 1952.580 4700.580 1952.860 4700.860 ;
        RECT 1953.200 4700.580 1953.480 4700.860 ;
        RECT 1953.820 4700.580 1954.100 4700.860 ;
        RECT 1944.520 4699.960 1944.800 4700.240 ;
        RECT 1945.140 4699.960 1945.420 4700.240 ;
        RECT 1945.760 4699.960 1946.040 4700.240 ;
        RECT 1946.380 4699.960 1946.660 4700.240 ;
        RECT 1947.000 4699.960 1947.280 4700.240 ;
        RECT 1947.620 4699.960 1947.900 4700.240 ;
        RECT 1948.240 4699.960 1948.520 4700.240 ;
        RECT 1948.860 4699.960 1949.140 4700.240 ;
        RECT 1949.480 4699.960 1949.760 4700.240 ;
        RECT 1950.100 4699.960 1950.380 4700.240 ;
        RECT 1950.720 4699.960 1951.000 4700.240 ;
        RECT 1951.340 4699.960 1951.620 4700.240 ;
        RECT 1951.960 4699.960 1952.240 4700.240 ;
        RECT 1952.580 4699.960 1952.860 4700.240 ;
        RECT 1953.200 4699.960 1953.480 4700.240 ;
        RECT 1953.820 4699.960 1954.100 4700.240 ;
        RECT 1956.370 4703.680 1956.650 4703.960 ;
        RECT 1956.990 4703.680 1957.270 4703.960 ;
        RECT 1957.610 4703.680 1957.890 4703.960 ;
        RECT 1958.230 4703.680 1958.510 4703.960 ;
        RECT 1958.850 4703.680 1959.130 4703.960 ;
        RECT 1959.470 4703.680 1959.750 4703.960 ;
        RECT 1960.090 4703.680 1960.370 4703.960 ;
        RECT 1960.710 4703.680 1960.990 4703.960 ;
        RECT 1961.330 4703.680 1961.610 4703.960 ;
        RECT 1961.950 4703.680 1962.230 4703.960 ;
        RECT 1962.570 4703.680 1962.850 4703.960 ;
        RECT 1963.190 4703.680 1963.470 4703.960 ;
        RECT 1963.810 4703.680 1964.090 4703.960 ;
        RECT 1964.430 4703.680 1964.710 4703.960 ;
        RECT 1965.050 4703.680 1965.330 4703.960 ;
        RECT 1965.670 4703.680 1965.950 4703.960 ;
        RECT 1956.370 4703.060 1956.650 4703.340 ;
        RECT 1956.990 4703.060 1957.270 4703.340 ;
        RECT 1957.610 4703.060 1957.890 4703.340 ;
        RECT 1958.230 4703.060 1958.510 4703.340 ;
        RECT 1958.850 4703.060 1959.130 4703.340 ;
        RECT 1959.470 4703.060 1959.750 4703.340 ;
        RECT 1960.090 4703.060 1960.370 4703.340 ;
        RECT 1960.710 4703.060 1960.990 4703.340 ;
        RECT 1961.330 4703.060 1961.610 4703.340 ;
        RECT 1961.950 4703.060 1962.230 4703.340 ;
        RECT 1962.570 4703.060 1962.850 4703.340 ;
        RECT 1963.190 4703.060 1963.470 4703.340 ;
        RECT 1963.810 4703.060 1964.090 4703.340 ;
        RECT 1964.430 4703.060 1964.710 4703.340 ;
        RECT 1965.050 4703.060 1965.330 4703.340 ;
        RECT 1965.670 4703.060 1965.950 4703.340 ;
        RECT 1956.370 4702.440 1956.650 4702.720 ;
        RECT 1956.990 4702.440 1957.270 4702.720 ;
        RECT 1957.610 4702.440 1957.890 4702.720 ;
        RECT 1958.230 4702.440 1958.510 4702.720 ;
        RECT 1958.850 4702.440 1959.130 4702.720 ;
        RECT 1959.470 4702.440 1959.750 4702.720 ;
        RECT 1960.090 4702.440 1960.370 4702.720 ;
        RECT 1960.710 4702.440 1960.990 4702.720 ;
        RECT 1961.330 4702.440 1961.610 4702.720 ;
        RECT 1961.950 4702.440 1962.230 4702.720 ;
        RECT 1962.570 4702.440 1962.850 4702.720 ;
        RECT 1963.190 4702.440 1963.470 4702.720 ;
        RECT 1963.810 4702.440 1964.090 4702.720 ;
        RECT 1964.430 4702.440 1964.710 4702.720 ;
        RECT 1965.050 4702.440 1965.330 4702.720 ;
        RECT 1965.670 4702.440 1965.950 4702.720 ;
        RECT 1956.370 4701.820 1956.650 4702.100 ;
        RECT 1956.990 4701.820 1957.270 4702.100 ;
        RECT 1957.610 4701.820 1957.890 4702.100 ;
        RECT 1958.230 4701.820 1958.510 4702.100 ;
        RECT 1958.850 4701.820 1959.130 4702.100 ;
        RECT 1959.470 4701.820 1959.750 4702.100 ;
        RECT 1960.090 4701.820 1960.370 4702.100 ;
        RECT 1960.710 4701.820 1960.990 4702.100 ;
        RECT 1961.330 4701.820 1961.610 4702.100 ;
        RECT 1961.950 4701.820 1962.230 4702.100 ;
        RECT 1962.570 4701.820 1962.850 4702.100 ;
        RECT 1963.190 4701.820 1963.470 4702.100 ;
        RECT 1963.810 4701.820 1964.090 4702.100 ;
        RECT 1964.430 4701.820 1964.710 4702.100 ;
        RECT 1965.050 4701.820 1965.330 4702.100 ;
        RECT 1965.670 4701.820 1965.950 4702.100 ;
        RECT 1956.370 4701.200 1956.650 4701.480 ;
        RECT 1956.990 4701.200 1957.270 4701.480 ;
        RECT 1957.610 4701.200 1957.890 4701.480 ;
        RECT 1958.230 4701.200 1958.510 4701.480 ;
        RECT 1958.850 4701.200 1959.130 4701.480 ;
        RECT 1959.470 4701.200 1959.750 4701.480 ;
        RECT 1960.090 4701.200 1960.370 4701.480 ;
        RECT 1960.710 4701.200 1960.990 4701.480 ;
        RECT 1961.330 4701.200 1961.610 4701.480 ;
        RECT 1961.950 4701.200 1962.230 4701.480 ;
        RECT 1962.570 4701.200 1962.850 4701.480 ;
        RECT 1963.190 4701.200 1963.470 4701.480 ;
        RECT 1963.810 4701.200 1964.090 4701.480 ;
        RECT 1964.430 4701.200 1964.710 4701.480 ;
        RECT 1965.050 4701.200 1965.330 4701.480 ;
        RECT 1965.670 4701.200 1965.950 4701.480 ;
        RECT 1956.370 4700.580 1956.650 4700.860 ;
        RECT 1956.990 4700.580 1957.270 4700.860 ;
        RECT 1957.610 4700.580 1957.890 4700.860 ;
        RECT 1958.230 4700.580 1958.510 4700.860 ;
        RECT 1958.850 4700.580 1959.130 4700.860 ;
        RECT 1959.470 4700.580 1959.750 4700.860 ;
        RECT 1960.090 4700.580 1960.370 4700.860 ;
        RECT 1960.710 4700.580 1960.990 4700.860 ;
        RECT 1961.330 4700.580 1961.610 4700.860 ;
        RECT 1961.950 4700.580 1962.230 4700.860 ;
        RECT 1962.570 4700.580 1962.850 4700.860 ;
        RECT 1963.190 4700.580 1963.470 4700.860 ;
        RECT 1963.810 4700.580 1964.090 4700.860 ;
        RECT 1964.430 4700.580 1964.710 4700.860 ;
        RECT 1965.050 4700.580 1965.330 4700.860 ;
        RECT 1965.670 4700.580 1965.950 4700.860 ;
        RECT 1956.370 4699.960 1956.650 4700.240 ;
        RECT 1956.990 4699.960 1957.270 4700.240 ;
        RECT 1957.610 4699.960 1957.890 4700.240 ;
        RECT 1958.230 4699.960 1958.510 4700.240 ;
        RECT 1958.850 4699.960 1959.130 4700.240 ;
        RECT 1959.470 4699.960 1959.750 4700.240 ;
        RECT 1960.090 4699.960 1960.370 4700.240 ;
        RECT 1960.710 4699.960 1960.990 4700.240 ;
        RECT 1961.330 4699.960 1961.610 4700.240 ;
        RECT 1961.950 4699.960 1962.230 4700.240 ;
        RECT 1962.570 4699.960 1962.850 4700.240 ;
        RECT 1963.190 4699.960 1963.470 4700.240 ;
        RECT 1963.810 4699.960 1964.090 4700.240 ;
        RECT 1964.430 4699.960 1964.710 4700.240 ;
        RECT 1965.050 4699.960 1965.330 4700.240 ;
        RECT 1965.670 4699.960 1965.950 4700.240 ;
        RECT 2202.740 4716.895 2203.020 4717.175 ;
        RECT 1969.390 4703.680 1969.670 4703.960 ;
        RECT 1970.010 4703.680 1970.290 4703.960 ;
        RECT 1970.630 4703.680 1970.910 4703.960 ;
        RECT 1971.250 4703.680 1971.530 4703.960 ;
        RECT 1971.870 4703.680 1972.150 4703.960 ;
        RECT 1972.490 4703.680 1972.770 4703.960 ;
        RECT 1973.110 4703.680 1973.390 4703.960 ;
        RECT 1973.730 4703.680 1974.010 4703.960 ;
        RECT 1974.350 4703.680 1974.630 4703.960 ;
        RECT 1974.970 4703.680 1975.250 4703.960 ;
        RECT 1975.590 4703.680 1975.870 4703.960 ;
        RECT 1976.210 4703.680 1976.490 4703.960 ;
        RECT 1976.830 4703.680 1977.110 4703.960 ;
        RECT 1977.450 4703.680 1977.730 4703.960 ;
        RECT 1978.070 4703.680 1978.350 4703.960 ;
        RECT 1969.390 4703.060 1969.670 4703.340 ;
        RECT 1970.010 4703.060 1970.290 4703.340 ;
        RECT 1970.630 4703.060 1970.910 4703.340 ;
        RECT 1971.250 4703.060 1971.530 4703.340 ;
        RECT 1971.870 4703.060 1972.150 4703.340 ;
        RECT 1972.490 4703.060 1972.770 4703.340 ;
        RECT 1973.110 4703.060 1973.390 4703.340 ;
        RECT 1973.730 4703.060 1974.010 4703.340 ;
        RECT 1974.350 4703.060 1974.630 4703.340 ;
        RECT 1974.970 4703.060 1975.250 4703.340 ;
        RECT 1975.590 4703.060 1975.870 4703.340 ;
        RECT 1976.210 4703.060 1976.490 4703.340 ;
        RECT 1976.830 4703.060 1977.110 4703.340 ;
        RECT 1977.450 4703.060 1977.730 4703.340 ;
        RECT 1978.070 4703.060 1978.350 4703.340 ;
        RECT 1969.390 4702.440 1969.670 4702.720 ;
        RECT 1970.010 4702.440 1970.290 4702.720 ;
        RECT 1970.630 4702.440 1970.910 4702.720 ;
        RECT 1971.250 4702.440 1971.530 4702.720 ;
        RECT 1971.870 4702.440 1972.150 4702.720 ;
        RECT 1972.490 4702.440 1972.770 4702.720 ;
        RECT 1973.110 4702.440 1973.390 4702.720 ;
        RECT 1973.730 4702.440 1974.010 4702.720 ;
        RECT 1974.350 4702.440 1974.630 4702.720 ;
        RECT 1974.970 4702.440 1975.250 4702.720 ;
        RECT 1975.590 4702.440 1975.870 4702.720 ;
        RECT 1976.210 4702.440 1976.490 4702.720 ;
        RECT 1976.830 4702.440 1977.110 4702.720 ;
        RECT 1977.450 4702.440 1977.730 4702.720 ;
        RECT 1978.070 4702.440 1978.350 4702.720 ;
        RECT 1969.390 4701.820 1969.670 4702.100 ;
        RECT 1970.010 4701.820 1970.290 4702.100 ;
        RECT 1970.630 4701.820 1970.910 4702.100 ;
        RECT 1971.250 4701.820 1971.530 4702.100 ;
        RECT 1971.870 4701.820 1972.150 4702.100 ;
        RECT 1972.490 4701.820 1972.770 4702.100 ;
        RECT 1973.110 4701.820 1973.390 4702.100 ;
        RECT 1973.730 4701.820 1974.010 4702.100 ;
        RECT 1974.350 4701.820 1974.630 4702.100 ;
        RECT 1974.970 4701.820 1975.250 4702.100 ;
        RECT 1975.590 4701.820 1975.870 4702.100 ;
        RECT 1976.210 4701.820 1976.490 4702.100 ;
        RECT 1976.830 4701.820 1977.110 4702.100 ;
        RECT 1977.450 4701.820 1977.730 4702.100 ;
        RECT 1978.070 4701.820 1978.350 4702.100 ;
        RECT 1969.390 4701.200 1969.670 4701.480 ;
        RECT 1970.010 4701.200 1970.290 4701.480 ;
        RECT 1970.630 4701.200 1970.910 4701.480 ;
        RECT 1971.250 4701.200 1971.530 4701.480 ;
        RECT 1971.870 4701.200 1972.150 4701.480 ;
        RECT 1972.490 4701.200 1972.770 4701.480 ;
        RECT 1973.110 4701.200 1973.390 4701.480 ;
        RECT 1973.730 4701.200 1974.010 4701.480 ;
        RECT 1974.350 4701.200 1974.630 4701.480 ;
        RECT 1974.970 4701.200 1975.250 4701.480 ;
        RECT 1975.590 4701.200 1975.870 4701.480 ;
        RECT 1976.210 4701.200 1976.490 4701.480 ;
        RECT 1976.830 4701.200 1977.110 4701.480 ;
        RECT 1977.450 4701.200 1977.730 4701.480 ;
        RECT 1978.070 4701.200 1978.350 4701.480 ;
        RECT 1969.390 4700.580 1969.670 4700.860 ;
        RECT 1970.010 4700.580 1970.290 4700.860 ;
        RECT 1970.630 4700.580 1970.910 4700.860 ;
        RECT 1971.250 4700.580 1971.530 4700.860 ;
        RECT 1971.870 4700.580 1972.150 4700.860 ;
        RECT 1972.490 4700.580 1972.770 4700.860 ;
        RECT 1973.110 4700.580 1973.390 4700.860 ;
        RECT 1973.730 4700.580 1974.010 4700.860 ;
        RECT 1974.350 4700.580 1974.630 4700.860 ;
        RECT 1974.970 4700.580 1975.250 4700.860 ;
        RECT 1975.590 4700.580 1975.870 4700.860 ;
        RECT 1976.210 4700.580 1976.490 4700.860 ;
        RECT 1976.830 4700.580 1977.110 4700.860 ;
        RECT 1977.450 4700.580 1977.730 4700.860 ;
        RECT 1978.070 4700.580 1978.350 4700.860 ;
        RECT 1969.390 4699.960 1969.670 4700.240 ;
        RECT 1970.010 4699.960 1970.290 4700.240 ;
        RECT 1970.630 4699.960 1970.910 4700.240 ;
        RECT 1971.250 4699.960 1971.530 4700.240 ;
        RECT 1971.870 4699.960 1972.150 4700.240 ;
        RECT 1972.490 4699.960 1972.770 4700.240 ;
        RECT 1973.110 4699.960 1973.390 4700.240 ;
        RECT 1973.730 4699.960 1974.010 4700.240 ;
        RECT 1974.350 4699.960 1974.630 4700.240 ;
        RECT 1974.970 4699.960 1975.250 4700.240 ;
        RECT 1975.590 4699.960 1975.870 4700.240 ;
        RECT 1976.210 4699.960 1976.490 4700.240 ;
        RECT 1976.830 4699.960 1977.110 4700.240 ;
        RECT 1977.450 4699.960 1977.730 4700.240 ;
        RECT 1978.070 4699.960 1978.350 4700.240 ;
        RECT 2061.035 4710.720 2061.315 4711.000 ;
        RECT 2062.035 4710.720 2062.315 4711.000 ;
        RECT 2061.035 4709.220 2061.315 4709.500 ;
        RECT 2062.035 4709.220 2062.315 4709.500 ;
        RECT 2061.035 4707.720 2061.315 4708.000 ;
        RECT 2062.035 4707.720 2062.315 4708.000 ;
        RECT 2151.035 4703.720 2151.315 4704.000 ;
        RECT 2152.035 4703.720 2152.315 4704.000 ;
        RECT 2151.035 4702.220 2151.315 4702.500 ;
        RECT 2152.035 4702.220 2152.315 4702.500 ;
        RECT 2151.035 4700.720 2151.315 4701.000 ;
        RECT 2152.035 4700.720 2152.315 4701.000 ;
        RECT 2202.730 4703.270 2203.010 4703.550 ;
        RECT 2202.730 4701.770 2203.010 4702.050 ;
        RECT 2202.730 4700.270 2203.010 4700.550 ;
        RECT 2237.740 4716.895 2238.020 4717.175 ;
        RECT 2272.740 4716.895 2273.020 4717.175 ;
        RECT 2237.730 4703.270 2238.010 4703.550 ;
        RECT 2237.730 4701.770 2238.010 4702.050 ;
        RECT 2237.730 4700.270 2238.010 4700.550 ;
        RECT 2241.035 4710.720 2241.315 4711.000 ;
        RECT 2242.035 4710.720 2242.315 4711.000 ;
        RECT 2241.035 4709.220 2241.315 4709.500 ;
        RECT 2242.035 4709.220 2242.315 4709.500 ;
        RECT 2241.035 4707.720 2241.315 4708.000 ;
        RECT 2242.035 4707.720 2242.315 4708.000 ;
        RECT 2352.030 4710.485 2352.310 4710.765 ;
        RECT 2352.030 4708.985 2352.310 4709.265 ;
        RECT 2352.030 4707.485 2352.310 4707.765 ;
        RECT 2272.730 4703.270 2273.010 4703.550 ;
        RECT 2272.730 4701.770 2273.010 4702.050 ;
        RECT 2272.730 4700.270 2273.010 4700.550 ;
        RECT 2331.035 4703.720 2331.315 4704.000 ;
        RECT 2332.035 4703.720 2332.315 4704.000 ;
        RECT 2331.035 4702.220 2331.315 4702.500 ;
        RECT 2332.035 4702.220 2332.315 4702.500 ;
        RECT 2331.035 4700.720 2331.315 4701.000 ;
        RECT 2332.035 4700.720 2332.315 4701.000 ;
        RECT 2477.740 4716.895 2478.020 4717.175 ;
        RECT 2354.105 4703.300 2354.385 4703.580 ;
        RECT 2354.105 4701.800 2354.385 4702.080 ;
        RECT 2354.105 4700.300 2354.385 4700.580 ;
        RECT 2421.035 4710.720 2421.315 4711.000 ;
        RECT 2422.035 4710.720 2422.315 4711.000 ;
        RECT 2421.035 4709.220 2421.315 4709.500 ;
        RECT 2422.035 4709.220 2422.315 4709.500 ;
        RECT 2421.035 4707.720 2421.315 4708.000 ;
        RECT 2422.035 4707.720 2422.315 4708.000 ;
        RECT 2512.740 4716.895 2513.020 4717.175 ;
        RECT 2477.730 4703.270 2478.010 4703.550 ;
        RECT 2477.730 4701.770 2478.010 4702.050 ;
        RECT 2477.730 4700.270 2478.010 4700.550 ;
        RECT 2511.035 4703.720 2511.315 4704.000 ;
        RECT 2512.035 4703.720 2512.315 4704.000 ;
        RECT 2512.730 4703.270 2513.010 4703.550 ;
        RECT 2511.035 4702.220 2511.315 4702.500 ;
        RECT 2512.035 4702.220 2512.315 4702.500 ;
        RECT 2512.730 4701.770 2513.010 4702.050 ;
        RECT 2511.035 4700.720 2511.315 4701.000 ;
        RECT 2512.035 4700.720 2512.315 4701.000 ;
        RECT 2512.730 4700.270 2513.010 4700.550 ;
        RECT 2547.740 4716.895 2548.020 4717.175 ;
        RECT 2547.730 4703.270 2548.010 4703.550 ;
        RECT 2547.730 4701.770 2548.010 4702.050 ;
        RECT 2547.730 4700.270 2548.010 4700.550 ;
        RECT 2601.035 4710.720 2601.315 4711.000 ;
        RECT 2602.035 4710.720 2602.315 4711.000 ;
        RECT 2601.035 4709.220 2601.315 4709.500 ;
        RECT 2602.035 4709.220 2602.315 4709.500 ;
        RECT 2601.035 4707.720 2601.315 4708.000 ;
        RECT 2602.035 4707.720 2602.315 4708.000 ;
        RECT 2627.030 4710.485 2627.310 4710.765 ;
        RECT 2627.030 4708.985 2627.310 4709.265 ;
        RECT 2627.030 4707.485 2627.310 4707.765 ;
        RECT 2752.740 4716.895 2753.020 4717.175 ;
        RECT 2629.105 4703.300 2629.385 4703.580 ;
        RECT 2629.105 4701.800 2629.385 4702.080 ;
        RECT 2629.105 4700.300 2629.385 4700.580 ;
        RECT 2691.035 4703.720 2691.315 4704.000 ;
        RECT 2692.035 4703.720 2692.315 4704.000 ;
        RECT 2691.035 4702.220 2691.315 4702.500 ;
        RECT 2692.035 4702.220 2692.315 4702.500 ;
        RECT 2691.035 4700.720 2691.315 4701.000 ;
        RECT 2692.035 4700.720 2692.315 4701.000 ;
        RECT 2787.740 4716.895 2788.020 4717.175 ;
        RECT 2752.730 4703.270 2753.010 4703.550 ;
        RECT 2752.730 4701.770 2753.010 4702.050 ;
        RECT 2752.730 4700.270 2753.010 4700.550 ;
        RECT 2781.035 4710.720 2781.315 4711.000 ;
        RECT 2782.035 4710.720 2782.315 4711.000 ;
        RECT 2781.035 4709.220 2781.315 4709.500 ;
        RECT 2782.035 4709.220 2782.315 4709.500 ;
        RECT 2781.035 4707.720 2781.315 4708.000 ;
        RECT 2782.035 4707.720 2782.315 4708.000 ;
        RECT 2787.730 4703.270 2788.010 4703.550 ;
        RECT 2787.730 4701.770 2788.010 4702.050 ;
        RECT 2787.730 4700.270 2788.010 4700.550 ;
        RECT 2822.740 4716.895 2823.020 4717.175 ;
        RECT 2902.030 4710.485 2902.310 4710.765 ;
        RECT 2902.030 4708.985 2902.310 4709.265 ;
        RECT 2902.030 4707.485 2902.310 4707.765 ;
        RECT 2822.730 4703.270 2823.010 4703.550 ;
        RECT 2822.730 4701.770 2823.010 4702.050 ;
        RECT 2822.730 4700.270 2823.010 4700.550 ;
        RECT 2871.035 4703.720 2871.315 4704.000 ;
        RECT 2872.035 4703.720 2872.315 4704.000 ;
        RECT 2871.035 4702.220 2871.315 4702.500 ;
        RECT 2872.035 4702.220 2872.315 4702.500 ;
        RECT 2871.035 4700.720 2871.315 4701.000 ;
        RECT 2872.035 4700.720 2872.315 4701.000 ;
        RECT 2904.105 4703.300 2904.385 4703.580 ;
        RECT 2904.105 4701.800 2904.385 4702.080 ;
        RECT 2904.105 4700.300 2904.385 4700.580 ;
        RECT 2961.035 4710.720 2961.315 4711.000 ;
        RECT 2962.035 4710.720 2962.315 4711.000 ;
        RECT 2961.035 4709.220 2961.315 4709.500 ;
        RECT 2962.035 4709.220 2962.315 4709.500 ;
        RECT 2961.035 4707.720 2961.315 4708.000 ;
        RECT 2962.035 4707.720 2962.315 4708.000 ;
        RECT 3006.740 4703.680 3007.020 4703.960 ;
        RECT 3007.360 4703.680 3007.640 4703.960 ;
        RECT 3007.980 4703.680 3008.260 4703.960 ;
        RECT 3008.600 4703.680 3008.880 4703.960 ;
        RECT 3009.220 4703.680 3009.500 4703.960 ;
        RECT 3009.840 4703.680 3010.120 4703.960 ;
        RECT 3010.460 4703.680 3010.740 4703.960 ;
        RECT 3011.080 4703.680 3011.360 4703.960 ;
        RECT 3011.700 4703.680 3011.980 4703.960 ;
        RECT 3012.320 4703.680 3012.600 4703.960 ;
        RECT 3012.940 4703.680 3013.220 4703.960 ;
        RECT 3013.560 4703.680 3013.840 4703.960 ;
        RECT 3014.180 4703.680 3014.460 4703.960 ;
        RECT 3014.800 4703.680 3015.080 4703.960 ;
        RECT 3015.420 4703.680 3015.700 4703.960 ;
        RECT 3006.740 4703.060 3007.020 4703.340 ;
        RECT 3007.360 4703.060 3007.640 4703.340 ;
        RECT 3007.980 4703.060 3008.260 4703.340 ;
        RECT 3008.600 4703.060 3008.880 4703.340 ;
        RECT 3009.220 4703.060 3009.500 4703.340 ;
        RECT 3009.840 4703.060 3010.120 4703.340 ;
        RECT 3010.460 4703.060 3010.740 4703.340 ;
        RECT 3011.080 4703.060 3011.360 4703.340 ;
        RECT 3011.700 4703.060 3011.980 4703.340 ;
        RECT 3012.320 4703.060 3012.600 4703.340 ;
        RECT 3012.940 4703.060 3013.220 4703.340 ;
        RECT 3013.560 4703.060 3013.840 4703.340 ;
        RECT 3014.180 4703.060 3014.460 4703.340 ;
        RECT 3014.800 4703.060 3015.080 4703.340 ;
        RECT 3015.420 4703.060 3015.700 4703.340 ;
        RECT 3006.740 4702.440 3007.020 4702.720 ;
        RECT 3007.360 4702.440 3007.640 4702.720 ;
        RECT 3007.980 4702.440 3008.260 4702.720 ;
        RECT 3008.600 4702.440 3008.880 4702.720 ;
        RECT 3009.220 4702.440 3009.500 4702.720 ;
        RECT 3009.840 4702.440 3010.120 4702.720 ;
        RECT 3010.460 4702.440 3010.740 4702.720 ;
        RECT 3011.080 4702.440 3011.360 4702.720 ;
        RECT 3011.700 4702.440 3011.980 4702.720 ;
        RECT 3012.320 4702.440 3012.600 4702.720 ;
        RECT 3012.940 4702.440 3013.220 4702.720 ;
        RECT 3013.560 4702.440 3013.840 4702.720 ;
        RECT 3014.180 4702.440 3014.460 4702.720 ;
        RECT 3014.800 4702.440 3015.080 4702.720 ;
        RECT 3015.420 4702.440 3015.700 4702.720 ;
        RECT 3006.740 4701.820 3007.020 4702.100 ;
        RECT 3007.360 4701.820 3007.640 4702.100 ;
        RECT 3007.980 4701.820 3008.260 4702.100 ;
        RECT 3008.600 4701.820 3008.880 4702.100 ;
        RECT 3009.220 4701.820 3009.500 4702.100 ;
        RECT 3009.840 4701.820 3010.120 4702.100 ;
        RECT 3010.460 4701.820 3010.740 4702.100 ;
        RECT 3011.080 4701.820 3011.360 4702.100 ;
        RECT 3011.700 4701.820 3011.980 4702.100 ;
        RECT 3012.320 4701.820 3012.600 4702.100 ;
        RECT 3012.940 4701.820 3013.220 4702.100 ;
        RECT 3013.560 4701.820 3013.840 4702.100 ;
        RECT 3014.180 4701.820 3014.460 4702.100 ;
        RECT 3014.800 4701.820 3015.080 4702.100 ;
        RECT 3015.420 4701.820 3015.700 4702.100 ;
        RECT 3006.740 4701.200 3007.020 4701.480 ;
        RECT 3007.360 4701.200 3007.640 4701.480 ;
        RECT 3007.980 4701.200 3008.260 4701.480 ;
        RECT 3008.600 4701.200 3008.880 4701.480 ;
        RECT 3009.220 4701.200 3009.500 4701.480 ;
        RECT 3009.840 4701.200 3010.120 4701.480 ;
        RECT 3010.460 4701.200 3010.740 4701.480 ;
        RECT 3011.080 4701.200 3011.360 4701.480 ;
        RECT 3011.700 4701.200 3011.980 4701.480 ;
        RECT 3012.320 4701.200 3012.600 4701.480 ;
        RECT 3012.940 4701.200 3013.220 4701.480 ;
        RECT 3013.560 4701.200 3013.840 4701.480 ;
        RECT 3014.180 4701.200 3014.460 4701.480 ;
        RECT 3014.800 4701.200 3015.080 4701.480 ;
        RECT 3015.420 4701.200 3015.700 4701.480 ;
        RECT 3006.740 4700.580 3007.020 4700.860 ;
        RECT 3007.360 4700.580 3007.640 4700.860 ;
        RECT 3007.980 4700.580 3008.260 4700.860 ;
        RECT 3008.600 4700.580 3008.880 4700.860 ;
        RECT 3009.220 4700.580 3009.500 4700.860 ;
        RECT 3009.840 4700.580 3010.120 4700.860 ;
        RECT 3010.460 4700.580 3010.740 4700.860 ;
        RECT 3011.080 4700.580 3011.360 4700.860 ;
        RECT 3011.700 4700.580 3011.980 4700.860 ;
        RECT 3012.320 4700.580 3012.600 4700.860 ;
        RECT 3012.940 4700.580 3013.220 4700.860 ;
        RECT 3013.560 4700.580 3013.840 4700.860 ;
        RECT 3014.180 4700.580 3014.460 4700.860 ;
        RECT 3014.800 4700.580 3015.080 4700.860 ;
        RECT 3015.420 4700.580 3015.700 4700.860 ;
        RECT 3006.740 4699.960 3007.020 4700.240 ;
        RECT 3007.360 4699.960 3007.640 4700.240 ;
        RECT 3007.980 4699.960 3008.260 4700.240 ;
        RECT 3008.600 4699.960 3008.880 4700.240 ;
        RECT 3009.220 4699.960 3009.500 4700.240 ;
        RECT 3009.840 4699.960 3010.120 4700.240 ;
        RECT 3010.460 4699.960 3010.740 4700.240 ;
        RECT 3011.080 4699.960 3011.360 4700.240 ;
        RECT 3011.700 4699.960 3011.980 4700.240 ;
        RECT 3012.320 4699.960 3012.600 4700.240 ;
        RECT 3012.940 4699.960 3013.220 4700.240 ;
        RECT 3013.560 4699.960 3013.840 4700.240 ;
        RECT 3014.180 4699.960 3014.460 4700.240 ;
        RECT 3014.800 4699.960 3015.080 4700.240 ;
        RECT 3015.420 4699.960 3015.700 4700.240 ;
        RECT 3019.140 4703.680 3019.420 4703.960 ;
        RECT 3019.760 4703.680 3020.040 4703.960 ;
        RECT 3020.380 4703.680 3020.660 4703.960 ;
        RECT 3021.000 4703.680 3021.280 4703.960 ;
        RECT 3021.620 4703.680 3021.900 4703.960 ;
        RECT 3022.240 4703.680 3022.520 4703.960 ;
        RECT 3022.860 4703.680 3023.140 4703.960 ;
        RECT 3023.480 4703.680 3023.760 4703.960 ;
        RECT 3024.100 4703.680 3024.380 4703.960 ;
        RECT 3024.720 4703.680 3025.000 4703.960 ;
        RECT 3025.340 4703.680 3025.620 4703.960 ;
        RECT 3025.960 4703.680 3026.240 4703.960 ;
        RECT 3026.580 4703.680 3026.860 4703.960 ;
        RECT 3027.200 4703.680 3027.480 4703.960 ;
        RECT 3027.820 4703.680 3028.100 4703.960 ;
        RECT 3028.440 4703.680 3028.720 4703.960 ;
        RECT 3019.140 4703.060 3019.420 4703.340 ;
        RECT 3019.760 4703.060 3020.040 4703.340 ;
        RECT 3020.380 4703.060 3020.660 4703.340 ;
        RECT 3021.000 4703.060 3021.280 4703.340 ;
        RECT 3021.620 4703.060 3021.900 4703.340 ;
        RECT 3022.240 4703.060 3022.520 4703.340 ;
        RECT 3022.860 4703.060 3023.140 4703.340 ;
        RECT 3023.480 4703.060 3023.760 4703.340 ;
        RECT 3024.100 4703.060 3024.380 4703.340 ;
        RECT 3024.720 4703.060 3025.000 4703.340 ;
        RECT 3025.340 4703.060 3025.620 4703.340 ;
        RECT 3025.960 4703.060 3026.240 4703.340 ;
        RECT 3026.580 4703.060 3026.860 4703.340 ;
        RECT 3027.200 4703.060 3027.480 4703.340 ;
        RECT 3027.820 4703.060 3028.100 4703.340 ;
        RECT 3028.440 4703.060 3028.720 4703.340 ;
        RECT 3019.140 4702.440 3019.420 4702.720 ;
        RECT 3019.760 4702.440 3020.040 4702.720 ;
        RECT 3020.380 4702.440 3020.660 4702.720 ;
        RECT 3021.000 4702.440 3021.280 4702.720 ;
        RECT 3021.620 4702.440 3021.900 4702.720 ;
        RECT 3022.240 4702.440 3022.520 4702.720 ;
        RECT 3022.860 4702.440 3023.140 4702.720 ;
        RECT 3023.480 4702.440 3023.760 4702.720 ;
        RECT 3024.100 4702.440 3024.380 4702.720 ;
        RECT 3024.720 4702.440 3025.000 4702.720 ;
        RECT 3025.340 4702.440 3025.620 4702.720 ;
        RECT 3025.960 4702.440 3026.240 4702.720 ;
        RECT 3026.580 4702.440 3026.860 4702.720 ;
        RECT 3027.200 4702.440 3027.480 4702.720 ;
        RECT 3027.820 4702.440 3028.100 4702.720 ;
        RECT 3028.440 4702.440 3028.720 4702.720 ;
        RECT 3019.140 4701.820 3019.420 4702.100 ;
        RECT 3019.760 4701.820 3020.040 4702.100 ;
        RECT 3020.380 4701.820 3020.660 4702.100 ;
        RECT 3021.000 4701.820 3021.280 4702.100 ;
        RECT 3021.620 4701.820 3021.900 4702.100 ;
        RECT 3022.240 4701.820 3022.520 4702.100 ;
        RECT 3022.860 4701.820 3023.140 4702.100 ;
        RECT 3023.480 4701.820 3023.760 4702.100 ;
        RECT 3024.100 4701.820 3024.380 4702.100 ;
        RECT 3024.720 4701.820 3025.000 4702.100 ;
        RECT 3025.340 4701.820 3025.620 4702.100 ;
        RECT 3025.960 4701.820 3026.240 4702.100 ;
        RECT 3026.580 4701.820 3026.860 4702.100 ;
        RECT 3027.200 4701.820 3027.480 4702.100 ;
        RECT 3027.820 4701.820 3028.100 4702.100 ;
        RECT 3028.440 4701.820 3028.720 4702.100 ;
        RECT 3019.140 4701.200 3019.420 4701.480 ;
        RECT 3019.760 4701.200 3020.040 4701.480 ;
        RECT 3020.380 4701.200 3020.660 4701.480 ;
        RECT 3021.000 4701.200 3021.280 4701.480 ;
        RECT 3021.620 4701.200 3021.900 4701.480 ;
        RECT 3022.240 4701.200 3022.520 4701.480 ;
        RECT 3022.860 4701.200 3023.140 4701.480 ;
        RECT 3023.480 4701.200 3023.760 4701.480 ;
        RECT 3024.100 4701.200 3024.380 4701.480 ;
        RECT 3024.720 4701.200 3025.000 4701.480 ;
        RECT 3025.340 4701.200 3025.620 4701.480 ;
        RECT 3025.960 4701.200 3026.240 4701.480 ;
        RECT 3026.580 4701.200 3026.860 4701.480 ;
        RECT 3027.200 4701.200 3027.480 4701.480 ;
        RECT 3027.820 4701.200 3028.100 4701.480 ;
        RECT 3028.440 4701.200 3028.720 4701.480 ;
        RECT 3019.140 4700.580 3019.420 4700.860 ;
        RECT 3019.760 4700.580 3020.040 4700.860 ;
        RECT 3020.380 4700.580 3020.660 4700.860 ;
        RECT 3021.000 4700.580 3021.280 4700.860 ;
        RECT 3021.620 4700.580 3021.900 4700.860 ;
        RECT 3022.240 4700.580 3022.520 4700.860 ;
        RECT 3022.860 4700.580 3023.140 4700.860 ;
        RECT 3023.480 4700.580 3023.760 4700.860 ;
        RECT 3024.100 4700.580 3024.380 4700.860 ;
        RECT 3024.720 4700.580 3025.000 4700.860 ;
        RECT 3025.340 4700.580 3025.620 4700.860 ;
        RECT 3025.960 4700.580 3026.240 4700.860 ;
        RECT 3026.580 4700.580 3026.860 4700.860 ;
        RECT 3027.200 4700.580 3027.480 4700.860 ;
        RECT 3027.820 4700.580 3028.100 4700.860 ;
        RECT 3028.440 4700.580 3028.720 4700.860 ;
        RECT 3019.140 4699.960 3019.420 4700.240 ;
        RECT 3019.760 4699.960 3020.040 4700.240 ;
        RECT 3020.380 4699.960 3020.660 4700.240 ;
        RECT 3021.000 4699.960 3021.280 4700.240 ;
        RECT 3021.620 4699.960 3021.900 4700.240 ;
        RECT 3022.240 4699.960 3022.520 4700.240 ;
        RECT 3022.860 4699.960 3023.140 4700.240 ;
        RECT 3023.480 4699.960 3023.760 4700.240 ;
        RECT 3024.100 4699.960 3024.380 4700.240 ;
        RECT 3024.720 4699.960 3025.000 4700.240 ;
        RECT 3025.340 4699.960 3025.620 4700.240 ;
        RECT 3025.960 4699.960 3026.240 4700.240 ;
        RECT 3026.580 4699.960 3026.860 4700.240 ;
        RECT 3027.200 4699.960 3027.480 4700.240 ;
        RECT 3027.820 4699.960 3028.100 4700.240 ;
        RECT 3028.440 4699.960 3028.720 4700.240 ;
        RECT 3030.990 4703.680 3031.270 4703.960 ;
        RECT 3031.610 4703.680 3031.890 4703.960 ;
        RECT 3032.230 4703.680 3032.510 4703.960 ;
        RECT 3032.850 4703.680 3033.130 4703.960 ;
        RECT 3033.470 4703.680 3033.750 4703.960 ;
        RECT 3034.090 4703.680 3034.370 4703.960 ;
        RECT 3034.710 4703.680 3034.990 4703.960 ;
        RECT 3035.330 4703.680 3035.610 4703.960 ;
        RECT 3035.950 4703.680 3036.230 4703.960 ;
        RECT 3036.570 4703.680 3036.850 4703.960 ;
        RECT 3037.190 4703.680 3037.470 4703.960 ;
        RECT 3037.810 4703.680 3038.090 4703.960 ;
        RECT 3038.430 4703.680 3038.710 4703.960 ;
        RECT 3039.050 4703.680 3039.330 4703.960 ;
        RECT 3039.670 4703.680 3039.950 4703.960 ;
        RECT 3040.290 4703.680 3040.570 4703.960 ;
        RECT 3030.990 4703.060 3031.270 4703.340 ;
        RECT 3031.610 4703.060 3031.890 4703.340 ;
        RECT 3032.230 4703.060 3032.510 4703.340 ;
        RECT 3032.850 4703.060 3033.130 4703.340 ;
        RECT 3033.470 4703.060 3033.750 4703.340 ;
        RECT 3034.090 4703.060 3034.370 4703.340 ;
        RECT 3034.710 4703.060 3034.990 4703.340 ;
        RECT 3035.330 4703.060 3035.610 4703.340 ;
        RECT 3035.950 4703.060 3036.230 4703.340 ;
        RECT 3036.570 4703.060 3036.850 4703.340 ;
        RECT 3037.190 4703.060 3037.470 4703.340 ;
        RECT 3037.810 4703.060 3038.090 4703.340 ;
        RECT 3038.430 4703.060 3038.710 4703.340 ;
        RECT 3039.050 4703.060 3039.330 4703.340 ;
        RECT 3039.670 4703.060 3039.950 4703.340 ;
        RECT 3040.290 4703.060 3040.570 4703.340 ;
        RECT 3030.990 4702.440 3031.270 4702.720 ;
        RECT 3031.610 4702.440 3031.890 4702.720 ;
        RECT 3032.230 4702.440 3032.510 4702.720 ;
        RECT 3032.850 4702.440 3033.130 4702.720 ;
        RECT 3033.470 4702.440 3033.750 4702.720 ;
        RECT 3034.090 4702.440 3034.370 4702.720 ;
        RECT 3034.710 4702.440 3034.990 4702.720 ;
        RECT 3035.330 4702.440 3035.610 4702.720 ;
        RECT 3035.950 4702.440 3036.230 4702.720 ;
        RECT 3036.570 4702.440 3036.850 4702.720 ;
        RECT 3037.190 4702.440 3037.470 4702.720 ;
        RECT 3037.810 4702.440 3038.090 4702.720 ;
        RECT 3038.430 4702.440 3038.710 4702.720 ;
        RECT 3039.050 4702.440 3039.330 4702.720 ;
        RECT 3039.670 4702.440 3039.950 4702.720 ;
        RECT 3040.290 4702.440 3040.570 4702.720 ;
        RECT 3030.990 4701.820 3031.270 4702.100 ;
        RECT 3031.610 4701.820 3031.890 4702.100 ;
        RECT 3032.230 4701.820 3032.510 4702.100 ;
        RECT 3032.850 4701.820 3033.130 4702.100 ;
        RECT 3033.470 4701.820 3033.750 4702.100 ;
        RECT 3034.090 4701.820 3034.370 4702.100 ;
        RECT 3034.710 4701.820 3034.990 4702.100 ;
        RECT 3035.330 4701.820 3035.610 4702.100 ;
        RECT 3035.950 4701.820 3036.230 4702.100 ;
        RECT 3036.570 4701.820 3036.850 4702.100 ;
        RECT 3037.190 4701.820 3037.470 4702.100 ;
        RECT 3037.810 4701.820 3038.090 4702.100 ;
        RECT 3038.430 4701.820 3038.710 4702.100 ;
        RECT 3039.050 4701.820 3039.330 4702.100 ;
        RECT 3039.670 4701.820 3039.950 4702.100 ;
        RECT 3040.290 4701.820 3040.570 4702.100 ;
        RECT 3030.990 4701.200 3031.270 4701.480 ;
        RECT 3031.610 4701.200 3031.890 4701.480 ;
        RECT 3032.230 4701.200 3032.510 4701.480 ;
        RECT 3032.850 4701.200 3033.130 4701.480 ;
        RECT 3033.470 4701.200 3033.750 4701.480 ;
        RECT 3034.090 4701.200 3034.370 4701.480 ;
        RECT 3034.710 4701.200 3034.990 4701.480 ;
        RECT 3035.330 4701.200 3035.610 4701.480 ;
        RECT 3035.950 4701.200 3036.230 4701.480 ;
        RECT 3036.570 4701.200 3036.850 4701.480 ;
        RECT 3037.190 4701.200 3037.470 4701.480 ;
        RECT 3037.810 4701.200 3038.090 4701.480 ;
        RECT 3038.430 4701.200 3038.710 4701.480 ;
        RECT 3039.050 4701.200 3039.330 4701.480 ;
        RECT 3039.670 4701.200 3039.950 4701.480 ;
        RECT 3040.290 4701.200 3040.570 4701.480 ;
        RECT 3030.990 4700.580 3031.270 4700.860 ;
        RECT 3031.610 4700.580 3031.890 4700.860 ;
        RECT 3032.230 4700.580 3032.510 4700.860 ;
        RECT 3032.850 4700.580 3033.130 4700.860 ;
        RECT 3033.470 4700.580 3033.750 4700.860 ;
        RECT 3034.090 4700.580 3034.370 4700.860 ;
        RECT 3034.710 4700.580 3034.990 4700.860 ;
        RECT 3035.330 4700.580 3035.610 4700.860 ;
        RECT 3035.950 4700.580 3036.230 4700.860 ;
        RECT 3036.570 4700.580 3036.850 4700.860 ;
        RECT 3037.190 4700.580 3037.470 4700.860 ;
        RECT 3037.810 4700.580 3038.090 4700.860 ;
        RECT 3038.430 4700.580 3038.710 4700.860 ;
        RECT 3039.050 4700.580 3039.330 4700.860 ;
        RECT 3039.670 4700.580 3039.950 4700.860 ;
        RECT 3040.290 4700.580 3040.570 4700.860 ;
        RECT 3030.990 4699.960 3031.270 4700.240 ;
        RECT 3031.610 4699.960 3031.890 4700.240 ;
        RECT 3032.230 4699.960 3032.510 4700.240 ;
        RECT 3032.850 4699.960 3033.130 4700.240 ;
        RECT 3033.470 4699.960 3033.750 4700.240 ;
        RECT 3034.090 4699.960 3034.370 4700.240 ;
        RECT 3034.710 4699.960 3034.990 4700.240 ;
        RECT 3035.330 4699.960 3035.610 4700.240 ;
        RECT 3035.950 4699.960 3036.230 4700.240 ;
        RECT 3036.570 4699.960 3036.850 4700.240 ;
        RECT 3037.190 4699.960 3037.470 4700.240 ;
        RECT 3037.810 4699.960 3038.090 4700.240 ;
        RECT 3038.430 4699.960 3038.710 4700.240 ;
        RECT 3039.050 4699.960 3039.330 4700.240 ;
        RECT 3039.670 4699.960 3039.950 4700.240 ;
        RECT 3040.290 4699.960 3040.570 4700.240 ;
        RECT 3044.520 4703.680 3044.800 4703.960 ;
        RECT 3045.140 4703.680 3045.420 4703.960 ;
        RECT 3045.760 4703.680 3046.040 4703.960 ;
        RECT 3046.380 4703.680 3046.660 4703.960 ;
        RECT 3047.000 4703.680 3047.280 4703.960 ;
        RECT 3047.620 4703.680 3047.900 4703.960 ;
        RECT 3048.240 4703.680 3048.520 4703.960 ;
        RECT 3048.860 4703.680 3049.140 4703.960 ;
        RECT 3049.480 4703.680 3049.760 4703.960 ;
        RECT 3050.100 4703.680 3050.380 4703.960 ;
        RECT 3050.720 4703.680 3051.000 4703.960 ;
        RECT 3051.340 4703.680 3051.620 4703.960 ;
        RECT 3051.960 4703.680 3052.240 4703.960 ;
        RECT 3052.580 4703.680 3052.860 4703.960 ;
        RECT 3053.200 4703.680 3053.480 4703.960 ;
        RECT 3053.820 4703.680 3054.100 4703.960 ;
        RECT 3044.520 4703.060 3044.800 4703.340 ;
        RECT 3045.140 4703.060 3045.420 4703.340 ;
        RECT 3045.760 4703.060 3046.040 4703.340 ;
        RECT 3046.380 4703.060 3046.660 4703.340 ;
        RECT 3047.000 4703.060 3047.280 4703.340 ;
        RECT 3047.620 4703.060 3047.900 4703.340 ;
        RECT 3048.240 4703.060 3048.520 4703.340 ;
        RECT 3048.860 4703.060 3049.140 4703.340 ;
        RECT 3049.480 4703.060 3049.760 4703.340 ;
        RECT 3050.100 4703.060 3050.380 4703.340 ;
        RECT 3050.720 4703.060 3051.000 4703.340 ;
        RECT 3051.340 4703.060 3051.620 4703.340 ;
        RECT 3051.960 4703.060 3052.240 4703.340 ;
        RECT 3052.580 4703.060 3052.860 4703.340 ;
        RECT 3053.200 4703.060 3053.480 4703.340 ;
        RECT 3053.820 4703.060 3054.100 4703.340 ;
        RECT 3044.520 4702.440 3044.800 4702.720 ;
        RECT 3045.140 4702.440 3045.420 4702.720 ;
        RECT 3045.760 4702.440 3046.040 4702.720 ;
        RECT 3046.380 4702.440 3046.660 4702.720 ;
        RECT 3047.000 4702.440 3047.280 4702.720 ;
        RECT 3047.620 4702.440 3047.900 4702.720 ;
        RECT 3048.240 4702.440 3048.520 4702.720 ;
        RECT 3048.860 4702.440 3049.140 4702.720 ;
        RECT 3049.480 4702.440 3049.760 4702.720 ;
        RECT 3050.100 4702.440 3050.380 4702.720 ;
        RECT 3050.720 4702.440 3051.000 4702.720 ;
        RECT 3051.340 4702.440 3051.620 4702.720 ;
        RECT 3051.960 4702.440 3052.240 4702.720 ;
        RECT 3052.580 4702.440 3052.860 4702.720 ;
        RECT 3053.200 4702.440 3053.480 4702.720 ;
        RECT 3053.820 4702.440 3054.100 4702.720 ;
        RECT 3044.520 4701.820 3044.800 4702.100 ;
        RECT 3045.140 4701.820 3045.420 4702.100 ;
        RECT 3045.760 4701.820 3046.040 4702.100 ;
        RECT 3046.380 4701.820 3046.660 4702.100 ;
        RECT 3047.000 4701.820 3047.280 4702.100 ;
        RECT 3047.620 4701.820 3047.900 4702.100 ;
        RECT 3048.240 4701.820 3048.520 4702.100 ;
        RECT 3048.860 4701.820 3049.140 4702.100 ;
        RECT 3049.480 4701.820 3049.760 4702.100 ;
        RECT 3050.100 4701.820 3050.380 4702.100 ;
        RECT 3050.720 4701.820 3051.000 4702.100 ;
        RECT 3051.340 4701.820 3051.620 4702.100 ;
        RECT 3051.960 4701.820 3052.240 4702.100 ;
        RECT 3052.580 4701.820 3052.860 4702.100 ;
        RECT 3053.200 4701.820 3053.480 4702.100 ;
        RECT 3053.820 4701.820 3054.100 4702.100 ;
        RECT 3044.520 4701.200 3044.800 4701.480 ;
        RECT 3045.140 4701.200 3045.420 4701.480 ;
        RECT 3045.760 4701.200 3046.040 4701.480 ;
        RECT 3046.380 4701.200 3046.660 4701.480 ;
        RECT 3047.000 4701.200 3047.280 4701.480 ;
        RECT 3047.620 4701.200 3047.900 4701.480 ;
        RECT 3048.240 4701.200 3048.520 4701.480 ;
        RECT 3048.860 4701.200 3049.140 4701.480 ;
        RECT 3049.480 4701.200 3049.760 4701.480 ;
        RECT 3050.100 4701.200 3050.380 4701.480 ;
        RECT 3050.720 4701.200 3051.000 4701.480 ;
        RECT 3051.340 4701.200 3051.620 4701.480 ;
        RECT 3051.960 4701.200 3052.240 4701.480 ;
        RECT 3052.580 4701.200 3052.860 4701.480 ;
        RECT 3053.200 4701.200 3053.480 4701.480 ;
        RECT 3053.820 4701.200 3054.100 4701.480 ;
        RECT 3044.520 4700.580 3044.800 4700.860 ;
        RECT 3045.140 4700.580 3045.420 4700.860 ;
        RECT 3045.760 4700.580 3046.040 4700.860 ;
        RECT 3046.380 4700.580 3046.660 4700.860 ;
        RECT 3047.000 4700.580 3047.280 4700.860 ;
        RECT 3047.620 4700.580 3047.900 4700.860 ;
        RECT 3048.240 4700.580 3048.520 4700.860 ;
        RECT 3048.860 4700.580 3049.140 4700.860 ;
        RECT 3049.480 4700.580 3049.760 4700.860 ;
        RECT 3050.100 4700.580 3050.380 4700.860 ;
        RECT 3050.720 4700.580 3051.000 4700.860 ;
        RECT 3051.340 4700.580 3051.620 4700.860 ;
        RECT 3051.960 4700.580 3052.240 4700.860 ;
        RECT 3052.580 4700.580 3052.860 4700.860 ;
        RECT 3053.200 4700.580 3053.480 4700.860 ;
        RECT 3053.820 4700.580 3054.100 4700.860 ;
        RECT 3044.520 4699.960 3044.800 4700.240 ;
        RECT 3045.140 4699.960 3045.420 4700.240 ;
        RECT 3045.760 4699.960 3046.040 4700.240 ;
        RECT 3046.380 4699.960 3046.660 4700.240 ;
        RECT 3047.000 4699.960 3047.280 4700.240 ;
        RECT 3047.620 4699.960 3047.900 4700.240 ;
        RECT 3048.240 4699.960 3048.520 4700.240 ;
        RECT 3048.860 4699.960 3049.140 4700.240 ;
        RECT 3049.480 4699.960 3049.760 4700.240 ;
        RECT 3050.100 4699.960 3050.380 4700.240 ;
        RECT 3050.720 4699.960 3051.000 4700.240 ;
        RECT 3051.340 4699.960 3051.620 4700.240 ;
        RECT 3051.960 4699.960 3052.240 4700.240 ;
        RECT 3052.580 4699.960 3052.860 4700.240 ;
        RECT 3053.200 4699.960 3053.480 4700.240 ;
        RECT 3053.820 4699.960 3054.100 4700.240 ;
        RECT 3056.370 4703.680 3056.650 4703.960 ;
        RECT 3056.990 4703.680 3057.270 4703.960 ;
        RECT 3057.610 4703.680 3057.890 4703.960 ;
        RECT 3058.230 4703.680 3058.510 4703.960 ;
        RECT 3058.850 4703.680 3059.130 4703.960 ;
        RECT 3059.470 4703.680 3059.750 4703.960 ;
        RECT 3060.090 4703.680 3060.370 4703.960 ;
        RECT 3060.710 4703.680 3060.990 4703.960 ;
        RECT 3061.330 4703.680 3061.610 4703.960 ;
        RECT 3061.950 4703.680 3062.230 4703.960 ;
        RECT 3062.570 4703.680 3062.850 4703.960 ;
        RECT 3063.190 4703.680 3063.470 4703.960 ;
        RECT 3063.810 4703.680 3064.090 4703.960 ;
        RECT 3064.430 4703.680 3064.710 4703.960 ;
        RECT 3065.050 4703.680 3065.330 4703.960 ;
        RECT 3065.670 4703.680 3065.950 4703.960 ;
        RECT 3056.370 4703.060 3056.650 4703.340 ;
        RECT 3056.990 4703.060 3057.270 4703.340 ;
        RECT 3057.610 4703.060 3057.890 4703.340 ;
        RECT 3058.230 4703.060 3058.510 4703.340 ;
        RECT 3058.850 4703.060 3059.130 4703.340 ;
        RECT 3059.470 4703.060 3059.750 4703.340 ;
        RECT 3060.090 4703.060 3060.370 4703.340 ;
        RECT 3060.710 4703.060 3060.990 4703.340 ;
        RECT 3061.330 4703.060 3061.610 4703.340 ;
        RECT 3061.950 4703.060 3062.230 4703.340 ;
        RECT 3062.570 4703.060 3062.850 4703.340 ;
        RECT 3063.190 4703.060 3063.470 4703.340 ;
        RECT 3063.810 4703.060 3064.090 4703.340 ;
        RECT 3064.430 4703.060 3064.710 4703.340 ;
        RECT 3065.050 4703.060 3065.330 4703.340 ;
        RECT 3065.670 4703.060 3065.950 4703.340 ;
        RECT 3056.370 4702.440 3056.650 4702.720 ;
        RECT 3056.990 4702.440 3057.270 4702.720 ;
        RECT 3057.610 4702.440 3057.890 4702.720 ;
        RECT 3058.230 4702.440 3058.510 4702.720 ;
        RECT 3058.850 4702.440 3059.130 4702.720 ;
        RECT 3059.470 4702.440 3059.750 4702.720 ;
        RECT 3060.090 4702.440 3060.370 4702.720 ;
        RECT 3060.710 4702.440 3060.990 4702.720 ;
        RECT 3061.330 4702.440 3061.610 4702.720 ;
        RECT 3061.950 4702.440 3062.230 4702.720 ;
        RECT 3062.570 4702.440 3062.850 4702.720 ;
        RECT 3063.190 4702.440 3063.470 4702.720 ;
        RECT 3063.810 4702.440 3064.090 4702.720 ;
        RECT 3064.430 4702.440 3064.710 4702.720 ;
        RECT 3065.050 4702.440 3065.330 4702.720 ;
        RECT 3065.670 4702.440 3065.950 4702.720 ;
        RECT 3056.370 4701.820 3056.650 4702.100 ;
        RECT 3056.990 4701.820 3057.270 4702.100 ;
        RECT 3057.610 4701.820 3057.890 4702.100 ;
        RECT 3058.230 4701.820 3058.510 4702.100 ;
        RECT 3058.850 4701.820 3059.130 4702.100 ;
        RECT 3059.470 4701.820 3059.750 4702.100 ;
        RECT 3060.090 4701.820 3060.370 4702.100 ;
        RECT 3060.710 4701.820 3060.990 4702.100 ;
        RECT 3061.330 4701.820 3061.610 4702.100 ;
        RECT 3061.950 4701.820 3062.230 4702.100 ;
        RECT 3062.570 4701.820 3062.850 4702.100 ;
        RECT 3063.190 4701.820 3063.470 4702.100 ;
        RECT 3063.810 4701.820 3064.090 4702.100 ;
        RECT 3064.430 4701.820 3064.710 4702.100 ;
        RECT 3065.050 4701.820 3065.330 4702.100 ;
        RECT 3065.670 4701.820 3065.950 4702.100 ;
        RECT 3056.370 4701.200 3056.650 4701.480 ;
        RECT 3056.990 4701.200 3057.270 4701.480 ;
        RECT 3057.610 4701.200 3057.890 4701.480 ;
        RECT 3058.230 4701.200 3058.510 4701.480 ;
        RECT 3058.850 4701.200 3059.130 4701.480 ;
        RECT 3059.470 4701.200 3059.750 4701.480 ;
        RECT 3060.090 4701.200 3060.370 4701.480 ;
        RECT 3060.710 4701.200 3060.990 4701.480 ;
        RECT 3061.330 4701.200 3061.610 4701.480 ;
        RECT 3061.950 4701.200 3062.230 4701.480 ;
        RECT 3062.570 4701.200 3062.850 4701.480 ;
        RECT 3063.190 4701.200 3063.470 4701.480 ;
        RECT 3063.810 4701.200 3064.090 4701.480 ;
        RECT 3064.430 4701.200 3064.710 4701.480 ;
        RECT 3065.050 4701.200 3065.330 4701.480 ;
        RECT 3065.670 4701.200 3065.950 4701.480 ;
        RECT 3056.370 4700.580 3056.650 4700.860 ;
        RECT 3056.990 4700.580 3057.270 4700.860 ;
        RECT 3057.610 4700.580 3057.890 4700.860 ;
        RECT 3058.230 4700.580 3058.510 4700.860 ;
        RECT 3058.850 4700.580 3059.130 4700.860 ;
        RECT 3059.470 4700.580 3059.750 4700.860 ;
        RECT 3060.090 4700.580 3060.370 4700.860 ;
        RECT 3060.710 4700.580 3060.990 4700.860 ;
        RECT 3061.330 4700.580 3061.610 4700.860 ;
        RECT 3061.950 4700.580 3062.230 4700.860 ;
        RECT 3062.570 4700.580 3062.850 4700.860 ;
        RECT 3063.190 4700.580 3063.470 4700.860 ;
        RECT 3063.810 4700.580 3064.090 4700.860 ;
        RECT 3064.430 4700.580 3064.710 4700.860 ;
        RECT 3065.050 4700.580 3065.330 4700.860 ;
        RECT 3065.670 4700.580 3065.950 4700.860 ;
        RECT 3056.370 4699.960 3056.650 4700.240 ;
        RECT 3056.990 4699.960 3057.270 4700.240 ;
        RECT 3057.610 4699.960 3057.890 4700.240 ;
        RECT 3058.230 4699.960 3058.510 4700.240 ;
        RECT 3058.850 4699.960 3059.130 4700.240 ;
        RECT 3059.470 4699.960 3059.750 4700.240 ;
        RECT 3060.090 4699.960 3060.370 4700.240 ;
        RECT 3060.710 4699.960 3060.990 4700.240 ;
        RECT 3061.330 4699.960 3061.610 4700.240 ;
        RECT 3061.950 4699.960 3062.230 4700.240 ;
        RECT 3062.570 4699.960 3062.850 4700.240 ;
        RECT 3063.190 4699.960 3063.470 4700.240 ;
        RECT 3063.810 4699.960 3064.090 4700.240 ;
        RECT 3064.430 4699.960 3064.710 4700.240 ;
        RECT 3065.050 4699.960 3065.330 4700.240 ;
        RECT 3065.670 4699.960 3065.950 4700.240 ;
        RECT 3302.740 4716.895 3303.020 4717.175 ;
        RECT 3069.390 4703.680 3069.670 4703.960 ;
        RECT 3070.010 4703.680 3070.290 4703.960 ;
        RECT 3070.630 4703.680 3070.910 4703.960 ;
        RECT 3071.250 4703.680 3071.530 4703.960 ;
        RECT 3071.870 4703.680 3072.150 4703.960 ;
        RECT 3072.490 4703.680 3072.770 4703.960 ;
        RECT 3073.110 4703.680 3073.390 4703.960 ;
        RECT 3073.730 4703.680 3074.010 4703.960 ;
        RECT 3074.350 4703.680 3074.630 4703.960 ;
        RECT 3074.970 4703.680 3075.250 4703.960 ;
        RECT 3075.590 4703.680 3075.870 4703.960 ;
        RECT 3076.210 4703.680 3076.490 4703.960 ;
        RECT 3076.830 4703.680 3077.110 4703.960 ;
        RECT 3077.450 4703.680 3077.730 4703.960 ;
        RECT 3078.070 4703.680 3078.350 4703.960 ;
        RECT 3069.390 4703.060 3069.670 4703.340 ;
        RECT 3070.010 4703.060 3070.290 4703.340 ;
        RECT 3070.630 4703.060 3070.910 4703.340 ;
        RECT 3071.250 4703.060 3071.530 4703.340 ;
        RECT 3071.870 4703.060 3072.150 4703.340 ;
        RECT 3072.490 4703.060 3072.770 4703.340 ;
        RECT 3073.110 4703.060 3073.390 4703.340 ;
        RECT 3073.730 4703.060 3074.010 4703.340 ;
        RECT 3074.350 4703.060 3074.630 4703.340 ;
        RECT 3074.970 4703.060 3075.250 4703.340 ;
        RECT 3075.590 4703.060 3075.870 4703.340 ;
        RECT 3076.210 4703.060 3076.490 4703.340 ;
        RECT 3076.830 4703.060 3077.110 4703.340 ;
        RECT 3077.450 4703.060 3077.730 4703.340 ;
        RECT 3078.070 4703.060 3078.350 4703.340 ;
        RECT 3069.390 4702.440 3069.670 4702.720 ;
        RECT 3070.010 4702.440 3070.290 4702.720 ;
        RECT 3070.630 4702.440 3070.910 4702.720 ;
        RECT 3071.250 4702.440 3071.530 4702.720 ;
        RECT 3071.870 4702.440 3072.150 4702.720 ;
        RECT 3072.490 4702.440 3072.770 4702.720 ;
        RECT 3073.110 4702.440 3073.390 4702.720 ;
        RECT 3073.730 4702.440 3074.010 4702.720 ;
        RECT 3074.350 4702.440 3074.630 4702.720 ;
        RECT 3074.970 4702.440 3075.250 4702.720 ;
        RECT 3075.590 4702.440 3075.870 4702.720 ;
        RECT 3076.210 4702.440 3076.490 4702.720 ;
        RECT 3076.830 4702.440 3077.110 4702.720 ;
        RECT 3077.450 4702.440 3077.730 4702.720 ;
        RECT 3078.070 4702.440 3078.350 4702.720 ;
        RECT 3069.390 4701.820 3069.670 4702.100 ;
        RECT 3070.010 4701.820 3070.290 4702.100 ;
        RECT 3070.630 4701.820 3070.910 4702.100 ;
        RECT 3071.250 4701.820 3071.530 4702.100 ;
        RECT 3071.870 4701.820 3072.150 4702.100 ;
        RECT 3072.490 4701.820 3072.770 4702.100 ;
        RECT 3073.110 4701.820 3073.390 4702.100 ;
        RECT 3073.730 4701.820 3074.010 4702.100 ;
        RECT 3074.350 4701.820 3074.630 4702.100 ;
        RECT 3074.970 4701.820 3075.250 4702.100 ;
        RECT 3075.590 4701.820 3075.870 4702.100 ;
        RECT 3076.210 4701.820 3076.490 4702.100 ;
        RECT 3076.830 4701.820 3077.110 4702.100 ;
        RECT 3077.450 4701.820 3077.730 4702.100 ;
        RECT 3078.070 4701.820 3078.350 4702.100 ;
        RECT 3069.390 4701.200 3069.670 4701.480 ;
        RECT 3070.010 4701.200 3070.290 4701.480 ;
        RECT 3070.630 4701.200 3070.910 4701.480 ;
        RECT 3071.250 4701.200 3071.530 4701.480 ;
        RECT 3071.870 4701.200 3072.150 4701.480 ;
        RECT 3072.490 4701.200 3072.770 4701.480 ;
        RECT 3073.110 4701.200 3073.390 4701.480 ;
        RECT 3073.730 4701.200 3074.010 4701.480 ;
        RECT 3074.350 4701.200 3074.630 4701.480 ;
        RECT 3074.970 4701.200 3075.250 4701.480 ;
        RECT 3075.590 4701.200 3075.870 4701.480 ;
        RECT 3076.210 4701.200 3076.490 4701.480 ;
        RECT 3076.830 4701.200 3077.110 4701.480 ;
        RECT 3077.450 4701.200 3077.730 4701.480 ;
        RECT 3078.070 4701.200 3078.350 4701.480 ;
        RECT 3069.390 4700.580 3069.670 4700.860 ;
        RECT 3070.010 4700.580 3070.290 4700.860 ;
        RECT 3070.630 4700.580 3070.910 4700.860 ;
        RECT 3071.250 4700.580 3071.530 4700.860 ;
        RECT 3071.870 4700.580 3072.150 4700.860 ;
        RECT 3072.490 4700.580 3072.770 4700.860 ;
        RECT 3073.110 4700.580 3073.390 4700.860 ;
        RECT 3073.730 4700.580 3074.010 4700.860 ;
        RECT 3074.350 4700.580 3074.630 4700.860 ;
        RECT 3074.970 4700.580 3075.250 4700.860 ;
        RECT 3075.590 4700.580 3075.870 4700.860 ;
        RECT 3076.210 4700.580 3076.490 4700.860 ;
        RECT 3076.830 4700.580 3077.110 4700.860 ;
        RECT 3077.450 4700.580 3077.730 4700.860 ;
        RECT 3078.070 4700.580 3078.350 4700.860 ;
        RECT 3069.390 4699.960 3069.670 4700.240 ;
        RECT 3070.010 4699.960 3070.290 4700.240 ;
        RECT 3070.630 4699.960 3070.910 4700.240 ;
        RECT 3071.250 4699.960 3071.530 4700.240 ;
        RECT 3071.870 4699.960 3072.150 4700.240 ;
        RECT 3072.490 4699.960 3072.770 4700.240 ;
        RECT 3073.110 4699.960 3073.390 4700.240 ;
        RECT 3073.730 4699.960 3074.010 4700.240 ;
        RECT 3074.350 4699.960 3074.630 4700.240 ;
        RECT 3074.970 4699.960 3075.250 4700.240 ;
        RECT 3075.590 4699.960 3075.870 4700.240 ;
        RECT 3076.210 4699.960 3076.490 4700.240 ;
        RECT 3076.830 4699.960 3077.110 4700.240 ;
        RECT 3077.450 4699.960 3077.730 4700.240 ;
        RECT 3078.070 4699.960 3078.350 4700.240 ;
        RECT 3141.035 4710.720 3141.315 4711.000 ;
        RECT 3142.035 4710.720 3142.315 4711.000 ;
        RECT 3141.035 4709.220 3141.315 4709.500 ;
        RECT 3142.035 4709.220 3142.315 4709.500 ;
        RECT 3141.035 4707.720 3141.315 4708.000 ;
        RECT 3142.035 4707.720 3142.315 4708.000 ;
        RECT 3231.035 4703.720 3231.315 4704.000 ;
        RECT 3232.035 4703.720 3232.315 4704.000 ;
        RECT 3231.035 4702.220 3231.315 4702.500 ;
        RECT 3232.035 4702.220 3232.315 4702.500 ;
        RECT 3231.035 4700.720 3231.315 4701.000 ;
        RECT 3232.035 4700.720 3232.315 4701.000 ;
        RECT 3337.740 4716.895 3338.020 4717.175 ;
        RECT 3302.730 4703.270 3303.010 4703.550 ;
        RECT 3302.730 4701.770 3303.010 4702.050 ;
        RECT 3302.730 4700.270 3303.010 4700.550 ;
        RECT 3321.035 4710.720 3321.315 4711.000 ;
        RECT 3322.035 4710.720 3322.315 4711.000 ;
        RECT 3321.035 4709.220 3321.315 4709.500 ;
        RECT 3322.035 4709.220 3322.315 4709.500 ;
        RECT 3321.035 4707.720 3321.315 4708.000 ;
        RECT 3322.035 4707.720 3322.315 4708.000 ;
        RECT 3337.730 4703.270 3338.010 4703.550 ;
        RECT 3337.730 4701.770 3338.010 4702.050 ;
        RECT 3337.730 4700.270 3338.010 4700.550 ;
        RECT 3372.740 4716.895 3373.020 4717.175 ;
        RECT 3452.030 4710.485 3452.310 4710.765 ;
        RECT 3452.030 4708.985 3452.310 4709.265 ;
        RECT 3452.030 4707.485 3452.310 4707.765 ;
        RECT 3372.730 4703.270 3373.010 4703.550 ;
        RECT 3372.730 4701.770 3373.010 4702.050 ;
        RECT 3372.730 4700.270 3373.010 4700.550 ;
        RECT 3411.035 4703.720 3411.315 4704.000 ;
        RECT 3412.035 4703.720 3412.315 4704.000 ;
        RECT 3411.035 4702.220 3411.315 4702.500 ;
        RECT 3412.035 4702.220 3412.315 4702.500 ;
        RECT 3411.035 4700.720 3411.315 4701.000 ;
        RECT 3412.035 4700.720 3412.315 4701.000 ;
        RECT 3497.260 4710.680 3497.540 4710.960 ;
        RECT 3497.880 4710.680 3498.160 4710.960 ;
        RECT 3498.500 4710.680 3498.780 4710.960 ;
        RECT 3499.120 4710.680 3499.400 4710.960 ;
        RECT 3499.740 4710.680 3500.020 4710.960 ;
        RECT 3500.360 4710.680 3500.640 4710.960 ;
        RECT 3500.980 4710.680 3501.260 4710.960 ;
        RECT 3497.260 4710.060 3497.540 4710.340 ;
        RECT 3497.880 4710.060 3498.160 4710.340 ;
        RECT 3498.500 4710.060 3498.780 4710.340 ;
        RECT 3499.120 4710.060 3499.400 4710.340 ;
        RECT 3499.740 4710.060 3500.020 4710.340 ;
        RECT 3500.360 4710.060 3500.640 4710.340 ;
        RECT 3500.980 4710.060 3501.260 4710.340 ;
        RECT 3497.260 4709.440 3497.540 4709.720 ;
        RECT 3497.880 4709.440 3498.160 4709.720 ;
        RECT 3498.500 4709.440 3498.780 4709.720 ;
        RECT 3499.120 4709.440 3499.400 4709.720 ;
        RECT 3499.740 4709.440 3500.020 4709.720 ;
        RECT 3500.360 4709.440 3500.640 4709.720 ;
        RECT 3500.980 4709.440 3501.260 4709.720 ;
        RECT 3497.260 4708.820 3497.540 4709.100 ;
        RECT 3497.880 4708.820 3498.160 4709.100 ;
        RECT 3498.500 4708.820 3498.780 4709.100 ;
        RECT 3499.120 4708.820 3499.400 4709.100 ;
        RECT 3499.740 4708.820 3500.020 4709.100 ;
        RECT 3500.360 4708.820 3500.640 4709.100 ;
        RECT 3500.980 4708.820 3501.260 4709.100 ;
        RECT 3497.260 4708.200 3497.540 4708.480 ;
        RECT 3497.880 4708.200 3498.160 4708.480 ;
        RECT 3498.500 4708.200 3498.780 4708.480 ;
        RECT 3499.120 4708.200 3499.400 4708.480 ;
        RECT 3499.740 4708.200 3500.020 4708.480 ;
        RECT 3500.360 4708.200 3500.640 4708.480 ;
        RECT 3500.980 4708.200 3501.260 4708.480 ;
        RECT 3497.260 4707.580 3497.540 4707.860 ;
        RECT 3497.880 4707.580 3498.160 4707.860 ;
        RECT 3498.500 4707.580 3498.780 4707.860 ;
        RECT 3499.120 4707.580 3499.400 4707.860 ;
        RECT 3499.740 4707.580 3500.020 4707.860 ;
        RECT 3500.360 4707.580 3500.640 4707.860 ;
        RECT 3500.980 4707.580 3501.260 4707.860 ;
        RECT 3497.260 4706.960 3497.540 4707.240 ;
        RECT 3497.880 4706.960 3498.160 4707.240 ;
        RECT 3498.500 4706.960 3498.780 4707.240 ;
        RECT 3499.120 4706.960 3499.400 4707.240 ;
        RECT 3499.740 4706.960 3500.020 4707.240 ;
        RECT 3500.360 4706.960 3500.640 4707.240 ;
        RECT 3500.980 4706.960 3501.260 4707.240 ;
        RECT 3454.105 4703.300 3454.385 4703.580 ;
        RECT 3454.105 4701.800 3454.385 4702.080 ;
        RECT 3454.105 4700.300 3454.385 4700.580 ;
        RECT 3490.260 4703.680 3490.540 4703.960 ;
        RECT 3490.880 4703.680 3491.160 4703.960 ;
        RECT 3491.500 4703.680 3491.780 4703.960 ;
        RECT 3492.120 4703.680 3492.400 4703.960 ;
        RECT 3492.740 4703.680 3493.020 4703.960 ;
        RECT 3493.360 4703.680 3493.640 4703.960 ;
        RECT 3493.980 4703.680 3494.260 4703.960 ;
        RECT 3490.260 4703.060 3490.540 4703.340 ;
        RECT 3490.880 4703.060 3491.160 4703.340 ;
        RECT 3491.500 4703.060 3491.780 4703.340 ;
        RECT 3492.120 4703.060 3492.400 4703.340 ;
        RECT 3492.740 4703.060 3493.020 4703.340 ;
        RECT 3493.360 4703.060 3493.640 4703.340 ;
        RECT 3493.980 4703.060 3494.260 4703.340 ;
        RECT 3490.260 4702.440 3490.540 4702.720 ;
        RECT 3490.880 4702.440 3491.160 4702.720 ;
        RECT 3491.500 4702.440 3491.780 4702.720 ;
        RECT 3492.120 4702.440 3492.400 4702.720 ;
        RECT 3492.740 4702.440 3493.020 4702.720 ;
        RECT 3493.360 4702.440 3493.640 4702.720 ;
        RECT 3493.980 4702.440 3494.260 4702.720 ;
        RECT 3490.260 4701.820 3490.540 4702.100 ;
        RECT 3490.880 4701.820 3491.160 4702.100 ;
        RECT 3491.500 4701.820 3491.780 4702.100 ;
        RECT 3492.120 4701.820 3492.400 4702.100 ;
        RECT 3492.740 4701.820 3493.020 4702.100 ;
        RECT 3493.360 4701.820 3493.640 4702.100 ;
        RECT 3493.980 4701.820 3494.260 4702.100 ;
        RECT 3490.260 4701.200 3490.540 4701.480 ;
        RECT 3490.880 4701.200 3491.160 4701.480 ;
        RECT 3491.500 4701.200 3491.780 4701.480 ;
        RECT 3492.120 4701.200 3492.400 4701.480 ;
        RECT 3492.740 4701.200 3493.020 4701.480 ;
        RECT 3493.360 4701.200 3493.640 4701.480 ;
        RECT 3493.980 4701.200 3494.260 4701.480 ;
        RECT 3490.260 4700.580 3490.540 4700.860 ;
        RECT 3490.880 4700.580 3491.160 4700.860 ;
        RECT 3491.500 4700.580 3491.780 4700.860 ;
        RECT 3492.120 4700.580 3492.400 4700.860 ;
        RECT 3492.740 4700.580 3493.020 4700.860 ;
        RECT 3493.360 4700.580 3493.640 4700.860 ;
        RECT 3493.980 4700.580 3494.260 4700.860 ;
        RECT 3490.260 4699.960 3490.540 4700.240 ;
        RECT 3490.880 4699.960 3491.160 4700.240 ;
        RECT 3491.500 4699.960 3491.780 4700.240 ;
        RECT 3492.120 4699.960 3492.400 4700.240 ;
        RECT 3492.740 4699.960 3493.020 4700.240 ;
        RECT 3493.360 4699.960 3493.640 4700.240 ;
        RECT 3493.980 4699.960 3494.260 4700.240 ;
        RECT 395.965 4648.090 396.245 4648.370 ;
        RECT 396.585 4648.090 396.865 4648.370 ;
        RECT 397.205 4648.090 397.485 4648.370 ;
        RECT 397.825 4648.090 398.105 4648.370 ;
        RECT 398.445 4648.090 398.725 4648.370 ;
        RECT 399.065 4648.090 399.345 4648.370 ;
        RECT 399.685 4648.090 399.965 4648.370 ;
        RECT 395.965 4647.470 396.245 4647.750 ;
        RECT 396.585 4647.470 396.865 4647.750 ;
        RECT 397.205 4647.470 397.485 4647.750 ;
        RECT 397.825 4647.470 398.105 4647.750 ;
        RECT 398.445 4647.470 398.725 4647.750 ;
        RECT 399.065 4647.470 399.345 4647.750 ;
        RECT 399.685 4647.470 399.965 4647.750 ;
        RECT 395.965 4613.090 396.245 4613.370 ;
        RECT 396.585 4613.090 396.865 4613.370 ;
        RECT 397.205 4613.090 397.485 4613.370 ;
        RECT 397.825 4613.090 398.105 4613.370 ;
        RECT 398.445 4613.090 398.725 4613.370 ;
        RECT 399.065 4613.090 399.345 4613.370 ;
        RECT 399.685 4613.090 399.965 4613.370 ;
        RECT 395.965 4612.470 396.245 4612.750 ;
        RECT 396.585 4612.470 396.865 4612.750 ;
        RECT 397.205 4612.470 397.485 4612.750 ;
        RECT 397.825 4612.470 398.105 4612.750 ;
        RECT 398.445 4612.470 398.725 4612.750 ;
        RECT 399.065 4612.470 399.345 4612.750 ;
        RECT 399.685 4612.470 399.965 4612.750 ;
        RECT 395.965 4578.090 396.245 4578.370 ;
        RECT 396.585 4578.090 396.865 4578.370 ;
        RECT 397.205 4578.090 397.485 4578.370 ;
        RECT 397.825 4578.090 398.105 4578.370 ;
        RECT 398.445 4578.090 398.725 4578.370 ;
        RECT 399.065 4578.090 399.345 4578.370 ;
        RECT 399.685 4578.090 399.965 4578.370 ;
        RECT 395.965 4577.470 396.245 4577.750 ;
        RECT 396.585 4577.470 396.865 4577.750 ;
        RECT 397.205 4577.470 397.485 4577.750 ;
        RECT 397.825 4577.470 398.105 4577.750 ;
        RECT 398.445 4577.470 398.725 4577.750 ;
        RECT 399.065 4577.470 399.345 4577.750 ;
        RECT 399.685 4577.470 399.965 4577.750 ;
        RECT 395.740 4482.670 396.020 4482.950 ;
        RECT 396.360 4482.670 396.640 4482.950 ;
        RECT 396.980 4482.670 397.260 4482.950 ;
        RECT 397.600 4482.670 397.880 4482.950 ;
        RECT 398.220 4482.670 398.500 4482.950 ;
        RECT 398.840 4482.670 399.120 4482.950 ;
        RECT 399.460 4482.670 399.740 4482.950 ;
        RECT 395.740 4482.050 396.020 4482.330 ;
        RECT 396.360 4482.050 396.640 4482.330 ;
        RECT 396.980 4482.050 397.260 4482.330 ;
        RECT 397.600 4482.050 397.880 4482.330 ;
        RECT 398.220 4482.050 398.500 4482.330 ;
        RECT 398.840 4482.050 399.120 4482.330 ;
        RECT 399.460 4482.050 399.740 4482.330 ;
        RECT 395.740 4481.430 396.020 4481.710 ;
        RECT 396.360 4481.430 396.640 4481.710 ;
        RECT 396.980 4481.430 397.260 4481.710 ;
        RECT 397.600 4481.430 397.880 4481.710 ;
        RECT 398.220 4481.430 398.500 4481.710 ;
        RECT 398.840 4481.430 399.120 4481.710 ;
        RECT 399.460 4481.430 399.740 4481.710 ;
        RECT 395.740 4480.810 396.020 4481.090 ;
        RECT 396.360 4480.810 396.640 4481.090 ;
        RECT 396.980 4480.810 397.260 4481.090 ;
        RECT 397.600 4480.810 397.880 4481.090 ;
        RECT 398.220 4480.810 398.500 4481.090 ;
        RECT 398.840 4480.810 399.120 4481.090 ;
        RECT 399.460 4480.810 399.740 4481.090 ;
        RECT 395.740 4480.190 396.020 4480.470 ;
        RECT 396.360 4480.190 396.640 4480.470 ;
        RECT 396.980 4480.190 397.260 4480.470 ;
        RECT 397.600 4480.190 397.880 4480.470 ;
        RECT 398.220 4480.190 398.500 4480.470 ;
        RECT 398.840 4480.190 399.120 4480.470 ;
        RECT 399.460 4480.190 399.740 4480.470 ;
        RECT 395.740 4302.670 396.020 4302.950 ;
        RECT 396.360 4302.670 396.640 4302.950 ;
        RECT 396.980 4302.670 397.260 4302.950 ;
        RECT 397.600 4302.670 397.880 4302.950 ;
        RECT 398.220 4302.670 398.500 4302.950 ;
        RECT 398.840 4302.670 399.120 4302.950 ;
        RECT 399.460 4302.670 399.740 4302.950 ;
        RECT 395.740 4302.050 396.020 4302.330 ;
        RECT 396.360 4302.050 396.640 4302.330 ;
        RECT 396.980 4302.050 397.260 4302.330 ;
        RECT 397.600 4302.050 397.880 4302.330 ;
        RECT 398.220 4302.050 398.500 4302.330 ;
        RECT 398.840 4302.050 399.120 4302.330 ;
        RECT 399.460 4302.050 399.740 4302.330 ;
        RECT 395.740 4301.430 396.020 4301.710 ;
        RECT 396.360 4301.430 396.640 4301.710 ;
        RECT 396.980 4301.430 397.260 4301.710 ;
        RECT 397.600 4301.430 397.880 4301.710 ;
        RECT 398.220 4301.430 398.500 4301.710 ;
        RECT 398.840 4301.430 399.120 4301.710 ;
        RECT 399.460 4301.430 399.740 4301.710 ;
        RECT 395.740 4300.810 396.020 4301.090 ;
        RECT 396.360 4300.810 396.640 4301.090 ;
        RECT 396.980 4300.810 397.260 4301.090 ;
        RECT 397.600 4300.810 397.880 4301.090 ;
        RECT 398.220 4300.810 398.500 4301.090 ;
        RECT 398.840 4300.810 399.120 4301.090 ;
        RECT 399.460 4300.810 399.740 4301.090 ;
        RECT 395.740 4300.190 396.020 4300.470 ;
        RECT 396.360 4300.190 396.640 4300.470 ;
        RECT 396.980 4300.190 397.260 4300.470 ;
        RECT 397.600 4300.190 397.880 4300.470 ;
        RECT 398.220 4300.190 398.500 4300.470 ;
        RECT 398.840 4300.190 399.120 4300.470 ;
        RECT 399.460 4300.190 399.740 4300.470 ;
        RECT 395.740 4122.670 396.020 4122.950 ;
        RECT 396.360 4122.670 396.640 4122.950 ;
        RECT 396.980 4122.670 397.260 4122.950 ;
        RECT 397.600 4122.670 397.880 4122.950 ;
        RECT 398.220 4122.670 398.500 4122.950 ;
        RECT 398.840 4122.670 399.120 4122.950 ;
        RECT 399.460 4122.670 399.740 4122.950 ;
        RECT 395.740 4122.050 396.020 4122.330 ;
        RECT 396.360 4122.050 396.640 4122.330 ;
        RECT 396.980 4122.050 397.260 4122.330 ;
        RECT 397.600 4122.050 397.880 4122.330 ;
        RECT 398.220 4122.050 398.500 4122.330 ;
        RECT 398.840 4122.050 399.120 4122.330 ;
        RECT 399.460 4122.050 399.740 4122.330 ;
        RECT 395.740 4121.430 396.020 4121.710 ;
        RECT 396.360 4121.430 396.640 4121.710 ;
        RECT 396.980 4121.430 397.260 4121.710 ;
        RECT 397.600 4121.430 397.880 4121.710 ;
        RECT 398.220 4121.430 398.500 4121.710 ;
        RECT 398.840 4121.430 399.120 4121.710 ;
        RECT 399.460 4121.430 399.740 4121.710 ;
        RECT 395.740 4120.810 396.020 4121.090 ;
        RECT 396.360 4120.810 396.640 4121.090 ;
        RECT 396.980 4120.810 397.260 4121.090 ;
        RECT 397.600 4120.810 397.880 4121.090 ;
        RECT 398.220 4120.810 398.500 4121.090 ;
        RECT 398.840 4120.810 399.120 4121.090 ;
        RECT 399.460 4120.810 399.740 4121.090 ;
        RECT 395.740 4120.190 396.020 4120.470 ;
        RECT 396.360 4120.190 396.640 4120.470 ;
        RECT 396.980 4120.190 397.260 4120.470 ;
        RECT 397.600 4120.190 397.880 4120.470 ;
        RECT 398.220 4120.190 398.500 4120.470 ;
        RECT 398.840 4120.190 399.120 4120.470 ;
        RECT 399.460 4120.190 399.740 4120.470 ;
        RECT 396.040 4013.070 396.320 4013.350 ;
        RECT 396.660 4013.070 396.940 4013.350 ;
        RECT 397.280 4013.070 397.560 4013.350 ;
        RECT 397.900 4013.070 398.180 4013.350 ;
        RECT 398.520 4013.070 398.800 4013.350 ;
        RECT 399.140 4013.070 399.420 4013.350 ;
        RECT 399.760 4013.070 400.040 4013.350 ;
        RECT 396.040 4012.450 396.320 4012.730 ;
        RECT 396.660 4012.450 396.940 4012.730 ;
        RECT 397.280 4012.450 397.560 4012.730 ;
        RECT 397.900 4012.450 398.180 4012.730 ;
        RECT 398.520 4012.450 398.800 4012.730 ;
        RECT 399.140 4012.450 399.420 4012.730 ;
        RECT 399.760 4012.450 400.040 4012.730 ;
        RECT 396.040 4011.830 396.320 4012.110 ;
        RECT 396.660 4011.830 396.940 4012.110 ;
        RECT 397.280 4011.830 397.560 4012.110 ;
        RECT 397.900 4011.830 398.180 4012.110 ;
        RECT 398.520 4011.830 398.800 4012.110 ;
        RECT 399.140 4011.830 399.420 4012.110 ;
        RECT 399.760 4011.830 400.040 4012.110 ;
        RECT 396.040 4011.210 396.320 4011.490 ;
        RECT 396.660 4011.210 396.940 4011.490 ;
        RECT 397.280 4011.210 397.560 4011.490 ;
        RECT 397.900 4011.210 398.180 4011.490 ;
        RECT 398.520 4011.210 398.800 4011.490 ;
        RECT 399.140 4011.210 399.420 4011.490 ;
        RECT 399.760 4011.210 400.040 4011.490 ;
        RECT 396.040 4010.590 396.320 4010.870 ;
        RECT 396.660 4010.590 396.940 4010.870 ;
        RECT 397.280 4010.590 397.560 4010.870 ;
        RECT 397.900 4010.590 398.180 4010.870 ;
        RECT 398.520 4010.590 398.800 4010.870 ;
        RECT 399.140 4010.590 399.420 4010.870 ;
        RECT 399.760 4010.590 400.040 4010.870 ;
        RECT 396.040 4009.970 396.320 4010.250 ;
        RECT 396.660 4009.970 396.940 4010.250 ;
        RECT 397.280 4009.970 397.560 4010.250 ;
        RECT 397.900 4009.970 398.180 4010.250 ;
        RECT 398.520 4009.970 398.800 4010.250 ;
        RECT 399.140 4009.970 399.420 4010.250 ;
        RECT 399.760 4009.970 400.040 4010.250 ;
        RECT 396.040 4009.350 396.320 4009.630 ;
        RECT 396.660 4009.350 396.940 4009.630 ;
        RECT 397.280 4009.350 397.560 4009.630 ;
        RECT 397.900 4009.350 398.180 4009.630 ;
        RECT 398.520 4009.350 398.800 4009.630 ;
        RECT 399.140 4009.350 399.420 4009.630 ;
        RECT 399.760 4009.350 400.040 4009.630 ;
        RECT 396.040 4008.730 396.320 4009.010 ;
        RECT 396.660 4008.730 396.940 4009.010 ;
        RECT 397.280 4008.730 397.560 4009.010 ;
        RECT 397.900 4008.730 398.180 4009.010 ;
        RECT 398.520 4008.730 398.800 4009.010 ;
        RECT 399.140 4008.730 399.420 4009.010 ;
        RECT 399.760 4008.730 400.040 4009.010 ;
        RECT 396.040 4008.110 396.320 4008.390 ;
        RECT 396.660 4008.110 396.940 4008.390 ;
        RECT 397.280 4008.110 397.560 4008.390 ;
        RECT 397.900 4008.110 398.180 4008.390 ;
        RECT 398.520 4008.110 398.800 4008.390 ;
        RECT 399.140 4008.110 399.420 4008.390 ;
        RECT 399.760 4008.110 400.040 4008.390 ;
        RECT 396.040 4007.490 396.320 4007.770 ;
        RECT 396.660 4007.490 396.940 4007.770 ;
        RECT 397.280 4007.490 397.560 4007.770 ;
        RECT 397.900 4007.490 398.180 4007.770 ;
        RECT 398.520 4007.490 398.800 4007.770 ;
        RECT 399.140 4007.490 399.420 4007.770 ;
        RECT 399.760 4007.490 400.040 4007.770 ;
        RECT 396.040 4006.870 396.320 4007.150 ;
        RECT 396.660 4006.870 396.940 4007.150 ;
        RECT 397.280 4006.870 397.560 4007.150 ;
        RECT 397.900 4006.870 398.180 4007.150 ;
        RECT 398.520 4006.870 398.800 4007.150 ;
        RECT 399.140 4006.870 399.420 4007.150 ;
        RECT 399.760 4006.870 400.040 4007.150 ;
        RECT 396.040 4006.250 396.320 4006.530 ;
        RECT 396.660 4006.250 396.940 4006.530 ;
        RECT 397.280 4006.250 397.560 4006.530 ;
        RECT 397.900 4006.250 398.180 4006.530 ;
        RECT 398.520 4006.250 398.800 4006.530 ;
        RECT 399.140 4006.250 399.420 4006.530 ;
        RECT 399.760 4006.250 400.040 4006.530 ;
        RECT 396.040 4005.630 396.320 4005.910 ;
        RECT 396.660 4005.630 396.940 4005.910 ;
        RECT 397.280 4005.630 397.560 4005.910 ;
        RECT 397.900 4005.630 398.180 4005.910 ;
        RECT 398.520 4005.630 398.800 4005.910 ;
        RECT 399.140 4005.630 399.420 4005.910 ;
        RECT 399.760 4005.630 400.040 4005.910 ;
        RECT 396.040 4005.010 396.320 4005.290 ;
        RECT 396.660 4005.010 396.940 4005.290 ;
        RECT 397.280 4005.010 397.560 4005.290 ;
        RECT 397.900 4005.010 398.180 4005.290 ;
        RECT 398.520 4005.010 398.800 4005.290 ;
        RECT 399.140 4005.010 399.420 4005.290 ;
        RECT 399.760 4005.010 400.040 4005.290 ;
        RECT 396.040 4004.390 396.320 4004.670 ;
        RECT 396.660 4004.390 396.940 4004.670 ;
        RECT 397.280 4004.390 397.560 4004.670 ;
        RECT 397.900 4004.390 398.180 4004.670 ;
        RECT 398.520 4004.390 398.800 4004.670 ;
        RECT 399.140 4004.390 399.420 4004.670 ;
        RECT 399.760 4004.390 400.040 4004.670 ;
        RECT 396.040 4000.670 396.320 4000.950 ;
        RECT 396.660 4000.670 396.940 4000.950 ;
        RECT 397.280 4000.670 397.560 4000.950 ;
        RECT 397.900 4000.670 398.180 4000.950 ;
        RECT 398.520 4000.670 398.800 4000.950 ;
        RECT 399.140 4000.670 399.420 4000.950 ;
        RECT 399.760 4000.670 400.040 4000.950 ;
        RECT 396.040 4000.050 396.320 4000.330 ;
        RECT 396.660 4000.050 396.940 4000.330 ;
        RECT 397.280 4000.050 397.560 4000.330 ;
        RECT 397.900 4000.050 398.180 4000.330 ;
        RECT 398.520 4000.050 398.800 4000.330 ;
        RECT 399.140 4000.050 399.420 4000.330 ;
        RECT 399.760 4000.050 400.040 4000.330 ;
        RECT 396.040 3999.430 396.320 3999.710 ;
        RECT 396.660 3999.430 396.940 3999.710 ;
        RECT 397.280 3999.430 397.560 3999.710 ;
        RECT 397.900 3999.430 398.180 3999.710 ;
        RECT 398.520 3999.430 398.800 3999.710 ;
        RECT 399.140 3999.430 399.420 3999.710 ;
        RECT 399.760 3999.430 400.040 3999.710 ;
        RECT 396.040 3998.810 396.320 3999.090 ;
        RECT 396.660 3998.810 396.940 3999.090 ;
        RECT 397.280 3998.810 397.560 3999.090 ;
        RECT 397.900 3998.810 398.180 3999.090 ;
        RECT 398.520 3998.810 398.800 3999.090 ;
        RECT 399.140 3998.810 399.420 3999.090 ;
        RECT 399.760 3998.810 400.040 3999.090 ;
        RECT 396.040 3998.190 396.320 3998.470 ;
        RECT 396.660 3998.190 396.940 3998.470 ;
        RECT 397.280 3998.190 397.560 3998.470 ;
        RECT 397.900 3998.190 398.180 3998.470 ;
        RECT 398.520 3998.190 398.800 3998.470 ;
        RECT 399.140 3998.190 399.420 3998.470 ;
        RECT 399.760 3998.190 400.040 3998.470 ;
        RECT 396.040 3997.570 396.320 3997.850 ;
        RECT 396.660 3997.570 396.940 3997.850 ;
        RECT 397.280 3997.570 397.560 3997.850 ;
        RECT 397.900 3997.570 398.180 3997.850 ;
        RECT 398.520 3997.570 398.800 3997.850 ;
        RECT 399.140 3997.570 399.420 3997.850 ;
        RECT 399.760 3997.570 400.040 3997.850 ;
        RECT 396.040 3996.950 396.320 3997.230 ;
        RECT 396.660 3996.950 396.940 3997.230 ;
        RECT 397.280 3996.950 397.560 3997.230 ;
        RECT 397.900 3996.950 398.180 3997.230 ;
        RECT 398.520 3996.950 398.800 3997.230 ;
        RECT 399.140 3996.950 399.420 3997.230 ;
        RECT 399.760 3996.950 400.040 3997.230 ;
        RECT 396.040 3996.330 396.320 3996.610 ;
        RECT 396.660 3996.330 396.940 3996.610 ;
        RECT 397.280 3996.330 397.560 3996.610 ;
        RECT 397.900 3996.330 398.180 3996.610 ;
        RECT 398.520 3996.330 398.800 3996.610 ;
        RECT 399.140 3996.330 399.420 3996.610 ;
        RECT 399.760 3996.330 400.040 3996.610 ;
        RECT 396.040 3995.710 396.320 3995.990 ;
        RECT 396.660 3995.710 396.940 3995.990 ;
        RECT 397.280 3995.710 397.560 3995.990 ;
        RECT 397.900 3995.710 398.180 3995.990 ;
        RECT 398.520 3995.710 398.800 3995.990 ;
        RECT 399.140 3995.710 399.420 3995.990 ;
        RECT 399.760 3995.710 400.040 3995.990 ;
        RECT 396.040 3995.090 396.320 3995.370 ;
        RECT 396.660 3995.090 396.940 3995.370 ;
        RECT 397.280 3995.090 397.560 3995.370 ;
        RECT 397.900 3995.090 398.180 3995.370 ;
        RECT 398.520 3995.090 398.800 3995.370 ;
        RECT 399.140 3995.090 399.420 3995.370 ;
        RECT 399.760 3995.090 400.040 3995.370 ;
        RECT 396.040 3994.470 396.320 3994.750 ;
        RECT 396.660 3994.470 396.940 3994.750 ;
        RECT 397.280 3994.470 397.560 3994.750 ;
        RECT 397.900 3994.470 398.180 3994.750 ;
        RECT 398.520 3994.470 398.800 3994.750 ;
        RECT 399.140 3994.470 399.420 3994.750 ;
        RECT 399.760 3994.470 400.040 3994.750 ;
        RECT 396.040 3993.850 396.320 3994.130 ;
        RECT 396.660 3993.850 396.940 3994.130 ;
        RECT 397.280 3993.850 397.560 3994.130 ;
        RECT 397.900 3993.850 398.180 3994.130 ;
        RECT 398.520 3993.850 398.800 3994.130 ;
        RECT 399.140 3993.850 399.420 3994.130 ;
        RECT 399.760 3993.850 400.040 3994.130 ;
        RECT 396.040 3993.230 396.320 3993.510 ;
        RECT 396.660 3993.230 396.940 3993.510 ;
        RECT 397.280 3993.230 397.560 3993.510 ;
        RECT 397.900 3993.230 398.180 3993.510 ;
        RECT 398.520 3993.230 398.800 3993.510 ;
        RECT 399.140 3993.230 399.420 3993.510 ;
        RECT 399.760 3993.230 400.040 3993.510 ;
        RECT 396.040 3992.610 396.320 3992.890 ;
        RECT 396.660 3992.610 396.940 3992.890 ;
        RECT 397.280 3992.610 397.560 3992.890 ;
        RECT 397.900 3992.610 398.180 3992.890 ;
        RECT 398.520 3992.610 398.800 3992.890 ;
        RECT 399.140 3992.610 399.420 3992.890 ;
        RECT 399.760 3992.610 400.040 3992.890 ;
        RECT 396.040 3991.990 396.320 3992.270 ;
        RECT 396.660 3991.990 396.940 3992.270 ;
        RECT 397.280 3991.990 397.560 3992.270 ;
        RECT 397.900 3991.990 398.180 3992.270 ;
        RECT 398.520 3991.990 398.800 3992.270 ;
        RECT 399.140 3991.990 399.420 3992.270 ;
        RECT 399.760 3991.990 400.040 3992.270 ;
        RECT 396.040 3991.370 396.320 3991.650 ;
        RECT 396.660 3991.370 396.940 3991.650 ;
        RECT 397.280 3991.370 397.560 3991.650 ;
        RECT 397.900 3991.370 398.180 3991.650 ;
        RECT 398.520 3991.370 398.800 3991.650 ;
        RECT 399.140 3991.370 399.420 3991.650 ;
        RECT 399.760 3991.370 400.040 3991.650 ;
        RECT 396.040 3988.820 396.320 3989.100 ;
        RECT 396.660 3988.820 396.940 3989.100 ;
        RECT 397.280 3988.820 397.560 3989.100 ;
        RECT 397.900 3988.820 398.180 3989.100 ;
        RECT 398.520 3988.820 398.800 3989.100 ;
        RECT 399.140 3988.820 399.420 3989.100 ;
        RECT 399.760 3988.820 400.040 3989.100 ;
        RECT 396.040 3988.200 396.320 3988.480 ;
        RECT 396.660 3988.200 396.940 3988.480 ;
        RECT 397.280 3988.200 397.560 3988.480 ;
        RECT 397.900 3988.200 398.180 3988.480 ;
        RECT 398.520 3988.200 398.800 3988.480 ;
        RECT 399.140 3988.200 399.420 3988.480 ;
        RECT 399.760 3988.200 400.040 3988.480 ;
        RECT 396.040 3987.580 396.320 3987.860 ;
        RECT 396.660 3987.580 396.940 3987.860 ;
        RECT 397.280 3987.580 397.560 3987.860 ;
        RECT 397.900 3987.580 398.180 3987.860 ;
        RECT 398.520 3987.580 398.800 3987.860 ;
        RECT 399.140 3987.580 399.420 3987.860 ;
        RECT 399.760 3987.580 400.040 3987.860 ;
        RECT 396.040 3986.960 396.320 3987.240 ;
        RECT 396.660 3986.960 396.940 3987.240 ;
        RECT 397.280 3986.960 397.560 3987.240 ;
        RECT 397.900 3986.960 398.180 3987.240 ;
        RECT 398.520 3986.960 398.800 3987.240 ;
        RECT 399.140 3986.960 399.420 3987.240 ;
        RECT 399.760 3986.960 400.040 3987.240 ;
        RECT 396.040 3986.340 396.320 3986.620 ;
        RECT 396.660 3986.340 396.940 3986.620 ;
        RECT 397.280 3986.340 397.560 3986.620 ;
        RECT 397.900 3986.340 398.180 3986.620 ;
        RECT 398.520 3986.340 398.800 3986.620 ;
        RECT 399.140 3986.340 399.420 3986.620 ;
        RECT 399.760 3986.340 400.040 3986.620 ;
        RECT 396.040 3985.720 396.320 3986.000 ;
        RECT 396.660 3985.720 396.940 3986.000 ;
        RECT 397.280 3985.720 397.560 3986.000 ;
        RECT 397.900 3985.720 398.180 3986.000 ;
        RECT 398.520 3985.720 398.800 3986.000 ;
        RECT 399.140 3985.720 399.420 3986.000 ;
        RECT 399.760 3985.720 400.040 3986.000 ;
        RECT 396.040 3985.100 396.320 3985.380 ;
        RECT 396.660 3985.100 396.940 3985.380 ;
        RECT 397.280 3985.100 397.560 3985.380 ;
        RECT 397.900 3985.100 398.180 3985.380 ;
        RECT 398.520 3985.100 398.800 3985.380 ;
        RECT 399.140 3985.100 399.420 3985.380 ;
        RECT 399.760 3985.100 400.040 3985.380 ;
        RECT 396.040 3984.480 396.320 3984.760 ;
        RECT 396.660 3984.480 396.940 3984.760 ;
        RECT 397.280 3984.480 397.560 3984.760 ;
        RECT 397.900 3984.480 398.180 3984.760 ;
        RECT 398.520 3984.480 398.800 3984.760 ;
        RECT 399.140 3984.480 399.420 3984.760 ;
        RECT 399.760 3984.480 400.040 3984.760 ;
        RECT 396.040 3983.860 396.320 3984.140 ;
        RECT 396.660 3983.860 396.940 3984.140 ;
        RECT 397.280 3983.860 397.560 3984.140 ;
        RECT 397.900 3983.860 398.180 3984.140 ;
        RECT 398.520 3983.860 398.800 3984.140 ;
        RECT 399.140 3983.860 399.420 3984.140 ;
        RECT 399.760 3983.860 400.040 3984.140 ;
        RECT 396.040 3983.240 396.320 3983.520 ;
        RECT 396.660 3983.240 396.940 3983.520 ;
        RECT 397.280 3983.240 397.560 3983.520 ;
        RECT 397.900 3983.240 398.180 3983.520 ;
        RECT 398.520 3983.240 398.800 3983.520 ;
        RECT 399.140 3983.240 399.420 3983.520 ;
        RECT 399.760 3983.240 400.040 3983.520 ;
        RECT 396.040 3982.620 396.320 3982.900 ;
        RECT 396.660 3982.620 396.940 3982.900 ;
        RECT 397.280 3982.620 397.560 3982.900 ;
        RECT 397.900 3982.620 398.180 3982.900 ;
        RECT 398.520 3982.620 398.800 3982.900 ;
        RECT 399.140 3982.620 399.420 3982.900 ;
        RECT 399.760 3982.620 400.040 3982.900 ;
        RECT 396.040 3982.000 396.320 3982.280 ;
        RECT 396.660 3982.000 396.940 3982.280 ;
        RECT 397.280 3982.000 397.560 3982.280 ;
        RECT 397.900 3982.000 398.180 3982.280 ;
        RECT 398.520 3982.000 398.800 3982.280 ;
        RECT 399.140 3982.000 399.420 3982.280 ;
        RECT 399.760 3982.000 400.040 3982.280 ;
        RECT 396.040 3981.380 396.320 3981.660 ;
        RECT 396.660 3981.380 396.940 3981.660 ;
        RECT 397.280 3981.380 397.560 3981.660 ;
        RECT 397.900 3981.380 398.180 3981.660 ;
        RECT 398.520 3981.380 398.800 3981.660 ;
        RECT 399.140 3981.380 399.420 3981.660 ;
        RECT 399.760 3981.380 400.040 3981.660 ;
        RECT 396.040 3980.760 396.320 3981.040 ;
        RECT 396.660 3980.760 396.940 3981.040 ;
        RECT 397.280 3980.760 397.560 3981.040 ;
        RECT 397.900 3980.760 398.180 3981.040 ;
        RECT 398.520 3980.760 398.800 3981.040 ;
        RECT 399.140 3980.760 399.420 3981.040 ;
        RECT 399.760 3980.760 400.040 3981.040 ;
        RECT 396.040 3980.140 396.320 3980.420 ;
        RECT 396.660 3980.140 396.940 3980.420 ;
        RECT 397.280 3980.140 397.560 3980.420 ;
        RECT 397.900 3980.140 398.180 3980.420 ;
        RECT 398.520 3980.140 398.800 3980.420 ;
        RECT 399.140 3980.140 399.420 3980.420 ;
        RECT 399.760 3980.140 400.040 3980.420 ;
        RECT 396.040 3979.520 396.320 3979.800 ;
        RECT 396.660 3979.520 396.940 3979.800 ;
        RECT 397.280 3979.520 397.560 3979.800 ;
        RECT 397.900 3979.520 398.180 3979.800 ;
        RECT 398.520 3979.520 398.800 3979.800 ;
        RECT 399.140 3979.520 399.420 3979.800 ;
        RECT 399.760 3979.520 400.040 3979.800 ;
        RECT 396.040 3975.290 396.320 3975.570 ;
        RECT 396.660 3975.290 396.940 3975.570 ;
        RECT 397.280 3975.290 397.560 3975.570 ;
        RECT 397.900 3975.290 398.180 3975.570 ;
        RECT 398.520 3975.290 398.800 3975.570 ;
        RECT 399.140 3975.290 399.420 3975.570 ;
        RECT 399.760 3975.290 400.040 3975.570 ;
        RECT 396.040 3974.670 396.320 3974.950 ;
        RECT 396.660 3974.670 396.940 3974.950 ;
        RECT 397.280 3974.670 397.560 3974.950 ;
        RECT 397.900 3974.670 398.180 3974.950 ;
        RECT 398.520 3974.670 398.800 3974.950 ;
        RECT 399.140 3974.670 399.420 3974.950 ;
        RECT 399.760 3974.670 400.040 3974.950 ;
        RECT 396.040 3974.050 396.320 3974.330 ;
        RECT 396.660 3974.050 396.940 3974.330 ;
        RECT 397.280 3974.050 397.560 3974.330 ;
        RECT 397.900 3974.050 398.180 3974.330 ;
        RECT 398.520 3974.050 398.800 3974.330 ;
        RECT 399.140 3974.050 399.420 3974.330 ;
        RECT 399.760 3974.050 400.040 3974.330 ;
        RECT 396.040 3973.430 396.320 3973.710 ;
        RECT 396.660 3973.430 396.940 3973.710 ;
        RECT 397.280 3973.430 397.560 3973.710 ;
        RECT 397.900 3973.430 398.180 3973.710 ;
        RECT 398.520 3973.430 398.800 3973.710 ;
        RECT 399.140 3973.430 399.420 3973.710 ;
        RECT 399.760 3973.430 400.040 3973.710 ;
        RECT 396.040 3972.810 396.320 3973.090 ;
        RECT 396.660 3972.810 396.940 3973.090 ;
        RECT 397.280 3972.810 397.560 3973.090 ;
        RECT 397.900 3972.810 398.180 3973.090 ;
        RECT 398.520 3972.810 398.800 3973.090 ;
        RECT 399.140 3972.810 399.420 3973.090 ;
        RECT 399.760 3972.810 400.040 3973.090 ;
        RECT 396.040 3972.190 396.320 3972.470 ;
        RECT 396.660 3972.190 396.940 3972.470 ;
        RECT 397.280 3972.190 397.560 3972.470 ;
        RECT 397.900 3972.190 398.180 3972.470 ;
        RECT 398.520 3972.190 398.800 3972.470 ;
        RECT 399.140 3972.190 399.420 3972.470 ;
        RECT 399.760 3972.190 400.040 3972.470 ;
        RECT 396.040 3971.570 396.320 3971.850 ;
        RECT 396.660 3971.570 396.940 3971.850 ;
        RECT 397.280 3971.570 397.560 3971.850 ;
        RECT 397.900 3971.570 398.180 3971.850 ;
        RECT 398.520 3971.570 398.800 3971.850 ;
        RECT 399.140 3971.570 399.420 3971.850 ;
        RECT 399.760 3971.570 400.040 3971.850 ;
        RECT 396.040 3970.950 396.320 3971.230 ;
        RECT 396.660 3970.950 396.940 3971.230 ;
        RECT 397.280 3970.950 397.560 3971.230 ;
        RECT 397.900 3970.950 398.180 3971.230 ;
        RECT 398.520 3970.950 398.800 3971.230 ;
        RECT 399.140 3970.950 399.420 3971.230 ;
        RECT 399.760 3970.950 400.040 3971.230 ;
        RECT 396.040 3970.330 396.320 3970.610 ;
        RECT 396.660 3970.330 396.940 3970.610 ;
        RECT 397.280 3970.330 397.560 3970.610 ;
        RECT 397.900 3970.330 398.180 3970.610 ;
        RECT 398.520 3970.330 398.800 3970.610 ;
        RECT 399.140 3970.330 399.420 3970.610 ;
        RECT 399.760 3970.330 400.040 3970.610 ;
        RECT 396.040 3969.710 396.320 3969.990 ;
        RECT 396.660 3969.710 396.940 3969.990 ;
        RECT 397.280 3969.710 397.560 3969.990 ;
        RECT 397.900 3969.710 398.180 3969.990 ;
        RECT 398.520 3969.710 398.800 3969.990 ;
        RECT 399.140 3969.710 399.420 3969.990 ;
        RECT 399.760 3969.710 400.040 3969.990 ;
        RECT 396.040 3969.090 396.320 3969.370 ;
        RECT 396.660 3969.090 396.940 3969.370 ;
        RECT 397.280 3969.090 397.560 3969.370 ;
        RECT 397.900 3969.090 398.180 3969.370 ;
        RECT 398.520 3969.090 398.800 3969.370 ;
        RECT 399.140 3969.090 399.420 3969.370 ;
        RECT 399.760 3969.090 400.040 3969.370 ;
        RECT 396.040 3968.470 396.320 3968.750 ;
        RECT 396.660 3968.470 396.940 3968.750 ;
        RECT 397.280 3968.470 397.560 3968.750 ;
        RECT 397.900 3968.470 398.180 3968.750 ;
        RECT 398.520 3968.470 398.800 3968.750 ;
        RECT 399.140 3968.470 399.420 3968.750 ;
        RECT 399.760 3968.470 400.040 3968.750 ;
        RECT 396.040 3967.850 396.320 3968.130 ;
        RECT 396.660 3967.850 396.940 3968.130 ;
        RECT 397.280 3967.850 397.560 3968.130 ;
        RECT 397.900 3967.850 398.180 3968.130 ;
        RECT 398.520 3967.850 398.800 3968.130 ;
        RECT 399.140 3967.850 399.420 3968.130 ;
        RECT 399.760 3967.850 400.040 3968.130 ;
        RECT 396.040 3967.230 396.320 3967.510 ;
        RECT 396.660 3967.230 396.940 3967.510 ;
        RECT 397.280 3967.230 397.560 3967.510 ;
        RECT 397.900 3967.230 398.180 3967.510 ;
        RECT 398.520 3967.230 398.800 3967.510 ;
        RECT 399.140 3967.230 399.420 3967.510 ;
        RECT 399.760 3967.230 400.040 3967.510 ;
        RECT 396.040 3966.610 396.320 3966.890 ;
        RECT 396.660 3966.610 396.940 3966.890 ;
        RECT 397.280 3966.610 397.560 3966.890 ;
        RECT 397.900 3966.610 398.180 3966.890 ;
        RECT 398.520 3966.610 398.800 3966.890 ;
        RECT 399.140 3966.610 399.420 3966.890 ;
        RECT 399.760 3966.610 400.040 3966.890 ;
        RECT 396.040 3965.990 396.320 3966.270 ;
        RECT 396.660 3965.990 396.940 3966.270 ;
        RECT 397.280 3965.990 397.560 3966.270 ;
        RECT 397.900 3965.990 398.180 3966.270 ;
        RECT 398.520 3965.990 398.800 3966.270 ;
        RECT 399.140 3965.990 399.420 3966.270 ;
        RECT 399.760 3965.990 400.040 3966.270 ;
        RECT 396.040 3963.440 396.320 3963.720 ;
        RECT 396.660 3963.440 396.940 3963.720 ;
        RECT 397.280 3963.440 397.560 3963.720 ;
        RECT 397.900 3963.440 398.180 3963.720 ;
        RECT 398.520 3963.440 398.800 3963.720 ;
        RECT 399.140 3963.440 399.420 3963.720 ;
        RECT 399.760 3963.440 400.040 3963.720 ;
        RECT 396.040 3962.820 396.320 3963.100 ;
        RECT 396.660 3962.820 396.940 3963.100 ;
        RECT 397.280 3962.820 397.560 3963.100 ;
        RECT 397.900 3962.820 398.180 3963.100 ;
        RECT 398.520 3962.820 398.800 3963.100 ;
        RECT 399.140 3962.820 399.420 3963.100 ;
        RECT 399.760 3962.820 400.040 3963.100 ;
        RECT 396.040 3962.200 396.320 3962.480 ;
        RECT 396.660 3962.200 396.940 3962.480 ;
        RECT 397.280 3962.200 397.560 3962.480 ;
        RECT 397.900 3962.200 398.180 3962.480 ;
        RECT 398.520 3962.200 398.800 3962.480 ;
        RECT 399.140 3962.200 399.420 3962.480 ;
        RECT 399.760 3962.200 400.040 3962.480 ;
        RECT 396.040 3961.580 396.320 3961.860 ;
        RECT 396.660 3961.580 396.940 3961.860 ;
        RECT 397.280 3961.580 397.560 3961.860 ;
        RECT 397.900 3961.580 398.180 3961.860 ;
        RECT 398.520 3961.580 398.800 3961.860 ;
        RECT 399.140 3961.580 399.420 3961.860 ;
        RECT 399.760 3961.580 400.040 3961.860 ;
        RECT 396.040 3960.960 396.320 3961.240 ;
        RECT 396.660 3960.960 396.940 3961.240 ;
        RECT 397.280 3960.960 397.560 3961.240 ;
        RECT 397.900 3960.960 398.180 3961.240 ;
        RECT 398.520 3960.960 398.800 3961.240 ;
        RECT 399.140 3960.960 399.420 3961.240 ;
        RECT 399.760 3960.960 400.040 3961.240 ;
        RECT 396.040 3960.340 396.320 3960.620 ;
        RECT 396.660 3960.340 396.940 3960.620 ;
        RECT 397.280 3960.340 397.560 3960.620 ;
        RECT 397.900 3960.340 398.180 3960.620 ;
        RECT 398.520 3960.340 398.800 3960.620 ;
        RECT 399.140 3960.340 399.420 3960.620 ;
        RECT 399.760 3960.340 400.040 3960.620 ;
        RECT 396.040 3959.720 396.320 3960.000 ;
        RECT 396.660 3959.720 396.940 3960.000 ;
        RECT 397.280 3959.720 397.560 3960.000 ;
        RECT 397.900 3959.720 398.180 3960.000 ;
        RECT 398.520 3959.720 398.800 3960.000 ;
        RECT 399.140 3959.720 399.420 3960.000 ;
        RECT 399.760 3959.720 400.040 3960.000 ;
        RECT 396.040 3959.100 396.320 3959.380 ;
        RECT 396.660 3959.100 396.940 3959.380 ;
        RECT 397.280 3959.100 397.560 3959.380 ;
        RECT 397.900 3959.100 398.180 3959.380 ;
        RECT 398.520 3959.100 398.800 3959.380 ;
        RECT 399.140 3959.100 399.420 3959.380 ;
        RECT 399.760 3959.100 400.040 3959.380 ;
        RECT 396.040 3958.480 396.320 3958.760 ;
        RECT 396.660 3958.480 396.940 3958.760 ;
        RECT 397.280 3958.480 397.560 3958.760 ;
        RECT 397.900 3958.480 398.180 3958.760 ;
        RECT 398.520 3958.480 398.800 3958.760 ;
        RECT 399.140 3958.480 399.420 3958.760 ;
        RECT 399.760 3958.480 400.040 3958.760 ;
        RECT 396.040 3957.860 396.320 3958.140 ;
        RECT 396.660 3957.860 396.940 3958.140 ;
        RECT 397.280 3957.860 397.560 3958.140 ;
        RECT 397.900 3957.860 398.180 3958.140 ;
        RECT 398.520 3957.860 398.800 3958.140 ;
        RECT 399.140 3957.860 399.420 3958.140 ;
        RECT 399.760 3957.860 400.040 3958.140 ;
        RECT 396.040 3957.240 396.320 3957.520 ;
        RECT 396.660 3957.240 396.940 3957.520 ;
        RECT 397.280 3957.240 397.560 3957.520 ;
        RECT 397.900 3957.240 398.180 3957.520 ;
        RECT 398.520 3957.240 398.800 3957.520 ;
        RECT 399.140 3957.240 399.420 3957.520 ;
        RECT 399.760 3957.240 400.040 3957.520 ;
        RECT 396.040 3956.620 396.320 3956.900 ;
        RECT 396.660 3956.620 396.940 3956.900 ;
        RECT 397.280 3956.620 397.560 3956.900 ;
        RECT 397.900 3956.620 398.180 3956.900 ;
        RECT 398.520 3956.620 398.800 3956.900 ;
        RECT 399.140 3956.620 399.420 3956.900 ;
        RECT 399.760 3956.620 400.040 3956.900 ;
        RECT 396.040 3956.000 396.320 3956.280 ;
        RECT 396.660 3956.000 396.940 3956.280 ;
        RECT 397.280 3956.000 397.560 3956.280 ;
        RECT 397.900 3956.000 398.180 3956.280 ;
        RECT 398.520 3956.000 398.800 3956.280 ;
        RECT 399.140 3956.000 399.420 3956.280 ;
        RECT 399.760 3956.000 400.040 3956.280 ;
        RECT 396.040 3955.380 396.320 3955.660 ;
        RECT 396.660 3955.380 396.940 3955.660 ;
        RECT 397.280 3955.380 397.560 3955.660 ;
        RECT 397.900 3955.380 398.180 3955.660 ;
        RECT 398.520 3955.380 398.800 3955.660 ;
        RECT 399.140 3955.380 399.420 3955.660 ;
        RECT 399.760 3955.380 400.040 3955.660 ;
        RECT 396.040 3954.760 396.320 3955.040 ;
        RECT 396.660 3954.760 396.940 3955.040 ;
        RECT 397.280 3954.760 397.560 3955.040 ;
        RECT 397.900 3954.760 398.180 3955.040 ;
        RECT 398.520 3954.760 398.800 3955.040 ;
        RECT 399.140 3954.760 399.420 3955.040 ;
        RECT 399.760 3954.760 400.040 3955.040 ;
        RECT 396.040 3954.140 396.320 3954.420 ;
        RECT 396.660 3954.140 396.940 3954.420 ;
        RECT 397.280 3954.140 397.560 3954.420 ;
        RECT 397.900 3954.140 398.180 3954.420 ;
        RECT 398.520 3954.140 398.800 3954.420 ;
        RECT 399.140 3954.140 399.420 3954.420 ;
        RECT 399.760 3954.140 400.040 3954.420 ;
        RECT 396.040 3950.420 396.320 3950.700 ;
        RECT 396.660 3950.420 396.940 3950.700 ;
        RECT 397.280 3950.420 397.560 3950.700 ;
        RECT 397.900 3950.420 398.180 3950.700 ;
        RECT 398.520 3950.420 398.800 3950.700 ;
        RECT 399.140 3950.420 399.420 3950.700 ;
        RECT 399.760 3950.420 400.040 3950.700 ;
        RECT 396.040 3949.800 396.320 3950.080 ;
        RECT 396.660 3949.800 396.940 3950.080 ;
        RECT 397.280 3949.800 397.560 3950.080 ;
        RECT 397.900 3949.800 398.180 3950.080 ;
        RECT 398.520 3949.800 398.800 3950.080 ;
        RECT 399.140 3949.800 399.420 3950.080 ;
        RECT 399.760 3949.800 400.040 3950.080 ;
        RECT 396.040 3949.180 396.320 3949.460 ;
        RECT 396.660 3949.180 396.940 3949.460 ;
        RECT 397.280 3949.180 397.560 3949.460 ;
        RECT 397.900 3949.180 398.180 3949.460 ;
        RECT 398.520 3949.180 398.800 3949.460 ;
        RECT 399.140 3949.180 399.420 3949.460 ;
        RECT 399.760 3949.180 400.040 3949.460 ;
        RECT 396.040 3948.560 396.320 3948.840 ;
        RECT 396.660 3948.560 396.940 3948.840 ;
        RECT 397.280 3948.560 397.560 3948.840 ;
        RECT 397.900 3948.560 398.180 3948.840 ;
        RECT 398.520 3948.560 398.800 3948.840 ;
        RECT 399.140 3948.560 399.420 3948.840 ;
        RECT 399.760 3948.560 400.040 3948.840 ;
        RECT 396.040 3947.940 396.320 3948.220 ;
        RECT 396.660 3947.940 396.940 3948.220 ;
        RECT 397.280 3947.940 397.560 3948.220 ;
        RECT 397.900 3947.940 398.180 3948.220 ;
        RECT 398.520 3947.940 398.800 3948.220 ;
        RECT 399.140 3947.940 399.420 3948.220 ;
        RECT 399.760 3947.940 400.040 3948.220 ;
        RECT 396.040 3947.320 396.320 3947.600 ;
        RECT 396.660 3947.320 396.940 3947.600 ;
        RECT 397.280 3947.320 397.560 3947.600 ;
        RECT 397.900 3947.320 398.180 3947.600 ;
        RECT 398.520 3947.320 398.800 3947.600 ;
        RECT 399.140 3947.320 399.420 3947.600 ;
        RECT 399.760 3947.320 400.040 3947.600 ;
        RECT 396.040 3946.700 396.320 3946.980 ;
        RECT 396.660 3946.700 396.940 3946.980 ;
        RECT 397.280 3946.700 397.560 3946.980 ;
        RECT 397.900 3946.700 398.180 3946.980 ;
        RECT 398.520 3946.700 398.800 3946.980 ;
        RECT 399.140 3946.700 399.420 3946.980 ;
        RECT 399.760 3946.700 400.040 3946.980 ;
        RECT 396.040 3946.080 396.320 3946.360 ;
        RECT 396.660 3946.080 396.940 3946.360 ;
        RECT 397.280 3946.080 397.560 3946.360 ;
        RECT 397.900 3946.080 398.180 3946.360 ;
        RECT 398.520 3946.080 398.800 3946.360 ;
        RECT 399.140 3946.080 399.420 3946.360 ;
        RECT 399.760 3946.080 400.040 3946.360 ;
        RECT 396.040 3945.460 396.320 3945.740 ;
        RECT 396.660 3945.460 396.940 3945.740 ;
        RECT 397.280 3945.460 397.560 3945.740 ;
        RECT 397.900 3945.460 398.180 3945.740 ;
        RECT 398.520 3945.460 398.800 3945.740 ;
        RECT 399.140 3945.460 399.420 3945.740 ;
        RECT 399.760 3945.460 400.040 3945.740 ;
        RECT 396.040 3944.840 396.320 3945.120 ;
        RECT 396.660 3944.840 396.940 3945.120 ;
        RECT 397.280 3944.840 397.560 3945.120 ;
        RECT 397.900 3944.840 398.180 3945.120 ;
        RECT 398.520 3944.840 398.800 3945.120 ;
        RECT 399.140 3944.840 399.420 3945.120 ;
        RECT 399.760 3944.840 400.040 3945.120 ;
        RECT 396.040 3944.220 396.320 3944.500 ;
        RECT 396.660 3944.220 396.940 3944.500 ;
        RECT 397.280 3944.220 397.560 3944.500 ;
        RECT 397.900 3944.220 398.180 3944.500 ;
        RECT 398.520 3944.220 398.800 3944.500 ;
        RECT 399.140 3944.220 399.420 3944.500 ;
        RECT 399.760 3944.220 400.040 3944.500 ;
        RECT 396.040 3943.600 396.320 3943.880 ;
        RECT 396.660 3943.600 396.940 3943.880 ;
        RECT 397.280 3943.600 397.560 3943.880 ;
        RECT 397.900 3943.600 398.180 3943.880 ;
        RECT 398.520 3943.600 398.800 3943.880 ;
        RECT 399.140 3943.600 399.420 3943.880 ;
        RECT 399.760 3943.600 400.040 3943.880 ;
        RECT 396.040 3942.980 396.320 3943.260 ;
        RECT 396.660 3942.980 396.940 3943.260 ;
        RECT 397.280 3942.980 397.560 3943.260 ;
        RECT 397.900 3942.980 398.180 3943.260 ;
        RECT 398.520 3942.980 398.800 3943.260 ;
        RECT 399.140 3942.980 399.420 3943.260 ;
        RECT 399.760 3942.980 400.040 3943.260 ;
        RECT 396.040 3942.360 396.320 3942.640 ;
        RECT 396.660 3942.360 396.940 3942.640 ;
        RECT 397.280 3942.360 397.560 3942.640 ;
        RECT 397.900 3942.360 398.180 3942.640 ;
        RECT 398.520 3942.360 398.800 3942.640 ;
        RECT 399.140 3942.360 399.420 3942.640 ;
        RECT 399.760 3942.360 400.040 3942.640 ;
        RECT 396.040 3941.740 396.320 3942.020 ;
        RECT 396.660 3941.740 396.940 3942.020 ;
        RECT 397.280 3941.740 397.560 3942.020 ;
        RECT 397.900 3941.740 398.180 3942.020 ;
        RECT 398.520 3941.740 398.800 3942.020 ;
        RECT 399.140 3941.740 399.420 3942.020 ;
        RECT 399.760 3941.740 400.040 3942.020 ;
        RECT 395.965 3909.920 396.245 3910.200 ;
        RECT 396.585 3909.920 396.865 3910.200 ;
        RECT 397.205 3909.920 397.485 3910.200 ;
        RECT 397.825 3909.920 398.105 3910.200 ;
        RECT 398.445 3909.920 398.725 3910.200 ;
        RECT 399.065 3909.920 399.345 3910.200 ;
        RECT 399.685 3909.920 399.965 3910.200 ;
        RECT 395.965 3828.090 396.245 3828.370 ;
        RECT 396.585 3828.090 396.865 3828.370 ;
        RECT 397.205 3828.090 397.485 3828.370 ;
        RECT 397.825 3828.090 398.105 3828.370 ;
        RECT 398.445 3828.090 398.725 3828.370 ;
        RECT 399.065 3828.090 399.345 3828.370 ;
        RECT 399.685 3828.090 399.965 3828.370 ;
        RECT 395.965 3827.470 396.245 3827.750 ;
        RECT 396.585 3827.470 396.865 3827.750 ;
        RECT 397.205 3827.470 397.485 3827.750 ;
        RECT 397.825 3827.470 398.105 3827.750 ;
        RECT 398.445 3827.470 398.725 3827.750 ;
        RECT 399.065 3827.470 399.345 3827.750 ;
        RECT 399.685 3827.470 399.965 3827.750 ;
        RECT 395.965 3793.090 396.245 3793.370 ;
        RECT 396.585 3793.090 396.865 3793.370 ;
        RECT 397.205 3793.090 397.485 3793.370 ;
        RECT 397.825 3793.090 398.105 3793.370 ;
        RECT 398.445 3793.090 398.725 3793.370 ;
        RECT 399.065 3793.090 399.345 3793.370 ;
        RECT 399.685 3793.090 399.965 3793.370 ;
        RECT 395.965 3792.470 396.245 3792.750 ;
        RECT 396.585 3792.470 396.865 3792.750 ;
        RECT 397.205 3792.470 397.485 3792.750 ;
        RECT 397.825 3792.470 398.105 3792.750 ;
        RECT 398.445 3792.470 398.725 3792.750 ;
        RECT 399.065 3792.470 399.345 3792.750 ;
        RECT 399.685 3792.470 399.965 3792.750 ;
        RECT 395.740 3762.670 396.020 3762.950 ;
        RECT 396.360 3762.670 396.640 3762.950 ;
        RECT 396.980 3762.670 397.260 3762.950 ;
        RECT 397.600 3762.670 397.880 3762.950 ;
        RECT 398.220 3762.670 398.500 3762.950 ;
        RECT 398.840 3762.670 399.120 3762.950 ;
        RECT 399.460 3762.670 399.740 3762.950 ;
        RECT 395.740 3762.050 396.020 3762.330 ;
        RECT 396.360 3762.050 396.640 3762.330 ;
        RECT 396.980 3762.050 397.260 3762.330 ;
        RECT 397.600 3762.050 397.880 3762.330 ;
        RECT 398.220 3762.050 398.500 3762.330 ;
        RECT 398.840 3762.050 399.120 3762.330 ;
        RECT 399.460 3762.050 399.740 3762.330 ;
        RECT 395.740 3761.430 396.020 3761.710 ;
        RECT 396.360 3761.430 396.640 3761.710 ;
        RECT 396.980 3761.430 397.260 3761.710 ;
        RECT 397.600 3761.430 397.880 3761.710 ;
        RECT 398.220 3761.430 398.500 3761.710 ;
        RECT 398.840 3761.430 399.120 3761.710 ;
        RECT 399.460 3761.430 399.740 3761.710 ;
        RECT 395.740 3760.810 396.020 3761.090 ;
        RECT 396.360 3760.810 396.640 3761.090 ;
        RECT 396.980 3760.810 397.260 3761.090 ;
        RECT 397.600 3760.810 397.880 3761.090 ;
        RECT 398.220 3760.810 398.500 3761.090 ;
        RECT 398.840 3760.810 399.120 3761.090 ;
        RECT 399.460 3760.810 399.740 3761.090 ;
        RECT 395.740 3760.190 396.020 3760.470 ;
        RECT 396.360 3760.190 396.640 3760.470 ;
        RECT 396.980 3760.190 397.260 3760.470 ;
        RECT 397.600 3760.190 397.880 3760.470 ;
        RECT 398.220 3760.190 398.500 3760.470 ;
        RECT 398.840 3760.190 399.120 3760.470 ;
        RECT 399.460 3760.190 399.740 3760.470 ;
        RECT 395.965 3758.090 396.245 3758.370 ;
        RECT 396.585 3758.090 396.865 3758.370 ;
        RECT 397.205 3758.090 397.485 3758.370 ;
        RECT 397.825 3758.090 398.105 3758.370 ;
        RECT 398.445 3758.090 398.725 3758.370 ;
        RECT 399.065 3758.090 399.345 3758.370 ;
        RECT 399.685 3758.090 399.965 3758.370 ;
        RECT 395.965 3757.470 396.245 3757.750 ;
        RECT 396.585 3757.470 396.865 3757.750 ;
        RECT 397.205 3757.470 397.485 3757.750 ;
        RECT 397.825 3757.470 398.105 3757.750 ;
        RECT 398.445 3757.470 398.725 3757.750 ;
        RECT 399.065 3757.470 399.345 3757.750 ;
        RECT 399.685 3757.470 399.965 3757.750 ;
        RECT 395.965 3704.920 396.245 3705.200 ;
        RECT 396.585 3704.920 396.865 3705.200 ;
        RECT 397.205 3704.920 397.485 3705.200 ;
        RECT 397.825 3704.920 398.105 3705.200 ;
        RECT 398.445 3704.920 398.725 3705.200 ;
        RECT 399.065 3704.920 399.345 3705.200 ;
        RECT 399.685 3704.920 399.965 3705.200 ;
        RECT 395.965 3623.090 396.245 3623.370 ;
        RECT 396.585 3623.090 396.865 3623.370 ;
        RECT 397.205 3623.090 397.485 3623.370 ;
        RECT 397.825 3623.090 398.105 3623.370 ;
        RECT 398.445 3623.090 398.725 3623.370 ;
        RECT 399.065 3623.090 399.345 3623.370 ;
        RECT 399.685 3623.090 399.965 3623.370 ;
        RECT 395.965 3622.470 396.245 3622.750 ;
        RECT 396.585 3622.470 396.865 3622.750 ;
        RECT 397.205 3622.470 397.485 3622.750 ;
        RECT 397.825 3622.470 398.105 3622.750 ;
        RECT 398.445 3622.470 398.725 3622.750 ;
        RECT 399.065 3622.470 399.345 3622.750 ;
        RECT 399.685 3622.470 399.965 3622.750 ;
        RECT 395.965 3588.090 396.245 3588.370 ;
        RECT 396.585 3588.090 396.865 3588.370 ;
        RECT 397.205 3588.090 397.485 3588.370 ;
        RECT 397.825 3588.090 398.105 3588.370 ;
        RECT 398.445 3588.090 398.725 3588.370 ;
        RECT 399.065 3588.090 399.345 3588.370 ;
        RECT 399.685 3588.090 399.965 3588.370 ;
        RECT 395.965 3587.470 396.245 3587.750 ;
        RECT 396.585 3587.470 396.865 3587.750 ;
        RECT 397.205 3587.470 397.485 3587.750 ;
        RECT 397.825 3587.470 398.105 3587.750 ;
        RECT 398.445 3587.470 398.725 3587.750 ;
        RECT 399.065 3587.470 399.345 3587.750 ;
        RECT 399.685 3587.470 399.965 3587.750 ;
        RECT 395.740 3582.670 396.020 3582.950 ;
        RECT 396.360 3582.670 396.640 3582.950 ;
        RECT 396.980 3582.670 397.260 3582.950 ;
        RECT 397.600 3582.670 397.880 3582.950 ;
        RECT 398.220 3582.670 398.500 3582.950 ;
        RECT 398.840 3582.670 399.120 3582.950 ;
        RECT 399.460 3582.670 399.740 3582.950 ;
        RECT 395.740 3582.050 396.020 3582.330 ;
        RECT 396.360 3582.050 396.640 3582.330 ;
        RECT 396.980 3582.050 397.260 3582.330 ;
        RECT 397.600 3582.050 397.880 3582.330 ;
        RECT 398.220 3582.050 398.500 3582.330 ;
        RECT 398.840 3582.050 399.120 3582.330 ;
        RECT 399.460 3582.050 399.740 3582.330 ;
        RECT 395.740 3581.430 396.020 3581.710 ;
        RECT 396.360 3581.430 396.640 3581.710 ;
        RECT 396.980 3581.430 397.260 3581.710 ;
        RECT 397.600 3581.430 397.880 3581.710 ;
        RECT 398.220 3581.430 398.500 3581.710 ;
        RECT 398.840 3581.430 399.120 3581.710 ;
        RECT 399.460 3581.430 399.740 3581.710 ;
        RECT 395.740 3580.810 396.020 3581.090 ;
        RECT 396.360 3580.810 396.640 3581.090 ;
        RECT 396.980 3580.810 397.260 3581.090 ;
        RECT 397.600 3580.810 397.880 3581.090 ;
        RECT 398.220 3580.810 398.500 3581.090 ;
        RECT 398.840 3580.810 399.120 3581.090 ;
        RECT 399.460 3580.810 399.740 3581.090 ;
        RECT 395.740 3580.190 396.020 3580.470 ;
        RECT 396.360 3580.190 396.640 3580.470 ;
        RECT 396.980 3580.190 397.260 3580.470 ;
        RECT 397.600 3580.190 397.880 3580.470 ;
        RECT 398.220 3580.190 398.500 3580.470 ;
        RECT 398.840 3580.190 399.120 3580.470 ;
        RECT 399.460 3580.190 399.740 3580.470 ;
        RECT 395.965 3553.090 396.245 3553.370 ;
        RECT 396.585 3553.090 396.865 3553.370 ;
        RECT 397.205 3553.090 397.485 3553.370 ;
        RECT 397.825 3553.090 398.105 3553.370 ;
        RECT 398.445 3553.090 398.725 3553.370 ;
        RECT 399.065 3553.090 399.345 3553.370 ;
        RECT 399.685 3553.090 399.965 3553.370 ;
        RECT 395.965 3552.470 396.245 3552.750 ;
        RECT 396.585 3552.470 396.865 3552.750 ;
        RECT 397.205 3552.470 397.485 3552.750 ;
        RECT 397.825 3552.470 398.105 3552.750 ;
        RECT 398.445 3552.470 398.725 3552.750 ;
        RECT 399.065 3552.470 399.345 3552.750 ;
        RECT 399.685 3552.470 399.965 3552.750 ;
        RECT 395.965 3499.920 396.245 3500.200 ;
        RECT 396.585 3499.920 396.865 3500.200 ;
        RECT 397.205 3499.920 397.485 3500.200 ;
        RECT 397.825 3499.920 398.105 3500.200 ;
        RECT 398.445 3499.920 398.725 3500.200 ;
        RECT 399.065 3499.920 399.345 3500.200 ;
        RECT 399.685 3499.920 399.965 3500.200 ;
        RECT 395.965 3418.090 396.245 3418.370 ;
        RECT 396.585 3418.090 396.865 3418.370 ;
        RECT 397.205 3418.090 397.485 3418.370 ;
        RECT 397.825 3418.090 398.105 3418.370 ;
        RECT 398.445 3418.090 398.725 3418.370 ;
        RECT 399.065 3418.090 399.345 3418.370 ;
        RECT 399.685 3418.090 399.965 3418.370 ;
        RECT 395.965 3417.470 396.245 3417.750 ;
        RECT 396.585 3417.470 396.865 3417.750 ;
        RECT 397.205 3417.470 397.485 3417.750 ;
        RECT 397.825 3417.470 398.105 3417.750 ;
        RECT 398.445 3417.470 398.725 3417.750 ;
        RECT 399.065 3417.470 399.345 3417.750 ;
        RECT 399.685 3417.470 399.965 3417.750 ;
        RECT 395.740 3402.670 396.020 3402.950 ;
        RECT 396.360 3402.670 396.640 3402.950 ;
        RECT 396.980 3402.670 397.260 3402.950 ;
        RECT 397.600 3402.670 397.880 3402.950 ;
        RECT 398.220 3402.670 398.500 3402.950 ;
        RECT 398.840 3402.670 399.120 3402.950 ;
        RECT 399.460 3402.670 399.740 3402.950 ;
        RECT 395.740 3402.050 396.020 3402.330 ;
        RECT 396.360 3402.050 396.640 3402.330 ;
        RECT 396.980 3402.050 397.260 3402.330 ;
        RECT 397.600 3402.050 397.880 3402.330 ;
        RECT 398.220 3402.050 398.500 3402.330 ;
        RECT 398.840 3402.050 399.120 3402.330 ;
        RECT 399.460 3402.050 399.740 3402.330 ;
        RECT 395.740 3401.430 396.020 3401.710 ;
        RECT 396.360 3401.430 396.640 3401.710 ;
        RECT 396.980 3401.430 397.260 3401.710 ;
        RECT 397.600 3401.430 397.880 3401.710 ;
        RECT 398.220 3401.430 398.500 3401.710 ;
        RECT 398.840 3401.430 399.120 3401.710 ;
        RECT 399.460 3401.430 399.740 3401.710 ;
        RECT 395.740 3400.810 396.020 3401.090 ;
        RECT 396.360 3400.810 396.640 3401.090 ;
        RECT 396.980 3400.810 397.260 3401.090 ;
        RECT 397.600 3400.810 397.880 3401.090 ;
        RECT 398.220 3400.810 398.500 3401.090 ;
        RECT 398.840 3400.810 399.120 3401.090 ;
        RECT 399.460 3400.810 399.740 3401.090 ;
        RECT 395.740 3400.190 396.020 3400.470 ;
        RECT 396.360 3400.190 396.640 3400.470 ;
        RECT 396.980 3400.190 397.260 3400.470 ;
        RECT 397.600 3400.190 397.880 3400.470 ;
        RECT 398.220 3400.190 398.500 3400.470 ;
        RECT 398.840 3400.190 399.120 3400.470 ;
        RECT 399.460 3400.190 399.740 3400.470 ;
        RECT 395.965 3383.090 396.245 3383.370 ;
        RECT 396.585 3383.090 396.865 3383.370 ;
        RECT 397.205 3383.090 397.485 3383.370 ;
        RECT 397.825 3383.090 398.105 3383.370 ;
        RECT 398.445 3383.090 398.725 3383.370 ;
        RECT 399.065 3383.090 399.345 3383.370 ;
        RECT 399.685 3383.090 399.965 3383.370 ;
        RECT 395.965 3382.470 396.245 3382.750 ;
        RECT 396.585 3382.470 396.865 3382.750 ;
        RECT 397.205 3382.470 397.485 3382.750 ;
        RECT 397.825 3382.470 398.105 3382.750 ;
        RECT 398.445 3382.470 398.725 3382.750 ;
        RECT 399.065 3382.470 399.345 3382.750 ;
        RECT 399.685 3382.470 399.965 3382.750 ;
        RECT 395.965 3348.090 396.245 3348.370 ;
        RECT 396.585 3348.090 396.865 3348.370 ;
        RECT 397.205 3348.090 397.485 3348.370 ;
        RECT 397.825 3348.090 398.105 3348.370 ;
        RECT 398.445 3348.090 398.725 3348.370 ;
        RECT 399.065 3348.090 399.345 3348.370 ;
        RECT 399.685 3348.090 399.965 3348.370 ;
        RECT 395.965 3347.470 396.245 3347.750 ;
        RECT 396.585 3347.470 396.865 3347.750 ;
        RECT 397.205 3347.470 397.485 3347.750 ;
        RECT 397.825 3347.470 398.105 3347.750 ;
        RECT 398.445 3347.470 398.725 3347.750 ;
        RECT 399.065 3347.470 399.345 3347.750 ;
        RECT 399.685 3347.470 399.965 3347.750 ;
        RECT 395.965 3294.920 396.245 3295.200 ;
        RECT 396.585 3294.920 396.865 3295.200 ;
        RECT 397.205 3294.920 397.485 3295.200 ;
        RECT 397.825 3294.920 398.105 3295.200 ;
        RECT 398.445 3294.920 398.725 3295.200 ;
        RECT 399.065 3294.920 399.345 3295.200 ;
        RECT 399.685 3294.920 399.965 3295.200 ;
        RECT 395.740 3222.670 396.020 3222.950 ;
        RECT 396.360 3222.670 396.640 3222.950 ;
        RECT 396.980 3222.670 397.260 3222.950 ;
        RECT 397.600 3222.670 397.880 3222.950 ;
        RECT 398.220 3222.670 398.500 3222.950 ;
        RECT 398.840 3222.670 399.120 3222.950 ;
        RECT 399.460 3222.670 399.740 3222.950 ;
        RECT 395.740 3222.050 396.020 3222.330 ;
        RECT 396.360 3222.050 396.640 3222.330 ;
        RECT 396.980 3222.050 397.260 3222.330 ;
        RECT 397.600 3222.050 397.880 3222.330 ;
        RECT 398.220 3222.050 398.500 3222.330 ;
        RECT 398.840 3222.050 399.120 3222.330 ;
        RECT 399.460 3222.050 399.740 3222.330 ;
        RECT 395.740 3221.430 396.020 3221.710 ;
        RECT 396.360 3221.430 396.640 3221.710 ;
        RECT 396.980 3221.430 397.260 3221.710 ;
        RECT 397.600 3221.430 397.880 3221.710 ;
        RECT 398.220 3221.430 398.500 3221.710 ;
        RECT 398.840 3221.430 399.120 3221.710 ;
        RECT 399.460 3221.430 399.740 3221.710 ;
        RECT 395.740 3220.810 396.020 3221.090 ;
        RECT 396.360 3220.810 396.640 3221.090 ;
        RECT 396.980 3220.810 397.260 3221.090 ;
        RECT 397.600 3220.810 397.880 3221.090 ;
        RECT 398.220 3220.810 398.500 3221.090 ;
        RECT 398.840 3220.810 399.120 3221.090 ;
        RECT 399.460 3220.810 399.740 3221.090 ;
        RECT 395.740 3220.190 396.020 3220.470 ;
        RECT 396.360 3220.190 396.640 3220.470 ;
        RECT 396.980 3220.190 397.260 3220.470 ;
        RECT 397.600 3220.190 397.880 3220.470 ;
        RECT 398.220 3220.190 398.500 3220.470 ;
        RECT 398.840 3220.190 399.120 3220.470 ;
        RECT 399.460 3220.190 399.740 3220.470 ;
        RECT 395.965 3213.090 396.245 3213.370 ;
        RECT 396.585 3213.090 396.865 3213.370 ;
        RECT 397.205 3213.090 397.485 3213.370 ;
        RECT 397.825 3213.090 398.105 3213.370 ;
        RECT 398.445 3213.090 398.725 3213.370 ;
        RECT 399.065 3213.090 399.345 3213.370 ;
        RECT 399.685 3213.090 399.965 3213.370 ;
        RECT 395.965 3212.470 396.245 3212.750 ;
        RECT 396.585 3212.470 396.865 3212.750 ;
        RECT 397.205 3212.470 397.485 3212.750 ;
        RECT 397.825 3212.470 398.105 3212.750 ;
        RECT 398.445 3212.470 398.725 3212.750 ;
        RECT 399.065 3212.470 399.345 3212.750 ;
        RECT 399.685 3212.470 399.965 3212.750 ;
        RECT 395.965 3178.090 396.245 3178.370 ;
        RECT 396.585 3178.090 396.865 3178.370 ;
        RECT 397.205 3178.090 397.485 3178.370 ;
        RECT 397.825 3178.090 398.105 3178.370 ;
        RECT 398.445 3178.090 398.725 3178.370 ;
        RECT 399.065 3178.090 399.345 3178.370 ;
        RECT 399.685 3178.090 399.965 3178.370 ;
        RECT 395.965 3177.470 396.245 3177.750 ;
        RECT 396.585 3177.470 396.865 3177.750 ;
        RECT 397.205 3177.470 397.485 3177.750 ;
        RECT 397.825 3177.470 398.105 3177.750 ;
        RECT 398.445 3177.470 398.725 3177.750 ;
        RECT 399.065 3177.470 399.345 3177.750 ;
        RECT 399.685 3177.470 399.965 3177.750 ;
        RECT 395.965 3143.090 396.245 3143.370 ;
        RECT 396.585 3143.090 396.865 3143.370 ;
        RECT 397.205 3143.090 397.485 3143.370 ;
        RECT 397.825 3143.090 398.105 3143.370 ;
        RECT 398.445 3143.090 398.725 3143.370 ;
        RECT 399.065 3143.090 399.345 3143.370 ;
        RECT 399.685 3143.090 399.965 3143.370 ;
        RECT 395.965 3142.470 396.245 3142.750 ;
        RECT 396.585 3142.470 396.865 3142.750 ;
        RECT 397.205 3142.470 397.485 3142.750 ;
        RECT 397.825 3142.470 398.105 3142.750 ;
        RECT 398.445 3142.470 398.725 3142.750 ;
        RECT 399.065 3142.470 399.345 3142.750 ;
        RECT 399.685 3142.470 399.965 3142.750 ;
        RECT 395.965 3089.920 396.245 3090.200 ;
        RECT 396.585 3089.920 396.865 3090.200 ;
        RECT 397.205 3089.920 397.485 3090.200 ;
        RECT 397.825 3089.920 398.105 3090.200 ;
        RECT 398.445 3089.920 398.725 3090.200 ;
        RECT 399.065 3089.920 399.345 3090.200 ;
        RECT 399.685 3089.920 399.965 3090.200 ;
        RECT 395.740 3042.670 396.020 3042.950 ;
        RECT 396.360 3042.670 396.640 3042.950 ;
        RECT 396.980 3042.670 397.260 3042.950 ;
        RECT 397.600 3042.670 397.880 3042.950 ;
        RECT 398.220 3042.670 398.500 3042.950 ;
        RECT 398.840 3042.670 399.120 3042.950 ;
        RECT 399.460 3042.670 399.740 3042.950 ;
        RECT 395.740 3042.050 396.020 3042.330 ;
        RECT 396.360 3042.050 396.640 3042.330 ;
        RECT 396.980 3042.050 397.260 3042.330 ;
        RECT 397.600 3042.050 397.880 3042.330 ;
        RECT 398.220 3042.050 398.500 3042.330 ;
        RECT 398.840 3042.050 399.120 3042.330 ;
        RECT 399.460 3042.050 399.740 3042.330 ;
        RECT 395.740 3041.430 396.020 3041.710 ;
        RECT 396.360 3041.430 396.640 3041.710 ;
        RECT 396.980 3041.430 397.260 3041.710 ;
        RECT 397.600 3041.430 397.880 3041.710 ;
        RECT 398.220 3041.430 398.500 3041.710 ;
        RECT 398.840 3041.430 399.120 3041.710 ;
        RECT 399.460 3041.430 399.740 3041.710 ;
        RECT 395.740 3040.810 396.020 3041.090 ;
        RECT 396.360 3040.810 396.640 3041.090 ;
        RECT 396.980 3040.810 397.260 3041.090 ;
        RECT 397.600 3040.810 397.880 3041.090 ;
        RECT 398.220 3040.810 398.500 3041.090 ;
        RECT 398.840 3040.810 399.120 3041.090 ;
        RECT 399.460 3040.810 399.740 3041.090 ;
        RECT 395.740 3040.190 396.020 3040.470 ;
        RECT 396.360 3040.190 396.640 3040.470 ;
        RECT 396.980 3040.190 397.260 3040.470 ;
        RECT 397.600 3040.190 397.880 3040.470 ;
        RECT 398.220 3040.190 398.500 3040.470 ;
        RECT 398.840 3040.190 399.120 3040.470 ;
        RECT 399.460 3040.190 399.740 3040.470 ;
        RECT 395.965 3008.090 396.245 3008.370 ;
        RECT 396.585 3008.090 396.865 3008.370 ;
        RECT 397.205 3008.090 397.485 3008.370 ;
        RECT 397.825 3008.090 398.105 3008.370 ;
        RECT 398.445 3008.090 398.725 3008.370 ;
        RECT 399.065 3008.090 399.345 3008.370 ;
        RECT 399.685 3008.090 399.965 3008.370 ;
        RECT 395.965 3007.470 396.245 3007.750 ;
        RECT 396.585 3007.470 396.865 3007.750 ;
        RECT 397.205 3007.470 397.485 3007.750 ;
        RECT 397.825 3007.470 398.105 3007.750 ;
        RECT 398.445 3007.470 398.725 3007.750 ;
        RECT 399.065 3007.470 399.345 3007.750 ;
        RECT 399.685 3007.470 399.965 3007.750 ;
        RECT 395.965 2973.090 396.245 2973.370 ;
        RECT 396.585 2973.090 396.865 2973.370 ;
        RECT 397.205 2973.090 397.485 2973.370 ;
        RECT 397.825 2973.090 398.105 2973.370 ;
        RECT 398.445 2973.090 398.725 2973.370 ;
        RECT 399.065 2973.090 399.345 2973.370 ;
        RECT 399.685 2973.090 399.965 2973.370 ;
        RECT 395.965 2972.470 396.245 2972.750 ;
        RECT 396.585 2972.470 396.865 2972.750 ;
        RECT 397.205 2972.470 397.485 2972.750 ;
        RECT 397.825 2972.470 398.105 2972.750 ;
        RECT 398.445 2972.470 398.725 2972.750 ;
        RECT 399.065 2972.470 399.345 2972.750 ;
        RECT 399.685 2972.470 399.965 2972.750 ;
        RECT 395.965 2938.090 396.245 2938.370 ;
        RECT 396.585 2938.090 396.865 2938.370 ;
        RECT 397.205 2938.090 397.485 2938.370 ;
        RECT 397.825 2938.090 398.105 2938.370 ;
        RECT 398.445 2938.090 398.725 2938.370 ;
        RECT 399.065 2938.090 399.345 2938.370 ;
        RECT 399.685 2938.090 399.965 2938.370 ;
        RECT 395.965 2937.470 396.245 2937.750 ;
        RECT 396.585 2937.470 396.865 2937.750 ;
        RECT 397.205 2937.470 397.485 2937.750 ;
        RECT 397.825 2937.470 398.105 2937.750 ;
        RECT 398.445 2937.470 398.725 2937.750 ;
        RECT 399.065 2937.470 399.345 2937.750 ;
        RECT 399.685 2937.470 399.965 2937.750 ;
        RECT 395.965 2884.920 396.245 2885.200 ;
        RECT 396.585 2884.920 396.865 2885.200 ;
        RECT 397.205 2884.920 397.485 2885.200 ;
        RECT 397.825 2884.920 398.105 2885.200 ;
        RECT 398.445 2884.920 398.725 2885.200 ;
        RECT 399.065 2884.920 399.345 2885.200 ;
        RECT 399.685 2884.920 399.965 2885.200 ;
        RECT 395.740 2862.670 396.020 2862.950 ;
        RECT 396.360 2862.670 396.640 2862.950 ;
        RECT 396.980 2862.670 397.260 2862.950 ;
        RECT 397.600 2862.670 397.880 2862.950 ;
        RECT 398.220 2862.670 398.500 2862.950 ;
        RECT 398.840 2862.670 399.120 2862.950 ;
        RECT 399.460 2862.670 399.740 2862.950 ;
        RECT 395.740 2862.050 396.020 2862.330 ;
        RECT 396.360 2862.050 396.640 2862.330 ;
        RECT 396.980 2862.050 397.260 2862.330 ;
        RECT 397.600 2862.050 397.880 2862.330 ;
        RECT 398.220 2862.050 398.500 2862.330 ;
        RECT 398.840 2862.050 399.120 2862.330 ;
        RECT 399.460 2862.050 399.740 2862.330 ;
        RECT 395.740 2861.430 396.020 2861.710 ;
        RECT 396.360 2861.430 396.640 2861.710 ;
        RECT 396.980 2861.430 397.260 2861.710 ;
        RECT 397.600 2861.430 397.880 2861.710 ;
        RECT 398.220 2861.430 398.500 2861.710 ;
        RECT 398.840 2861.430 399.120 2861.710 ;
        RECT 399.460 2861.430 399.740 2861.710 ;
        RECT 395.740 2860.810 396.020 2861.090 ;
        RECT 396.360 2860.810 396.640 2861.090 ;
        RECT 396.980 2860.810 397.260 2861.090 ;
        RECT 397.600 2860.810 397.880 2861.090 ;
        RECT 398.220 2860.810 398.500 2861.090 ;
        RECT 398.840 2860.810 399.120 2861.090 ;
        RECT 399.460 2860.810 399.740 2861.090 ;
        RECT 395.740 2860.190 396.020 2860.470 ;
        RECT 396.360 2860.190 396.640 2860.470 ;
        RECT 396.980 2860.190 397.260 2860.470 ;
        RECT 397.600 2860.190 397.880 2860.470 ;
        RECT 398.220 2860.190 398.500 2860.470 ;
        RECT 398.840 2860.190 399.120 2860.470 ;
        RECT 399.460 2860.190 399.740 2860.470 ;
        RECT 395.965 2803.090 396.245 2803.370 ;
        RECT 396.585 2803.090 396.865 2803.370 ;
        RECT 397.205 2803.090 397.485 2803.370 ;
        RECT 397.825 2803.090 398.105 2803.370 ;
        RECT 398.445 2803.090 398.725 2803.370 ;
        RECT 399.065 2803.090 399.345 2803.370 ;
        RECT 399.685 2803.090 399.965 2803.370 ;
        RECT 395.965 2802.470 396.245 2802.750 ;
        RECT 396.585 2802.470 396.865 2802.750 ;
        RECT 397.205 2802.470 397.485 2802.750 ;
        RECT 397.825 2802.470 398.105 2802.750 ;
        RECT 398.445 2802.470 398.725 2802.750 ;
        RECT 399.065 2802.470 399.345 2802.750 ;
        RECT 399.685 2802.470 399.965 2802.750 ;
        RECT 395.965 2768.090 396.245 2768.370 ;
        RECT 396.585 2768.090 396.865 2768.370 ;
        RECT 397.205 2768.090 397.485 2768.370 ;
        RECT 397.825 2768.090 398.105 2768.370 ;
        RECT 398.445 2768.090 398.725 2768.370 ;
        RECT 399.065 2768.090 399.345 2768.370 ;
        RECT 399.685 2768.090 399.965 2768.370 ;
        RECT 395.965 2767.470 396.245 2767.750 ;
        RECT 396.585 2767.470 396.865 2767.750 ;
        RECT 397.205 2767.470 397.485 2767.750 ;
        RECT 397.825 2767.470 398.105 2767.750 ;
        RECT 398.445 2767.470 398.725 2767.750 ;
        RECT 399.065 2767.470 399.345 2767.750 ;
        RECT 399.685 2767.470 399.965 2767.750 ;
        RECT 395.965 2733.090 396.245 2733.370 ;
        RECT 396.585 2733.090 396.865 2733.370 ;
        RECT 397.205 2733.090 397.485 2733.370 ;
        RECT 397.825 2733.090 398.105 2733.370 ;
        RECT 398.445 2733.090 398.725 2733.370 ;
        RECT 399.065 2733.090 399.345 2733.370 ;
        RECT 399.685 2733.090 399.965 2733.370 ;
        RECT 395.965 2732.470 396.245 2732.750 ;
        RECT 396.585 2732.470 396.865 2732.750 ;
        RECT 397.205 2732.470 397.485 2732.750 ;
        RECT 397.825 2732.470 398.105 2732.750 ;
        RECT 398.445 2732.470 398.725 2732.750 ;
        RECT 399.065 2732.470 399.345 2732.750 ;
        RECT 399.685 2732.470 399.965 2732.750 ;
        RECT 395.740 2682.670 396.020 2682.950 ;
        RECT 396.360 2682.670 396.640 2682.950 ;
        RECT 396.980 2682.670 397.260 2682.950 ;
        RECT 397.600 2682.670 397.880 2682.950 ;
        RECT 398.220 2682.670 398.500 2682.950 ;
        RECT 398.840 2682.670 399.120 2682.950 ;
        RECT 399.460 2682.670 399.740 2682.950 ;
        RECT 395.740 2682.050 396.020 2682.330 ;
        RECT 396.360 2682.050 396.640 2682.330 ;
        RECT 396.980 2682.050 397.260 2682.330 ;
        RECT 397.600 2682.050 397.880 2682.330 ;
        RECT 398.220 2682.050 398.500 2682.330 ;
        RECT 398.840 2682.050 399.120 2682.330 ;
        RECT 399.460 2682.050 399.740 2682.330 ;
        RECT 395.740 2681.430 396.020 2681.710 ;
        RECT 396.360 2681.430 396.640 2681.710 ;
        RECT 396.980 2681.430 397.260 2681.710 ;
        RECT 397.600 2681.430 397.880 2681.710 ;
        RECT 398.220 2681.430 398.500 2681.710 ;
        RECT 398.840 2681.430 399.120 2681.710 ;
        RECT 399.460 2681.430 399.740 2681.710 ;
        RECT 395.740 2680.810 396.020 2681.090 ;
        RECT 396.360 2680.810 396.640 2681.090 ;
        RECT 396.980 2680.810 397.260 2681.090 ;
        RECT 397.600 2680.810 397.880 2681.090 ;
        RECT 398.220 2680.810 398.500 2681.090 ;
        RECT 398.840 2680.810 399.120 2681.090 ;
        RECT 399.460 2680.810 399.740 2681.090 ;
        RECT 395.965 2598.090 396.245 2598.370 ;
        RECT 396.585 2598.090 396.865 2598.370 ;
        RECT 397.205 2598.090 397.485 2598.370 ;
        RECT 397.825 2598.090 398.105 2598.370 ;
        RECT 398.445 2598.090 398.725 2598.370 ;
        RECT 399.065 2598.090 399.345 2598.370 ;
        RECT 399.685 2598.090 399.965 2598.370 ;
        RECT 395.965 2597.470 396.245 2597.750 ;
        RECT 396.585 2597.470 396.865 2597.750 ;
        RECT 397.205 2597.470 397.485 2597.750 ;
        RECT 397.825 2597.470 398.105 2597.750 ;
        RECT 398.445 2597.470 398.725 2597.750 ;
        RECT 399.065 2597.470 399.345 2597.750 ;
        RECT 399.685 2597.470 399.965 2597.750 ;
        RECT 395.965 2563.090 396.245 2563.370 ;
        RECT 396.585 2563.090 396.865 2563.370 ;
        RECT 397.205 2563.090 397.485 2563.370 ;
        RECT 397.825 2563.090 398.105 2563.370 ;
        RECT 398.445 2563.090 398.725 2563.370 ;
        RECT 399.065 2563.090 399.345 2563.370 ;
        RECT 399.685 2563.090 399.965 2563.370 ;
        RECT 395.965 2562.470 396.245 2562.750 ;
        RECT 396.585 2562.470 396.865 2562.750 ;
        RECT 397.205 2562.470 397.485 2562.750 ;
        RECT 397.825 2562.470 398.105 2562.750 ;
        RECT 398.445 2562.470 398.725 2562.750 ;
        RECT 399.065 2562.470 399.345 2562.750 ;
        RECT 399.685 2562.470 399.965 2562.750 ;
        RECT 395.965 2528.090 396.245 2528.370 ;
        RECT 396.585 2528.090 396.865 2528.370 ;
        RECT 397.205 2528.090 397.485 2528.370 ;
        RECT 397.825 2528.090 398.105 2528.370 ;
        RECT 398.445 2528.090 398.725 2528.370 ;
        RECT 399.065 2528.090 399.345 2528.370 ;
        RECT 399.685 2528.090 399.965 2528.370 ;
        RECT 395.965 2527.470 396.245 2527.750 ;
        RECT 396.585 2527.470 396.865 2527.750 ;
        RECT 397.205 2527.470 397.485 2527.750 ;
        RECT 397.825 2527.470 398.105 2527.750 ;
        RECT 398.445 2527.470 398.725 2527.750 ;
        RECT 399.065 2527.470 399.345 2527.750 ;
        RECT 399.685 2527.470 399.965 2527.750 ;
        RECT 395.740 2502.670 396.020 2502.950 ;
        RECT 396.360 2502.670 396.640 2502.950 ;
        RECT 396.980 2502.670 397.260 2502.950 ;
        RECT 397.600 2502.670 397.880 2502.950 ;
        RECT 398.220 2502.670 398.500 2502.950 ;
        RECT 398.840 2502.670 399.120 2502.950 ;
        RECT 399.460 2502.670 399.740 2502.950 ;
        RECT 395.740 2502.050 396.020 2502.330 ;
        RECT 396.360 2502.050 396.640 2502.330 ;
        RECT 396.980 2502.050 397.260 2502.330 ;
        RECT 397.600 2502.050 397.880 2502.330 ;
        RECT 398.220 2502.050 398.500 2502.330 ;
        RECT 398.840 2502.050 399.120 2502.330 ;
        RECT 399.460 2502.050 399.740 2502.330 ;
        RECT 395.740 2501.430 396.020 2501.710 ;
        RECT 396.360 2501.430 396.640 2501.710 ;
        RECT 396.980 2501.430 397.260 2501.710 ;
        RECT 397.600 2501.430 397.880 2501.710 ;
        RECT 398.220 2501.430 398.500 2501.710 ;
        RECT 398.840 2501.430 399.120 2501.710 ;
        RECT 399.460 2501.430 399.740 2501.710 ;
        RECT 395.740 2500.810 396.020 2501.090 ;
        RECT 396.360 2500.810 396.640 2501.090 ;
        RECT 396.980 2500.810 397.260 2501.090 ;
        RECT 397.600 2500.810 397.880 2501.090 ;
        RECT 398.220 2500.810 398.500 2501.090 ;
        RECT 398.840 2500.810 399.120 2501.090 ;
        RECT 399.460 2500.810 399.740 2501.090 ;
        RECT 395.740 2500.190 396.020 2500.470 ;
        RECT 396.360 2500.190 396.640 2500.470 ;
        RECT 396.980 2500.190 397.260 2500.470 ;
        RECT 397.600 2500.190 397.880 2500.470 ;
        RECT 398.220 2500.190 398.500 2500.470 ;
        RECT 398.840 2500.190 399.120 2500.470 ;
        RECT 399.460 2500.190 399.740 2500.470 ;
        RECT 396.040 2168.070 396.320 2168.350 ;
        RECT 396.660 2168.070 396.940 2168.350 ;
        RECT 397.280 2168.070 397.560 2168.350 ;
        RECT 397.900 2168.070 398.180 2168.350 ;
        RECT 398.520 2168.070 398.800 2168.350 ;
        RECT 399.140 2168.070 399.420 2168.350 ;
        RECT 399.760 2168.070 400.040 2168.350 ;
        RECT 396.040 2167.450 396.320 2167.730 ;
        RECT 396.660 2167.450 396.940 2167.730 ;
        RECT 397.280 2167.450 397.560 2167.730 ;
        RECT 397.900 2167.450 398.180 2167.730 ;
        RECT 398.520 2167.450 398.800 2167.730 ;
        RECT 399.140 2167.450 399.420 2167.730 ;
        RECT 399.760 2167.450 400.040 2167.730 ;
        RECT 396.040 2166.830 396.320 2167.110 ;
        RECT 396.660 2166.830 396.940 2167.110 ;
        RECT 397.280 2166.830 397.560 2167.110 ;
        RECT 397.900 2166.830 398.180 2167.110 ;
        RECT 398.520 2166.830 398.800 2167.110 ;
        RECT 399.140 2166.830 399.420 2167.110 ;
        RECT 399.760 2166.830 400.040 2167.110 ;
        RECT 396.040 2166.210 396.320 2166.490 ;
        RECT 396.660 2166.210 396.940 2166.490 ;
        RECT 397.280 2166.210 397.560 2166.490 ;
        RECT 397.900 2166.210 398.180 2166.490 ;
        RECT 398.520 2166.210 398.800 2166.490 ;
        RECT 399.140 2166.210 399.420 2166.490 ;
        RECT 399.760 2166.210 400.040 2166.490 ;
        RECT 396.040 2165.590 396.320 2165.870 ;
        RECT 396.660 2165.590 396.940 2165.870 ;
        RECT 397.280 2165.590 397.560 2165.870 ;
        RECT 397.900 2165.590 398.180 2165.870 ;
        RECT 398.520 2165.590 398.800 2165.870 ;
        RECT 399.140 2165.590 399.420 2165.870 ;
        RECT 399.760 2165.590 400.040 2165.870 ;
        RECT 396.040 2164.970 396.320 2165.250 ;
        RECT 396.660 2164.970 396.940 2165.250 ;
        RECT 397.280 2164.970 397.560 2165.250 ;
        RECT 397.900 2164.970 398.180 2165.250 ;
        RECT 398.520 2164.970 398.800 2165.250 ;
        RECT 399.140 2164.970 399.420 2165.250 ;
        RECT 399.760 2164.970 400.040 2165.250 ;
        RECT 396.040 2164.350 396.320 2164.630 ;
        RECT 396.660 2164.350 396.940 2164.630 ;
        RECT 397.280 2164.350 397.560 2164.630 ;
        RECT 397.900 2164.350 398.180 2164.630 ;
        RECT 398.520 2164.350 398.800 2164.630 ;
        RECT 399.140 2164.350 399.420 2164.630 ;
        RECT 399.760 2164.350 400.040 2164.630 ;
        RECT 396.040 2163.730 396.320 2164.010 ;
        RECT 396.660 2163.730 396.940 2164.010 ;
        RECT 397.280 2163.730 397.560 2164.010 ;
        RECT 397.900 2163.730 398.180 2164.010 ;
        RECT 398.520 2163.730 398.800 2164.010 ;
        RECT 399.140 2163.730 399.420 2164.010 ;
        RECT 399.760 2163.730 400.040 2164.010 ;
        RECT 396.040 2163.110 396.320 2163.390 ;
        RECT 396.660 2163.110 396.940 2163.390 ;
        RECT 397.280 2163.110 397.560 2163.390 ;
        RECT 397.900 2163.110 398.180 2163.390 ;
        RECT 398.520 2163.110 398.800 2163.390 ;
        RECT 399.140 2163.110 399.420 2163.390 ;
        RECT 399.760 2163.110 400.040 2163.390 ;
        RECT 396.040 2162.490 396.320 2162.770 ;
        RECT 396.660 2162.490 396.940 2162.770 ;
        RECT 397.280 2162.490 397.560 2162.770 ;
        RECT 397.900 2162.490 398.180 2162.770 ;
        RECT 398.520 2162.490 398.800 2162.770 ;
        RECT 399.140 2162.490 399.420 2162.770 ;
        RECT 399.760 2162.490 400.040 2162.770 ;
        RECT 396.040 2161.870 396.320 2162.150 ;
        RECT 396.660 2161.870 396.940 2162.150 ;
        RECT 397.280 2161.870 397.560 2162.150 ;
        RECT 397.900 2161.870 398.180 2162.150 ;
        RECT 398.520 2161.870 398.800 2162.150 ;
        RECT 399.140 2161.870 399.420 2162.150 ;
        RECT 399.760 2161.870 400.040 2162.150 ;
        RECT 396.040 2161.250 396.320 2161.530 ;
        RECT 396.660 2161.250 396.940 2161.530 ;
        RECT 397.280 2161.250 397.560 2161.530 ;
        RECT 397.900 2161.250 398.180 2161.530 ;
        RECT 398.520 2161.250 398.800 2161.530 ;
        RECT 399.140 2161.250 399.420 2161.530 ;
        RECT 399.760 2161.250 400.040 2161.530 ;
        RECT 396.040 2160.630 396.320 2160.910 ;
        RECT 396.660 2160.630 396.940 2160.910 ;
        RECT 397.280 2160.630 397.560 2160.910 ;
        RECT 397.900 2160.630 398.180 2160.910 ;
        RECT 398.520 2160.630 398.800 2160.910 ;
        RECT 399.140 2160.630 399.420 2160.910 ;
        RECT 399.760 2160.630 400.040 2160.910 ;
        RECT 396.040 2160.010 396.320 2160.290 ;
        RECT 396.660 2160.010 396.940 2160.290 ;
        RECT 397.280 2160.010 397.560 2160.290 ;
        RECT 397.900 2160.010 398.180 2160.290 ;
        RECT 398.520 2160.010 398.800 2160.290 ;
        RECT 399.140 2160.010 399.420 2160.290 ;
        RECT 399.760 2160.010 400.040 2160.290 ;
        RECT 396.040 2159.390 396.320 2159.670 ;
        RECT 396.660 2159.390 396.940 2159.670 ;
        RECT 397.280 2159.390 397.560 2159.670 ;
        RECT 397.900 2159.390 398.180 2159.670 ;
        RECT 398.520 2159.390 398.800 2159.670 ;
        RECT 399.140 2159.390 399.420 2159.670 ;
        RECT 399.760 2159.390 400.040 2159.670 ;
        RECT 396.040 2155.670 396.320 2155.950 ;
        RECT 396.660 2155.670 396.940 2155.950 ;
        RECT 397.280 2155.670 397.560 2155.950 ;
        RECT 397.900 2155.670 398.180 2155.950 ;
        RECT 398.520 2155.670 398.800 2155.950 ;
        RECT 399.140 2155.670 399.420 2155.950 ;
        RECT 399.760 2155.670 400.040 2155.950 ;
        RECT 396.040 2155.050 396.320 2155.330 ;
        RECT 396.660 2155.050 396.940 2155.330 ;
        RECT 397.280 2155.050 397.560 2155.330 ;
        RECT 397.900 2155.050 398.180 2155.330 ;
        RECT 398.520 2155.050 398.800 2155.330 ;
        RECT 399.140 2155.050 399.420 2155.330 ;
        RECT 399.760 2155.050 400.040 2155.330 ;
        RECT 396.040 2154.430 396.320 2154.710 ;
        RECT 396.660 2154.430 396.940 2154.710 ;
        RECT 397.280 2154.430 397.560 2154.710 ;
        RECT 397.900 2154.430 398.180 2154.710 ;
        RECT 398.520 2154.430 398.800 2154.710 ;
        RECT 399.140 2154.430 399.420 2154.710 ;
        RECT 399.760 2154.430 400.040 2154.710 ;
        RECT 396.040 2153.810 396.320 2154.090 ;
        RECT 396.660 2153.810 396.940 2154.090 ;
        RECT 397.280 2153.810 397.560 2154.090 ;
        RECT 397.900 2153.810 398.180 2154.090 ;
        RECT 398.520 2153.810 398.800 2154.090 ;
        RECT 399.140 2153.810 399.420 2154.090 ;
        RECT 399.760 2153.810 400.040 2154.090 ;
        RECT 396.040 2153.190 396.320 2153.470 ;
        RECT 396.660 2153.190 396.940 2153.470 ;
        RECT 397.280 2153.190 397.560 2153.470 ;
        RECT 397.900 2153.190 398.180 2153.470 ;
        RECT 398.520 2153.190 398.800 2153.470 ;
        RECT 399.140 2153.190 399.420 2153.470 ;
        RECT 399.760 2153.190 400.040 2153.470 ;
        RECT 396.040 2152.570 396.320 2152.850 ;
        RECT 396.660 2152.570 396.940 2152.850 ;
        RECT 397.280 2152.570 397.560 2152.850 ;
        RECT 397.900 2152.570 398.180 2152.850 ;
        RECT 398.520 2152.570 398.800 2152.850 ;
        RECT 399.140 2152.570 399.420 2152.850 ;
        RECT 399.760 2152.570 400.040 2152.850 ;
        RECT 396.040 2151.950 396.320 2152.230 ;
        RECT 396.660 2151.950 396.940 2152.230 ;
        RECT 397.280 2151.950 397.560 2152.230 ;
        RECT 397.900 2151.950 398.180 2152.230 ;
        RECT 398.520 2151.950 398.800 2152.230 ;
        RECT 399.140 2151.950 399.420 2152.230 ;
        RECT 399.760 2151.950 400.040 2152.230 ;
        RECT 396.040 2151.330 396.320 2151.610 ;
        RECT 396.660 2151.330 396.940 2151.610 ;
        RECT 397.280 2151.330 397.560 2151.610 ;
        RECT 397.900 2151.330 398.180 2151.610 ;
        RECT 398.520 2151.330 398.800 2151.610 ;
        RECT 399.140 2151.330 399.420 2151.610 ;
        RECT 399.760 2151.330 400.040 2151.610 ;
        RECT 396.040 2150.710 396.320 2150.990 ;
        RECT 396.660 2150.710 396.940 2150.990 ;
        RECT 397.280 2150.710 397.560 2150.990 ;
        RECT 397.900 2150.710 398.180 2150.990 ;
        RECT 398.520 2150.710 398.800 2150.990 ;
        RECT 399.140 2150.710 399.420 2150.990 ;
        RECT 399.760 2150.710 400.040 2150.990 ;
        RECT 396.040 2150.090 396.320 2150.370 ;
        RECT 396.660 2150.090 396.940 2150.370 ;
        RECT 397.280 2150.090 397.560 2150.370 ;
        RECT 397.900 2150.090 398.180 2150.370 ;
        RECT 398.520 2150.090 398.800 2150.370 ;
        RECT 399.140 2150.090 399.420 2150.370 ;
        RECT 399.760 2150.090 400.040 2150.370 ;
        RECT 396.040 2149.470 396.320 2149.750 ;
        RECT 396.660 2149.470 396.940 2149.750 ;
        RECT 397.280 2149.470 397.560 2149.750 ;
        RECT 397.900 2149.470 398.180 2149.750 ;
        RECT 398.520 2149.470 398.800 2149.750 ;
        RECT 399.140 2149.470 399.420 2149.750 ;
        RECT 399.760 2149.470 400.040 2149.750 ;
        RECT 396.040 2148.850 396.320 2149.130 ;
        RECT 396.660 2148.850 396.940 2149.130 ;
        RECT 397.280 2148.850 397.560 2149.130 ;
        RECT 397.900 2148.850 398.180 2149.130 ;
        RECT 398.520 2148.850 398.800 2149.130 ;
        RECT 399.140 2148.850 399.420 2149.130 ;
        RECT 399.760 2148.850 400.040 2149.130 ;
        RECT 396.040 2148.230 396.320 2148.510 ;
        RECT 396.660 2148.230 396.940 2148.510 ;
        RECT 397.280 2148.230 397.560 2148.510 ;
        RECT 397.900 2148.230 398.180 2148.510 ;
        RECT 398.520 2148.230 398.800 2148.510 ;
        RECT 399.140 2148.230 399.420 2148.510 ;
        RECT 399.760 2148.230 400.040 2148.510 ;
        RECT 396.040 2147.610 396.320 2147.890 ;
        RECT 396.660 2147.610 396.940 2147.890 ;
        RECT 397.280 2147.610 397.560 2147.890 ;
        RECT 397.900 2147.610 398.180 2147.890 ;
        RECT 398.520 2147.610 398.800 2147.890 ;
        RECT 399.140 2147.610 399.420 2147.890 ;
        RECT 399.760 2147.610 400.040 2147.890 ;
        RECT 396.040 2146.990 396.320 2147.270 ;
        RECT 396.660 2146.990 396.940 2147.270 ;
        RECT 397.280 2146.990 397.560 2147.270 ;
        RECT 397.900 2146.990 398.180 2147.270 ;
        RECT 398.520 2146.990 398.800 2147.270 ;
        RECT 399.140 2146.990 399.420 2147.270 ;
        RECT 399.760 2146.990 400.040 2147.270 ;
        RECT 396.040 2146.370 396.320 2146.650 ;
        RECT 396.660 2146.370 396.940 2146.650 ;
        RECT 397.280 2146.370 397.560 2146.650 ;
        RECT 397.900 2146.370 398.180 2146.650 ;
        RECT 398.520 2146.370 398.800 2146.650 ;
        RECT 399.140 2146.370 399.420 2146.650 ;
        RECT 399.760 2146.370 400.040 2146.650 ;
        RECT 396.040 2143.820 396.320 2144.100 ;
        RECT 396.660 2143.820 396.940 2144.100 ;
        RECT 397.280 2143.820 397.560 2144.100 ;
        RECT 397.900 2143.820 398.180 2144.100 ;
        RECT 398.520 2143.820 398.800 2144.100 ;
        RECT 399.140 2143.820 399.420 2144.100 ;
        RECT 399.760 2143.820 400.040 2144.100 ;
        RECT 396.040 2143.200 396.320 2143.480 ;
        RECT 396.660 2143.200 396.940 2143.480 ;
        RECT 397.280 2143.200 397.560 2143.480 ;
        RECT 397.900 2143.200 398.180 2143.480 ;
        RECT 398.520 2143.200 398.800 2143.480 ;
        RECT 399.140 2143.200 399.420 2143.480 ;
        RECT 399.760 2143.200 400.040 2143.480 ;
        RECT 396.040 2142.580 396.320 2142.860 ;
        RECT 396.660 2142.580 396.940 2142.860 ;
        RECT 397.280 2142.580 397.560 2142.860 ;
        RECT 397.900 2142.580 398.180 2142.860 ;
        RECT 398.520 2142.580 398.800 2142.860 ;
        RECT 399.140 2142.580 399.420 2142.860 ;
        RECT 399.760 2142.580 400.040 2142.860 ;
        RECT 396.040 2141.960 396.320 2142.240 ;
        RECT 396.660 2141.960 396.940 2142.240 ;
        RECT 397.280 2141.960 397.560 2142.240 ;
        RECT 397.900 2141.960 398.180 2142.240 ;
        RECT 398.520 2141.960 398.800 2142.240 ;
        RECT 399.140 2141.960 399.420 2142.240 ;
        RECT 399.760 2141.960 400.040 2142.240 ;
        RECT 396.040 2141.340 396.320 2141.620 ;
        RECT 396.660 2141.340 396.940 2141.620 ;
        RECT 397.280 2141.340 397.560 2141.620 ;
        RECT 397.900 2141.340 398.180 2141.620 ;
        RECT 398.520 2141.340 398.800 2141.620 ;
        RECT 399.140 2141.340 399.420 2141.620 ;
        RECT 399.760 2141.340 400.040 2141.620 ;
        RECT 396.040 2140.720 396.320 2141.000 ;
        RECT 396.660 2140.720 396.940 2141.000 ;
        RECT 397.280 2140.720 397.560 2141.000 ;
        RECT 397.900 2140.720 398.180 2141.000 ;
        RECT 398.520 2140.720 398.800 2141.000 ;
        RECT 399.140 2140.720 399.420 2141.000 ;
        RECT 399.760 2140.720 400.040 2141.000 ;
        RECT 396.040 2140.100 396.320 2140.380 ;
        RECT 396.660 2140.100 396.940 2140.380 ;
        RECT 397.280 2140.100 397.560 2140.380 ;
        RECT 397.900 2140.100 398.180 2140.380 ;
        RECT 398.520 2140.100 398.800 2140.380 ;
        RECT 399.140 2140.100 399.420 2140.380 ;
        RECT 399.760 2140.100 400.040 2140.380 ;
        RECT 396.040 2139.480 396.320 2139.760 ;
        RECT 396.660 2139.480 396.940 2139.760 ;
        RECT 397.280 2139.480 397.560 2139.760 ;
        RECT 397.900 2139.480 398.180 2139.760 ;
        RECT 398.520 2139.480 398.800 2139.760 ;
        RECT 399.140 2139.480 399.420 2139.760 ;
        RECT 399.760 2139.480 400.040 2139.760 ;
        RECT 396.040 2138.860 396.320 2139.140 ;
        RECT 396.660 2138.860 396.940 2139.140 ;
        RECT 397.280 2138.860 397.560 2139.140 ;
        RECT 397.900 2138.860 398.180 2139.140 ;
        RECT 398.520 2138.860 398.800 2139.140 ;
        RECT 399.140 2138.860 399.420 2139.140 ;
        RECT 399.760 2138.860 400.040 2139.140 ;
        RECT 396.040 2138.240 396.320 2138.520 ;
        RECT 396.660 2138.240 396.940 2138.520 ;
        RECT 397.280 2138.240 397.560 2138.520 ;
        RECT 397.900 2138.240 398.180 2138.520 ;
        RECT 398.520 2138.240 398.800 2138.520 ;
        RECT 399.140 2138.240 399.420 2138.520 ;
        RECT 399.760 2138.240 400.040 2138.520 ;
        RECT 396.040 2137.620 396.320 2137.900 ;
        RECT 396.660 2137.620 396.940 2137.900 ;
        RECT 397.280 2137.620 397.560 2137.900 ;
        RECT 397.900 2137.620 398.180 2137.900 ;
        RECT 398.520 2137.620 398.800 2137.900 ;
        RECT 399.140 2137.620 399.420 2137.900 ;
        RECT 399.760 2137.620 400.040 2137.900 ;
        RECT 396.040 2137.000 396.320 2137.280 ;
        RECT 396.660 2137.000 396.940 2137.280 ;
        RECT 397.280 2137.000 397.560 2137.280 ;
        RECT 397.900 2137.000 398.180 2137.280 ;
        RECT 398.520 2137.000 398.800 2137.280 ;
        RECT 399.140 2137.000 399.420 2137.280 ;
        RECT 399.760 2137.000 400.040 2137.280 ;
        RECT 396.040 2136.380 396.320 2136.660 ;
        RECT 396.660 2136.380 396.940 2136.660 ;
        RECT 397.280 2136.380 397.560 2136.660 ;
        RECT 397.900 2136.380 398.180 2136.660 ;
        RECT 398.520 2136.380 398.800 2136.660 ;
        RECT 399.140 2136.380 399.420 2136.660 ;
        RECT 399.760 2136.380 400.040 2136.660 ;
        RECT 396.040 2135.760 396.320 2136.040 ;
        RECT 396.660 2135.760 396.940 2136.040 ;
        RECT 397.280 2135.760 397.560 2136.040 ;
        RECT 397.900 2135.760 398.180 2136.040 ;
        RECT 398.520 2135.760 398.800 2136.040 ;
        RECT 399.140 2135.760 399.420 2136.040 ;
        RECT 399.760 2135.760 400.040 2136.040 ;
        RECT 396.040 2135.140 396.320 2135.420 ;
        RECT 396.660 2135.140 396.940 2135.420 ;
        RECT 397.280 2135.140 397.560 2135.420 ;
        RECT 397.900 2135.140 398.180 2135.420 ;
        RECT 398.520 2135.140 398.800 2135.420 ;
        RECT 399.140 2135.140 399.420 2135.420 ;
        RECT 399.760 2135.140 400.040 2135.420 ;
        RECT 396.040 2134.520 396.320 2134.800 ;
        RECT 396.660 2134.520 396.940 2134.800 ;
        RECT 397.280 2134.520 397.560 2134.800 ;
        RECT 397.900 2134.520 398.180 2134.800 ;
        RECT 398.520 2134.520 398.800 2134.800 ;
        RECT 399.140 2134.520 399.420 2134.800 ;
        RECT 399.760 2134.520 400.040 2134.800 ;
        RECT 396.040 2130.290 396.320 2130.570 ;
        RECT 396.660 2130.290 396.940 2130.570 ;
        RECT 397.280 2130.290 397.560 2130.570 ;
        RECT 397.900 2130.290 398.180 2130.570 ;
        RECT 398.520 2130.290 398.800 2130.570 ;
        RECT 399.140 2130.290 399.420 2130.570 ;
        RECT 399.760 2130.290 400.040 2130.570 ;
        RECT 396.040 2129.670 396.320 2129.950 ;
        RECT 396.660 2129.670 396.940 2129.950 ;
        RECT 397.280 2129.670 397.560 2129.950 ;
        RECT 397.900 2129.670 398.180 2129.950 ;
        RECT 398.520 2129.670 398.800 2129.950 ;
        RECT 399.140 2129.670 399.420 2129.950 ;
        RECT 399.760 2129.670 400.040 2129.950 ;
        RECT 396.040 2129.050 396.320 2129.330 ;
        RECT 396.660 2129.050 396.940 2129.330 ;
        RECT 397.280 2129.050 397.560 2129.330 ;
        RECT 397.900 2129.050 398.180 2129.330 ;
        RECT 398.520 2129.050 398.800 2129.330 ;
        RECT 399.140 2129.050 399.420 2129.330 ;
        RECT 399.760 2129.050 400.040 2129.330 ;
        RECT 396.040 2128.430 396.320 2128.710 ;
        RECT 396.660 2128.430 396.940 2128.710 ;
        RECT 397.280 2128.430 397.560 2128.710 ;
        RECT 397.900 2128.430 398.180 2128.710 ;
        RECT 398.520 2128.430 398.800 2128.710 ;
        RECT 399.140 2128.430 399.420 2128.710 ;
        RECT 399.760 2128.430 400.040 2128.710 ;
        RECT 396.040 2127.810 396.320 2128.090 ;
        RECT 396.660 2127.810 396.940 2128.090 ;
        RECT 397.280 2127.810 397.560 2128.090 ;
        RECT 397.900 2127.810 398.180 2128.090 ;
        RECT 398.520 2127.810 398.800 2128.090 ;
        RECT 399.140 2127.810 399.420 2128.090 ;
        RECT 399.760 2127.810 400.040 2128.090 ;
        RECT 396.040 2127.190 396.320 2127.470 ;
        RECT 396.660 2127.190 396.940 2127.470 ;
        RECT 397.280 2127.190 397.560 2127.470 ;
        RECT 397.900 2127.190 398.180 2127.470 ;
        RECT 398.520 2127.190 398.800 2127.470 ;
        RECT 399.140 2127.190 399.420 2127.470 ;
        RECT 399.760 2127.190 400.040 2127.470 ;
        RECT 396.040 2126.570 396.320 2126.850 ;
        RECT 396.660 2126.570 396.940 2126.850 ;
        RECT 397.280 2126.570 397.560 2126.850 ;
        RECT 397.900 2126.570 398.180 2126.850 ;
        RECT 398.520 2126.570 398.800 2126.850 ;
        RECT 399.140 2126.570 399.420 2126.850 ;
        RECT 399.760 2126.570 400.040 2126.850 ;
        RECT 396.040 2125.950 396.320 2126.230 ;
        RECT 396.660 2125.950 396.940 2126.230 ;
        RECT 397.280 2125.950 397.560 2126.230 ;
        RECT 397.900 2125.950 398.180 2126.230 ;
        RECT 398.520 2125.950 398.800 2126.230 ;
        RECT 399.140 2125.950 399.420 2126.230 ;
        RECT 399.760 2125.950 400.040 2126.230 ;
        RECT 396.040 2125.330 396.320 2125.610 ;
        RECT 396.660 2125.330 396.940 2125.610 ;
        RECT 397.280 2125.330 397.560 2125.610 ;
        RECT 397.900 2125.330 398.180 2125.610 ;
        RECT 398.520 2125.330 398.800 2125.610 ;
        RECT 399.140 2125.330 399.420 2125.610 ;
        RECT 399.760 2125.330 400.040 2125.610 ;
        RECT 396.040 2124.710 396.320 2124.990 ;
        RECT 396.660 2124.710 396.940 2124.990 ;
        RECT 397.280 2124.710 397.560 2124.990 ;
        RECT 397.900 2124.710 398.180 2124.990 ;
        RECT 398.520 2124.710 398.800 2124.990 ;
        RECT 399.140 2124.710 399.420 2124.990 ;
        RECT 399.760 2124.710 400.040 2124.990 ;
        RECT 396.040 2124.090 396.320 2124.370 ;
        RECT 396.660 2124.090 396.940 2124.370 ;
        RECT 397.280 2124.090 397.560 2124.370 ;
        RECT 397.900 2124.090 398.180 2124.370 ;
        RECT 398.520 2124.090 398.800 2124.370 ;
        RECT 399.140 2124.090 399.420 2124.370 ;
        RECT 399.760 2124.090 400.040 2124.370 ;
        RECT 396.040 2123.470 396.320 2123.750 ;
        RECT 396.660 2123.470 396.940 2123.750 ;
        RECT 397.280 2123.470 397.560 2123.750 ;
        RECT 397.900 2123.470 398.180 2123.750 ;
        RECT 398.520 2123.470 398.800 2123.750 ;
        RECT 399.140 2123.470 399.420 2123.750 ;
        RECT 399.760 2123.470 400.040 2123.750 ;
        RECT 396.040 2122.850 396.320 2123.130 ;
        RECT 396.660 2122.850 396.940 2123.130 ;
        RECT 397.280 2122.850 397.560 2123.130 ;
        RECT 397.900 2122.850 398.180 2123.130 ;
        RECT 398.520 2122.850 398.800 2123.130 ;
        RECT 399.140 2122.850 399.420 2123.130 ;
        RECT 399.760 2122.850 400.040 2123.130 ;
        RECT 396.040 2122.230 396.320 2122.510 ;
        RECT 396.660 2122.230 396.940 2122.510 ;
        RECT 397.280 2122.230 397.560 2122.510 ;
        RECT 397.900 2122.230 398.180 2122.510 ;
        RECT 398.520 2122.230 398.800 2122.510 ;
        RECT 399.140 2122.230 399.420 2122.510 ;
        RECT 399.760 2122.230 400.040 2122.510 ;
        RECT 396.040 2121.610 396.320 2121.890 ;
        RECT 396.660 2121.610 396.940 2121.890 ;
        RECT 397.280 2121.610 397.560 2121.890 ;
        RECT 397.900 2121.610 398.180 2121.890 ;
        RECT 398.520 2121.610 398.800 2121.890 ;
        RECT 399.140 2121.610 399.420 2121.890 ;
        RECT 399.760 2121.610 400.040 2121.890 ;
        RECT 396.040 2120.990 396.320 2121.270 ;
        RECT 396.660 2120.990 396.940 2121.270 ;
        RECT 397.280 2120.990 397.560 2121.270 ;
        RECT 397.900 2120.990 398.180 2121.270 ;
        RECT 398.520 2120.990 398.800 2121.270 ;
        RECT 399.140 2120.990 399.420 2121.270 ;
        RECT 399.760 2120.990 400.040 2121.270 ;
        RECT 396.040 2118.440 396.320 2118.720 ;
        RECT 396.660 2118.440 396.940 2118.720 ;
        RECT 397.280 2118.440 397.560 2118.720 ;
        RECT 397.900 2118.440 398.180 2118.720 ;
        RECT 398.520 2118.440 398.800 2118.720 ;
        RECT 399.140 2118.440 399.420 2118.720 ;
        RECT 399.760 2118.440 400.040 2118.720 ;
        RECT 396.040 2117.820 396.320 2118.100 ;
        RECT 396.660 2117.820 396.940 2118.100 ;
        RECT 397.280 2117.820 397.560 2118.100 ;
        RECT 397.900 2117.820 398.180 2118.100 ;
        RECT 398.520 2117.820 398.800 2118.100 ;
        RECT 399.140 2117.820 399.420 2118.100 ;
        RECT 399.760 2117.820 400.040 2118.100 ;
        RECT 396.040 2117.200 396.320 2117.480 ;
        RECT 396.660 2117.200 396.940 2117.480 ;
        RECT 397.280 2117.200 397.560 2117.480 ;
        RECT 397.900 2117.200 398.180 2117.480 ;
        RECT 398.520 2117.200 398.800 2117.480 ;
        RECT 399.140 2117.200 399.420 2117.480 ;
        RECT 399.760 2117.200 400.040 2117.480 ;
        RECT 396.040 2116.580 396.320 2116.860 ;
        RECT 396.660 2116.580 396.940 2116.860 ;
        RECT 397.280 2116.580 397.560 2116.860 ;
        RECT 397.900 2116.580 398.180 2116.860 ;
        RECT 398.520 2116.580 398.800 2116.860 ;
        RECT 399.140 2116.580 399.420 2116.860 ;
        RECT 399.760 2116.580 400.040 2116.860 ;
        RECT 396.040 2115.960 396.320 2116.240 ;
        RECT 396.660 2115.960 396.940 2116.240 ;
        RECT 397.280 2115.960 397.560 2116.240 ;
        RECT 397.900 2115.960 398.180 2116.240 ;
        RECT 398.520 2115.960 398.800 2116.240 ;
        RECT 399.140 2115.960 399.420 2116.240 ;
        RECT 399.760 2115.960 400.040 2116.240 ;
        RECT 396.040 2115.340 396.320 2115.620 ;
        RECT 396.660 2115.340 396.940 2115.620 ;
        RECT 397.280 2115.340 397.560 2115.620 ;
        RECT 397.900 2115.340 398.180 2115.620 ;
        RECT 398.520 2115.340 398.800 2115.620 ;
        RECT 399.140 2115.340 399.420 2115.620 ;
        RECT 399.760 2115.340 400.040 2115.620 ;
        RECT 396.040 2114.720 396.320 2115.000 ;
        RECT 396.660 2114.720 396.940 2115.000 ;
        RECT 397.280 2114.720 397.560 2115.000 ;
        RECT 397.900 2114.720 398.180 2115.000 ;
        RECT 398.520 2114.720 398.800 2115.000 ;
        RECT 399.140 2114.720 399.420 2115.000 ;
        RECT 399.760 2114.720 400.040 2115.000 ;
        RECT 396.040 2114.100 396.320 2114.380 ;
        RECT 396.660 2114.100 396.940 2114.380 ;
        RECT 397.280 2114.100 397.560 2114.380 ;
        RECT 397.900 2114.100 398.180 2114.380 ;
        RECT 398.520 2114.100 398.800 2114.380 ;
        RECT 399.140 2114.100 399.420 2114.380 ;
        RECT 399.760 2114.100 400.040 2114.380 ;
        RECT 396.040 2113.480 396.320 2113.760 ;
        RECT 396.660 2113.480 396.940 2113.760 ;
        RECT 397.280 2113.480 397.560 2113.760 ;
        RECT 397.900 2113.480 398.180 2113.760 ;
        RECT 398.520 2113.480 398.800 2113.760 ;
        RECT 399.140 2113.480 399.420 2113.760 ;
        RECT 399.760 2113.480 400.040 2113.760 ;
        RECT 396.040 2112.860 396.320 2113.140 ;
        RECT 396.660 2112.860 396.940 2113.140 ;
        RECT 397.280 2112.860 397.560 2113.140 ;
        RECT 397.900 2112.860 398.180 2113.140 ;
        RECT 398.520 2112.860 398.800 2113.140 ;
        RECT 399.140 2112.860 399.420 2113.140 ;
        RECT 399.760 2112.860 400.040 2113.140 ;
        RECT 396.040 2112.240 396.320 2112.520 ;
        RECT 396.660 2112.240 396.940 2112.520 ;
        RECT 397.280 2112.240 397.560 2112.520 ;
        RECT 397.900 2112.240 398.180 2112.520 ;
        RECT 398.520 2112.240 398.800 2112.520 ;
        RECT 399.140 2112.240 399.420 2112.520 ;
        RECT 399.760 2112.240 400.040 2112.520 ;
        RECT 396.040 2111.620 396.320 2111.900 ;
        RECT 396.660 2111.620 396.940 2111.900 ;
        RECT 397.280 2111.620 397.560 2111.900 ;
        RECT 397.900 2111.620 398.180 2111.900 ;
        RECT 398.520 2111.620 398.800 2111.900 ;
        RECT 399.140 2111.620 399.420 2111.900 ;
        RECT 399.760 2111.620 400.040 2111.900 ;
        RECT 396.040 2111.000 396.320 2111.280 ;
        RECT 396.660 2111.000 396.940 2111.280 ;
        RECT 397.280 2111.000 397.560 2111.280 ;
        RECT 397.900 2111.000 398.180 2111.280 ;
        RECT 398.520 2111.000 398.800 2111.280 ;
        RECT 399.140 2111.000 399.420 2111.280 ;
        RECT 399.760 2111.000 400.040 2111.280 ;
        RECT 396.040 2110.380 396.320 2110.660 ;
        RECT 396.660 2110.380 396.940 2110.660 ;
        RECT 397.280 2110.380 397.560 2110.660 ;
        RECT 397.900 2110.380 398.180 2110.660 ;
        RECT 398.520 2110.380 398.800 2110.660 ;
        RECT 399.140 2110.380 399.420 2110.660 ;
        RECT 399.760 2110.380 400.040 2110.660 ;
        RECT 396.040 2109.760 396.320 2110.040 ;
        RECT 396.660 2109.760 396.940 2110.040 ;
        RECT 397.280 2109.760 397.560 2110.040 ;
        RECT 397.900 2109.760 398.180 2110.040 ;
        RECT 398.520 2109.760 398.800 2110.040 ;
        RECT 399.140 2109.760 399.420 2110.040 ;
        RECT 399.760 2109.760 400.040 2110.040 ;
        RECT 396.040 2109.140 396.320 2109.420 ;
        RECT 396.660 2109.140 396.940 2109.420 ;
        RECT 397.280 2109.140 397.560 2109.420 ;
        RECT 397.900 2109.140 398.180 2109.420 ;
        RECT 398.520 2109.140 398.800 2109.420 ;
        RECT 399.140 2109.140 399.420 2109.420 ;
        RECT 399.760 2109.140 400.040 2109.420 ;
        RECT 396.040 2105.420 396.320 2105.700 ;
        RECT 396.660 2105.420 396.940 2105.700 ;
        RECT 397.280 2105.420 397.560 2105.700 ;
        RECT 397.900 2105.420 398.180 2105.700 ;
        RECT 398.520 2105.420 398.800 2105.700 ;
        RECT 399.140 2105.420 399.420 2105.700 ;
        RECT 399.760 2105.420 400.040 2105.700 ;
        RECT 396.040 2104.800 396.320 2105.080 ;
        RECT 396.660 2104.800 396.940 2105.080 ;
        RECT 397.280 2104.800 397.560 2105.080 ;
        RECT 397.900 2104.800 398.180 2105.080 ;
        RECT 398.520 2104.800 398.800 2105.080 ;
        RECT 399.140 2104.800 399.420 2105.080 ;
        RECT 399.760 2104.800 400.040 2105.080 ;
        RECT 396.040 2104.180 396.320 2104.460 ;
        RECT 396.660 2104.180 396.940 2104.460 ;
        RECT 397.280 2104.180 397.560 2104.460 ;
        RECT 397.900 2104.180 398.180 2104.460 ;
        RECT 398.520 2104.180 398.800 2104.460 ;
        RECT 399.140 2104.180 399.420 2104.460 ;
        RECT 399.760 2104.180 400.040 2104.460 ;
        RECT 396.040 2103.560 396.320 2103.840 ;
        RECT 396.660 2103.560 396.940 2103.840 ;
        RECT 397.280 2103.560 397.560 2103.840 ;
        RECT 397.900 2103.560 398.180 2103.840 ;
        RECT 398.520 2103.560 398.800 2103.840 ;
        RECT 399.140 2103.560 399.420 2103.840 ;
        RECT 399.760 2103.560 400.040 2103.840 ;
        RECT 396.040 2102.940 396.320 2103.220 ;
        RECT 396.660 2102.940 396.940 2103.220 ;
        RECT 397.280 2102.940 397.560 2103.220 ;
        RECT 397.900 2102.940 398.180 2103.220 ;
        RECT 398.520 2102.940 398.800 2103.220 ;
        RECT 399.140 2102.940 399.420 2103.220 ;
        RECT 399.760 2102.940 400.040 2103.220 ;
        RECT 396.040 2102.320 396.320 2102.600 ;
        RECT 396.660 2102.320 396.940 2102.600 ;
        RECT 397.280 2102.320 397.560 2102.600 ;
        RECT 397.900 2102.320 398.180 2102.600 ;
        RECT 398.520 2102.320 398.800 2102.600 ;
        RECT 399.140 2102.320 399.420 2102.600 ;
        RECT 399.760 2102.320 400.040 2102.600 ;
        RECT 396.040 2101.700 396.320 2101.980 ;
        RECT 396.660 2101.700 396.940 2101.980 ;
        RECT 397.280 2101.700 397.560 2101.980 ;
        RECT 397.900 2101.700 398.180 2101.980 ;
        RECT 398.520 2101.700 398.800 2101.980 ;
        RECT 399.140 2101.700 399.420 2101.980 ;
        RECT 399.760 2101.700 400.040 2101.980 ;
        RECT 396.040 2101.080 396.320 2101.360 ;
        RECT 396.660 2101.080 396.940 2101.360 ;
        RECT 397.280 2101.080 397.560 2101.360 ;
        RECT 397.900 2101.080 398.180 2101.360 ;
        RECT 398.520 2101.080 398.800 2101.360 ;
        RECT 399.140 2101.080 399.420 2101.360 ;
        RECT 399.760 2101.080 400.040 2101.360 ;
        RECT 396.040 2100.460 396.320 2100.740 ;
        RECT 396.660 2100.460 396.940 2100.740 ;
        RECT 397.280 2100.460 397.560 2100.740 ;
        RECT 397.900 2100.460 398.180 2100.740 ;
        RECT 398.520 2100.460 398.800 2100.740 ;
        RECT 399.140 2100.460 399.420 2100.740 ;
        RECT 399.760 2100.460 400.040 2100.740 ;
        RECT 396.040 2099.840 396.320 2100.120 ;
        RECT 396.660 2099.840 396.940 2100.120 ;
        RECT 397.280 2099.840 397.560 2100.120 ;
        RECT 397.900 2099.840 398.180 2100.120 ;
        RECT 398.520 2099.840 398.800 2100.120 ;
        RECT 399.140 2099.840 399.420 2100.120 ;
        RECT 399.760 2099.840 400.040 2100.120 ;
        RECT 396.040 2099.220 396.320 2099.500 ;
        RECT 396.660 2099.220 396.940 2099.500 ;
        RECT 397.280 2099.220 397.560 2099.500 ;
        RECT 397.900 2099.220 398.180 2099.500 ;
        RECT 398.520 2099.220 398.800 2099.500 ;
        RECT 399.140 2099.220 399.420 2099.500 ;
        RECT 399.760 2099.220 400.040 2099.500 ;
        RECT 396.040 2098.600 396.320 2098.880 ;
        RECT 396.660 2098.600 396.940 2098.880 ;
        RECT 397.280 2098.600 397.560 2098.880 ;
        RECT 397.900 2098.600 398.180 2098.880 ;
        RECT 398.520 2098.600 398.800 2098.880 ;
        RECT 399.140 2098.600 399.420 2098.880 ;
        RECT 399.760 2098.600 400.040 2098.880 ;
        RECT 396.040 2097.980 396.320 2098.260 ;
        RECT 396.660 2097.980 396.940 2098.260 ;
        RECT 397.280 2097.980 397.560 2098.260 ;
        RECT 397.900 2097.980 398.180 2098.260 ;
        RECT 398.520 2097.980 398.800 2098.260 ;
        RECT 399.140 2097.980 399.420 2098.260 ;
        RECT 399.760 2097.980 400.040 2098.260 ;
        RECT 396.040 2097.360 396.320 2097.640 ;
        RECT 396.660 2097.360 396.940 2097.640 ;
        RECT 397.280 2097.360 397.560 2097.640 ;
        RECT 397.900 2097.360 398.180 2097.640 ;
        RECT 398.520 2097.360 398.800 2097.640 ;
        RECT 399.140 2097.360 399.420 2097.640 ;
        RECT 399.760 2097.360 400.040 2097.640 ;
        RECT 396.040 2096.740 396.320 2097.020 ;
        RECT 396.660 2096.740 396.940 2097.020 ;
        RECT 397.280 2096.740 397.560 2097.020 ;
        RECT 397.900 2096.740 398.180 2097.020 ;
        RECT 398.520 2096.740 398.800 2097.020 ;
        RECT 399.140 2096.740 399.420 2097.020 ;
        RECT 399.760 2096.740 400.040 2097.020 ;
        RECT 396.420 2064.960 396.700 2065.240 ;
        RECT 397.920 2064.960 398.200 2065.240 ;
        RECT 399.420 2064.960 399.700 2065.240 ;
        RECT 396.500 1982.830 396.780 1983.110 ;
        RECT 398.000 1982.830 398.280 1983.110 ;
        RECT 399.500 1982.830 399.780 1983.110 ;
        RECT 396.000 1961.865 396.280 1962.145 ;
        RECT 397.500 1961.865 397.780 1962.145 ;
        RECT 399.000 1961.865 399.280 1962.145 ;
        RECT 396.000 1960.865 396.280 1961.145 ;
        RECT 397.500 1960.865 397.780 1961.145 ;
        RECT 399.000 1960.865 399.280 1961.145 ;
        RECT 396.500 1947.830 396.780 1948.110 ;
        RECT 398.000 1947.830 398.280 1948.110 ;
        RECT 399.500 1947.830 399.780 1948.110 ;
        RECT 396.500 1912.830 396.780 1913.110 ;
        RECT 398.000 1912.830 398.280 1913.110 ;
        RECT 399.500 1912.830 399.780 1913.110 ;
        RECT 396.420 1859.960 396.700 1860.240 ;
        RECT 397.920 1859.960 398.200 1860.240 ;
        RECT 399.420 1859.960 399.700 1860.240 ;
        RECT 396.000 1781.865 396.280 1782.145 ;
        RECT 397.500 1781.865 397.780 1782.145 ;
        RECT 399.000 1781.865 399.280 1782.145 ;
        RECT 396.000 1780.865 396.280 1781.145 ;
        RECT 397.500 1780.865 397.780 1781.145 ;
        RECT 399.000 1780.865 399.280 1781.145 ;
        RECT 396.500 1777.830 396.780 1778.110 ;
        RECT 398.000 1777.830 398.280 1778.110 ;
        RECT 399.500 1777.830 399.780 1778.110 ;
        RECT 396.500 1742.830 396.780 1743.110 ;
        RECT 398.000 1742.830 398.280 1743.110 ;
        RECT 399.500 1742.830 399.780 1743.110 ;
        RECT 396.500 1707.830 396.780 1708.110 ;
        RECT 398.000 1707.830 398.280 1708.110 ;
        RECT 399.500 1707.830 399.780 1708.110 ;
        RECT 3490.220 4611.890 3490.500 4612.170 ;
        RECT 3491.720 4611.890 3492.000 4612.170 ;
        RECT 3493.220 4611.890 3493.500 4612.170 ;
        RECT 3490.220 4576.890 3490.500 4577.170 ;
        RECT 3491.720 4576.890 3492.000 4577.170 ;
        RECT 3493.220 4576.890 3493.500 4577.170 ;
        RECT 3490.220 4541.890 3490.500 4542.170 ;
        RECT 3491.720 4541.890 3492.000 4542.170 ;
        RECT 3493.220 4541.890 3493.500 4542.170 ;
        RECT 3490.720 4481.865 3491.000 4482.145 ;
        RECT 3492.220 4481.865 3492.500 4482.145 ;
        RECT 3493.720 4481.865 3494.000 4482.145 ;
        RECT 3490.720 4480.865 3491.000 4481.145 ;
        RECT 3492.220 4480.865 3492.500 4481.145 ;
        RECT 3493.720 4480.865 3494.000 4481.145 ;
        RECT 3490.300 4459.760 3490.580 4460.040 ;
        RECT 3491.800 4459.760 3492.080 4460.040 ;
        RECT 3493.300 4459.760 3493.580 4460.040 ;
        RECT 3490.720 4301.865 3491.000 4302.145 ;
        RECT 3492.220 4301.865 3492.500 4302.145 ;
        RECT 3493.720 4301.865 3494.000 4302.145 ;
        RECT 3490.720 4300.865 3491.000 4301.145 ;
        RECT 3492.220 4300.865 3492.500 4301.145 ;
        RECT 3493.720 4300.865 3494.000 4301.145 ;
        RECT 3490.220 4181.890 3490.500 4182.170 ;
        RECT 3491.720 4181.890 3492.000 4182.170 ;
        RECT 3493.220 4181.890 3493.500 4182.170 ;
        RECT 3490.220 4146.890 3490.500 4147.170 ;
        RECT 3491.720 4146.890 3492.000 4147.170 ;
        RECT 3493.220 4146.890 3493.500 4147.170 ;
        RECT 3490.720 4121.865 3491.000 4122.145 ;
        RECT 3492.220 4121.865 3492.500 4122.145 ;
        RECT 3493.720 4121.865 3494.000 4122.145 ;
        RECT 3490.720 4120.865 3491.000 4121.145 ;
        RECT 3492.220 4120.865 3492.500 4121.145 ;
        RECT 3493.720 4120.865 3494.000 4121.145 ;
        RECT 3490.220 4111.890 3490.500 4112.170 ;
        RECT 3491.720 4111.890 3492.000 4112.170 ;
        RECT 3493.220 4111.890 3493.500 4112.170 ;
        RECT 3490.300 4029.760 3490.580 4030.040 ;
        RECT 3491.800 4029.760 3492.080 4030.040 ;
        RECT 3493.300 4029.760 3493.580 4030.040 ;
        RECT 3490.720 3761.865 3491.000 3762.145 ;
        RECT 3492.220 3761.865 3492.500 3762.145 ;
        RECT 3493.720 3761.865 3494.000 3762.145 ;
        RECT 3490.720 3760.865 3491.000 3761.145 ;
        RECT 3492.220 3760.865 3492.500 3761.145 ;
        RECT 3493.720 3760.865 3494.000 3761.145 ;
        RECT 3490.220 3751.890 3490.500 3752.170 ;
        RECT 3491.720 3751.890 3492.000 3752.170 ;
        RECT 3493.220 3751.890 3493.500 3752.170 ;
        RECT 3490.220 3716.890 3490.500 3717.170 ;
        RECT 3491.720 3716.890 3492.000 3717.170 ;
        RECT 3493.220 3716.890 3493.500 3717.170 ;
        RECT 3490.220 3681.890 3490.500 3682.170 ;
        RECT 3491.720 3681.890 3492.000 3682.170 ;
        RECT 3493.220 3681.890 3493.500 3682.170 ;
        RECT 3490.300 3599.760 3490.580 3600.040 ;
        RECT 3491.800 3599.760 3492.080 3600.040 ;
        RECT 3493.300 3599.760 3493.580 3600.040 ;
        RECT 3490.720 3581.865 3491.000 3582.145 ;
        RECT 3492.220 3581.865 3492.500 3582.145 ;
        RECT 3493.720 3581.865 3494.000 3582.145 ;
        RECT 3490.720 3580.865 3491.000 3581.145 ;
        RECT 3492.220 3580.865 3492.500 3581.145 ;
        RECT 3493.720 3580.865 3494.000 3581.145 ;
        RECT 3490.220 3536.890 3490.500 3537.170 ;
        RECT 3491.720 3536.890 3492.000 3537.170 ;
        RECT 3493.220 3536.890 3493.500 3537.170 ;
        RECT 3490.220 3501.890 3490.500 3502.170 ;
        RECT 3491.720 3501.890 3492.000 3502.170 ;
        RECT 3493.220 3501.890 3493.500 3502.170 ;
        RECT 3490.220 3466.890 3490.500 3467.170 ;
        RECT 3491.720 3466.890 3492.000 3467.170 ;
        RECT 3493.220 3466.890 3493.500 3467.170 ;
        RECT 3490.720 3401.865 3491.000 3402.145 ;
        RECT 3492.220 3401.865 3492.500 3402.145 ;
        RECT 3493.720 3401.865 3494.000 3402.145 ;
        RECT 3490.720 3400.865 3491.000 3401.145 ;
        RECT 3492.220 3400.865 3492.500 3401.145 ;
        RECT 3493.720 3400.865 3494.000 3401.145 ;
        RECT 3490.300 3384.760 3490.580 3385.040 ;
        RECT 3491.800 3384.760 3492.080 3385.040 ;
        RECT 3493.300 3384.760 3493.580 3385.040 ;
        RECT 3490.220 3321.890 3490.500 3322.170 ;
        RECT 3491.720 3321.890 3492.000 3322.170 ;
        RECT 3493.220 3321.890 3493.500 3322.170 ;
        RECT 3490.220 3286.890 3490.500 3287.170 ;
        RECT 3491.720 3286.890 3492.000 3287.170 ;
        RECT 3493.220 3286.890 3493.500 3287.170 ;
        RECT 3490.220 3251.890 3490.500 3252.170 ;
        RECT 3491.720 3251.890 3492.000 3252.170 ;
        RECT 3493.220 3251.890 3493.500 3252.170 ;
        RECT 3490.720 3221.865 3491.000 3222.145 ;
        RECT 3492.220 3221.865 3492.500 3222.145 ;
        RECT 3493.720 3221.865 3494.000 3222.145 ;
        RECT 3490.720 3220.865 3491.000 3221.145 ;
        RECT 3492.220 3220.865 3492.500 3221.145 ;
        RECT 3493.720 3220.865 3494.000 3221.145 ;
        RECT 3490.300 3169.760 3490.580 3170.040 ;
        RECT 3491.800 3169.760 3492.080 3170.040 ;
        RECT 3493.300 3169.760 3493.580 3170.040 ;
        RECT 3490.220 3106.890 3490.500 3107.170 ;
        RECT 3491.720 3106.890 3492.000 3107.170 ;
        RECT 3493.220 3106.890 3493.500 3107.170 ;
        RECT 3490.220 3071.890 3490.500 3072.170 ;
        RECT 3491.720 3071.890 3492.000 3072.170 ;
        RECT 3493.220 3071.890 3493.500 3072.170 ;
        RECT 3490.720 3041.865 3491.000 3042.145 ;
        RECT 3492.220 3041.865 3492.500 3042.145 ;
        RECT 3493.720 3041.865 3494.000 3042.145 ;
        RECT 3490.720 3040.865 3491.000 3041.145 ;
        RECT 3492.220 3040.865 3492.500 3041.145 ;
        RECT 3493.720 3040.865 3494.000 3041.145 ;
        RECT 3490.220 3036.890 3490.500 3037.170 ;
        RECT 3491.720 3036.890 3492.000 3037.170 ;
        RECT 3493.220 3036.890 3493.500 3037.170 ;
        RECT 3490.300 2954.760 3490.580 2955.040 ;
        RECT 3491.800 2954.760 3492.080 2955.040 ;
        RECT 3493.300 2954.760 3493.580 2955.040 ;
        RECT 3490.220 2891.890 3490.500 2892.170 ;
        RECT 3491.720 2891.890 3492.000 2892.170 ;
        RECT 3493.220 2891.890 3493.500 2892.170 ;
        RECT 3490.720 2861.865 3491.000 2862.145 ;
        RECT 3492.220 2861.865 3492.500 2862.145 ;
        RECT 3493.720 2861.865 3494.000 2862.145 ;
        RECT 3490.720 2860.865 3491.000 2861.145 ;
        RECT 3492.220 2860.865 3492.500 2861.145 ;
        RECT 3493.720 2860.865 3494.000 2861.145 ;
        RECT 3490.220 2856.890 3490.500 2857.170 ;
        RECT 3491.720 2856.890 3492.000 2857.170 ;
        RECT 3493.220 2856.890 3493.500 2857.170 ;
        RECT 3490.220 2821.890 3490.500 2822.170 ;
        RECT 3491.720 2821.890 3492.000 2822.170 ;
        RECT 3493.220 2821.890 3493.500 2822.170 ;
        RECT 3490.300 2739.760 3490.580 2740.040 ;
        RECT 3491.800 2739.760 3492.080 2740.040 ;
        RECT 3493.300 2739.760 3493.580 2740.040 ;
        RECT 3490.720 2681.865 3491.000 2682.145 ;
        RECT 3492.220 2681.865 3492.500 2682.145 ;
        RECT 3493.720 2681.865 3494.000 2682.145 ;
        RECT 3490.720 2680.865 3491.000 2681.145 ;
        RECT 3492.220 2680.865 3492.500 2681.145 ;
        RECT 3493.720 2680.865 3494.000 2681.145 ;
        RECT 3490.220 2676.890 3490.500 2677.170 ;
        RECT 3491.720 2676.890 3492.000 2677.170 ;
        RECT 3493.220 2676.890 3493.500 2677.170 ;
        RECT 3490.220 2641.890 3490.500 2642.170 ;
        RECT 3491.720 2641.890 3492.000 2642.170 ;
        RECT 3493.220 2641.890 3493.500 2642.170 ;
        RECT 3490.220 2606.890 3490.500 2607.170 ;
        RECT 3491.720 2606.890 3492.000 2607.170 ;
        RECT 3493.220 2606.890 3493.500 2607.170 ;
        RECT 3490.300 2524.760 3490.580 2525.040 ;
        RECT 3491.800 2524.760 3492.080 2525.040 ;
        RECT 3493.300 2524.760 3493.580 2525.040 ;
        RECT 3490.720 2501.865 3491.000 2502.145 ;
        RECT 3492.220 2501.865 3492.500 2502.145 ;
        RECT 3493.720 2501.865 3494.000 2502.145 ;
        RECT 3490.720 2500.865 3491.000 2501.145 ;
        RECT 3492.220 2500.865 3492.500 2501.145 ;
        RECT 3493.720 2500.865 3494.000 2501.145 ;
        RECT 3490.720 2321.865 3491.000 2322.145 ;
        RECT 3492.220 2321.865 3492.500 2322.145 ;
        RECT 3493.720 2321.865 3494.000 2322.145 ;
        RECT 3490.720 2320.865 3491.000 2321.145 ;
        RECT 3492.220 2320.865 3492.500 2321.145 ;
        RECT 3493.720 2320.865 3494.000 2321.145 ;
        RECT 3489.960 2267.980 3490.240 2268.260 ;
        RECT 3490.580 2267.980 3490.860 2268.260 ;
        RECT 3491.200 2267.980 3491.480 2268.260 ;
        RECT 3491.820 2267.980 3492.100 2268.260 ;
        RECT 3492.440 2267.980 3492.720 2268.260 ;
        RECT 3493.060 2267.980 3493.340 2268.260 ;
        RECT 3493.680 2267.980 3493.960 2268.260 ;
        RECT 3489.960 2267.360 3490.240 2267.640 ;
        RECT 3490.580 2267.360 3490.860 2267.640 ;
        RECT 3491.200 2267.360 3491.480 2267.640 ;
        RECT 3491.820 2267.360 3492.100 2267.640 ;
        RECT 3492.440 2267.360 3492.720 2267.640 ;
        RECT 3493.060 2267.360 3493.340 2267.640 ;
        RECT 3493.680 2267.360 3493.960 2267.640 ;
        RECT 3489.960 2266.740 3490.240 2267.020 ;
        RECT 3490.580 2266.740 3490.860 2267.020 ;
        RECT 3491.200 2266.740 3491.480 2267.020 ;
        RECT 3491.820 2266.740 3492.100 2267.020 ;
        RECT 3492.440 2266.740 3492.720 2267.020 ;
        RECT 3493.060 2266.740 3493.340 2267.020 ;
        RECT 3493.680 2266.740 3493.960 2267.020 ;
        RECT 3489.960 2266.120 3490.240 2266.400 ;
        RECT 3490.580 2266.120 3490.860 2266.400 ;
        RECT 3491.200 2266.120 3491.480 2266.400 ;
        RECT 3491.820 2266.120 3492.100 2266.400 ;
        RECT 3492.440 2266.120 3492.720 2266.400 ;
        RECT 3493.060 2266.120 3493.340 2266.400 ;
        RECT 3493.680 2266.120 3493.960 2266.400 ;
        RECT 3489.960 2265.500 3490.240 2265.780 ;
        RECT 3490.580 2265.500 3490.860 2265.780 ;
        RECT 3491.200 2265.500 3491.480 2265.780 ;
        RECT 3491.820 2265.500 3492.100 2265.780 ;
        RECT 3492.440 2265.500 3492.720 2265.780 ;
        RECT 3493.060 2265.500 3493.340 2265.780 ;
        RECT 3493.680 2265.500 3493.960 2265.780 ;
        RECT 3489.960 2264.880 3490.240 2265.160 ;
        RECT 3490.580 2264.880 3490.860 2265.160 ;
        RECT 3491.200 2264.880 3491.480 2265.160 ;
        RECT 3491.820 2264.880 3492.100 2265.160 ;
        RECT 3492.440 2264.880 3492.720 2265.160 ;
        RECT 3493.060 2264.880 3493.340 2265.160 ;
        RECT 3493.680 2264.880 3493.960 2265.160 ;
        RECT 3489.960 2264.260 3490.240 2264.540 ;
        RECT 3490.580 2264.260 3490.860 2264.540 ;
        RECT 3491.200 2264.260 3491.480 2264.540 ;
        RECT 3491.820 2264.260 3492.100 2264.540 ;
        RECT 3492.440 2264.260 3492.720 2264.540 ;
        RECT 3493.060 2264.260 3493.340 2264.540 ;
        RECT 3493.680 2264.260 3493.960 2264.540 ;
        RECT 3489.960 2263.640 3490.240 2263.920 ;
        RECT 3490.580 2263.640 3490.860 2263.920 ;
        RECT 3491.200 2263.640 3491.480 2263.920 ;
        RECT 3491.820 2263.640 3492.100 2263.920 ;
        RECT 3492.440 2263.640 3492.720 2263.920 ;
        RECT 3493.060 2263.640 3493.340 2263.920 ;
        RECT 3493.680 2263.640 3493.960 2263.920 ;
        RECT 3489.960 2263.020 3490.240 2263.300 ;
        RECT 3490.580 2263.020 3490.860 2263.300 ;
        RECT 3491.200 2263.020 3491.480 2263.300 ;
        RECT 3491.820 2263.020 3492.100 2263.300 ;
        RECT 3492.440 2263.020 3492.720 2263.300 ;
        RECT 3493.060 2263.020 3493.340 2263.300 ;
        RECT 3493.680 2263.020 3493.960 2263.300 ;
        RECT 3489.960 2262.400 3490.240 2262.680 ;
        RECT 3490.580 2262.400 3490.860 2262.680 ;
        RECT 3491.200 2262.400 3491.480 2262.680 ;
        RECT 3491.820 2262.400 3492.100 2262.680 ;
        RECT 3492.440 2262.400 3492.720 2262.680 ;
        RECT 3493.060 2262.400 3493.340 2262.680 ;
        RECT 3493.680 2262.400 3493.960 2262.680 ;
        RECT 3489.960 2261.780 3490.240 2262.060 ;
        RECT 3490.580 2261.780 3490.860 2262.060 ;
        RECT 3491.200 2261.780 3491.480 2262.060 ;
        RECT 3491.820 2261.780 3492.100 2262.060 ;
        RECT 3492.440 2261.780 3492.720 2262.060 ;
        RECT 3493.060 2261.780 3493.340 2262.060 ;
        RECT 3493.680 2261.780 3493.960 2262.060 ;
        RECT 3489.960 2261.160 3490.240 2261.440 ;
        RECT 3490.580 2261.160 3490.860 2261.440 ;
        RECT 3491.200 2261.160 3491.480 2261.440 ;
        RECT 3491.820 2261.160 3492.100 2261.440 ;
        RECT 3492.440 2261.160 3492.720 2261.440 ;
        RECT 3493.060 2261.160 3493.340 2261.440 ;
        RECT 3493.680 2261.160 3493.960 2261.440 ;
        RECT 3489.960 2260.540 3490.240 2260.820 ;
        RECT 3490.580 2260.540 3490.860 2260.820 ;
        RECT 3491.200 2260.540 3491.480 2260.820 ;
        RECT 3491.820 2260.540 3492.100 2260.820 ;
        RECT 3492.440 2260.540 3492.720 2260.820 ;
        RECT 3493.060 2260.540 3493.340 2260.820 ;
        RECT 3493.680 2260.540 3493.960 2260.820 ;
        RECT 3489.960 2259.920 3490.240 2260.200 ;
        RECT 3490.580 2259.920 3490.860 2260.200 ;
        RECT 3491.200 2259.920 3491.480 2260.200 ;
        RECT 3491.820 2259.920 3492.100 2260.200 ;
        RECT 3492.440 2259.920 3492.720 2260.200 ;
        RECT 3493.060 2259.920 3493.340 2260.200 ;
        RECT 3493.680 2259.920 3493.960 2260.200 ;
        RECT 3489.960 2259.300 3490.240 2259.580 ;
        RECT 3490.580 2259.300 3490.860 2259.580 ;
        RECT 3491.200 2259.300 3491.480 2259.580 ;
        RECT 3491.820 2259.300 3492.100 2259.580 ;
        RECT 3492.440 2259.300 3492.720 2259.580 ;
        RECT 3493.060 2259.300 3493.340 2259.580 ;
        RECT 3493.680 2259.300 3493.960 2259.580 ;
        RECT 3489.960 2255.580 3490.240 2255.860 ;
        RECT 3490.580 2255.580 3490.860 2255.860 ;
        RECT 3491.200 2255.580 3491.480 2255.860 ;
        RECT 3491.820 2255.580 3492.100 2255.860 ;
        RECT 3492.440 2255.580 3492.720 2255.860 ;
        RECT 3493.060 2255.580 3493.340 2255.860 ;
        RECT 3493.680 2255.580 3493.960 2255.860 ;
        RECT 3489.960 2254.960 3490.240 2255.240 ;
        RECT 3490.580 2254.960 3490.860 2255.240 ;
        RECT 3491.200 2254.960 3491.480 2255.240 ;
        RECT 3491.820 2254.960 3492.100 2255.240 ;
        RECT 3492.440 2254.960 3492.720 2255.240 ;
        RECT 3493.060 2254.960 3493.340 2255.240 ;
        RECT 3493.680 2254.960 3493.960 2255.240 ;
        RECT 3489.960 2254.340 3490.240 2254.620 ;
        RECT 3490.580 2254.340 3490.860 2254.620 ;
        RECT 3491.200 2254.340 3491.480 2254.620 ;
        RECT 3491.820 2254.340 3492.100 2254.620 ;
        RECT 3492.440 2254.340 3492.720 2254.620 ;
        RECT 3493.060 2254.340 3493.340 2254.620 ;
        RECT 3493.680 2254.340 3493.960 2254.620 ;
        RECT 3489.960 2253.720 3490.240 2254.000 ;
        RECT 3490.580 2253.720 3490.860 2254.000 ;
        RECT 3491.200 2253.720 3491.480 2254.000 ;
        RECT 3491.820 2253.720 3492.100 2254.000 ;
        RECT 3492.440 2253.720 3492.720 2254.000 ;
        RECT 3493.060 2253.720 3493.340 2254.000 ;
        RECT 3493.680 2253.720 3493.960 2254.000 ;
        RECT 3489.960 2253.100 3490.240 2253.380 ;
        RECT 3490.580 2253.100 3490.860 2253.380 ;
        RECT 3491.200 2253.100 3491.480 2253.380 ;
        RECT 3491.820 2253.100 3492.100 2253.380 ;
        RECT 3492.440 2253.100 3492.720 2253.380 ;
        RECT 3493.060 2253.100 3493.340 2253.380 ;
        RECT 3493.680 2253.100 3493.960 2253.380 ;
        RECT 3489.960 2252.480 3490.240 2252.760 ;
        RECT 3490.580 2252.480 3490.860 2252.760 ;
        RECT 3491.200 2252.480 3491.480 2252.760 ;
        RECT 3491.820 2252.480 3492.100 2252.760 ;
        RECT 3492.440 2252.480 3492.720 2252.760 ;
        RECT 3493.060 2252.480 3493.340 2252.760 ;
        RECT 3493.680 2252.480 3493.960 2252.760 ;
        RECT 3489.960 2251.860 3490.240 2252.140 ;
        RECT 3490.580 2251.860 3490.860 2252.140 ;
        RECT 3491.200 2251.860 3491.480 2252.140 ;
        RECT 3491.820 2251.860 3492.100 2252.140 ;
        RECT 3492.440 2251.860 3492.720 2252.140 ;
        RECT 3493.060 2251.860 3493.340 2252.140 ;
        RECT 3493.680 2251.860 3493.960 2252.140 ;
        RECT 3489.960 2251.240 3490.240 2251.520 ;
        RECT 3490.580 2251.240 3490.860 2251.520 ;
        RECT 3491.200 2251.240 3491.480 2251.520 ;
        RECT 3491.820 2251.240 3492.100 2251.520 ;
        RECT 3492.440 2251.240 3492.720 2251.520 ;
        RECT 3493.060 2251.240 3493.340 2251.520 ;
        RECT 3493.680 2251.240 3493.960 2251.520 ;
        RECT 3489.960 2250.620 3490.240 2250.900 ;
        RECT 3490.580 2250.620 3490.860 2250.900 ;
        RECT 3491.200 2250.620 3491.480 2250.900 ;
        RECT 3491.820 2250.620 3492.100 2250.900 ;
        RECT 3492.440 2250.620 3492.720 2250.900 ;
        RECT 3493.060 2250.620 3493.340 2250.900 ;
        RECT 3493.680 2250.620 3493.960 2250.900 ;
        RECT 3489.960 2250.000 3490.240 2250.280 ;
        RECT 3490.580 2250.000 3490.860 2250.280 ;
        RECT 3491.200 2250.000 3491.480 2250.280 ;
        RECT 3491.820 2250.000 3492.100 2250.280 ;
        RECT 3492.440 2250.000 3492.720 2250.280 ;
        RECT 3493.060 2250.000 3493.340 2250.280 ;
        RECT 3493.680 2250.000 3493.960 2250.280 ;
        RECT 3489.960 2249.380 3490.240 2249.660 ;
        RECT 3490.580 2249.380 3490.860 2249.660 ;
        RECT 3491.200 2249.380 3491.480 2249.660 ;
        RECT 3491.820 2249.380 3492.100 2249.660 ;
        RECT 3492.440 2249.380 3492.720 2249.660 ;
        RECT 3493.060 2249.380 3493.340 2249.660 ;
        RECT 3493.680 2249.380 3493.960 2249.660 ;
        RECT 3489.960 2248.760 3490.240 2249.040 ;
        RECT 3490.580 2248.760 3490.860 2249.040 ;
        RECT 3491.200 2248.760 3491.480 2249.040 ;
        RECT 3491.820 2248.760 3492.100 2249.040 ;
        RECT 3492.440 2248.760 3492.720 2249.040 ;
        RECT 3493.060 2248.760 3493.340 2249.040 ;
        RECT 3493.680 2248.760 3493.960 2249.040 ;
        RECT 3489.960 2248.140 3490.240 2248.420 ;
        RECT 3490.580 2248.140 3490.860 2248.420 ;
        RECT 3491.200 2248.140 3491.480 2248.420 ;
        RECT 3491.820 2248.140 3492.100 2248.420 ;
        RECT 3492.440 2248.140 3492.720 2248.420 ;
        RECT 3493.060 2248.140 3493.340 2248.420 ;
        RECT 3493.680 2248.140 3493.960 2248.420 ;
        RECT 3489.960 2247.520 3490.240 2247.800 ;
        RECT 3490.580 2247.520 3490.860 2247.800 ;
        RECT 3491.200 2247.520 3491.480 2247.800 ;
        RECT 3491.820 2247.520 3492.100 2247.800 ;
        RECT 3492.440 2247.520 3492.720 2247.800 ;
        RECT 3493.060 2247.520 3493.340 2247.800 ;
        RECT 3493.680 2247.520 3493.960 2247.800 ;
        RECT 3489.960 2246.900 3490.240 2247.180 ;
        RECT 3490.580 2246.900 3490.860 2247.180 ;
        RECT 3491.200 2246.900 3491.480 2247.180 ;
        RECT 3491.820 2246.900 3492.100 2247.180 ;
        RECT 3492.440 2246.900 3492.720 2247.180 ;
        RECT 3493.060 2246.900 3493.340 2247.180 ;
        RECT 3493.680 2246.900 3493.960 2247.180 ;
        RECT 3489.960 2246.280 3490.240 2246.560 ;
        RECT 3490.580 2246.280 3490.860 2246.560 ;
        RECT 3491.200 2246.280 3491.480 2246.560 ;
        RECT 3491.820 2246.280 3492.100 2246.560 ;
        RECT 3492.440 2246.280 3492.720 2246.560 ;
        RECT 3493.060 2246.280 3493.340 2246.560 ;
        RECT 3493.680 2246.280 3493.960 2246.560 ;
        RECT 3489.960 2243.730 3490.240 2244.010 ;
        RECT 3490.580 2243.730 3490.860 2244.010 ;
        RECT 3491.200 2243.730 3491.480 2244.010 ;
        RECT 3491.820 2243.730 3492.100 2244.010 ;
        RECT 3492.440 2243.730 3492.720 2244.010 ;
        RECT 3493.060 2243.730 3493.340 2244.010 ;
        RECT 3493.680 2243.730 3493.960 2244.010 ;
        RECT 3489.960 2243.110 3490.240 2243.390 ;
        RECT 3490.580 2243.110 3490.860 2243.390 ;
        RECT 3491.200 2243.110 3491.480 2243.390 ;
        RECT 3491.820 2243.110 3492.100 2243.390 ;
        RECT 3492.440 2243.110 3492.720 2243.390 ;
        RECT 3493.060 2243.110 3493.340 2243.390 ;
        RECT 3493.680 2243.110 3493.960 2243.390 ;
        RECT 3489.960 2242.490 3490.240 2242.770 ;
        RECT 3490.580 2242.490 3490.860 2242.770 ;
        RECT 3491.200 2242.490 3491.480 2242.770 ;
        RECT 3491.820 2242.490 3492.100 2242.770 ;
        RECT 3492.440 2242.490 3492.720 2242.770 ;
        RECT 3493.060 2242.490 3493.340 2242.770 ;
        RECT 3493.680 2242.490 3493.960 2242.770 ;
        RECT 3489.960 2241.870 3490.240 2242.150 ;
        RECT 3490.580 2241.870 3490.860 2242.150 ;
        RECT 3491.200 2241.870 3491.480 2242.150 ;
        RECT 3491.820 2241.870 3492.100 2242.150 ;
        RECT 3492.440 2241.870 3492.720 2242.150 ;
        RECT 3493.060 2241.870 3493.340 2242.150 ;
        RECT 3493.680 2241.870 3493.960 2242.150 ;
        RECT 3489.960 2241.250 3490.240 2241.530 ;
        RECT 3490.580 2241.250 3490.860 2241.530 ;
        RECT 3491.200 2241.250 3491.480 2241.530 ;
        RECT 3491.820 2241.250 3492.100 2241.530 ;
        RECT 3492.440 2241.250 3492.720 2241.530 ;
        RECT 3493.060 2241.250 3493.340 2241.530 ;
        RECT 3493.680 2241.250 3493.960 2241.530 ;
        RECT 3489.960 2240.630 3490.240 2240.910 ;
        RECT 3490.580 2240.630 3490.860 2240.910 ;
        RECT 3491.200 2240.630 3491.480 2240.910 ;
        RECT 3491.820 2240.630 3492.100 2240.910 ;
        RECT 3492.440 2240.630 3492.720 2240.910 ;
        RECT 3493.060 2240.630 3493.340 2240.910 ;
        RECT 3493.680 2240.630 3493.960 2240.910 ;
        RECT 3489.960 2240.010 3490.240 2240.290 ;
        RECT 3490.580 2240.010 3490.860 2240.290 ;
        RECT 3491.200 2240.010 3491.480 2240.290 ;
        RECT 3491.820 2240.010 3492.100 2240.290 ;
        RECT 3492.440 2240.010 3492.720 2240.290 ;
        RECT 3493.060 2240.010 3493.340 2240.290 ;
        RECT 3493.680 2240.010 3493.960 2240.290 ;
        RECT 3489.960 2239.390 3490.240 2239.670 ;
        RECT 3490.580 2239.390 3490.860 2239.670 ;
        RECT 3491.200 2239.390 3491.480 2239.670 ;
        RECT 3491.820 2239.390 3492.100 2239.670 ;
        RECT 3492.440 2239.390 3492.720 2239.670 ;
        RECT 3493.060 2239.390 3493.340 2239.670 ;
        RECT 3493.680 2239.390 3493.960 2239.670 ;
        RECT 3489.960 2238.770 3490.240 2239.050 ;
        RECT 3490.580 2238.770 3490.860 2239.050 ;
        RECT 3491.200 2238.770 3491.480 2239.050 ;
        RECT 3491.820 2238.770 3492.100 2239.050 ;
        RECT 3492.440 2238.770 3492.720 2239.050 ;
        RECT 3493.060 2238.770 3493.340 2239.050 ;
        RECT 3493.680 2238.770 3493.960 2239.050 ;
        RECT 3489.960 2238.150 3490.240 2238.430 ;
        RECT 3490.580 2238.150 3490.860 2238.430 ;
        RECT 3491.200 2238.150 3491.480 2238.430 ;
        RECT 3491.820 2238.150 3492.100 2238.430 ;
        RECT 3492.440 2238.150 3492.720 2238.430 ;
        RECT 3493.060 2238.150 3493.340 2238.430 ;
        RECT 3493.680 2238.150 3493.960 2238.430 ;
        RECT 3489.960 2237.530 3490.240 2237.810 ;
        RECT 3490.580 2237.530 3490.860 2237.810 ;
        RECT 3491.200 2237.530 3491.480 2237.810 ;
        RECT 3491.820 2237.530 3492.100 2237.810 ;
        RECT 3492.440 2237.530 3492.720 2237.810 ;
        RECT 3493.060 2237.530 3493.340 2237.810 ;
        RECT 3493.680 2237.530 3493.960 2237.810 ;
        RECT 3489.960 2236.910 3490.240 2237.190 ;
        RECT 3490.580 2236.910 3490.860 2237.190 ;
        RECT 3491.200 2236.910 3491.480 2237.190 ;
        RECT 3491.820 2236.910 3492.100 2237.190 ;
        RECT 3492.440 2236.910 3492.720 2237.190 ;
        RECT 3493.060 2236.910 3493.340 2237.190 ;
        RECT 3493.680 2236.910 3493.960 2237.190 ;
        RECT 3489.960 2236.290 3490.240 2236.570 ;
        RECT 3490.580 2236.290 3490.860 2236.570 ;
        RECT 3491.200 2236.290 3491.480 2236.570 ;
        RECT 3491.820 2236.290 3492.100 2236.570 ;
        RECT 3492.440 2236.290 3492.720 2236.570 ;
        RECT 3493.060 2236.290 3493.340 2236.570 ;
        RECT 3493.680 2236.290 3493.960 2236.570 ;
        RECT 3489.960 2235.670 3490.240 2235.950 ;
        RECT 3490.580 2235.670 3490.860 2235.950 ;
        RECT 3491.200 2235.670 3491.480 2235.950 ;
        RECT 3491.820 2235.670 3492.100 2235.950 ;
        RECT 3492.440 2235.670 3492.720 2235.950 ;
        RECT 3493.060 2235.670 3493.340 2235.950 ;
        RECT 3493.680 2235.670 3493.960 2235.950 ;
        RECT 3489.960 2235.050 3490.240 2235.330 ;
        RECT 3490.580 2235.050 3490.860 2235.330 ;
        RECT 3491.200 2235.050 3491.480 2235.330 ;
        RECT 3491.820 2235.050 3492.100 2235.330 ;
        RECT 3492.440 2235.050 3492.720 2235.330 ;
        RECT 3493.060 2235.050 3493.340 2235.330 ;
        RECT 3493.680 2235.050 3493.960 2235.330 ;
        RECT 3489.960 2234.430 3490.240 2234.710 ;
        RECT 3490.580 2234.430 3490.860 2234.710 ;
        RECT 3491.200 2234.430 3491.480 2234.710 ;
        RECT 3491.820 2234.430 3492.100 2234.710 ;
        RECT 3492.440 2234.430 3492.720 2234.710 ;
        RECT 3493.060 2234.430 3493.340 2234.710 ;
        RECT 3493.680 2234.430 3493.960 2234.710 ;
        RECT 3489.960 2230.200 3490.240 2230.480 ;
        RECT 3490.580 2230.200 3490.860 2230.480 ;
        RECT 3491.200 2230.200 3491.480 2230.480 ;
        RECT 3491.820 2230.200 3492.100 2230.480 ;
        RECT 3492.440 2230.200 3492.720 2230.480 ;
        RECT 3493.060 2230.200 3493.340 2230.480 ;
        RECT 3493.680 2230.200 3493.960 2230.480 ;
        RECT 3489.960 2229.580 3490.240 2229.860 ;
        RECT 3490.580 2229.580 3490.860 2229.860 ;
        RECT 3491.200 2229.580 3491.480 2229.860 ;
        RECT 3491.820 2229.580 3492.100 2229.860 ;
        RECT 3492.440 2229.580 3492.720 2229.860 ;
        RECT 3493.060 2229.580 3493.340 2229.860 ;
        RECT 3493.680 2229.580 3493.960 2229.860 ;
        RECT 3489.960 2228.960 3490.240 2229.240 ;
        RECT 3490.580 2228.960 3490.860 2229.240 ;
        RECT 3491.200 2228.960 3491.480 2229.240 ;
        RECT 3491.820 2228.960 3492.100 2229.240 ;
        RECT 3492.440 2228.960 3492.720 2229.240 ;
        RECT 3493.060 2228.960 3493.340 2229.240 ;
        RECT 3493.680 2228.960 3493.960 2229.240 ;
        RECT 3489.960 2228.340 3490.240 2228.620 ;
        RECT 3490.580 2228.340 3490.860 2228.620 ;
        RECT 3491.200 2228.340 3491.480 2228.620 ;
        RECT 3491.820 2228.340 3492.100 2228.620 ;
        RECT 3492.440 2228.340 3492.720 2228.620 ;
        RECT 3493.060 2228.340 3493.340 2228.620 ;
        RECT 3493.680 2228.340 3493.960 2228.620 ;
        RECT 3489.960 2227.720 3490.240 2228.000 ;
        RECT 3490.580 2227.720 3490.860 2228.000 ;
        RECT 3491.200 2227.720 3491.480 2228.000 ;
        RECT 3491.820 2227.720 3492.100 2228.000 ;
        RECT 3492.440 2227.720 3492.720 2228.000 ;
        RECT 3493.060 2227.720 3493.340 2228.000 ;
        RECT 3493.680 2227.720 3493.960 2228.000 ;
        RECT 3489.960 2227.100 3490.240 2227.380 ;
        RECT 3490.580 2227.100 3490.860 2227.380 ;
        RECT 3491.200 2227.100 3491.480 2227.380 ;
        RECT 3491.820 2227.100 3492.100 2227.380 ;
        RECT 3492.440 2227.100 3492.720 2227.380 ;
        RECT 3493.060 2227.100 3493.340 2227.380 ;
        RECT 3493.680 2227.100 3493.960 2227.380 ;
        RECT 3489.960 2226.480 3490.240 2226.760 ;
        RECT 3490.580 2226.480 3490.860 2226.760 ;
        RECT 3491.200 2226.480 3491.480 2226.760 ;
        RECT 3491.820 2226.480 3492.100 2226.760 ;
        RECT 3492.440 2226.480 3492.720 2226.760 ;
        RECT 3493.060 2226.480 3493.340 2226.760 ;
        RECT 3493.680 2226.480 3493.960 2226.760 ;
        RECT 3489.960 2225.860 3490.240 2226.140 ;
        RECT 3490.580 2225.860 3490.860 2226.140 ;
        RECT 3491.200 2225.860 3491.480 2226.140 ;
        RECT 3491.820 2225.860 3492.100 2226.140 ;
        RECT 3492.440 2225.860 3492.720 2226.140 ;
        RECT 3493.060 2225.860 3493.340 2226.140 ;
        RECT 3493.680 2225.860 3493.960 2226.140 ;
        RECT 3489.960 2225.240 3490.240 2225.520 ;
        RECT 3490.580 2225.240 3490.860 2225.520 ;
        RECT 3491.200 2225.240 3491.480 2225.520 ;
        RECT 3491.820 2225.240 3492.100 2225.520 ;
        RECT 3492.440 2225.240 3492.720 2225.520 ;
        RECT 3493.060 2225.240 3493.340 2225.520 ;
        RECT 3493.680 2225.240 3493.960 2225.520 ;
        RECT 3489.960 2224.620 3490.240 2224.900 ;
        RECT 3490.580 2224.620 3490.860 2224.900 ;
        RECT 3491.200 2224.620 3491.480 2224.900 ;
        RECT 3491.820 2224.620 3492.100 2224.900 ;
        RECT 3492.440 2224.620 3492.720 2224.900 ;
        RECT 3493.060 2224.620 3493.340 2224.900 ;
        RECT 3493.680 2224.620 3493.960 2224.900 ;
        RECT 3489.960 2224.000 3490.240 2224.280 ;
        RECT 3490.580 2224.000 3490.860 2224.280 ;
        RECT 3491.200 2224.000 3491.480 2224.280 ;
        RECT 3491.820 2224.000 3492.100 2224.280 ;
        RECT 3492.440 2224.000 3492.720 2224.280 ;
        RECT 3493.060 2224.000 3493.340 2224.280 ;
        RECT 3493.680 2224.000 3493.960 2224.280 ;
        RECT 3489.960 2223.380 3490.240 2223.660 ;
        RECT 3490.580 2223.380 3490.860 2223.660 ;
        RECT 3491.200 2223.380 3491.480 2223.660 ;
        RECT 3491.820 2223.380 3492.100 2223.660 ;
        RECT 3492.440 2223.380 3492.720 2223.660 ;
        RECT 3493.060 2223.380 3493.340 2223.660 ;
        RECT 3493.680 2223.380 3493.960 2223.660 ;
        RECT 3489.960 2222.760 3490.240 2223.040 ;
        RECT 3490.580 2222.760 3490.860 2223.040 ;
        RECT 3491.200 2222.760 3491.480 2223.040 ;
        RECT 3491.820 2222.760 3492.100 2223.040 ;
        RECT 3492.440 2222.760 3492.720 2223.040 ;
        RECT 3493.060 2222.760 3493.340 2223.040 ;
        RECT 3493.680 2222.760 3493.960 2223.040 ;
        RECT 3489.960 2222.140 3490.240 2222.420 ;
        RECT 3490.580 2222.140 3490.860 2222.420 ;
        RECT 3491.200 2222.140 3491.480 2222.420 ;
        RECT 3491.820 2222.140 3492.100 2222.420 ;
        RECT 3492.440 2222.140 3492.720 2222.420 ;
        RECT 3493.060 2222.140 3493.340 2222.420 ;
        RECT 3493.680 2222.140 3493.960 2222.420 ;
        RECT 3489.960 2221.520 3490.240 2221.800 ;
        RECT 3490.580 2221.520 3490.860 2221.800 ;
        RECT 3491.200 2221.520 3491.480 2221.800 ;
        RECT 3491.820 2221.520 3492.100 2221.800 ;
        RECT 3492.440 2221.520 3492.720 2221.800 ;
        RECT 3493.060 2221.520 3493.340 2221.800 ;
        RECT 3493.680 2221.520 3493.960 2221.800 ;
        RECT 3489.960 2220.900 3490.240 2221.180 ;
        RECT 3490.580 2220.900 3490.860 2221.180 ;
        RECT 3491.200 2220.900 3491.480 2221.180 ;
        RECT 3491.820 2220.900 3492.100 2221.180 ;
        RECT 3492.440 2220.900 3492.720 2221.180 ;
        RECT 3493.060 2220.900 3493.340 2221.180 ;
        RECT 3493.680 2220.900 3493.960 2221.180 ;
        RECT 3489.960 2218.350 3490.240 2218.630 ;
        RECT 3490.580 2218.350 3490.860 2218.630 ;
        RECT 3491.200 2218.350 3491.480 2218.630 ;
        RECT 3491.820 2218.350 3492.100 2218.630 ;
        RECT 3492.440 2218.350 3492.720 2218.630 ;
        RECT 3493.060 2218.350 3493.340 2218.630 ;
        RECT 3493.680 2218.350 3493.960 2218.630 ;
        RECT 3489.960 2217.730 3490.240 2218.010 ;
        RECT 3490.580 2217.730 3490.860 2218.010 ;
        RECT 3491.200 2217.730 3491.480 2218.010 ;
        RECT 3491.820 2217.730 3492.100 2218.010 ;
        RECT 3492.440 2217.730 3492.720 2218.010 ;
        RECT 3493.060 2217.730 3493.340 2218.010 ;
        RECT 3493.680 2217.730 3493.960 2218.010 ;
        RECT 3489.960 2217.110 3490.240 2217.390 ;
        RECT 3490.580 2217.110 3490.860 2217.390 ;
        RECT 3491.200 2217.110 3491.480 2217.390 ;
        RECT 3491.820 2217.110 3492.100 2217.390 ;
        RECT 3492.440 2217.110 3492.720 2217.390 ;
        RECT 3493.060 2217.110 3493.340 2217.390 ;
        RECT 3493.680 2217.110 3493.960 2217.390 ;
        RECT 3489.960 2216.490 3490.240 2216.770 ;
        RECT 3490.580 2216.490 3490.860 2216.770 ;
        RECT 3491.200 2216.490 3491.480 2216.770 ;
        RECT 3491.820 2216.490 3492.100 2216.770 ;
        RECT 3492.440 2216.490 3492.720 2216.770 ;
        RECT 3493.060 2216.490 3493.340 2216.770 ;
        RECT 3493.680 2216.490 3493.960 2216.770 ;
        RECT 3489.960 2215.870 3490.240 2216.150 ;
        RECT 3490.580 2215.870 3490.860 2216.150 ;
        RECT 3491.200 2215.870 3491.480 2216.150 ;
        RECT 3491.820 2215.870 3492.100 2216.150 ;
        RECT 3492.440 2215.870 3492.720 2216.150 ;
        RECT 3493.060 2215.870 3493.340 2216.150 ;
        RECT 3493.680 2215.870 3493.960 2216.150 ;
        RECT 3489.960 2215.250 3490.240 2215.530 ;
        RECT 3490.580 2215.250 3490.860 2215.530 ;
        RECT 3491.200 2215.250 3491.480 2215.530 ;
        RECT 3491.820 2215.250 3492.100 2215.530 ;
        RECT 3492.440 2215.250 3492.720 2215.530 ;
        RECT 3493.060 2215.250 3493.340 2215.530 ;
        RECT 3493.680 2215.250 3493.960 2215.530 ;
        RECT 3489.960 2214.630 3490.240 2214.910 ;
        RECT 3490.580 2214.630 3490.860 2214.910 ;
        RECT 3491.200 2214.630 3491.480 2214.910 ;
        RECT 3491.820 2214.630 3492.100 2214.910 ;
        RECT 3492.440 2214.630 3492.720 2214.910 ;
        RECT 3493.060 2214.630 3493.340 2214.910 ;
        RECT 3493.680 2214.630 3493.960 2214.910 ;
        RECT 3489.960 2214.010 3490.240 2214.290 ;
        RECT 3490.580 2214.010 3490.860 2214.290 ;
        RECT 3491.200 2214.010 3491.480 2214.290 ;
        RECT 3491.820 2214.010 3492.100 2214.290 ;
        RECT 3492.440 2214.010 3492.720 2214.290 ;
        RECT 3493.060 2214.010 3493.340 2214.290 ;
        RECT 3493.680 2214.010 3493.960 2214.290 ;
        RECT 3489.960 2213.390 3490.240 2213.670 ;
        RECT 3490.580 2213.390 3490.860 2213.670 ;
        RECT 3491.200 2213.390 3491.480 2213.670 ;
        RECT 3491.820 2213.390 3492.100 2213.670 ;
        RECT 3492.440 2213.390 3492.720 2213.670 ;
        RECT 3493.060 2213.390 3493.340 2213.670 ;
        RECT 3493.680 2213.390 3493.960 2213.670 ;
        RECT 3489.960 2212.770 3490.240 2213.050 ;
        RECT 3490.580 2212.770 3490.860 2213.050 ;
        RECT 3491.200 2212.770 3491.480 2213.050 ;
        RECT 3491.820 2212.770 3492.100 2213.050 ;
        RECT 3492.440 2212.770 3492.720 2213.050 ;
        RECT 3493.060 2212.770 3493.340 2213.050 ;
        RECT 3493.680 2212.770 3493.960 2213.050 ;
        RECT 3489.960 2212.150 3490.240 2212.430 ;
        RECT 3490.580 2212.150 3490.860 2212.430 ;
        RECT 3491.200 2212.150 3491.480 2212.430 ;
        RECT 3491.820 2212.150 3492.100 2212.430 ;
        RECT 3492.440 2212.150 3492.720 2212.430 ;
        RECT 3493.060 2212.150 3493.340 2212.430 ;
        RECT 3493.680 2212.150 3493.960 2212.430 ;
        RECT 3489.960 2211.530 3490.240 2211.810 ;
        RECT 3490.580 2211.530 3490.860 2211.810 ;
        RECT 3491.200 2211.530 3491.480 2211.810 ;
        RECT 3491.820 2211.530 3492.100 2211.810 ;
        RECT 3492.440 2211.530 3492.720 2211.810 ;
        RECT 3493.060 2211.530 3493.340 2211.810 ;
        RECT 3493.680 2211.530 3493.960 2211.810 ;
        RECT 3489.960 2210.910 3490.240 2211.190 ;
        RECT 3490.580 2210.910 3490.860 2211.190 ;
        RECT 3491.200 2210.910 3491.480 2211.190 ;
        RECT 3491.820 2210.910 3492.100 2211.190 ;
        RECT 3492.440 2210.910 3492.720 2211.190 ;
        RECT 3493.060 2210.910 3493.340 2211.190 ;
        RECT 3493.680 2210.910 3493.960 2211.190 ;
        RECT 3489.960 2210.290 3490.240 2210.570 ;
        RECT 3490.580 2210.290 3490.860 2210.570 ;
        RECT 3491.200 2210.290 3491.480 2210.570 ;
        RECT 3491.820 2210.290 3492.100 2210.570 ;
        RECT 3492.440 2210.290 3492.720 2210.570 ;
        RECT 3493.060 2210.290 3493.340 2210.570 ;
        RECT 3493.680 2210.290 3493.960 2210.570 ;
        RECT 3489.960 2209.670 3490.240 2209.950 ;
        RECT 3490.580 2209.670 3490.860 2209.950 ;
        RECT 3491.200 2209.670 3491.480 2209.950 ;
        RECT 3491.820 2209.670 3492.100 2209.950 ;
        RECT 3492.440 2209.670 3492.720 2209.950 ;
        RECT 3493.060 2209.670 3493.340 2209.950 ;
        RECT 3493.680 2209.670 3493.960 2209.950 ;
        RECT 3489.960 2209.050 3490.240 2209.330 ;
        RECT 3490.580 2209.050 3490.860 2209.330 ;
        RECT 3491.200 2209.050 3491.480 2209.330 ;
        RECT 3491.820 2209.050 3492.100 2209.330 ;
        RECT 3492.440 2209.050 3492.720 2209.330 ;
        RECT 3493.060 2209.050 3493.340 2209.330 ;
        RECT 3493.680 2209.050 3493.960 2209.330 ;
        RECT 3489.960 2205.330 3490.240 2205.610 ;
        RECT 3490.580 2205.330 3490.860 2205.610 ;
        RECT 3491.200 2205.330 3491.480 2205.610 ;
        RECT 3491.820 2205.330 3492.100 2205.610 ;
        RECT 3492.440 2205.330 3492.720 2205.610 ;
        RECT 3493.060 2205.330 3493.340 2205.610 ;
        RECT 3493.680 2205.330 3493.960 2205.610 ;
        RECT 3489.960 2204.710 3490.240 2204.990 ;
        RECT 3490.580 2204.710 3490.860 2204.990 ;
        RECT 3491.200 2204.710 3491.480 2204.990 ;
        RECT 3491.820 2204.710 3492.100 2204.990 ;
        RECT 3492.440 2204.710 3492.720 2204.990 ;
        RECT 3493.060 2204.710 3493.340 2204.990 ;
        RECT 3493.680 2204.710 3493.960 2204.990 ;
        RECT 3489.960 2204.090 3490.240 2204.370 ;
        RECT 3490.580 2204.090 3490.860 2204.370 ;
        RECT 3491.200 2204.090 3491.480 2204.370 ;
        RECT 3491.820 2204.090 3492.100 2204.370 ;
        RECT 3492.440 2204.090 3492.720 2204.370 ;
        RECT 3493.060 2204.090 3493.340 2204.370 ;
        RECT 3493.680 2204.090 3493.960 2204.370 ;
        RECT 3489.960 2203.470 3490.240 2203.750 ;
        RECT 3490.580 2203.470 3490.860 2203.750 ;
        RECT 3491.200 2203.470 3491.480 2203.750 ;
        RECT 3491.820 2203.470 3492.100 2203.750 ;
        RECT 3492.440 2203.470 3492.720 2203.750 ;
        RECT 3493.060 2203.470 3493.340 2203.750 ;
        RECT 3493.680 2203.470 3493.960 2203.750 ;
        RECT 3489.960 2202.850 3490.240 2203.130 ;
        RECT 3490.580 2202.850 3490.860 2203.130 ;
        RECT 3491.200 2202.850 3491.480 2203.130 ;
        RECT 3491.820 2202.850 3492.100 2203.130 ;
        RECT 3492.440 2202.850 3492.720 2203.130 ;
        RECT 3493.060 2202.850 3493.340 2203.130 ;
        RECT 3493.680 2202.850 3493.960 2203.130 ;
        RECT 3489.960 2202.230 3490.240 2202.510 ;
        RECT 3490.580 2202.230 3490.860 2202.510 ;
        RECT 3491.200 2202.230 3491.480 2202.510 ;
        RECT 3491.820 2202.230 3492.100 2202.510 ;
        RECT 3492.440 2202.230 3492.720 2202.510 ;
        RECT 3493.060 2202.230 3493.340 2202.510 ;
        RECT 3493.680 2202.230 3493.960 2202.510 ;
        RECT 3489.960 2201.610 3490.240 2201.890 ;
        RECT 3490.580 2201.610 3490.860 2201.890 ;
        RECT 3491.200 2201.610 3491.480 2201.890 ;
        RECT 3491.820 2201.610 3492.100 2201.890 ;
        RECT 3492.440 2201.610 3492.720 2201.890 ;
        RECT 3493.060 2201.610 3493.340 2201.890 ;
        RECT 3493.680 2201.610 3493.960 2201.890 ;
        RECT 3489.960 2200.990 3490.240 2201.270 ;
        RECT 3490.580 2200.990 3490.860 2201.270 ;
        RECT 3491.200 2200.990 3491.480 2201.270 ;
        RECT 3491.820 2200.990 3492.100 2201.270 ;
        RECT 3492.440 2200.990 3492.720 2201.270 ;
        RECT 3493.060 2200.990 3493.340 2201.270 ;
        RECT 3493.680 2200.990 3493.960 2201.270 ;
        RECT 3489.960 2200.370 3490.240 2200.650 ;
        RECT 3490.580 2200.370 3490.860 2200.650 ;
        RECT 3491.200 2200.370 3491.480 2200.650 ;
        RECT 3491.820 2200.370 3492.100 2200.650 ;
        RECT 3492.440 2200.370 3492.720 2200.650 ;
        RECT 3493.060 2200.370 3493.340 2200.650 ;
        RECT 3493.680 2200.370 3493.960 2200.650 ;
        RECT 3489.960 2199.750 3490.240 2200.030 ;
        RECT 3490.580 2199.750 3490.860 2200.030 ;
        RECT 3491.200 2199.750 3491.480 2200.030 ;
        RECT 3491.820 2199.750 3492.100 2200.030 ;
        RECT 3492.440 2199.750 3492.720 2200.030 ;
        RECT 3493.060 2199.750 3493.340 2200.030 ;
        RECT 3493.680 2199.750 3493.960 2200.030 ;
        RECT 3489.960 2199.130 3490.240 2199.410 ;
        RECT 3490.580 2199.130 3490.860 2199.410 ;
        RECT 3491.200 2199.130 3491.480 2199.410 ;
        RECT 3491.820 2199.130 3492.100 2199.410 ;
        RECT 3492.440 2199.130 3492.720 2199.410 ;
        RECT 3493.060 2199.130 3493.340 2199.410 ;
        RECT 3493.680 2199.130 3493.960 2199.410 ;
        RECT 3489.960 2198.510 3490.240 2198.790 ;
        RECT 3490.580 2198.510 3490.860 2198.790 ;
        RECT 3491.200 2198.510 3491.480 2198.790 ;
        RECT 3491.820 2198.510 3492.100 2198.790 ;
        RECT 3492.440 2198.510 3492.720 2198.790 ;
        RECT 3493.060 2198.510 3493.340 2198.790 ;
        RECT 3493.680 2198.510 3493.960 2198.790 ;
        RECT 3489.960 2197.890 3490.240 2198.170 ;
        RECT 3490.580 2197.890 3490.860 2198.170 ;
        RECT 3491.200 2197.890 3491.480 2198.170 ;
        RECT 3491.820 2197.890 3492.100 2198.170 ;
        RECT 3492.440 2197.890 3492.720 2198.170 ;
        RECT 3493.060 2197.890 3493.340 2198.170 ;
        RECT 3493.680 2197.890 3493.960 2198.170 ;
        RECT 3489.960 2197.270 3490.240 2197.550 ;
        RECT 3490.580 2197.270 3490.860 2197.550 ;
        RECT 3491.200 2197.270 3491.480 2197.550 ;
        RECT 3491.820 2197.270 3492.100 2197.550 ;
        RECT 3492.440 2197.270 3492.720 2197.550 ;
        RECT 3493.060 2197.270 3493.340 2197.550 ;
        RECT 3493.680 2197.270 3493.960 2197.550 ;
        RECT 3489.960 2196.650 3490.240 2196.930 ;
        RECT 3490.580 2196.650 3490.860 2196.930 ;
        RECT 3491.200 2196.650 3491.480 2196.930 ;
        RECT 3491.820 2196.650 3492.100 2196.930 ;
        RECT 3492.440 2196.650 3492.720 2196.930 ;
        RECT 3493.060 2196.650 3493.340 2196.930 ;
        RECT 3493.680 2196.650 3493.960 2196.930 ;
        RECT 3490.720 2141.865 3491.000 2142.145 ;
        RECT 3492.220 2141.865 3492.500 2142.145 ;
        RECT 3493.720 2141.865 3494.000 2142.145 ;
        RECT 3490.720 2140.865 3491.000 2141.145 ;
        RECT 3492.220 2140.865 3492.500 2141.145 ;
        RECT 3493.720 2140.865 3494.000 2141.145 ;
        RECT 3489.960 2052.980 3490.240 2053.260 ;
        RECT 3490.580 2052.980 3490.860 2053.260 ;
        RECT 3491.200 2052.980 3491.480 2053.260 ;
        RECT 3491.820 2052.980 3492.100 2053.260 ;
        RECT 3492.440 2052.980 3492.720 2053.260 ;
        RECT 3493.060 2052.980 3493.340 2053.260 ;
        RECT 3493.680 2052.980 3493.960 2053.260 ;
        RECT 3489.960 2052.360 3490.240 2052.640 ;
        RECT 3490.580 2052.360 3490.860 2052.640 ;
        RECT 3491.200 2052.360 3491.480 2052.640 ;
        RECT 3491.820 2052.360 3492.100 2052.640 ;
        RECT 3492.440 2052.360 3492.720 2052.640 ;
        RECT 3493.060 2052.360 3493.340 2052.640 ;
        RECT 3493.680 2052.360 3493.960 2052.640 ;
        RECT 3489.960 2051.740 3490.240 2052.020 ;
        RECT 3490.580 2051.740 3490.860 2052.020 ;
        RECT 3491.200 2051.740 3491.480 2052.020 ;
        RECT 3491.820 2051.740 3492.100 2052.020 ;
        RECT 3492.440 2051.740 3492.720 2052.020 ;
        RECT 3493.060 2051.740 3493.340 2052.020 ;
        RECT 3493.680 2051.740 3493.960 2052.020 ;
        RECT 3489.960 2051.120 3490.240 2051.400 ;
        RECT 3490.580 2051.120 3490.860 2051.400 ;
        RECT 3491.200 2051.120 3491.480 2051.400 ;
        RECT 3491.820 2051.120 3492.100 2051.400 ;
        RECT 3492.440 2051.120 3492.720 2051.400 ;
        RECT 3493.060 2051.120 3493.340 2051.400 ;
        RECT 3493.680 2051.120 3493.960 2051.400 ;
        RECT 3489.960 2050.500 3490.240 2050.780 ;
        RECT 3490.580 2050.500 3490.860 2050.780 ;
        RECT 3491.200 2050.500 3491.480 2050.780 ;
        RECT 3491.820 2050.500 3492.100 2050.780 ;
        RECT 3492.440 2050.500 3492.720 2050.780 ;
        RECT 3493.060 2050.500 3493.340 2050.780 ;
        RECT 3493.680 2050.500 3493.960 2050.780 ;
        RECT 3489.960 2049.880 3490.240 2050.160 ;
        RECT 3490.580 2049.880 3490.860 2050.160 ;
        RECT 3491.200 2049.880 3491.480 2050.160 ;
        RECT 3491.820 2049.880 3492.100 2050.160 ;
        RECT 3492.440 2049.880 3492.720 2050.160 ;
        RECT 3493.060 2049.880 3493.340 2050.160 ;
        RECT 3493.680 2049.880 3493.960 2050.160 ;
        RECT 3489.960 2049.260 3490.240 2049.540 ;
        RECT 3490.580 2049.260 3490.860 2049.540 ;
        RECT 3491.200 2049.260 3491.480 2049.540 ;
        RECT 3491.820 2049.260 3492.100 2049.540 ;
        RECT 3492.440 2049.260 3492.720 2049.540 ;
        RECT 3493.060 2049.260 3493.340 2049.540 ;
        RECT 3493.680 2049.260 3493.960 2049.540 ;
        RECT 3489.960 2048.640 3490.240 2048.920 ;
        RECT 3490.580 2048.640 3490.860 2048.920 ;
        RECT 3491.200 2048.640 3491.480 2048.920 ;
        RECT 3491.820 2048.640 3492.100 2048.920 ;
        RECT 3492.440 2048.640 3492.720 2048.920 ;
        RECT 3493.060 2048.640 3493.340 2048.920 ;
        RECT 3493.680 2048.640 3493.960 2048.920 ;
        RECT 3489.960 2048.020 3490.240 2048.300 ;
        RECT 3490.580 2048.020 3490.860 2048.300 ;
        RECT 3491.200 2048.020 3491.480 2048.300 ;
        RECT 3491.820 2048.020 3492.100 2048.300 ;
        RECT 3492.440 2048.020 3492.720 2048.300 ;
        RECT 3493.060 2048.020 3493.340 2048.300 ;
        RECT 3493.680 2048.020 3493.960 2048.300 ;
        RECT 3489.960 2047.400 3490.240 2047.680 ;
        RECT 3490.580 2047.400 3490.860 2047.680 ;
        RECT 3491.200 2047.400 3491.480 2047.680 ;
        RECT 3491.820 2047.400 3492.100 2047.680 ;
        RECT 3492.440 2047.400 3492.720 2047.680 ;
        RECT 3493.060 2047.400 3493.340 2047.680 ;
        RECT 3493.680 2047.400 3493.960 2047.680 ;
        RECT 3489.960 2046.780 3490.240 2047.060 ;
        RECT 3490.580 2046.780 3490.860 2047.060 ;
        RECT 3491.200 2046.780 3491.480 2047.060 ;
        RECT 3491.820 2046.780 3492.100 2047.060 ;
        RECT 3492.440 2046.780 3492.720 2047.060 ;
        RECT 3493.060 2046.780 3493.340 2047.060 ;
        RECT 3493.680 2046.780 3493.960 2047.060 ;
        RECT 3489.960 2046.160 3490.240 2046.440 ;
        RECT 3490.580 2046.160 3490.860 2046.440 ;
        RECT 3491.200 2046.160 3491.480 2046.440 ;
        RECT 3491.820 2046.160 3492.100 2046.440 ;
        RECT 3492.440 2046.160 3492.720 2046.440 ;
        RECT 3493.060 2046.160 3493.340 2046.440 ;
        RECT 3493.680 2046.160 3493.960 2046.440 ;
        RECT 3489.960 2045.540 3490.240 2045.820 ;
        RECT 3490.580 2045.540 3490.860 2045.820 ;
        RECT 3491.200 2045.540 3491.480 2045.820 ;
        RECT 3491.820 2045.540 3492.100 2045.820 ;
        RECT 3492.440 2045.540 3492.720 2045.820 ;
        RECT 3493.060 2045.540 3493.340 2045.820 ;
        RECT 3493.680 2045.540 3493.960 2045.820 ;
        RECT 3489.960 2044.920 3490.240 2045.200 ;
        RECT 3490.580 2044.920 3490.860 2045.200 ;
        RECT 3491.200 2044.920 3491.480 2045.200 ;
        RECT 3491.820 2044.920 3492.100 2045.200 ;
        RECT 3492.440 2044.920 3492.720 2045.200 ;
        RECT 3493.060 2044.920 3493.340 2045.200 ;
        RECT 3493.680 2044.920 3493.960 2045.200 ;
        RECT 3489.960 2044.300 3490.240 2044.580 ;
        RECT 3490.580 2044.300 3490.860 2044.580 ;
        RECT 3491.200 2044.300 3491.480 2044.580 ;
        RECT 3491.820 2044.300 3492.100 2044.580 ;
        RECT 3492.440 2044.300 3492.720 2044.580 ;
        RECT 3493.060 2044.300 3493.340 2044.580 ;
        RECT 3493.680 2044.300 3493.960 2044.580 ;
        RECT 3489.960 2040.580 3490.240 2040.860 ;
        RECT 3490.580 2040.580 3490.860 2040.860 ;
        RECT 3491.200 2040.580 3491.480 2040.860 ;
        RECT 3491.820 2040.580 3492.100 2040.860 ;
        RECT 3492.440 2040.580 3492.720 2040.860 ;
        RECT 3493.060 2040.580 3493.340 2040.860 ;
        RECT 3493.680 2040.580 3493.960 2040.860 ;
        RECT 3489.960 2039.960 3490.240 2040.240 ;
        RECT 3490.580 2039.960 3490.860 2040.240 ;
        RECT 3491.200 2039.960 3491.480 2040.240 ;
        RECT 3491.820 2039.960 3492.100 2040.240 ;
        RECT 3492.440 2039.960 3492.720 2040.240 ;
        RECT 3493.060 2039.960 3493.340 2040.240 ;
        RECT 3493.680 2039.960 3493.960 2040.240 ;
        RECT 3489.960 2039.340 3490.240 2039.620 ;
        RECT 3490.580 2039.340 3490.860 2039.620 ;
        RECT 3491.200 2039.340 3491.480 2039.620 ;
        RECT 3491.820 2039.340 3492.100 2039.620 ;
        RECT 3492.440 2039.340 3492.720 2039.620 ;
        RECT 3493.060 2039.340 3493.340 2039.620 ;
        RECT 3493.680 2039.340 3493.960 2039.620 ;
        RECT 3489.960 2038.720 3490.240 2039.000 ;
        RECT 3490.580 2038.720 3490.860 2039.000 ;
        RECT 3491.200 2038.720 3491.480 2039.000 ;
        RECT 3491.820 2038.720 3492.100 2039.000 ;
        RECT 3492.440 2038.720 3492.720 2039.000 ;
        RECT 3493.060 2038.720 3493.340 2039.000 ;
        RECT 3493.680 2038.720 3493.960 2039.000 ;
        RECT 3489.960 2038.100 3490.240 2038.380 ;
        RECT 3490.580 2038.100 3490.860 2038.380 ;
        RECT 3491.200 2038.100 3491.480 2038.380 ;
        RECT 3491.820 2038.100 3492.100 2038.380 ;
        RECT 3492.440 2038.100 3492.720 2038.380 ;
        RECT 3493.060 2038.100 3493.340 2038.380 ;
        RECT 3493.680 2038.100 3493.960 2038.380 ;
        RECT 3489.960 2037.480 3490.240 2037.760 ;
        RECT 3490.580 2037.480 3490.860 2037.760 ;
        RECT 3491.200 2037.480 3491.480 2037.760 ;
        RECT 3491.820 2037.480 3492.100 2037.760 ;
        RECT 3492.440 2037.480 3492.720 2037.760 ;
        RECT 3493.060 2037.480 3493.340 2037.760 ;
        RECT 3493.680 2037.480 3493.960 2037.760 ;
        RECT 3489.960 2036.860 3490.240 2037.140 ;
        RECT 3490.580 2036.860 3490.860 2037.140 ;
        RECT 3491.200 2036.860 3491.480 2037.140 ;
        RECT 3491.820 2036.860 3492.100 2037.140 ;
        RECT 3492.440 2036.860 3492.720 2037.140 ;
        RECT 3493.060 2036.860 3493.340 2037.140 ;
        RECT 3493.680 2036.860 3493.960 2037.140 ;
        RECT 3489.960 2036.240 3490.240 2036.520 ;
        RECT 3490.580 2036.240 3490.860 2036.520 ;
        RECT 3491.200 2036.240 3491.480 2036.520 ;
        RECT 3491.820 2036.240 3492.100 2036.520 ;
        RECT 3492.440 2036.240 3492.720 2036.520 ;
        RECT 3493.060 2036.240 3493.340 2036.520 ;
        RECT 3493.680 2036.240 3493.960 2036.520 ;
        RECT 3489.960 2035.620 3490.240 2035.900 ;
        RECT 3490.580 2035.620 3490.860 2035.900 ;
        RECT 3491.200 2035.620 3491.480 2035.900 ;
        RECT 3491.820 2035.620 3492.100 2035.900 ;
        RECT 3492.440 2035.620 3492.720 2035.900 ;
        RECT 3493.060 2035.620 3493.340 2035.900 ;
        RECT 3493.680 2035.620 3493.960 2035.900 ;
        RECT 3489.960 2035.000 3490.240 2035.280 ;
        RECT 3490.580 2035.000 3490.860 2035.280 ;
        RECT 3491.200 2035.000 3491.480 2035.280 ;
        RECT 3491.820 2035.000 3492.100 2035.280 ;
        RECT 3492.440 2035.000 3492.720 2035.280 ;
        RECT 3493.060 2035.000 3493.340 2035.280 ;
        RECT 3493.680 2035.000 3493.960 2035.280 ;
        RECT 3489.960 2034.380 3490.240 2034.660 ;
        RECT 3490.580 2034.380 3490.860 2034.660 ;
        RECT 3491.200 2034.380 3491.480 2034.660 ;
        RECT 3491.820 2034.380 3492.100 2034.660 ;
        RECT 3492.440 2034.380 3492.720 2034.660 ;
        RECT 3493.060 2034.380 3493.340 2034.660 ;
        RECT 3493.680 2034.380 3493.960 2034.660 ;
        RECT 3489.960 2033.760 3490.240 2034.040 ;
        RECT 3490.580 2033.760 3490.860 2034.040 ;
        RECT 3491.200 2033.760 3491.480 2034.040 ;
        RECT 3491.820 2033.760 3492.100 2034.040 ;
        RECT 3492.440 2033.760 3492.720 2034.040 ;
        RECT 3493.060 2033.760 3493.340 2034.040 ;
        RECT 3493.680 2033.760 3493.960 2034.040 ;
        RECT 3489.960 2033.140 3490.240 2033.420 ;
        RECT 3490.580 2033.140 3490.860 2033.420 ;
        RECT 3491.200 2033.140 3491.480 2033.420 ;
        RECT 3491.820 2033.140 3492.100 2033.420 ;
        RECT 3492.440 2033.140 3492.720 2033.420 ;
        RECT 3493.060 2033.140 3493.340 2033.420 ;
        RECT 3493.680 2033.140 3493.960 2033.420 ;
        RECT 3489.960 2032.520 3490.240 2032.800 ;
        RECT 3490.580 2032.520 3490.860 2032.800 ;
        RECT 3491.200 2032.520 3491.480 2032.800 ;
        RECT 3491.820 2032.520 3492.100 2032.800 ;
        RECT 3492.440 2032.520 3492.720 2032.800 ;
        RECT 3493.060 2032.520 3493.340 2032.800 ;
        RECT 3493.680 2032.520 3493.960 2032.800 ;
        RECT 3489.960 2031.900 3490.240 2032.180 ;
        RECT 3490.580 2031.900 3490.860 2032.180 ;
        RECT 3491.200 2031.900 3491.480 2032.180 ;
        RECT 3491.820 2031.900 3492.100 2032.180 ;
        RECT 3492.440 2031.900 3492.720 2032.180 ;
        RECT 3493.060 2031.900 3493.340 2032.180 ;
        RECT 3493.680 2031.900 3493.960 2032.180 ;
        RECT 3489.960 2031.280 3490.240 2031.560 ;
        RECT 3490.580 2031.280 3490.860 2031.560 ;
        RECT 3491.200 2031.280 3491.480 2031.560 ;
        RECT 3491.820 2031.280 3492.100 2031.560 ;
        RECT 3492.440 2031.280 3492.720 2031.560 ;
        RECT 3493.060 2031.280 3493.340 2031.560 ;
        RECT 3493.680 2031.280 3493.960 2031.560 ;
        RECT 3489.960 2028.730 3490.240 2029.010 ;
        RECT 3490.580 2028.730 3490.860 2029.010 ;
        RECT 3491.200 2028.730 3491.480 2029.010 ;
        RECT 3491.820 2028.730 3492.100 2029.010 ;
        RECT 3492.440 2028.730 3492.720 2029.010 ;
        RECT 3493.060 2028.730 3493.340 2029.010 ;
        RECT 3493.680 2028.730 3493.960 2029.010 ;
        RECT 3489.960 2028.110 3490.240 2028.390 ;
        RECT 3490.580 2028.110 3490.860 2028.390 ;
        RECT 3491.200 2028.110 3491.480 2028.390 ;
        RECT 3491.820 2028.110 3492.100 2028.390 ;
        RECT 3492.440 2028.110 3492.720 2028.390 ;
        RECT 3493.060 2028.110 3493.340 2028.390 ;
        RECT 3493.680 2028.110 3493.960 2028.390 ;
        RECT 3489.960 2027.490 3490.240 2027.770 ;
        RECT 3490.580 2027.490 3490.860 2027.770 ;
        RECT 3491.200 2027.490 3491.480 2027.770 ;
        RECT 3491.820 2027.490 3492.100 2027.770 ;
        RECT 3492.440 2027.490 3492.720 2027.770 ;
        RECT 3493.060 2027.490 3493.340 2027.770 ;
        RECT 3493.680 2027.490 3493.960 2027.770 ;
        RECT 3489.960 2026.870 3490.240 2027.150 ;
        RECT 3490.580 2026.870 3490.860 2027.150 ;
        RECT 3491.200 2026.870 3491.480 2027.150 ;
        RECT 3491.820 2026.870 3492.100 2027.150 ;
        RECT 3492.440 2026.870 3492.720 2027.150 ;
        RECT 3493.060 2026.870 3493.340 2027.150 ;
        RECT 3493.680 2026.870 3493.960 2027.150 ;
        RECT 3489.960 2026.250 3490.240 2026.530 ;
        RECT 3490.580 2026.250 3490.860 2026.530 ;
        RECT 3491.200 2026.250 3491.480 2026.530 ;
        RECT 3491.820 2026.250 3492.100 2026.530 ;
        RECT 3492.440 2026.250 3492.720 2026.530 ;
        RECT 3493.060 2026.250 3493.340 2026.530 ;
        RECT 3493.680 2026.250 3493.960 2026.530 ;
        RECT 3489.960 2025.630 3490.240 2025.910 ;
        RECT 3490.580 2025.630 3490.860 2025.910 ;
        RECT 3491.200 2025.630 3491.480 2025.910 ;
        RECT 3491.820 2025.630 3492.100 2025.910 ;
        RECT 3492.440 2025.630 3492.720 2025.910 ;
        RECT 3493.060 2025.630 3493.340 2025.910 ;
        RECT 3493.680 2025.630 3493.960 2025.910 ;
        RECT 3489.960 2025.010 3490.240 2025.290 ;
        RECT 3490.580 2025.010 3490.860 2025.290 ;
        RECT 3491.200 2025.010 3491.480 2025.290 ;
        RECT 3491.820 2025.010 3492.100 2025.290 ;
        RECT 3492.440 2025.010 3492.720 2025.290 ;
        RECT 3493.060 2025.010 3493.340 2025.290 ;
        RECT 3493.680 2025.010 3493.960 2025.290 ;
        RECT 3489.960 2024.390 3490.240 2024.670 ;
        RECT 3490.580 2024.390 3490.860 2024.670 ;
        RECT 3491.200 2024.390 3491.480 2024.670 ;
        RECT 3491.820 2024.390 3492.100 2024.670 ;
        RECT 3492.440 2024.390 3492.720 2024.670 ;
        RECT 3493.060 2024.390 3493.340 2024.670 ;
        RECT 3493.680 2024.390 3493.960 2024.670 ;
        RECT 3489.960 2023.770 3490.240 2024.050 ;
        RECT 3490.580 2023.770 3490.860 2024.050 ;
        RECT 3491.200 2023.770 3491.480 2024.050 ;
        RECT 3491.820 2023.770 3492.100 2024.050 ;
        RECT 3492.440 2023.770 3492.720 2024.050 ;
        RECT 3493.060 2023.770 3493.340 2024.050 ;
        RECT 3493.680 2023.770 3493.960 2024.050 ;
        RECT 3489.960 2023.150 3490.240 2023.430 ;
        RECT 3490.580 2023.150 3490.860 2023.430 ;
        RECT 3491.200 2023.150 3491.480 2023.430 ;
        RECT 3491.820 2023.150 3492.100 2023.430 ;
        RECT 3492.440 2023.150 3492.720 2023.430 ;
        RECT 3493.060 2023.150 3493.340 2023.430 ;
        RECT 3493.680 2023.150 3493.960 2023.430 ;
        RECT 3489.960 2022.530 3490.240 2022.810 ;
        RECT 3490.580 2022.530 3490.860 2022.810 ;
        RECT 3491.200 2022.530 3491.480 2022.810 ;
        RECT 3491.820 2022.530 3492.100 2022.810 ;
        RECT 3492.440 2022.530 3492.720 2022.810 ;
        RECT 3493.060 2022.530 3493.340 2022.810 ;
        RECT 3493.680 2022.530 3493.960 2022.810 ;
        RECT 3489.960 2021.910 3490.240 2022.190 ;
        RECT 3490.580 2021.910 3490.860 2022.190 ;
        RECT 3491.200 2021.910 3491.480 2022.190 ;
        RECT 3491.820 2021.910 3492.100 2022.190 ;
        RECT 3492.440 2021.910 3492.720 2022.190 ;
        RECT 3493.060 2021.910 3493.340 2022.190 ;
        RECT 3493.680 2021.910 3493.960 2022.190 ;
        RECT 3489.960 2021.290 3490.240 2021.570 ;
        RECT 3490.580 2021.290 3490.860 2021.570 ;
        RECT 3491.200 2021.290 3491.480 2021.570 ;
        RECT 3491.820 2021.290 3492.100 2021.570 ;
        RECT 3492.440 2021.290 3492.720 2021.570 ;
        RECT 3493.060 2021.290 3493.340 2021.570 ;
        RECT 3493.680 2021.290 3493.960 2021.570 ;
        RECT 3489.960 2020.670 3490.240 2020.950 ;
        RECT 3490.580 2020.670 3490.860 2020.950 ;
        RECT 3491.200 2020.670 3491.480 2020.950 ;
        RECT 3491.820 2020.670 3492.100 2020.950 ;
        RECT 3492.440 2020.670 3492.720 2020.950 ;
        RECT 3493.060 2020.670 3493.340 2020.950 ;
        RECT 3493.680 2020.670 3493.960 2020.950 ;
        RECT 3489.960 2020.050 3490.240 2020.330 ;
        RECT 3490.580 2020.050 3490.860 2020.330 ;
        RECT 3491.200 2020.050 3491.480 2020.330 ;
        RECT 3491.820 2020.050 3492.100 2020.330 ;
        RECT 3492.440 2020.050 3492.720 2020.330 ;
        RECT 3493.060 2020.050 3493.340 2020.330 ;
        RECT 3493.680 2020.050 3493.960 2020.330 ;
        RECT 3489.960 2019.430 3490.240 2019.710 ;
        RECT 3490.580 2019.430 3490.860 2019.710 ;
        RECT 3491.200 2019.430 3491.480 2019.710 ;
        RECT 3491.820 2019.430 3492.100 2019.710 ;
        RECT 3492.440 2019.430 3492.720 2019.710 ;
        RECT 3493.060 2019.430 3493.340 2019.710 ;
        RECT 3493.680 2019.430 3493.960 2019.710 ;
        RECT 3489.960 2015.200 3490.240 2015.480 ;
        RECT 3490.580 2015.200 3490.860 2015.480 ;
        RECT 3491.200 2015.200 3491.480 2015.480 ;
        RECT 3491.820 2015.200 3492.100 2015.480 ;
        RECT 3492.440 2015.200 3492.720 2015.480 ;
        RECT 3493.060 2015.200 3493.340 2015.480 ;
        RECT 3493.680 2015.200 3493.960 2015.480 ;
        RECT 3489.960 2014.580 3490.240 2014.860 ;
        RECT 3490.580 2014.580 3490.860 2014.860 ;
        RECT 3491.200 2014.580 3491.480 2014.860 ;
        RECT 3491.820 2014.580 3492.100 2014.860 ;
        RECT 3492.440 2014.580 3492.720 2014.860 ;
        RECT 3493.060 2014.580 3493.340 2014.860 ;
        RECT 3493.680 2014.580 3493.960 2014.860 ;
        RECT 3489.960 2013.960 3490.240 2014.240 ;
        RECT 3490.580 2013.960 3490.860 2014.240 ;
        RECT 3491.200 2013.960 3491.480 2014.240 ;
        RECT 3491.820 2013.960 3492.100 2014.240 ;
        RECT 3492.440 2013.960 3492.720 2014.240 ;
        RECT 3493.060 2013.960 3493.340 2014.240 ;
        RECT 3493.680 2013.960 3493.960 2014.240 ;
        RECT 3489.960 2013.340 3490.240 2013.620 ;
        RECT 3490.580 2013.340 3490.860 2013.620 ;
        RECT 3491.200 2013.340 3491.480 2013.620 ;
        RECT 3491.820 2013.340 3492.100 2013.620 ;
        RECT 3492.440 2013.340 3492.720 2013.620 ;
        RECT 3493.060 2013.340 3493.340 2013.620 ;
        RECT 3493.680 2013.340 3493.960 2013.620 ;
        RECT 3489.960 2012.720 3490.240 2013.000 ;
        RECT 3490.580 2012.720 3490.860 2013.000 ;
        RECT 3491.200 2012.720 3491.480 2013.000 ;
        RECT 3491.820 2012.720 3492.100 2013.000 ;
        RECT 3492.440 2012.720 3492.720 2013.000 ;
        RECT 3493.060 2012.720 3493.340 2013.000 ;
        RECT 3493.680 2012.720 3493.960 2013.000 ;
        RECT 3489.960 2012.100 3490.240 2012.380 ;
        RECT 3490.580 2012.100 3490.860 2012.380 ;
        RECT 3491.200 2012.100 3491.480 2012.380 ;
        RECT 3491.820 2012.100 3492.100 2012.380 ;
        RECT 3492.440 2012.100 3492.720 2012.380 ;
        RECT 3493.060 2012.100 3493.340 2012.380 ;
        RECT 3493.680 2012.100 3493.960 2012.380 ;
        RECT 3489.960 2011.480 3490.240 2011.760 ;
        RECT 3490.580 2011.480 3490.860 2011.760 ;
        RECT 3491.200 2011.480 3491.480 2011.760 ;
        RECT 3491.820 2011.480 3492.100 2011.760 ;
        RECT 3492.440 2011.480 3492.720 2011.760 ;
        RECT 3493.060 2011.480 3493.340 2011.760 ;
        RECT 3493.680 2011.480 3493.960 2011.760 ;
        RECT 3489.960 2010.860 3490.240 2011.140 ;
        RECT 3490.580 2010.860 3490.860 2011.140 ;
        RECT 3491.200 2010.860 3491.480 2011.140 ;
        RECT 3491.820 2010.860 3492.100 2011.140 ;
        RECT 3492.440 2010.860 3492.720 2011.140 ;
        RECT 3493.060 2010.860 3493.340 2011.140 ;
        RECT 3493.680 2010.860 3493.960 2011.140 ;
        RECT 3489.960 2010.240 3490.240 2010.520 ;
        RECT 3490.580 2010.240 3490.860 2010.520 ;
        RECT 3491.200 2010.240 3491.480 2010.520 ;
        RECT 3491.820 2010.240 3492.100 2010.520 ;
        RECT 3492.440 2010.240 3492.720 2010.520 ;
        RECT 3493.060 2010.240 3493.340 2010.520 ;
        RECT 3493.680 2010.240 3493.960 2010.520 ;
        RECT 3489.960 2009.620 3490.240 2009.900 ;
        RECT 3490.580 2009.620 3490.860 2009.900 ;
        RECT 3491.200 2009.620 3491.480 2009.900 ;
        RECT 3491.820 2009.620 3492.100 2009.900 ;
        RECT 3492.440 2009.620 3492.720 2009.900 ;
        RECT 3493.060 2009.620 3493.340 2009.900 ;
        RECT 3493.680 2009.620 3493.960 2009.900 ;
        RECT 3489.960 2009.000 3490.240 2009.280 ;
        RECT 3490.580 2009.000 3490.860 2009.280 ;
        RECT 3491.200 2009.000 3491.480 2009.280 ;
        RECT 3491.820 2009.000 3492.100 2009.280 ;
        RECT 3492.440 2009.000 3492.720 2009.280 ;
        RECT 3493.060 2009.000 3493.340 2009.280 ;
        RECT 3493.680 2009.000 3493.960 2009.280 ;
        RECT 3489.960 2008.380 3490.240 2008.660 ;
        RECT 3490.580 2008.380 3490.860 2008.660 ;
        RECT 3491.200 2008.380 3491.480 2008.660 ;
        RECT 3491.820 2008.380 3492.100 2008.660 ;
        RECT 3492.440 2008.380 3492.720 2008.660 ;
        RECT 3493.060 2008.380 3493.340 2008.660 ;
        RECT 3493.680 2008.380 3493.960 2008.660 ;
        RECT 3489.960 2007.760 3490.240 2008.040 ;
        RECT 3490.580 2007.760 3490.860 2008.040 ;
        RECT 3491.200 2007.760 3491.480 2008.040 ;
        RECT 3491.820 2007.760 3492.100 2008.040 ;
        RECT 3492.440 2007.760 3492.720 2008.040 ;
        RECT 3493.060 2007.760 3493.340 2008.040 ;
        RECT 3493.680 2007.760 3493.960 2008.040 ;
        RECT 3489.960 2007.140 3490.240 2007.420 ;
        RECT 3490.580 2007.140 3490.860 2007.420 ;
        RECT 3491.200 2007.140 3491.480 2007.420 ;
        RECT 3491.820 2007.140 3492.100 2007.420 ;
        RECT 3492.440 2007.140 3492.720 2007.420 ;
        RECT 3493.060 2007.140 3493.340 2007.420 ;
        RECT 3493.680 2007.140 3493.960 2007.420 ;
        RECT 3489.960 2006.520 3490.240 2006.800 ;
        RECT 3490.580 2006.520 3490.860 2006.800 ;
        RECT 3491.200 2006.520 3491.480 2006.800 ;
        RECT 3491.820 2006.520 3492.100 2006.800 ;
        RECT 3492.440 2006.520 3492.720 2006.800 ;
        RECT 3493.060 2006.520 3493.340 2006.800 ;
        RECT 3493.680 2006.520 3493.960 2006.800 ;
        RECT 3489.960 2005.900 3490.240 2006.180 ;
        RECT 3490.580 2005.900 3490.860 2006.180 ;
        RECT 3491.200 2005.900 3491.480 2006.180 ;
        RECT 3491.820 2005.900 3492.100 2006.180 ;
        RECT 3492.440 2005.900 3492.720 2006.180 ;
        RECT 3493.060 2005.900 3493.340 2006.180 ;
        RECT 3493.680 2005.900 3493.960 2006.180 ;
        RECT 3489.960 2003.350 3490.240 2003.630 ;
        RECT 3490.580 2003.350 3490.860 2003.630 ;
        RECT 3491.200 2003.350 3491.480 2003.630 ;
        RECT 3491.820 2003.350 3492.100 2003.630 ;
        RECT 3492.440 2003.350 3492.720 2003.630 ;
        RECT 3493.060 2003.350 3493.340 2003.630 ;
        RECT 3493.680 2003.350 3493.960 2003.630 ;
        RECT 3489.960 2002.730 3490.240 2003.010 ;
        RECT 3490.580 2002.730 3490.860 2003.010 ;
        RECT 3491.200 2002.730 3491.480 2003.010 ;
        RECT 3491.820 2002.730 3492.100 2003.010 ;
        RECT 3492.440 2002.730 3492.720 2003.010 ;
        RECT 3493.060 2002.730 3493.340 2003.010 ;
        RECT 3493.680 2002.730 3493.960 2003.010 ;
        RECT 3489.960 2002.110 3490.240 2002.390 ;
        RECT 3490.580 2002.110 3490.860 2002.390 ;
        RECT 3491.200 2002.110 3491.480 2002.390 ;
        RECT 3491.820 2002.110 3492.100 2002.390 ;
        RECT 3492.440 2002.110 3492.720 2002.390 ;
        RECT 3493.060 2002.110 3493.340 2002.390 ;
        RECT 3493.680 2002.110 3493.960 2002.390 ;
        RECT 3489.960 2001.490 3490.240 2001.770 ;
        RECT 3490.580 2001.490 3490.860 2001.770 ;
        RECT 3491.200 2001.490 3491.480 2001.770 ;
        RECT 3491.820 2001.490 3492.100 2001.770 ;
        RECT 3492.440 2001.490 3492.720 2001.770 ;
        RECT 3493.060 2001.490 3493.340 2001.770 ;
        RECT 3493.680 2001.490 3493.960 2001.770 ;
        RECT 3489.960 2000.870 3490.240 2001.150 ;
        RECT 3490.580 2000.870 3490.860 2001.150 ;
        RECT 3491.200 2000.870 3491.480 2001.150 ;
        RECT 3491.820 2000.870 3492.100 2001.150 ;
        RECT 3492.440 2000.870 3492.720 2001.150 ;
        RECT 3493.060 2000.870 3493.340 2001.150 ;
        RECT 3493.680 2000.870 3493.960 2001.150 ;
        RECT 3489.960 2000.250 3490.240 2000.530 ;
        RECT 3490.580 2000.250 3490.860 2000.530 ;
        RECT 3491.200 2000.250 3491.480 2000.530 ;
        RECT 3491.820 2000.250 3492.100 2000.530 ;
        RECT 3492.440 2000.250 3492.720 2000.530 ;
        RECT 3493.060 2000.250 3493.340 2000.530 ;
        RECT 3493.680 2000.250 3493.960 2000.530 ;
        RECT 3489.960 1999.630 3490.240 1999.910 ;
        RECT 3490.580 1999.630 3490.860 1999.910 ;
        RECT 3491.200 1999.630 3491.480 1999.910 ;
        RECT 3491.820 1999.630 3492.100 1999.910 ;
        RECT 3492.440 1999.630 3492.720 1999.910 ;
        RECT 3493.060 1999.630 3493.340 1999.910 ;
        RECT 3493.680 1999.630 3493.960 1999.910 ;
        RECT 3489.960 1999.010 3490.240 1999.290 ;
        RECT 3490.580 1999.010 3490.860 1999.290 ;
        RECT 3491.200 1999.010 3491.480 1999.290 ;
        RECT 3491.820 1999.010 3492.100 1999.290 ;
        RECT 3492.440 1999.010 3492.720 1999.290 ;
        RECT 3493.060 1999.010 3493.340 1999.290 ;
        RECT 3493.680 1999.010 3493.960 1999.290 ;
        RECT 3489.960 1998.390 3490.240 1998.670 ;
        RECT 3490.580 1998.390 3490.860 1998.670 ;
        RECT 3491.200 1998.390 3491.480 1998.670 ;
        RECT 3491.820 1998.390 3492.100 1998.670 ;
        RECT 3492.440 1998.390 3492.720 1998.670 ;
        RECT 3493.060 1998.390 3493.340 1998.670 ;
        RECT 3493.680 1998.390 3493.960 1998.670 ;
        RECT 3489.960 1997.770 3490.240 1998.050 ;
        RECT 3490.580 1997.770 3490.860 1998.050 ;
        RECT 3491.200 1997.770 3491.480 1998.050 ;
        RECT 3491.820 1997.770 3492.100 1998.050 ;
        RECT 3492.440 1997.770 3492.720 1998.050 ;
        RECT 3493.060 1997.770 3493.340 1998.050 ;
        RECT 3493.680 1997.770 3493.960 1998.050 ;
        RECT 3489.960 1997.150 3490.240 1997.430 ;
        RECT 3490.580 1997.150 3490.860 1997.430 ;
        RECT 3491.200 1997.150 3491.480 1997.430 ;
        RECT 3491.820 1997.150 3492.100 1997.430 ;
        RECT 3492.440 1997.150 3492.720 1997.430 ;
        RECT 3493.060 1997.150 3493.340 1997.430 ;
        RECT 3493.680 1997.150 3493.960 1997.430 ;
        RECT 3489.960 1996.530 3490.240 1996.810 ;
        RECT 3490.580 1996.530 3490.860 1996.810 ;
        RECT 3491.200 1996.530 3491.480 1996.810 ;
        RECT 3491.820 1996.530 3492.100 1996.810 ;
        RECT 3492.440 1996.530 3492.720 1996.810 ;
        RECT 3493.060 1996.530 3493.340 1996.810 ;
        RECT 3493.680 1996.530 3493.960 1996.810 ;
        RECT 3489.960 1995.910 3490.240 1996.190 ;
        RECT 3490.580 1995.910 3490.860 1996.190 ;
        RECT 3491.200 1995.910 3491.480 1996.190 ;
        RECT 3491.820 1995.910 3492.100 1996.190 ;
        RECT 3492.440 1995.910 3492.720 1996.190 ;
        RECT 3493.060 1995.910 3493.340 1996.190 ;
        RECT 3493.680 1995.910 3493.960 1996.190 ;
        RECT 3489.960 1995.290 3490.240 1995.570 ;
        RECT 3490.580 1995.290 3490.860 1995.570 ;
        RECT 3491.200 1995.290 3491.480 1995.570 ;
        RECT 3491.820 1995.290 3492.100 1995.570 ;
        RECT 3492.440 1995.290 3492.720 1995.570 ;
        RECT 3493.060 1995.290 3493.340 1995.570 ;
        RECT 3493.680 1995.290 3493.960 1995.570 ;
        RECT 3489.960 1994.670 3490.240 1994.950 ;
        RECT 3490.580 1994.670 3490.860 1994.950 ;
        RECT 3491.200 1994.670 3491.480 1994.950 ;
        RECT 3491.820 1994.670 3492.100 1994.950 ;
        RECT 3492.440 1994.670 3492.720 1994.950 ;
        RECT 3493.060 1994.670 3493.340 1994.950 ;
        RECT 3493.680 1994.670 3493.960 1994.950 ;
        RECT 3489.960 1994.050 3490.240 1994.330 ;
        RECT 3490.580 1994.050 3490.860 1994.330 ;
        RECT 3491.200 1994.050 3491.480 1994.330 ;
        RECT 3491.820 1994.050 3492.100 1994.330 ;
        RECT 3492.440 1994.050 3492.720 1994.330 ;
        RECT 3493.060 1994.050 3493.340 1994.330 ;
        RECT 3493.680 1994.050 3493.960 1994.330 ;
        RECT 3489.960 1990.330 3490.240 1990.610 ;
        RECT 3490.580 1990.330 3490.860 1990.610 ;
        RECT 3491.200 1990.330 3491.480 1990.610 ;
        RECT 3491.820 1990.330 3492.100 1990.610 ;
        RECT 3492.440 1990.330 3492.720 1990.610 ;
        RECT 3493.060 1990.330 3493.340 1990.610 ;
        RECT 3493.680 1990.330 3493.960 1990.610 ;
        RECT 3489.960 1989.710 3490.240 1989.990 ;
        RECT 3490.580 1989.710 3490.860 1989.990 ;
        RECT 3491.200 1989.710 3491.480 1989.990 ;
        RECT 3491.820 1989.710 3492.100 1989.990 ;
        RECT 3492.440 1989.710 3492.720 1989.990 ;
        RECT 3493.060 1989.710 3493.340 1989.990 ;
        RECT 3493.680 1989.710 3493.960 1989.990 ;
        RECT 3489.960 1989.090 3490.240 1989.370 ;
        RECT 3490.580 1989.090 3490.860 1989.370 ;
        RECT 3491.200 1989.090 3491.480 1989.370 ;
        RECT 3491.820 1989.090 3492.100 1989.370 ;
        RECT 3492.440 1989.090 3492.720 1989.370 ;
        RECT 3493.060 1989.090 3493.340 1989.370 ;
        RECT 3493.680 1989.090 3493.960 1989.370 ;
        RECT 3489.960 1988.470 3490.240 1988.750 ;
        RECT 3490.580 1988.470 3490.860 1988.750 ;
        RECT 3491.200 1988.470 3491.480 1988.750 ;
        RECT 3491.820 1988.470 3492.100 1988.750 ;
        RECT 3492.440 1988.470 3492.720 1988.750 ;
        RECT 3493.060 1988.470 3493.340 1988.750 ;
        RECT 3493.680 1988.470 3493.960 1988.750 ;
        RECT 3489.960 1987.850 3490.240 1988.130 ;
        RECT 3490.580 1987.850 3490.860 1988.130 ;
        RECT 3491.200 1987.850 3491.480 1988.130 ;
        RECT 3491.820 1987.850 3492.100 1988.130 ;
        RECT 3492.440 1987.850 3492.720 1988.130 ;
        RECT 3493.060 1987.850 3493.340 1988.130 ;
        RECT 3493.680 1987.850 3493.960 1988.130 ;
        RECT 3489.960 1987.230 3490.240 1987.510 ;
        RECT 3490.580 1987.230 3490.860 1987.510 ;
        RECT 3491.200 1987.230 3491.480 1987.510 ;
        RECT 3491.820 1987.230 3492.100 1987.510 ;
        RECT 3492.440 1987.230 3492.720 1987.510 ;
        RECT 3493.060 1987.230 3493.340 1987.510 ;
        RECT 3493.680 1987.230 3493.960 1987.510 ;
        RECT 3489.960 1986.610 3490.240 1986.890 ;
        RECT 3490.580 1986.610 3490.860 1986.890 ;
        RECT 3491.200 1986.610 3491.480 1986.890 ;
        RECT 3491.820 1986.610 3492.100 1986.890 ;
        RECT 3492.440 1986.610 3492.720 1986.890 ;
        RECT 3493.060 1986.610 3493.340 1986.890 ;
        RECT 3493.680 1986.610 3493.960 1986.890 ;
        RECT 3489.960 1985.990 3490.240 1986.270 ;
        RECT 3490.580 1985.990 3490.860 1986.270 ;
        RECT 3491.200 1985.990 3491.480 1986.270 ;
        RECT 3491.820 1985.990 3492.100 1986.270 ;
        RECT 3492.440 1985.990 3492.720 1986.270 ;
        RECT 3493.060 1985.990 3493.340 1986.270 ;
        RECT 3493.680 1985.990 3493.960 1986.270 ;
        RECT 3489.960 1985.370 3490.240 1985.650 ;
        RECT 3490.580 1985.370 3490.860 1985.650 ;
        RECT 3491.200 1985.370 3491.480 1985.650 ;
        RECT 3491.820 1985.370 3492.100 1985.650 ;
        RECT 3492.440 1985.370 3492.720 1985.650 ;
        RECT 3493.060 1985.370 3493.340 1985.650 ;
        RECT 3493.680 1985.370 3493.960 1985.650 ;
        RECT 3489.960 1984.750 3490.240 1985.030 ;
        RECT 3490.580 1984.750 3490.860 1985.030 ;
        RECT 3491.200 1984.750 3491.480 1985.030 ;
        RECT 3491.820 1984.750 3492.100 1985.030 ;
        RECT 3492.440 1984.750 3492.720 1985.030 ;
        RECT 3493.060 1984.750 3493.340 1985.030 ;
        RECT 3493.680 1984.750 3493.960 1985.030 ;
        RECT 3489.960 1984.130 3490.240 1984.410 ;
        RECT 3490.580 1984.130 3490.860 1984.410 ;
        RECT 3491.200 1984.130 3491.480 1984.410 ;
        RECT 3491.820 1984.130 3492.100 1984.410 ;
        RECT 3492.440 1984.130 3492.720 1984.410 ;
        RECT 3493.060 1984.130 3493.340 1984.410 ;
        RECT 3493.680 1984.130 3493.960 1984.410 ;
        RECT 3489.960 1983.510 3490.240 1983.790 ;
        RECT 3490.580 1983.510 3490.860 1983.790 ;
        RECT 3491.200 1983.510 3491.480 1983.790 ;
        RECT 3491.820 1983.510 3492.100 1983.790 ;
        RECT 3492.440 1983.510 3492.720 1983.790 ;
        RECT 3493.060 1983.510 3493.340 1983.790 ;
        RECT 3493.680 1983.510 3493.960 1983.790 ;
        RECT 3489.960 1982.890 3490.240 1983.170 ;
        RECT 3490.580 1982.890 3490.860 1983.170 ;
        RECT 3491.200 1982.890 3491.480 1983.170 ;
        RECT 3491.820 1982.890 3492.100 1983.170 ;
        RECT 3492.440 1982.890 3492.720 1983.170 ;
        RECT 3493.060 1982.890 3493.340 1983.170 ;
        RECT 3493.680 1982.890 3493.960 1983.170 ;
        RECT 3489.960 1982.270 3490.240 1982.550 ;
        RECT 3490.580 1982.270 3490.860 1982.550 ;
        RECT 3491.200 1982.270 3491.480 1982.550 ;
        RECT 3491.820 1982.270 3492.100 1982.550 ;
        RECT 3492.440 1982.270 3492.720 1982.550 ;
        RECT 3493.060 1982.270 3493.340 1982.550 ;
        RECT 3493.680 1982.270 3493.960 1982.550 ;
        RECT 3489.960 1981.650 3490.240 1981.930 ;
        RECT 3490.580 1981.650 3490.860 1981.930 ;
        RECT 3491.200 1981.650 3491.480 1981.930 ;
        RECT 3491.820 1981.650 3492.100 1981.930 ;
        RECT 3492.440 1981.650 3492.720 1981.930 ;
        RECT 3493.060 1981.650 3493.340 1981.930 ;
        RECT 3493.680 1981.650 3493.960 1981.930 ;
        RECT 3490.720 1961.865 3491.000 1962.145 ;
        RECT 3492.220 1961.865 3492.500 1962.145 ;
        RECT 3493.720 1961.865 3494.000 1962.145 ;
        RECT 3490.720 1960.865 3491.000 1961.145 ;
        RECT 3492.220 1960.865 3492.500 1961.145 ;
        RECT 3493.720 1960.865 3494.000 1961.145 ;
        RECT 3490.220 1816.890 3490.500 1817.170 ;
        RECT 3491.720 1816.890 3492.000 1817.170 ;
        RECT 3493.220 1816.890 3493.500 1817.170 ;
        RECT 3490.720 1781.865 3491.000 1782.145 ;
        RECT 3492.220 1781.865 3492.500 1782.145 ;
        RECT 3493.720 1781.865 3494.000 1782.145 ;
        RECT 3490.720 1780.865 3491.000 1781.145 ;
        RECT 3492.220 1780.865 3492.500 1781.145 ;
        RECT 3493.720 1780.865 3494.000 1781.145 ;
        RECT 3490.220 1746.890 3490.500 1747.170 ;
        RECT 3491.720 1746.890 3492.000 1747.170 ;
        RECT 3493.220 1746.890 3493.500 1747.170 ;
        RECT 396.040 1654.920 396.320 1655.200 ;
        RECT 396.660 1654.920 396.940 1655.200 ;
        RECT 397.280 1654.920 397.560 1655.200 ;
        RECT 397.900 1654.920 398.180 1655.200 ;
        RECT 398.520 1654.920 398.800 1655.200 ;
        RECT 399.140 1654.920 399.420 1655.200 ;
        RECT 399.760 1654.920 400.040 1655.200 ;
        RECT 396.040 1654.300 396.320 1654.580 ;
        RECT 396.660 1654.300 396.940 1654.580 ;
        RECT 397.280 1654.300 397.560 1654.580 ;
        RECT 397.900 1654.300 398.180 1654.580 ;
        RECT 398.520 1654.300 398.800 1654.580 ;
        RECT 399.140 1654.300 399.420 1654.580 ;
        RECT 399.760 1654.300 400.040 1654.580 ;
        RECT 396.040 1653.680 396.320 1653.960 ;
        RECT 396.660 1653.680 396.940 1653.960 ;
        RECT 397.280 1653.680 397.560 1653.960 ;
        RECT 397.900 1653.680 398.180 1653.960 ;
        RECT 398.520 1653.680 398.800 1653.960 ;
        RECT 399.140 1653.680 399.420 1653.960 ;
        RECT 399.760 1653.680 400.040 1653.960 ;
        RECT 396.040 1653.060 396.320 1653.340 ;
        RECT 396.660 1653.060 396.940 1653.340 ;
        RECT 397.280 1653.060 397.560 1653.340 ;
        RECT 397.900 1653.060 398.180 1653.340 ;
        RECT 398.520 1653.060 398.800 1653.340 ;
        RECT 399.140 1653.060 399.420 1653.340 ;
        RECT 399.760 1653.060 400.040 1653.340 ;
        RECT 396.040 1652.440 396.320 1652.720 ;
        RECT 396.660 1652.440 396.940 1652.720 ;
        RECT 397.280 1652.440 397.560 1652.720 ;
        RECT 397.900 1652.440 398.180 1652.720 ;
        RECT 398.520 1652.440 398.800 1652.720 ;
        RECT 399.140 1652.440 399.420 1652.720 ;
        RECT 399.760 1652.440 400.040 1652.720 ;
        RECT 396.040 1651.820 396.320 1652.100 ;
        RECT 396.660 1651.820 396.940 1652.100 ;
        RECT 397.280 1651.820 397.560 1652.100 ;
        RECT 397.900 1651.820 398.180 1652.100 ;
        RECT 398.520 1651.820 398.800 1652.100 ;
        RECT 399.140 1651.820 399.420 1652.100 ;
        RECT 399.760 1651.820 400.040 1652.100 ;
        RECT 396.040 1651.200 396.320 1651.480 ;
        RECT 396.660 1651.200 396.940 1651.480 ;
        RECT 397.280 1651.200 397.560 1651.480 ;
        RECT 397.900 1651.200 398.180 1651.480 ;
        RECT 398.520 1651.200 398.800 1651.480 ;
        RECT 399.140 1651.200 399.420 1651.480 ;
        RECT 399.760 1651.200 400.040 1651.480 ;
        RECT 531.035 1654.160 531.315 1654.440 ;
        RECT 532.035 1654.160 532.315 1654.440 ;
        RECT 531.035 1652.660 531.315 1652.940 ;
        RECT 532.035 1652.660 532.315 1652.940 ;
        RECT 531.035 1651.160 531.315 1651.440 ;
        RECT 532.035 1651.160 532.315 1651.440 ;
        RECT 441.035 1647.160 441.315 1647.440 ;
        RECT 442.035 1647.160 442.315 1647.440 ;
        RECT 441.035 1645.660 441.315 1645.940 ;
        RECT 442.035 1645.660 442.315 1645.940 ;
        RECT 441.035 1644.160 441.315 1644.440 ;
        RECT 442.035 1644.160 442.315 1644.440 ;
        RECT 711.035 1654.160 711.315 1654.440 ;
        RECT 712.035 1654.160 712.315 1654.440 ;
        RECT 711.035 1652.660 711.315 1652.940 ;
        RECT 712.035 1652.660 712.315 1652.940 ;
        RECT 711.035 1651.160 711.315 1651.440 ;
        RECT 712.035 1651.160 712.315 1651.440 ;
        RECT 790.890 1654.920 791.170 1655.200 ;
        RECT 791.510 1654.920 791.790 1655.200 ;
        RECT 792.130 1654.920 792.410 1655.200 ;
        RECT 792.750 1654.920 793.030 1655.200 ;
        RECT 790.890 1654.300 791.170 1654.580 ;
        RECT 791.510 1654.300 791.790 1654.580 ;
        RECT 792.130 1654.300 792.410 1654.580 ;
        RECT 792.750 1654.300 793.030 1654.580 ;
        RECT 790.890 1653.680 791.170 1653.960 ;
        RECT 791.510 1653.680 791.790 1653.960 ;
        RECT 792.130 1653.680 792.410 1653.960 ;
        RECT 792.750 1653.680 793.030 1653.960 ;
        RECT 790.890 1653.060 791.170 1653.340 ;
        RECT 791.510 1653.060 791.790 1653.340 ;
        RECT 792.130 1653.060 792.410 1653.340 ;
        RECT 792.750 1653.060 793.030 1653.340 ;
        RECT 790.890 1652.440 791.170 1652.720 ;
        RECT 791.510 1652.440 791.790 1652.720 ;
        RECT 792.130 1652.440 792.410 1652.720 ;
        RECT 792.750 1652.440 793.030 1652.720 ;
        RECT 790.890 1651.820 791.170 1652.100 ;
        RECT 791.510 1651.820 791.790 1652.100 ;
        RECT 792.130 1651.820 792.410 1652.100 ;
        RECT 792.750 1651.820 793.030 1652.100 ;
        RECT 790.890 1651.200 791.170 1651.480 ;
        RECT 791.510 1651.200 791.790 1651.480 ;
        RECT 792.130 1651.200 792.410 1651.480 ;
        RECT 792.750 1651.200 793.030 1651.480 ;
        RECT 621.035 1647.160 621.315 1647.440 ;
        RECT 622.035 1647.160 622.315 1647.440 ;
        RECT 621.035 1645.660 621.315 1645.940 ;
        RECT 622.035 1645.660 622.315 1645.940 ;
        RECT 621.035 1644.160 621.315 1644.440 ;
        RECT 622.035 1644.160 622.315 1644.440 ;
        RECT 785.790 1647.920 786.070 1648.200 ;
        RECT 786.410 1647.920 786.690 1648.200 ;
        RECT 787.030 1647.920 787.310 1648.200 ;
        RECT 787.650 1647.920 787.930 1648.200 ;
        RECT 785.790 1647.300 786.070 1647.580 ;
        RECT 786.410 1647.300 786.690 1647.580 ;
        RECT 787.030 1647.300 787.310 1647.580 ;
        RECT 787.650 1647.300 787.930 1647.580 ;
        RECT 785.790 1646.680 786.070 1646.960 ;
        RECT 786.410 1646.680 786.690 1646.960 ;
        RECT 787.030 1646.680 787.310 1646.960 ;
        RECT 787.650 1646.680 787.930 1646.960 ;
        RECT 785.790 1646.060 786.070 1646.340 ;
        RECT 786.410 1646.060 786.690 1646.340 ;
        RECT 787.030 1646.060 787.310 1646.340 ;
        RECT 787.650 1646.060 787.930 1646.340 ;
        RECT 785.790 1645.440 786.070 1645.720 ;
        RECT 786.410 1645.440 786.690 1645.720 ;
        RECT 787.030 1645.440 787.310 1645.720 ;
        RECT 787.650 1645.440 787.930 1645.720 ;
        RECT 785.790 1644.820 786.070 1645.100 ;
        RECT 786.410 1644.820 786.690 1645.100 ;
        RECT 787.030 1644.820 787.310 1645.100 ;
        RECT 787.650 1644.820 787.930 1645.100 ;
        RECT 785.790 1644.200 786.070 1644.480 ;
        RECT 786.410 1644.200 786.690 1644.480 ;
        RECT 787.030 1644.200 787.310 1644.480 ;
        RECT 787.650 1644.200 787.930 1644.480 ;
        RECT 396.500 1572.830 396.780 1573.110 ;
        RECT 398.000 1572.830 398.280 1573.110 ;
        RECT 399.500 1572.830 399.780 1573.110 ;
        RECT 786.050 1591.840 786.330 1592.120 ;
        RECT 787.550 1591.840 787.830 1592.120 ;
        RECT 786.050 1584.850 786.330 1585.130 ;
        RECT 787.550 1584.850 787.830 1585.130 ;
        RECT 786.050 1577.860 786.330 1578.140 ;
        RECT 787.550 1577.860 787.830 1578.140 ;
        RECT 396.500 1537.830 396.780 1538.110 ;
        RECT 398.000 1537.830 398.280 1538.110 ;
        RECT 399.500 1537.830 399.780 1538.110 ;
        RECT 396.040 1535.650 396.320 1535.930 ;
        RECT 396.660 1535.650 396.940 1535.930 ;
        RECT 397.280 1535.650 397.560 1535.930 ;
        RECT 397.900 1535.650 398.180 1535.930 ;
        RECT 398.520 1535.650 398.800 1535.930 ;
        RECT 399.140 1535.650 399.420 1535.930 ;
        RECT 399.760 1535.650 400.040 1535.930 ;
        RECT 396.040 1535.030 396.320 1535.310 ;
        RECT 396.660 1535.030 396.940 1535.310 ;
        RECT 397.280 1535.030 397.560 1535.310 ;
        RECT 397.900 1535.030 398.180 1535.310 ;
        RECT 398.520 1535.030 398.800 1535.310 ;
        RECT 399.140 1535.030 399.420 1535.310 ;
        RECT 399.760 1535.030 400.040 1535.310 ;
        RECT 396.040 1534.410 396.320 1534.690 ;
        RECT 396.660 1534.410 396.940 1534.690 ;
        RECT 397.280 1534.410 397.560 1534.690 ;
        RECT 397.900 1534.410 398.180 1534.690 ;
        RECT 398.520 1534.410 398.800 1534.690 ;
        RECT 399.140 1534.410 399.420 1534.690 ;
        RECT 399.760 1534.410 400.040 1534.690 ;
        RECT 396.040 1533.790 396.320 1534.070 ;
        RECT 396.660 1533.790 396.940 1534.070 ;
        RECT 397.280 1533.790 397.560 1534.070 ;
        RECT 397.900 1533.790 398.180 1534.070 ;
        RECT 398.520 1533.790 398.800 1534.070 ;
        RECT 399.140 1533.790 399.420 1534.070 ;
        RECT 399.760 1533.790 400.040 1534.070 ;
        RECT 396.040 1533.170 396.320 1533.450 ;
        RECT 396.660 1533.170 396.940 1533.450 ;
        RECT 397.280 1533.170 397.560 1533.450 ;
        RECT 397.900 1533.170 398.180 1533.450 ;
        RECT 398.520 1533.170 398.800 1533.450 ;
        RECT 399.140 1533.170 399.420 1533.450 ;
        RECT 399.760 1533.170 400.040 1533.450 ;
        RECT 396.040 1532.550 396.320 1532.830 ;
        RECT 396.660 1532.550 396.940 1532.830 ;
        RECT 397.280 1532.550 397.560 1532.830 ;
        RECT 397.900 1532.550 398.180 1532.830 ;
        RECT 398.520 1532.550 398.800 1532.830 ;
        RECT 399.140 1532.550 399.420 1532.830 ;
        RECT 399.760 1532.550 400.040 1532.830 ;
        RECT 396.040 1531.930 396.320 1532.210 ;
        RECT 396.660 1531.930 396.940 1532.210 ;
        RECT 397.280 1531.930 397.560 1532.210 ;
        RECT 397.900 1531.930 398.180 1532.210 ;
        RECT 398.520 1531.930 398.800 1532.210 ;
        RECT 399.140 1531.930 399.420 1532.210 ;
        RECT 399.760 1531.930 400.040 1532.210 ;
        RECT 581.100 1535.650 581.380 1535.930 ;
        RECT 581.720 1535.650 582.000 1535.930 ;
        RECT 581.100 1535.030 581.380 1535.310 ;
        RECT 581.720 1535.030 582.000 1535.310 ;
        RECT 581.100 1534.410 581.380 1534.690 ;
        RECT 581.720 1534.410 582.000 1534.690 ;
        RECT 581.100 1533.790 581.380 1534.070 ;
        RECT 581.720 1533.790 582.000 1534.070 ;
        RECT 581.100 1533.170 581.380 1533.450 ;
        RECT 581.720 1533.170 582.000 1533.450 ;
        RECT 581.100 1532.550 581.380 1532.830 ;
        RECT 581.720 1532.550 582.000 1532.830 ;
        RECT 581.100 1531.930 581.380 1532.210 ;
        RECT 581.720 1531.930 582.000 1532.210 ;
        RECT 573.125 1528.650 573.405 1528.930 ;
        RECT 573.745 1528.650 574.025 1528.930 ;
        RECT 573.125 1528.030 573.405 1528.310 ;
        RECT 573.745 1528.030 574.025 1528.310 ;
        RECT 573.125 1527.410 573.405 1527.690 ;
        RECT 573.745 1527.410 574.025 1527.690 ;
        RECT 573.125 1526.790 573.405 1527.070 ;
        RECT 573.745 1526.790 574.025 1527.070 ;
        RECT 573.125 1526.170 573.405 1526.450 ;
        RECT 573.745 1526.170 574.025 1526.450 ;
        RECT 573.125 1525.550 573.405 1525.830 ;
        RECT 573.745 1525.550 574.025 1525.830 ;
        RECT 573.125 1524.930 573.405 1525.210 ;
        RECT 573.745 1524.930 574.025 1525.210 ;
        RECT 597.050 1535.650 597.330 1535.930 ;
        RECT 597.670 1535.650 597.950 1535.930 ;
        RECT 597.050 1535.030 597.330 1535.310 ;
        RECT 597.670 1535.030 597.950 1535.310 ;
        RECT 597.050 1534.410 597.330 1534.690 ;
        RECT 597.670 1534.410 597.950 1534.690 ;
        RECT 597.050 1533.790 597.330 1534.070 ;
        RECT 597.670 1533.790 597.950 1534.070 ;
        RECT 597.050 1533.170 597.330 1533.450 ;
        RECT 597.670 1533.170 597.950 1533.450 ;
        RECT 597.050 1532.550 597.330 1532.830 ;
        RECT 597.670 1532.550 597.950 1532.830 ;
        RECT 597.050 1531.930 597.330 1532.210 ;
        RECT 597.670 1531.930 597.950 1532.210 ;
        RECT 589.075 1528.650 589.355 1528.930 ;
        RECT 589.695 1528.650 589.975 1528.930 ;
        RECT 589.075 1528.030 589.355 1528.310 ;
        RECT 589.695 1528.030 589.975 1528.310 ;
        RECT 589.075 1527.410 589.355 1527.690 ;
        RECT 589.695 1527.410 589.975 1527.690 ;
        RECT 589.075 1526.790 589.355 1527.070 ;
        RECT 589.695 1526.790 589.975 1527.070 ;
        RECT 589.075 1526.170 589.355 1526.450 ;
        RECT 589.695 1526.170 589.975 1526.450 ;
        RECT 589.075 1525.550 589.355 1525.830 ;
        RECT 589.695 1525.550 589.975 1525.830 ;
        RECT 589.075 1524.930 589.355 1525.210 ;
        RECT 589.695 1524.930 589.975 1525.210 ;
        RECT 613.000 1535.650 613.280 1535.930 ;
        RECT 613.620 1535.650 613.900 1535.930 ;
        RECT 613.000 1535.030 613.280 1535.310 ;
        RECT 613.620 1535.030 613.900 1535.310 ;
        RECT 613.000 1534.410 613.280 1534.690 ;
        RECT 613.620 1534.410 613.900 1534.690 ;
        RECT 613.000 1533.790 613.280 1534.070 ;
        RECT 613.620 1533.790 613.900 1534.070 ;
        RECT 613.000 1533.170 613.280 1533.450 ;
        RECT 613.620 1533.170 613.900 1533.450 ;
        RECT 613.000 1532.550 613.280 1532.830 ;
        RECT 613.620 1532.550 613.900 1532.830 ;
        RECT 613.000 1531.930 613.280 1532.210 ;
        RECT 613.620 1531.930 613.900 1532.210 ;
        RECT 605.025 1528.650 605.305 1528.930 ;
        RECT 605.645 1528.650 605.925 1528.930 ;
        RECT 605.025 1528.030 605.305 1528.310 ;
        RECT 605.645 1528.030 605.925 1528.310 ;
        RECT 605.025 1527.410 605.305 1527.690 ;
        RECT 605.645 1527.410 605.925 1527.690 ;
        RECT 605.025 1526.790 605.305 1527.070 ;
        RECT 605.645 1526.790 605.925 1527.070 ;
        RECT 605.025 1526.170 605.305 1526.450 ;
        RECT 605.645 1526.170 605.925 1526.450 ;
        RECT 605.025 1525.550 605.305 1525.830 ;
        RECT 605.645 1525.550 605.925 1525.830 ;
        RECT 605.025 1524.930 605.305 1525.210 ;
        RECT 605.645 1524.930 605.925 1525.210 ;
        RECT 620.975 1528.650 621.255 1528.930 ;
        RECT 621.595 1528.650 621.875 1528.930 ;
        RECT 620.975 1528.030 621.255 1528.310 ;
        RECT 621.595 1528.030 621.875 1528.310 ;
        RECT 620.975 1527.410 621.255 1527.690 ;
        RECT 621.595 1527.410 621.875 1527.690 ;
        RECT 620.975 1526.790 621.255 1527.070 ;
        RECT 621.595 1526.790 621.875 1527.070 ;
        RECT 620.975 1526.170 621.255 1526.450 ;
        RECT 621.595 1526.170 621.875 1526.450 ;
        RECT 620.975 1525.550 621.255 1525.830 ;
        RECT 621.595 1525.550 621.875 1525.830 ;
        RECT 620.975 1524.930 621.255 1525.210 ;
        RECT 621.595 1524.930 621.875 1525.210 ;
        RECT 786.050 1570.870 786.330 1571.150 ;
        RECT 787.550 1570.870 787.830 1571.150 ;
        RECT 891.035 1654.160 891.315 1654.440 ;
        RECT 892.035 1654.160 892.315 1654.440 ;
        RECT 891.035 1652.660 891.315 1652.940 ;
        RECT 892.035 1652.660 892.315 1652.940 ;
        RECT 891.035 1651.160 891.315 1651.440 ;
        RECT 892.035 1651.160 892.315 1651.440 ;
        RECT 801.035 1647.160 801.315 1647.440 ;
        RECT 802.035 1647.160 802.315 1647.440 ;
        RECT 801.035 1645.660 801.315 1645.940 ;
        RECT 802.035 1645.660 802.315 1645.940 ;
        RECT 801.035 1644.160 801.315 1644.440 ;
        RECT 802.035 1644.160 802.315 1644.440 ;
        RECT 1071.035 1654.160 1071.315 1654.440 ;
        RECT 1072.035 1654.160 1072.315 1654.440 ;
        RECT 1071.035 1652.660 1071.315 1652.940 ;
        RECT 1072.035 1652.660 1072.315 1652.940 ;
        RECT 1071.035 1651.160 1071.315 1651.440 ;
        RECT 1072.035 1651.160 1072.315 1651.440 ;
        RECT 981.035 1647.160 981.315 1647.440 ;
        RECT 982.035 1647.160 982.315 1647.440 ;
        RECT 981.035 1645.660 981.315 1645.940 ;
        RECT 982.035 1645.660 982.315 1645.940 ;
        RECT 981.035 1644.160 981.315 1644.440 ;
        RECT 982.035 1644.160 982.315 1644.440 ;
        RECT 1251.035 1654.160 1251.315 1654.440 ;
        RECT 1252.035 1654.160 1252.315 1654.440 ;
        RECT 1251.035 1652.660 1251.315 1652.940 ;
        RECT 1252.035 1652.660 1252.315 1652.940 ;
        RECT 1251.035 1651.160 1251.315 1651.440 ;
        RECT 1252.035 1651.160 1252.315 1651.440 ;
        RECT 1161.035 1647.160 1161.315 1647.440 ;
        RECT 1162.035 1647.160 1162.315 1647.440 ;
        RECT 1161.035 1645.660 1161.315 1645.940 ;
        RECT 1162.035 1645.660 1162.315 1645.940 ;
        RECT 1161.035 1644.160 1161.315 1644.440 ;
        RECT 1162.035 1644.160 1162.315 1644.440 ;
        RECT 1431.035 1654.160 1431.315 1654.440 ;
        RECT 1432.035 1654.160 1432.315 1654.440 ;
        RECT 1431.035 1652.660 1431.315 1652.940 ;
        RECT 1432.035 1652.660 1432.315 1652.940 ;
        RECT 1431.035 1651.160 1431.315 1651.440 ;
        RECT 1432.035 1651.160 1432.315 1651.440 ;
        RECT 1341.035 1647.160 1341.315 1647.440 ;
        RECT 1342.035 1647.160 1342.315 1647.440 ;
        RECT 1341.035 1645.660 1341.315 1645.940 ;
        RECT 1342.035 1645.660 1342.315 1645.940 ;
        RECT 1341.035 1644.160 1341.315 1644.440 ;
        RECT 1342.035 1644.160 1342.315 1644.440 ;
        RECT 1611.035 1654.160 1611.315 1654.440 ;
        RECT 1612.035 1654.160 1612.315 1654.440 ;
        RECT 1611.035 1652.660 1611.315 1652.940 ;
        RECT 1612.035 1652.660 1612.315 1652.940 ;
        RECT 1611.035 1651.160 1611.315 1651.440 ;
        RECT 1612.035 1651.160 1612.315 1651.440 ;
        RECT 1521.035 1647.160 1521.315 1647.440 ;
        RECT 1522.035 1647.160 1522.315 1647.440 ;
        RECT 1521.035 1645.660 1521.315 1645.940 ;
        RECT 1522.035 1645.660 1522.315 1645.940 ;
        RECT 1521.035 1644.160 1521.315 1644.440 ;
        RECT 1522.035 1644.160 1522.315 1644.440 ;
        RECT 1791.035 1654.160 1791.315 1654.440 ;
        RECT 1792.035 1654.160 1792.315 1654.440 ;
        RECT 1791.035 1652.660 1791.315 1652.940 ;
        RECT 1792.035 1652.660 1792.315 1652.940 ;
        RECT 1791.035 1651.160 1791.315 1651.440 ;
        RECT 1792.035 1651.160 1792.315 1651.440 ;
        RECT 1701.035 1647.160 1701.315 1647.440 ;
        RECT 1702.035 1647.160 1702.315 1647.440 ;
        RECT 1701.035 1645.660 1701.315 1645.940 ;
        RECT 1702.035 1645.660 1702.315 1645.940 ;
        RECT 1701.035 1644.160 1701.315 1644.440 ;
        RECT 1702.035 1644.160 1702.315 1644.440 ;
        RECT 1881.035 1647.160 1881.315 1647.440 ;
        RECT 1882.035 1647.160 1882.315 1647.440 ;
        RECT 1881.035 1645.660 1881.315 1645.940 ;
        RECT 1882.035 1645.660 1882.315 1645.940 ;
        RECT 1881.035 1644.160 1881.315 1644.440 ;
        RECT 1882.035 1644.160 1882.315 1644.440 ;
        RECT 1906.550 1654.920 1906.830 1655.200 ;
        RECT 1907.170 1654.920 1907.450 1655.200 ;
        RECT 1907.790 1654.920 1908.070 1655.200 ;
        RECT 1908.410 1654.920 1908.690 1655.200 ;
        RECT 1906.550 1654.300 1906.830 1654.580 ;
        RECT 1907.170 1654.300 1907.450 1654.580 ;
        RECT 1907.790 1654.300 1908.070 1654.580 ;
        RECT 1908.410 1654.300 1908.690 1654.580 ;
        RECT 1906.550 1653.680 1906.830 1653.960 ;
        RECT 1907.170 1653.680 1907.450 1653.960 ;
        RECT 1907.790 1653.680 1908.070 1653.960 ;
        RECT 1908.410 1653.680 1908.690 1653.960 ;
        RECT 1906.550 1653.060 1906.830 1653.340 ;
        RECT 1907.170 1653.060 1907.450 1653.340 ;
        RECT 1907.790 1653.060 1908.070 1653.340 ;
        RECT 1908.410 1653.060 1908.690 1653.340 ;
        RECT 1906.550 1652.440 1906.830 1652.720 ;
        RECT 1907.170 1652.440 1907.450 1652.720 ;
        RECT 1907.790 1652.440 1908.070 1652.720 ;
        RECT 1908.410 1652.440 1908.690 1652.720 ;
        RECT 1906.550 1651.820 1906.830 1652.100 ;
        RECT 1907.170 1651.820 1907.450 1652.100 ;
        RECT 1907.790 1651.820 1908.070 1652.100 ;
        RECT 1908.410 1651.820 1908.690 1652.100 ;
        RECT 1906.550 1651.200 1906.830 1651.480 ;
        RECT 1907.170 1651.200 1907.450 1651.480 ;
        RECT 1907.790 1651.200 1908.070 1651.480 ;
        RECT 1908.410 1651.200 1908.690 1651.480 ;
        RECT 791.150 1588.345 791.430 1588.625 ;
        RECT 792.650 1588.345 792.930 1588.625 ;
        RECT 791.150 1581.355 791.430 1581.635 ;
        RECT 792.650 1581.355 792.930 1581.635 ;
        RECT 791.150 1574.365 791.430 1574.645 ;
        RECT 792.650 1574.365 792.930 1574.645 ;
        RECT 790.890 1535.350 791.170 1535.630 ;
        RECT 791.510 1535.350 791.790 1535.630 ;
        RECT 792.130 1535.350 792.410 1535.630 ;
        RECT 792.750 1535.350 793.030 1535.630 ;
        RECT 790.890 1534.730 791.170 1535.010 ;
        RECT 791.510 1534.730 791.790 1535.010 ;
        RECT 792.130 1534.730 792.410 1535.010 ;
        RECT 792.750 1534.730 793.030 1535.010 ;
        RECT 790.890 1534.110 791.170 1534.390 ;
        RECT 791.510 1534.110 791.790 1534.390 ;
        RECT 792.130 1534.110 792.410 1534.390 ;
        RECT 792.750 1534.110 793.030 1534.390 ;
        RECT 790.890 1533.490 791.170 1533.770 ;
        RECT 791.510 1533.490 791.790 1533.770 ;
        RECT 792.130 1533.490 792.410 1533.770 ;
        RECT 792.750 1533.490 793.030 1533.770 ;
        RECT 790.890 1532.870 791.170 1533.150 ;
        RECT 791.510 1532.870 791.790 1533.150 ;
        RECT 792.130 1532.870 792.410 1533.150 ;
        RECT 792.750 1532.870 793.030 1533.150 ;
        RECT 790.890 1532.250 791.170 1532.530 ;
        RECT 791.510 1532.250 791.790 1532.530 ;
        RECT 792.130 1532.250 792.410 1532.530 ;
        RECT 792.750 1532.250 793.030 1532.530 ;
        RECT 790.890 1531.630 791.170 1531.910 ;
        RECT 791.510 1531.630 791.790 1531.910 ;
        RECT 792.130 1531.630 792.410 1531.910 ;
        RECT 792.750 1531.630 793.030 1531.910 ;
        RECT 1971.035 1654.160 1971.315 1654.440 ;
        RECT 1972.035 1654.160 1972.315 1654.440 ;
        RECT 1971.035 1652.660 1971.315 1652.940 ;
        RECT 1972.035 1652.660 1972.315 1652.940 ;
        RECT 1971.035 1651.160 1971.315 1651.440 ;
        RECT 1972.035 1651.160 1972.315 1651.440 ;
        RECT 1906.910 1588.355 1907.190 1588.635 ;
        RECT 1908.410 1588.355 1908.690 1588.635 ;
        RECT 1906.910 1581.365 1907.190 1581.645 ;
        RECT 1908.410 1581.365 1908.690 1581.645 ;
        RECT 1906.910 1574.375 1907.190 1574.655 ;
        RECT 1908.410 1574.375 1908.690 1574.655 ;
        RECT 1906.550 1535.350 1906.830 1535.630 ;
        RECT 1907.170 1535.350 1907.450 1535.630 ;
        RECT 1907.790 1535.350 1908.070 1535.630 ;
        RECT 1908.410 1535.350 1908.690 1535.630 ;
        RECT 1906.550 1534.730 1906.830 1535.010 ;
        RECT 1907.170 1534.730 1907.450 1535.010 ;
        RECT 1907.790 1534.730 1908.070 1535.010 ;
        RECT 1908.410 1534.730 1908.690 1535.010 ;
        RECT 1906.550 1534.110 1906.830 1534.390 ;
        RECT 1907.170 1534.110 1907.450 1534.390 ;
        RECT 1907.790 1534.110 1908.070 1534.390 ;
        RECT 1908.410 1534.110 1908.690 1534.390 ;
        RECT 1906.550 1533.490 1906.830 1533.770 ;
        RECT 1907.170 1533.490 1907.450 1533.770 ;
        RECT 1907.790 1533.490 1908.070 1533.770 ;
        RECT 1908.410 1533.490 1908.690 1533.770 ;
        RECT 1906.550 1532.870 1906.830 1533.150 ;
        RECT 1907.170 1532.870 1907.450 1533.150 ;
        RECT 1907.790 1532.870 1908.070 1533.150 ;
        RECT 1908.410 1532.870 1908.690 1533.150 ;
        RECT 1906.550 1532.250 1906.830 1532.530 ;
        RECT 1907.170 1532.250 1907.450 1532.530 ;
        RECT 1907.790 1532.250 1908.070 1532.530 ;
        RECT 1908.410 1532.250 1908.690 1532.530 ;
        RECT 1906.550 1531.630 1906.830 1531.910 ;
        RECT 1907.170 1531.630 1907.450 1531.910 ;
        RECT 1907.790 1531.630 1908.070 1531.910 ;
        RECT 1908.410 1531.630 1908.690 1531.910 ;
        RECT 1911.650 1647.920 1911.930 1648.200 ;
        RECT 1912.270 1647.920 1912.550 1648.200 ;
        RECT 1912.890 1647.920 1913.170 1648.200 ;
        RECT 1913.510 1647.920 1913.790 1648.200 ;
        RECT 1911.650 1647.300 1911.930 1647.580 ;
        RECT 1912.270 1647.300 1912.550 1647.580 ;
        RECT 1912.890 1647.300 1913.170 1647.580 ;
        RECT 1913.510 1647.300 1913.790 1647.580 ;
        RECT 1911.650 1646.680 1911.930 1646.960 ;
        RECT 1912.270 1646.680 1912.550 1646.960 ;
        RECT 1912.890 1646.680 1913.170 1646.960 ;
        RECT 1913.510 1646.680 1913.790 1646.960 ;
        RECT 1911.650 1646.060 1911.930 1646.340 ;
        RECT 1912.270 1646.060 1912.550 1646.340 ;
        RECT 1912.890 1646.060 1913.170 1646.340 ;
        RECT 1913.510 1646.060 1913.790 1646.340 ;
        RECT 1911.650 1645.440 1911.930 1645.720 ;
        RECT 1912.270 1645.440 1912.550 1645.720 ;
        RECT 1912.890 1645.440 1913.170 1645.720 ;
        RECT 1913.510 1645.440 1913.790 1645.720 ;
        RECT 1911.650 1644.820 1911.930 1645.100 ;
        RECT 1912.270 1644.820 1912.550 1645.100 ;
        RECT 1912.890 1644.820 1913.170 1645.100 ;
        RECT 1913.510 1644.820 1913.790 1645.100 ;
        RECT 1911.650 1644.200 1911.930 1644.480 ;
        RECT 1912.270 1644.200 1912.550 1644.480 ;
        RECT 1912.890 1644.200 1913.170 1644.480 ;
        RECT 1913.510 1644.200 1913.790 1644.480 ;
        RECT 2151.035 1654.160 2151.315 1654.440 ;
        RECT 2152.035 1654.160 2152.315 1654.440 ;
        RECT 2151.035 1652.660 2151.315 1652.940 ;
        RECT 2152.035 1652.660 2152.315 1652.940 ;
        RECT 2151.035 1651.160 2151.315 1651.440 ;
        RECT 2152.035 1651.160 2152.315 1651.440 ;
        RECT 2061.035 1647.160 2061.315 1647.440 ;
        RECT 2062.035 1647.160 2062.315 1647.440 ;
        RECT 2061.035 1645.660 2061.315 1645.940 ;
        RECT 2062.035 1645.660 2062.315 1645.940 ;
        RECT 2061.035 1644.160 2061.315 1644.440 ;
        RECT 2062.035 1644.160 2062.315 1644.440 ;
        RECT 2331.035 1654.160 2331.315 1654.440 ;
        RECT 2332.035 1654.160 2332.315 1654.440 ;
        RECT 2331.035 1652.660 2331.315 1652.940 ;
        RECT 2332.035 1652.660 2332.315 1652.940 ;
        RECT 2331.035 1651.160 2331.315 1651.440 ;
        RECT 2332.035 1651.160 2332.315 1651.440 ;
        RECT 2241.035 1647.160 2241.315 1647.440 ;
        RECT 2242.035 1647.160 2242.315 1647.440 ;
        RECT 2241.035 1645.660 2241.315 1645.940 ;
        RECT 2242.035 1645.660 2242.315 1645.940 ;
        RECT 2241.035 1644.160 2241.315 1644.440 ;
        RECT 2242.035 1644.160 2242.315 1644.440 ;
        RECT 2511.035 1654.160 2511.315 1654.440 ;
        RECT 2512.035 1654.160 2512.315 1654.440 ;
        RECT 2511.035 1652.660 2511.315 1652.940 ;
        RECT 2512.035 1652.660 2512.315 1652.940 ;
        RECT 2511.035 1651.160 2511.315 1651.440 ;
        RECT 2512.035 1651.160 2512.315 1651.440 ;
        RECT 2421.035 1647.160 2421.315 1647.440 ;
        RECT 2422.035 1647.160 2422.315 1647.440 ;
        RECT 2421.035 1645.660 2421.315 1645.940 ;
        RECT 2422.035 1645.660 2422.315 1645.940 ;
        RECT 2421.035 1644.160 2421.315 1644.440 ;
        RECT 2422.035 1644.160 2422.315 1644.440 ;
        RECT 2691.035 1654.160 2691.315 1654.440 ;
        RECT 2692.035 1654.160 2692.315 1654.440 ;
        RECT 2691.035 1652.660 2691.315 1652.940 ;
        RECT 2692.035 1652.660 2692.315 1652.940 ;
        RECT 2691.035 1651.160 2691.315 1651.440 ;
        RECT 2692.035 1651.160 2692.315 1651.440 ;
        RECT 2601.035 1647.160 2601.315 1647.440 ;
        RECT 2602.035 1647.160 2602.315 1647.440 ;
        RECT 2601.035 1645.660 2601.315 1645.940 ;
        RECT 2602.035 1645.660 2602.315 1645.940 ;
        RECT 2601.035 1644.160 2601.315 1644.440 ;
        RECT 2602.035 1644.160 2602.315 1644.440 ;
        RECT 2871.035 1654.160 2871.315 1654.440 ;
        RECT 2872.035 1654.160 2872.315 1654.440 ;
        RECT 2871.035 1652.660 2871.315 1652.940 ;
        RECT 2872.035 1652.660 2872.315 1652.940 ;
        RECT 2871.035 1651.160 2871.315 1651.440 ;
        RECT 2872.035 1651.160 2872.315 1651.440 ;
        RECT 2781.035 1647.160 2781.315 1647.440 ;
        RECT 2782.035 1647.160 2782.315 1647.440 ;
        RECT 2781.035 1645.660 2781.315 1645.940 ;
        RECT 2782.035 1645.660 2782.315 1645.940 ;
        RECT 2781.035 1644.160 2781.315 1644.440 ;
        RECT 2782.035 1644.160 2782.315 1644.440 ;
        RECT 3051.035 1654.160 3051.315 1654.440 ;
        RECT 3052.035 1654.160 3052.315 1654.440 ;
        RECT 3051.035 1652.660 3051.315 1652.940 ;
        RECT 3052.035 1652.660 3052.315 1652.940 ;
        RECT 3051.035 1651.160 3051.315 1651.440 ;
        RECT 3052.035 1651.160 3052.315 1651.440 ;
        RECT 2961.035 1647.160 2961.315 1647.440 ;
        RECT 2962.035 1647.160 2962.315 1647.440 ;
        RECT 2961.035 1645.660 2961.315 1645.940 ;
        RECT 2962.035 1645.660 2962.315 1645.940 ;
        RECT 2961.035 1644.160 2961.315 1644.440 ;
        RECT 2962.035 1644.160 2962.315 1644.440 ;
        RECT 3231.035 1654.160 3231.315 1654.440 ;
        RECT 3232.035 1654.160 3232.315 1654.440 ;
        RECT 3231.035 1652.660 3231.315 1652.940 ;
        RECT 3232.035 1652.660 3232.315 1652.940 ;
        RECT 3231.035 1651.160 3231.315 1651.440 ;
        RECT 3232.035 1651.160 3232.315 1651.440 ;
        RECT 3141.035 1647.160 3141.315 1647.440 ;
        RECT 3142.035 1647.160 3142.315 1647.440 ;
        RECT 3141.035 1645.660 3141.315 1645.940 ;
        RECT 3142.035 1645.660 3142.315 1645.940 ;
        RECT 3141.035 1644.160 3141.315 1644.440 ;
        RECT 3142.035 1644.160 3142.315 1644.440 ;
        RECT 3411.035 1654.160 3411.315 1654.440 ;
        RECT 3412.035 1654.160 3412.315 1654.440 ;
        RECT 3411.035 1652.660 3411.315 1652.940 ;
        RECT 3412.035 1652.660 3412.315 1652.940 ;
        RECT 3411.035 1651.160 3411.315 1651.440 ;
        RECT 3412.035 1651.160 3412.315 1651.440 ;
        RECT 3490.300 1664.760 3490.580 1665.040 ;
        RECT 3491.800 1664.760 3492.080 1665.040 ;
        RECT 3493.300 1664.760 3493.580 1665.040 ;
        RECT 3490.260 1654.920 3490.540 1655.200 ;
        RECT 3490.880 1654.920 3491.160 1655.200 ;
        RECT 3491.500 1654.920 3491.780 1655.200 ;
        RECT 3492.120 1654.920 3492.400 1655.200 ;
        RECT 3492.740 1654.920 3493.020 1655.200 ;
        RECT 3493.360 1654.920 3493.640 1655.200 ;
        RECT 3493.980 1654.920 3494.260 1655.200 ;
        RECT 3490.260 1654.300 3490.540 1654.580 ;
        RECT 3490.880 1654.300 3491.160 1654.580 ;
        RECT 3491.500 1654.300 3491.780 1654.580 ;
        RECT 3492.120 1654.300 3492.400 1654.580 ;
        RECT 3492.740 1654.300 3493.020 1654.580 ;
        RECT 3493.360 1654.300 3493.640 1654.580 ;
        RECT 3493.980 1654.300 3494.260 1654.580 ;
        RECT 3490.260 1653.680 3490.540 1653.960 ;
        RECT 3490.880 1653.680 3491.160 1653.960 ;
        RECT 3491.500 1653.680 3491.780 1653.960 ;
        RECT 3492.120 1653.680 3492.400 1653.960 ;
        RECT 3492.740 1653.680 3493.020 1653.960 ;
        RECT 3493.360 1653.680 3493.640 1653.960 ;
        RECT 3493.980 1653.680 3494.260 1653.960 ;
        RECT 3490.260 1653.060 3490.540 1653.340 ;
        RECT 3490.880 1653.060 3491.160 1653.340 ;
        RECT 3491.500 1653.060 3491.780 1653.340 ;
        RECT 3492.120 1653.060 3492.400 1653.340 ;
        RECT 3492.740 1653.060 3493.020 1653.340 ;
        RECT 3493.360 1653.060 3493.640 1653.340 ;
        RECT 3493.980 1653.060 3494.260 1653.340 ;
        RECT 3490.260 1652.440 3490.540 1652.720 ;
        RECT 3490.880 1652.440 3491.160 1652.720 ;
        RECT 3491.500 1652.440 3491.780 1652.720 ;
        RECT 3492.120 1652.440 3492.400 1652.720 ;
        RECT 3492.740 1652.440 3493.020 1652.720 ;
        RECT 3493.360 1652.440 3493.640 1652.720 ;
        RECT 3493.980 1652.440 3494.260 1652.720 ;
        RECT 3490.260 1651.820 3490.540 1652.100 ;
        RECT 3490.880 1651.820 3491.160 1652.100 ;
        RECT 3491.500 1651.820 3491.780 1652.100 ;
        RECT 3492.120 1651.820 3492.400 1652.100 ;
        RECT 3492.740 1651.820 3493.020 1652.100 ;
        RECT 3493.360 1651.820 3493.640 1652.100 ;
        RECT 3493.980 1651.820 3494.260 1652.100 ;
        RECT 3490.260 1651.200 3490.540 1651.480 ;
        RECT 3490.880 1651.200 3491.160 1651.480 ;
        RECT 3491.500 1651.200 3491.780 1651.480 ;
        RECT 3492.120 1651.200 3492.400 1651.480 ;
        RECT 3492.740 1651.200 3493.020 1651.480 ;
        RECT 3493.360 1651.200 3493.640 1651.480 ;
        RECT 3493.980 1651.200 3494.260 1651.480 ;
        RECT 3321.035 1647.160 3321.315 1647.440 ;
        RECT 3322.035 1647.160 3322.315 1647.440 ;
        RECT 3321.035 1645.660 3321.315 1645.940 ;
        RECT 3322.035 1645.660 3322.315 1645.940 ;
        RECT 3321.035 1644.160 3321.315 1644.440 ;
        RECT 3322.035 1644.160 3322.315 1644.440 ;
        RECT 1912.010 1591.850 1912.290 1592.130 ;
        RECT 1913.510 1591.850 1913.790 1592.130 ;
        RECT 1912.010 1584.860 1912.290 1585.140 ;
        RECT 1913.510 1584.860 1913.790 1585.140 ;
        RECT 1912.010 1577.870 1912.290 1578.150 ;
        RECT 1913.510 1577.870 1913.790 1578.150 ;
        RECT 3490.220 1601.890 3490.500 1602.170 ;
        RECT 3491.720 1601.890 3492.000 1602.170 ;
        RECT 3493.220 1601.890 3493.500 1602.170 ;
        RECT 1912.010 1570.880 1912.290 1571.160 ;
        RECT 1913.510 1570.880 1913.790 1571.160 ;
        RECT 785.790 1528.350 786.070 1528.630 ;
        RECT 786.410 1528.350 786.690 1528.630 ;
        RECT 787.030 1528.350 787.310 1528.630 ;
        RECT 787.650 1528.350 787.930 1528.630 ;
        RECT 785.790 1527.730 786.070 1528.010 ;
        RECT 786.410 1527.730 786.690 1528.010 ;
        RECT 787.030 1527.730 787.310 1528.010 ;
        RECT 787.650 1527.730 787.930 1528.010 ;
        RECT 785.790 1527.110 786.070 1527.390 ;
        RECT 786.410 1527.110 786.690 1527.390 ;
        RECT 787.030 1527.110 787.310 1527.390 ;
        RECT 787.650 1527.110 787.930 1527.390 ;
        RECT 785.790 1526.490 786.070 1526.770 ;
        RECT 786.410 1526.490 786.690 1526.770 ;
        RECT 787.030 1526.490 787.310 1526.770 ;
        RECT 787.650 1526.490 787.930 1526.770 ;
        RECT 785.790 1525.870 786.070 1526.150 ;
        RECT 786.410 1525.870 786.690 1526.150 ;
        RECT 787.030 1525.870 787.310 1526.150 ;
        RECT 787.650 1525.870 787.930 1526.150 ;
        RECT 785.790 1525.250 786.070 1525.530 ;
        RECT 786.410 1525.250 786.690 1525.530 ;
        RECT 787.030 1525.250 787.310 1525.530 ;
        RECT 787.650 1525.250 787.930 1525.530 ;
        RECT 785.790 1524.630 786.070 1524.910 ;
        RECT 786.410 1524.630 786.690 1524.910 ;
        RECT 787.030 1524.630 787.310 1524.910 ;
        RECT 787.650 1524.630 787.930 1524.910 ;
        RECT 1911.650 1528.350 1911.930 1528.630 ;
        RECT 1912.270 1528.350 1912.550 1528.630 ;
        RECT 1912.890 1528.350 1913.170 1528.630 ;
        RECT 1913.510 1528.350 1913.790 1528.630 ;
        RECT 1911.650 1527.730 1911.930 1528.010 ;
        RECT 1912.270 1527.730 1912.550 1528.010 ;
        RECT 1912.890 1527.730 1913.170 1528.010 ;
        RECT 1913.510 1527.730 1913.790 1528.010 ;
        RECT 1911.650 1527.110 1911.930 1527.390 ;
        RECT 1912.270 1527.110 1912.550 1527.390 ;
        RECT 1912.890 1527.110 1913.170 1527.390 ;
        RECT 1913.510 1527.110 1913.790 1527.390 ;
        RECT 1911.650 1526.490 1911.930 1526.770 ;
        RECT 1912.270 1526.490 1912.550 1526.770 ;
        RECT 1912.890 1526.490 1913.170 1526.770 ;
        RECT 1913.510 1526.490 1913.790 1526.770 ;
        RECT 1911.650 1525.870 1911.930 1526.150 ;
        RECT 1912.270 1525.870 1912.550 1526.150 ;
        RECT 1912.890 1525.870 1913.170 1526.150 ;
        RECT 1913.510 1525.870 1913.790 1526.150 ;
        RECT 1911.650 1525.250 1911.930 1525.530 ;
        RECT 1912.270 1525.250 1912.550 1525.530 ;
        RECT 1912.890 1525.250 1913.170 1525.530 ;
        RECT 1913.510 1525.250 1913.790 1525.530 ;
        RECT 1911.650 1524.630 1911.930 1524.910 ;
        RECT 1912.270 1524.630 1912.550 1524.910 ;
        RECT 1912.890 1524.630 1913.170 1524.910 ;
        RECT 1913.510 1524.630 1913.790 1524.910 ;
        RECT 1951.100 1535.650 1951.380 1535.930 ;
        RECT 1951.720 1535.650 1952.000 1535.930 ;
        RECT 1951.100 1535.030 1951.380 1535.310 ;
        RECT 1951.720 1535.030 1952.000 1535.310 ;
        RECT 1951.100 1534.410 1951.380 1534.690 ;
        RECT 1951.720 1534.410 1952.000 1534.690 ;
        RECT 1951.100 1533.790 1951.380 1534.070 ;
        RECT 1951.720 1533.790 1952.000 1534.070 ;
        RECT 1951.100 1533.170 1951.380 1533.450 ;
        RECT 1951.720 1533.170 1952.000 1533.450 ;
        RECT 1951.100 1532.550 1951.380 1532.830 ;
        RECT 1951.720 1532.550 1952.000 1532.830 ;
        RECT 1951.100 1531.930 1951.380 1532.210 ;
        RECT 1951.720 1531.930 1952.000 1532.210 ;
        RECT 1943.125 1528.650 1943.405 1528.930 ;
        RECT 1943.745 1528.650 1944.025 1528.930 ;
        RECT 1943.125 1528.030 1943.405 1528.310 ;
        RECT 1943.745 1528.030 1944.025 1528.310 ;
        RECT 1943.125 1527.410 1943.405 1527.690 ;
        RECT 1943.745 1527.410 1944.025 1527.690 ;
        RECT 1943.125 1526.790 1943.405 1527.070 ;
        RECT 1943.745 1526.790 1944.025 1527.070 ;
        RECT 1943.125 1526.170 1943.405 1526.450 ;
        RECT 1943.745 1526.170 1944.025 1526.450 ;
        RECT 1943.125 1525.550 1943.405 1525.830 ;
        RECT 1943.745 1525.550 1944.025 1525.830 ;
        RECT 1943.125 1524.930 1943.405 1525.210 ;
        RECT 1943.745 1524.930 1944.025 1525.210 ;
        RECT 1967.050 1535.650 1967.330 1535.930 ;
        RECT 1967.670 1535.650 1967.950 1535.930 ;
        RECT 1967.050 1535.030 1967.330 1535.310 ;
        RECT 1967.670 1535.030 1967.950 1535.310 ;
        RECT 1967.050 1534.410 1967.330 1534.690 ;
        RECT 1967.670 1534.410 1967.950 1534.690 ;
        RECT 1967.050 1533.790 1967.330 1534.070 ;
        RECT 1967.670 1533.790 1967.950 1534.070 ;
        RECT 1967.050 1533.170 1967.330 1533.450 ;
        RECT 1967.670 1533.170 1967.950 1533.450 ;
        RECT 1967.050 1532.550 1967.330 1532.830 ;
        RECT 1967.670 1532.550 1967.950 1532.830 ;
        RECT 1967.050 1531.930 1967.330 1532.210 ;
        RECT 1967.670 1531.930 1967.950 1532.210 ;
        RECT 1959.075 1528.650 1959.355 1528.930 ;
        RECT 1959.695 1528.650 1959.975 1528.930 ;
        RECT 1959.075 1528.030 1959.355 1528.310 ;
        RECT 1959.695 1528.030 1959.975 1528.310 ;
        RECT 1959.075 1527.410 1959.355 1527.690 ;
        RECT 1959.695 1527.410 1959.975 1527.690 ;
        RECT 1959.075 1526.790 1959.355 1527.070 ;
        RECT 1959.695 1526.790 1959.975 1527.070 ;
        RECT 1959.075 1526.170 1959.355 1526.450 ;
        RECT 1959.695 1526.170 1959.975 1526.450 ;
        RECT 1959.075 1525.550 1959.355 1525.830 ;
        RECT 1959.695 1525.550 1959.975 1525.830 ;
        RECT 1959.075 1524.930 1959.355 1525.210 ;
        RECT 1959.695 1524.930 1959.975 1525.210 ;
        RECT 1983.000 1535.650 1983.280 1535.930 ;
        RECT 1983.620 1535.650 1983.900 1535.930 ;
        RECT 1983.000 1535.030 1983.280 1535.310 ;
        RECT 1983.620 1535.030 1983.900 1535.310 ;
        RECT 1983.000 1534.410 1983.280 1534.690 ;
        RECT 1983.620 1534.410 1983.900 1534.690 ;
        RECT 1983.000 1533.790 1983.280 1534.070 ;
        RECT 1983.620 1533.790 1983.900 1534.070 ;
        RECT 1983.000 1533.170 1983.280 1533.450 ;
        RECT 1983.620 1533.170 1983.900 1533.450 ;
        RECT 1983.000 1532.550 1983.280 1532.830 ;
        RECT 1983.620 1532.550 1983.900 1532.830 ;
        RECT 1983.000 1531.930 1983.280 1532.210 ;
        RECT 1983.620 1531.930 1983.900 1532.210 ;
        RECT 1975.025 1528.650 1975.305 1528.930 ;
        RECT 1975.645 1528.650 1975.925 1528.930 ;
        RECT 1975.025 1528.030 1975.305 1528.310 ;
        RECT 1975.645 1528.030 1975.925 1528.310 ;
        RECT 1975.025 1527.410 1975.305 1527.690 ;
        RECT 1975.645 1527.410 1975.925 1527.690 ;
        RECT 1975.025 1526.790 1975.305 1527.070 ;
        RECT 1975.645 1526.790 1975.925 1527.070 ;
        RECT 1975.025 1526.170 1975.305 1526.450 ;
        RECT 1975.645 1526.170 1975.925 1526.450 ;
        RECT 1975.025 1525.550 1975.305 1525.830 ;
        RECT 1975.645 1525.550 1975.925 1525.830 ;
        RECT 1975.025 1524.930 1975.305 1525.210 ;
        RECT 1975.645 1524.930 1975.925 1525.210 ;
        RECT 1990.975 1528.650 1991.255 1528.930 ;
        RECT 1991.595 1528.650 1991.875 1528.930 ;
        RECT 1990.975 1528.030 1991.255 1528.310 ;
        RECT 1991.595 1528.030 1991.875 1528.310 ;
        RECT 1990.975 1527.410 1991.255 1527.690 ;
        RECT 1991.595 1527.410 1991.875 1527.690 ;
        RECT 1990.975 1526.790 1991.255 1527.070 ;
        RECT 1991.595 1526.790 1991.875 1527.070 ;
        RECT 1990.975 1526.170 1991.255 1526.450 ;
        RECT 1991.595 1526.170 1991.875 1526.450 ;
        RECT 1990.975 1525.550 1991.255 1525.830 ;
        RECT 1991.595 1525.550 1991.875 1525.830 ;
        RECT 1990.975 1524.930 1991.255 1525.210 ;
        RECT 1991.595 1524.930 1991.875 1525.210 ;
        RECT 2451.100 1535.650 2451.380 1535.930 ;
        RECT 2451.720 1535.650 2452.000 1535.930 ;
        RECT 2451.100 1535.030 2451.380 1535.310 ;
        RECT 2451.720 1535.030 2452.000 1535.310 ;
        RECT 2451.100 1534.410 2451.380 1534.690 ;
        RECT 2451.720 1534.410 2452.000 1534.690 ;
        RECT 2451.100 1533.790 2451.380 1534.070 ;
        RECT 2451.720 1533.790 2452.000 1534.070 ;
        RECT 2451.100 1533.170 2451.380 1533.450 ;
        RECT 2451.720 1533.170 2452.000 1533.450 ;
        RECT 2451.100 1532.550 2451.380 1532.830 ;
        RECT 2451.720 1532.550 2452.000 1532.830 ;
        RECT 2451.100 1531.930 2451.380 1532.210 ;
        RECT 2451.720 1531.930 2452.000 1532.210 ;
        RECT 2443.125 1528.650 2443.405 1528.930 ;
        RECT 2443.745 1528.650 2444.025 1528.930 ;
        RECT 2443.125 1528.030 2443.405 1528.310 ;
        RECT 2443.745 1528.030 2444.025 1528.310 ;
        RECT 2443.125 1527.410 2443.405 1527.690 ;
        RECT 2443.745 1527.410 2444.025 1527.690 ;
        RECT 2443.125 1526.790 2443.405 1527.070 ;
        RECT 2443.745 1526.790 2444.025 1527.070 ;
        RECT 2443.125 1526.170 2443.405 1526.450 ;
        RECT 2443.745 1526.170 2444.025 1526.450 ;
        RECT 2443.125 1525.550 2443.405 1525.830 ;
        RECT 2443.745 1525.550 2444.025 1525.830 ;
        RECT 2443.125 1524.930 2443.405 1525.210 ;
        RECT 2443.745 1524.930 2444.025 1525.210 ;
        RECT 2467.050 1535.650 2467.330 1535.930 ;
        RECT 2467.670 1535.650 2467.950 1535.930 ;
        RECT 2467.050 1535.030 2467.330 1535.310 ;
        RECT 2467.670 1535.030 2467.950 1535.310 ;
        RECT 2467.050 1534.410 2467.330 1534.690 ;
        RECT 2467.670 1534.410 2467.950 1534.690 ;
        RECT 2467.050 1533.790 2467.330 1534.070 ;
        RECT 2467.670 1533.790 2467.950 1534.070 ;
        RECT 2467.050 1533.170 2467.330 1533.450 ;
        RECT 2467.670 1533.170 2467.950 1533.450 ;
        RECT 2467.050 1532.550 2467.330 1532.830 ;
        RECT 2467.670 1532.550 2467.950 1532.830 ;
        RECT 2467.050 1531.930 2467.330 1532.210 ;
        RECT 2467.670 1531.930 2467.950 1532.210 ;
        RECT 2459.075 1528.650 2459.355 1528.930 ;
        RECT 2459.695 1528.650 2459.975 1528.930 ;
        RECT 2459.075 1528.030 2459.355 1528.310 ;
        RECT 2459.695 1528.030 2459.975 1528.310 ;
        RECT 2459.075 1527.410 2459.355 1527.690 ;
        RECT 2459.695 1527.410 2459.975 1527.690 ;
        RECT 2459.075 1526.790 2459.355 1527.070 ;
        RECT 2459.695 1526.790 2459.975 1527.070 ;
        RECT 2459.075 1526.170 2459.355 1526.450 ;
        RECT 2459.695 1526.170 2459.975 1526.450 ;
        RECT 2459.075 1525.550 2459.355 1525.830 ;
        RECT 2459.695 1525.550 2459.975 1525.830 ;
        RECT 2459.075 1524.930 2459.355 1525.210 ;
        RECT 2459.695 1524.930 2459.975 1525.210 ;
        RECT 2483.000 1535.650 2483.280 1535.930 ;
        RECT 2483.620 1535.650 2483.900 1535.930 ;
        RECT 2483.000 1535.030 2483.280 1535.310 ;
        RECT 2483.620 1535.030 2483.900 1535.310 ;
        RECT 2483.000 1534.410 2483.280 1534.690 ;
        RECT 2483.620 1534.410 2483.900 1534.690 ;
        RECT 2483.000 1533.790 2483.280 1534.070 ;
        RECT 2483.620 1533.790 2483.900 1534.070 ;
        RECT 2483.000 1533.170 2483.280 1533.450 ;
        RECT 2483.620 1533.170 2483.900 1533.450 ;
        RECT 2483.000 1532.550 2483.280 1532.830 ;
        RECT 2483.620 1532.550 2483.900 1532.830 ;
        RECT 2483.000 1531.930 2483.280 1532.210 ;
        RECT 2483.620 1531.930 2483.900 1532.210 ;
        RECT 2475.025 1528.650 2475.305 1528.930 ;
        RECT 2475.645 1528.650 2475.925 1528.930 ;
        RECT 2475.025 1528.030 2475.305 1528.310 ;
        RECT 2475.645 1528.030 2475.925 1528.310 ;
        RECT 2475.025 1527.410 2475.305 1527.690 ;
        RECT 2475.645 1527.410 2475.925 1527.690 ;
        RECT 2475.025 1526.790 2475.305 1527.070 ;
        RECT 2475.645 1526.790 2475.925 1527.070 ;
        RECT 2475.025 1526.170 2475.305 1526.450 ;
        RECT 2475.645 1526.170 2475.925 1526.450 ;
        RECT 2475.025 1525.550 2475.305 1525.830 ;
        RECT 2475.645 1525.550 2475.925 1525.830 ;
        RECT 2475.025 1524.930 2475.305 1525.210 ;
        RECT 2475.645 1524.930 2475.925 1525.210 ;
        RECT 2490.975 1528.650 2491.255 1528.930 ;
        RECT 2491.595 1528.650 2491.875 1528.930 ;
        RECT 2490.975 1528.030 2491.255 1528.310 ;
        RECT 2491.595 1528.030 2491.875 1528.310 ;
        RECT 2490.975 1527.410 2491.255 1527.690 ;
        RECT 2491.595 1527.410 2491.875 1527.690 ;
        RECT 2490.975 1526.790 2491.255 1527.070 ;
        RECT 2491.595 1526.790 2491.875 1527.070 ;
        RECT 2490.975 1526.170 2491.255 1526.450 ;
        RECT 2491.595 1526.170 2491.875 1526.450 ;
        RECT 2490.975 1525.550 2491.255 1525.830 ;
        RECT 2491.595 1525.550 2491.875 1525.830 ;
        RECT 2490.975 1524.930 2491.255 1525.210 ;
        RECT 2491.595 1524.930 2491.875 1525.210 ;
        RECT 2954.550 1535.350 2954.830 1535.630 ;
        RECT 2955.170 1535.350 2955.450 1535.630 ;
        RECT 2955.790 1535.350 2956.070 1535.630 ;
        RECT 2956.410 1535.350 2956.690 1535.630 ;
        RECT 2957.030 1535.350 2957.310 1535.630 ;
        RECT 2957.650 1535.350 2957.930 1535.630 ;
        RECT 2958.270 1535.350 2958.550 1535.630 ;
        RECT 2954.550 1534.730 2954.830 1535.010 ;
        RECT 2955.170 1534.730 2955.450 1535.010 ;
        RECT 2955.790 1534.730 2956.070 1535.010 ;
        RECT 2956.410 1534.730 2956.690 1535.010 ;
        RECT 2957.030 1534.730 2957.310 1535.010 ;
        RECT 2957.650 1534.730 2957.930 1535.010 ;
        RECT 2958.270 1534.730 2958.550 1535.010 ;
        RECT 2954.550 1534.110 2954.830 1534.390 ;
        RECT 2955.170 1534.110 2955.450 1534.390 ;
        RECT 2955.790 1534.110 2956.070 1534.390 ;
        RECT 2956.410 1534.110 2956.690 1534.390 ;
        RECT 2957.030 1534.110 2957.310 1534.390 ;
        RECT 2957.650 1534.110 2957.930 1534.390 ;
        RECT 2958.270 1534.110 2958.550 1534.390 ;
        RECT 2954.550 1533.490 2954.830 1533.770 ;
        RECT 2955.170 1533.490 2955.450 1533.770 ;
        RECT 2955.790 1533.490 2956.070 1533.770 ;
        RECT 2956.410 1533.490 2956.690 1533.770 ;
        RECT 2957.030 1533.490 2957.310 1533.770 ;
        RECT 2957.650 1533.490 2957.930 1533.770 ;
        RECT 2958.270 1533.490 2958.550 1533.770 ;
        RECT 2954.550 1532.870 2954.830 1533.150 ;
        RECT 2955.170 1532.870 2955.450 1533.150 ;
        RECT 2955.790 1532.870 2956.070 1533.150 ;
        RECT 2956.410 1532.870 2956.690 1533.150 ;
        RECT 2957.030 1532.870 2957.310 1533.150 ;
        RECT 2957.650 1532.870 2957.930 1533.150 ;
        RECT 2958.270 1532.870 2958.550 1533.150 ;
        RECT 2954.550 1532.250 2954.830 1532.530 ;
        RECT 2955.170 1532.250 2955.450 1532.530 ;
        RECT 2955.790 1532.250 2956.070 1532.530 ;
        RECT 2956.410 1532.250 2956.690 1532.530 ;
        RECT 2957.030 1532.250 2957.310 1532.530 ;
        RECT 2957.650 1532.250 2957.930 1532.530 ;
        RECT 2958.270 1532.250 2958.550 1532.530 ;
        RECT 2954.550 1531.630 2954.830 1531.910 ;
        RECT 2955.170 1531.630 2955.450 1531.910 ;
        RECT 2955.790 1531.630 2956.070 1531.910 ;
        RECT 2956.410 1531.630 2956.690 1531.910 ;
        RECT 2957.030 1531.630 2957.310 1531.910 ;
        RECT 2957.650 1531.630 2957.930 1531.910 ;
        RECT 2958.270 1531.630 2958.550 1531.910 ;
        RECT 396.500 1502.830 396.780 1503.110 ;
        RECT 398.000 1502.830 398.280 1503.110 ;
        RECT 399.500 1502.830 399.780 1503.110 ;
        RECT 396.420 1449.960 396.700 1450.240 ;
        RECT 397.920 1449.960 398.200 1450.240 ;
        RECT 399.420 1449.960 399.700 1450.240 ;
        RECT 396.040 1416.580 396.320 1416.860 ;
        RECT 396.660 1416.580 396.940 1416.860 ;
        RECT 397.280 1416.580 397.560 1416.860 ;
        RECT 397.900 1416.580 398.180 1416.860 ;
        RECT 398.520 1416.580 398.800 1416.860 ;
        RECT 399.140 1416.580 399.420 1416.860 ;
        RECT 399.760 1416.580 400.040 1416.860 ;
        RECT 396.040 1415.960 396.320 1416.240 ;
        RECT 396.660 1415.960 396.940 1416.240 ;
        RECT 397.280 1415.960 397.560 1416.240 ;
        RECT 397.900 1415.960 398.180 1416.240 ;
        RECT 398.520 1415.960 398.800 1416.240 ;
        RECT 399.140 1415.960 399.420 1416.240 ;
        RECT 399.760 1415.960 400.040 1416.240 ;
        RECT 396.040 1415.340 396.320 1415.620 ;
        RECT 396.660 1415.340 396.940 1415.620 ;
        RECT 397.280 1415.340 397.560 1415.620 ;
        RECT 397.900 1415.340 398.180 1415.620 ;
        RECT 398.520 1415.340 398.800 1415.620 ;
        RECT 399.140 1415.340 399.420 1415.620 ;
        RECT 399.760 1415.340 400.040 1415.620 ;
        RECT 396.040 1414.720 396.320 1415.000 ;
        RECT 396.660 1414.720 396.940 1415.000 ;
        RECT 397.280 1414.720 397.560 1415.000 ;
        RECT 397.900 1414.720 398.180 1415.000 ;
        RECT 398.520 1414.720 398.800 1415.000 ;
        RECT 399.140 1414.720 399.420 1415.000 ;
        RECT 399.760 1414.720 400.040 1415.000 ;
        RECT 396.040 1414.100 396.320 1414.380 ;
        RECT 396.660 1414.100 396.940 1414.380 ;
        RECT 397.280 1414.100 397.560 1414.380 ;
        RECT 397.900 1414.100 398.180 1414.380 ;
        RECT 398.520 1414.100 398.800 1414.380 ;
        RECT 399.140 1414.100 399.420 1414.380 ;
        RECT 399.760 1414.100 400.040 1414.380 ;
        RECT 396.040 1413.480 396.320 1413.760 ;
        RECT 396.660 1413.480 396.940 1413.760 ;
        RECT 397.280 1413.480 397.560 1413.760 ;
        RECT 397.900 1413.480 398.180 1413.760 ;
        RECT 398.520 1413.480 398.800 1413.760 ;
        RECT 399.140 1413.480 399.420 1413.760 ;
        RECT 399.760 1413.480 400.040 1413.760 ;
        RECT 396.040 1412.860 396.320 1413.140 ;
        RECT 396.660 1412.860 396.940 1413.140 ;
        RECT 397.280 1412.860 397.560 1413.140 ;
        RECT 397.900 1412.860 398.180 1413.140 ;
        RECT 398.520 1412.860 398.800 1413.140 ;
        RECT 399.140 1412.860 399.420 1413.140 ;
        RECT 399.760 1412.860 400.040 1413.140 ;
        RECT 496.470 1416.280 496.750 1416.560 ;
        RECT 497.090 1416.280 497.370 1416.560 ;
        RECT 496.470 1415.660 496.750 1415.940 ;
        RECT 497.090 1415.660 497.370 1415.940 ;
        RECT 496.470 1415.040 496.750 1415.320 ;
        RECT 497.090 1415.040 497.370 1415.320 ;
        RECT 496.470 1414.420 496.750 1414.700 ;
        RECT 497.090 1414.420 497.370 1414.700 ;
        RECT 496.470 1413.800 496.750 1414.080 ;
        RECT 497.090 1413.800 497.370 1414.080 ;
        RECT 496.470 1413.180 496.750 1413.460 ;
        RECT 497.090 1413.180 497.370 1413.460 ;
        RECT 496.470 1412.560 496.750 1412.840 ;
        RECT 497.090 1412.560 497.370 1412.840 ;
        RECT 471.470 1409.280 471.750 1409.560 ;
        RECT 472.090 1409.280 472.370 1409.560 ;
        RECT 471.470 1408.660 471.750 1408.940 ;
        RECT 472.090 1408.660 472.370 1408.940 ;
        RECT 471.470 1408.040 471.750 1408.320 ;
        RECT 472.090 1408.040 472.370 1408.320 ;
        RECT 471.470 1407.420 471.750 1407.700 ;
        RECT 472.090 1407.420 472.370 1407.700 ;
        RECT 471.470 1406.800 471.750 1407.080 ;
        RECT 472.090 1406.800 472.370 1407.080 ;
        RECT 471.470 1406.180 471.750 1406.460 ;
        RECT 472.090 1406.180 472.370 1406.460 ;
        RECT 471.470 1405.560 471.750 1405.840 ;
        RECT 472.090 1405.560 472.370 1405.840 ;
        RECT 546.470 1416.280 546.750 1416.560 ;
        RECT 547.090 1416.280 547.370 1416.560 ;
        RECT 546.470 1415.660 546.750 1415.940 ;
        RECT 547.090 1415.660 547.370 1415.940 ;
        RECT 546.470 1415.040 546.750 1415.320 ;
        RECT 547.090 1415.040 547.370 1415.320 ;
        RECT 546.470 1414.420 546.750 1414.700 ;
        RECT 547.090 1414.420 547.370 1414.700 ;
        RECT 546.470 1413.800 546.750 1414.080 ;
        RECT 547.090 1413.800 547.370 1414.080 ;
        RECT 546.470 1413.180 546.750 1413.460 ;
        RECT 547.090 1413.180 547.370 1413.460 ;
        RECT 546.470 1412.560 546.750 1412.840 ;
        RECT 547.090 1412.560 547.370 1412.840 ;
        RECT 521.470 1409.280 521.750 1409.560 ;
        RECT 522.090 1409.280 522.370 1409.560 ;
        RECT 521.470 1408.660 521.750 1408.940 ;
        RECT 522.090 1408.660 522.370 1408.940 ;
        RECT 521.470 1408.040 521.750 1408.320 ;
        RECT 522.090 1408.040 522.370 1408.320 ;
        RECT 521.470 1407.420 521.750 1407.700 ;
        RECT 522.090 1407.420 522.370 1407.700 ;
        RECT 521.470 1406.800 521.750 1407.080 ;
        RECT 522.090 1406.800 522.370 1407.080 ;
        RECT 521.470 1406.180 521.750 1406.460 ;
        RECT 522.090 1406.180 522.370 1406.460 ;
        RECT 521.470 1405.560 521.750 1405.840 ;
        RECT 522.090 1405.560 522.370 1405.840 ;
        RECT 596.470 1416.280 596.750 1416.560 ;
        RECT 597.090 1416.280 597.370 1416.560 ;
        RECT 596.470 1415.660 596.750 1415.940 ;
        RECT 597.090 1415.660 597.370 1415.940 ;
        RECT 596.470 1415.040 596.750 1415.320 ;
        RECT 597.090 1415.040 597.370 1415.320 ;
        RECT 596.470 1414.420 596.750 1414.700 ;
        RECT 597.090 1414.420 597.370 1414.700 ;
        RECT 596.470 1413.800 596.750 1414.080 ;
        RECT 597.090 1413.800 597.370 1414.080 ;
        RECT 596.470 1413.180 596.750 1413.460 ;
        RECT 597.090 1413.180 597.370 1413.460 ;
        RECT 596.470 1412.560 596.750 1412.840 ;
        RECT 597.090 1412.560 597.370 1412.840 ;
        RECT 571.470 1409.280 571.750 1409.560 ;
        RECT 572.090 1409.280 572.370 1409.560 ;
        RECT 571.470 1408.660 571.750 1408.940 ;
        RECT 572.090 1408.660 572.370 1408.940 ;
        RECT 571.470 1408.040 571.750 1408.320 ;
        RECT 572.090 1408.040 572.370 1408.320 ;
        RECT 571.470 1407.420 571.750 1407.700 ;
        RECT 572.090 1407.420 572.370 1407.700 ;
        RECT 571.470 1406.800 571.750 1407.080 ;
        RECT 572.090 1406.800 572.370 1407.080 ;
        RECT 571.470 1406.180 571.750 1406.460 ;
        RECT 572.090 1406.180 572.370 1406.460 ;
        RECT 571.470 1405.560 571.750 1405.840 ;
        RECT 572.090 1405.560 572.370 1405.840 ;
        RECT 646.470 1416.280 646.750 1416.560 ;
        RECT 647.090 1416.280 647.370 1416.560 ;
        RECT 646.470 1415.660 646.750 1415.940 ;
        RECT 647.090 1415.660 647.370 1415.940 ;
        RECT 646.470 1415.040 646.750 1415.320 ;
        RECT 647.090 1415.040 647.370 1415.320 ;
        RECT 646.470 1414.420 646.750 1414.700 ;
        RECT 647.090 1414.420 647.370 1414.700 ;
        RECT 646.470 1413.800 646.750 1414.080 ;
        RECT 647.090 1413.800 647.370 1414.080 ;
        RECT 646.470 1413.180 646.750 1413.460 ;
        RECT 647.090 1413.180 647.370 1413.460 ;
        RECT 646.470 1412.560 646.750 1412.840 ;
        RECT 647.090 1412.560 647.370 1412.840 ;
        RECT 621.470 1409.280 621.750 1409.560 ;
        RECT 622.090 1409.280 622.370 1409.560 ;
        RECT 621.470 1408.660 621.750 1408.940 ;
        RECT 622.090 1408.660 622.370 1408.940 ;
        RECT 621.470 1408.040 621.750 1408.320 ;
        RECT 622.090 1408.040 622.370 1408.320 ;
        RECT 621.470 1407.420 621.750 1407.700 ;
        RECT 622.090 1407.420 622.370 1407.700 ;
        RECT 621.470 1406.800 621.750 1407.080 ;
        RECT 622.090 1406.800 622.370 1407.080 ;
        RECT 621.470 1406.180 621.750 1406.460 ;
        RECT 622.090 1406.180 622.370 1406.460 ;
        RECT 621.470 1405.560 621.750 1405.840 ;
        RECT 622.090 1405.560 622.370 1405.840 ;
        RECT 696.470 1416.280 696.750 1416.560 ;
        RECT 697.090 1416.280 697.370 1416.560 ;
        RECT 696.470 1415.660 696.750 1415.940 ;
        RECT 697.090 1415.660 697.370 1415.940 ;
        RECT 696.470 1415.040 696.750 1415.320 ;
        RECT 697.090 1415.040 697.370 1415.320 ;
        RECT 696.470 1414.420 696.750 1414.700 ;
        RECT 697.090 1414.420 697.370 1414.700 ;
        RECT 696.470 1413.800 696.750 1414.080 ;
        RECT 697.090 1413.800 697.370 1414.080 ;
        RECT 696.470 1413.180 696.750 1413.460 ;
        RECT 697.090 1413.180 697.370 1413.460 ;
        RECT 696.470 1412.560 696.750 1412.840 ;
        RECT 697.090 1412.560 697.370 1412.840 ;
        RECT 671.470 1409.280 671.750 1409.560 ;
        RECT 672.090 1409.280 672.370 1409.560 ;
        RECT 671.470 1408.660 671.750 1408.940 ;
        RECT 672.090 1408.660 672.370 1408.940 ;
        RECT 671.470 1408.040 671.750 1408.320 ;
        RECT 672.090 1408.040 672.370 1408.320 ;
        RECT 671.470 1407.420 671.750 1407.700 ;
        RECT 672.090 1407.420 672.370 1407.700 ;
        RECT 671.470 1406.800 671.750 1407.080 ;
        RECT 672.090 1406.800 672.370 1407.080 ;
        RECT 671.470 1406.180 671.750 1406.460 ;
        RECT 672.090 1406.180 672.370 1406.460 ;
        RECT 671.470 1405.560 671.750 1405.840 ;
        RECT 672.090 1405.560 672.370 1405.840 ;
        RECT 746.470 1416.280 746.750 1416.560 ;
        RECT 747.090 1416.280 747.370 1416.560 ;
        RECT 746.470 1415.660 746.750 1415.940 ;
        RECT 747.090 1415.660 747.370 1415.940 ;
        RECT 746.470 1415.040 746.750 1415.320 ;
        RECT 747.090 1415.040 747.370 1415.320 ;
        RECT 746.470 1414.420 746.750 1414.700 ;
        RECT 747.090 1414.420 747.370 1414.700 ;
        RECT 746.470 1413.800 746.750 1414.080 ;
        RECT 747.090 1413.800 747.370 1414.080 ;
        RECT 746.470 1413.180 746.750 1413.460 ;
        RECT 747.090 1413.180 747.370 1413.460 ;
        RECT 746.470 1412.560 746.750 1412.840 ;
        RECT 747.090 1412.560 747.370 1412.840 ;
        RECT 721.470 1409.280 721.750 1409.560 ;
        RECT 722.090 1409.280 722.370 1409.560 ;
        RECT 721.470 1408.660 721.750 1408.940 ;
        RECT 722.090 1408.660 722.370 1408.940 ;
        RECT 721.470 1408.040 721.750 1408.320 ;
        RECT 722.090 1408.040 722.370 1408.320 ;
        RECT 721.470 1407.420 721.750 1407.700 ;
        RECT 722.090 1407.420 722.370 1407.700 ;
        RECT 721.470 1406.800 721.750 1407.080 ;
        RECT 722.090 1406.800 722.370 1407.080 ;
        RECT 721.470 1406.180 721.750 1406.460 ;
        RECT 722.090 1406.180 722.370 1406.460 ;
        RECT 721.470 1405.560 721.750 1405.840 ;
        RECT 722.090 1405.560 722.370 1405.840 ;
        RECT 796.470 1416.280 796.750 1416.560 ;
        RECT 797.090 1416.280 797.370 1416.560 ;
        RECT 796.470 1415.660 796.750 1415.940 ;
        RECT 797.090 1415.660 797.370 1415.940 ;
        RECT 796.470 1415.040 796.750 1415.320 ;
        RECT 797.090 1415.040 797.370 1415.320 ;
        RECT 796.470 1414.420 796.750 1414.700 ;
        RECT 797.090 1414.420 797.370 1414.700 ;
        RECT 796.470 1413.800 796.750 1414.080 ;
        RECT 797.090 1413.800 797.370 1414.080 ;
        RECT 796.470 1413.180 796.750 1413.460 ;
        RECT 797.090 1413.180 797.370 1413.460 ;
        RECT 796.470 1412.560 796.750 1412.840 ;
        RECT 797.090 1412.560 797.370 1412.840 ;
        RECT 771.470 1409.280 771.750 1409.560 ;
        RECT 772.090 1409.280 772.370 1409.560 ;
        RECT 771.470 1408.660 771.750 1408.940 ;
        RECT 772.090 1408.660 772.370 1408.940 ;
        RECT 771.470 1408.040 771.750 1408.320 ;
        RECT 772.090 1408.040 772.370 1408.320 ;
        RECT 771.470 1407.420 771.750 1407.700 ;
        RECT 772.090 1407.420 772.370 1407.700 ;
        RECT 771.470 1406.800 771.750 1407.080 ;
        RECT 772.090 1406.800 772.370 1407.080 ;
        RECT 771.470 1406.180 771.750 1406.460 ;
        RECT 772.090 1406.180 772.370 1406.460 ;
        RECT 771.470 1405.560 771.750 1405.840 ;
        RECT 772.090 1405.560 772.370 1405.840 ;
        RECT 846.470 1416.280 846.750 1416.560 ;
        RECT 847.090 1416.280 847.370 1416.560 ;
        RECT 846.470 1415.660 846.750 1415.940 ;
        RECT 847.090 1415.660 847.370 1415.940 ;
        RECT 846.470 1415.040 846.750 1415.320 ;
        RECT 847.090 1415.040 847.370 1415.320 ;
        RECT 846.470 1414.420 846.750 1414.700 ;
        RECT 847.090 1414.420 847.370 1414.700 ;
        RECT 846.470 1413.800 846.750 1414.080 ;
        RECT 847.090 1413.800 847.370 1414.080 ;
        RECT 846.470 1413.180 846.750 1413.460 ;
        RECT 847.090 1413.180 847.370 1413.460 ;
        RECT 846.470 1412.560 846.750 1412.840 ;
        RECT 847.090 1412.560 847.370 1412.840 ;
        RECT 821.470 1409.280 821.750 1409.560 ;
        RECT 822.090 1409.280 822.370 1409.560 ;
        RECT 821.470 1408.660 821.750 1408.940 ;
        RECT 822.090 1408.660 822.370 1408.940 ;
        RECT 821.470 1408.040 821.750 1408.320 ;
        RECT 822.090 1408.040 822.370 1408.320 ;
        RECT 821.470 1407.420 821.750 1407.700 ;
        RECT 822.090 1407.420 822.370 1407.700 ;
        RECT 821.470 1406.800 821.750 1407.080 ;
        RECT 822.090 1406.800 822.370 1407.080 ;
        RECT 821.470 1406.180 821.750 1406.460 ;
        RECT 822.090 1406.180 822.370 1406.460 ;
        RECT 821.470 1405.560 821.750 1405.840 ;
        RECT 822.090 1405.560 822.370 1405.840 ;
        RECT 896.470 1416.280 896.750 1416.560 ;
        RECT 897.090 1416.280 897.370 1416.560 ;
        RECT 896.470 1415.660 896.750 1415.940 ;
        RECT 897.090 1415.660 897.370 1415.940 ;
        RECT 896.470 1415.040 896.750 1415.320 ;
        RECT 897.090 1415.040 897.370 1415.320 ;
        RECT 896.470 1414.420 896.750 1414.700 ;
        RECT 897.090 1414.420 897.370 1414.700 ;
        RECT 896.470 1413.800 896.750 1414.080 ;
        RECT 897.090 1413.800 897.370 1414.080 ;
        RECT 896.470 1413.180 896.750 1413.460 ;
        RECT 897.090 1413.180 897.370 1413.460 ;
        RECT 896.470 1412.560 896.750 1412.840 ;
        RECT 897.090 1412.560 897.370 1412.840 ;
        RECT 871.470 1409.280 871.750 1409.560 ;
        RECT 872.090 1409.280 872.370 1409.560 ;
        RECT 871.470 1408.660 871.750 1408.940 ;
        RECT 872.090 1408.660 872.370 1408.940 ;
        RECT 871.470 1408.040 871.750 1408.320 ;
        RECT 872.090 1408.040 872.370 1408.320 ;
        RECT 871.470 1407.420 871.750 1407.700 ;
        RECT 872.090 1407.420 872.370 1407.700 ;
        RECT 871.470 1406.800 871.750 1407.080 ;
        RECT 872.090 1406.800 872.370 1407.080 ;
        RECT 871.470 1406.180 871.750 1406.460 ;
        RECT 872.090 1406.180 872.370 1406.460 ;
        RECT 871.470 1405.560 871.750 1405.840 ;
        RECT 872.090 1405.560 872.370 1405.840 ;
        RECT 946.470 1416.280 946.750 1416.560 ;
        RECT 947.090 1416.280 947.370 1416.560 ;
        RECT 946.470 1415.660 946.750 1415.940 ;
        RECT 947.090 1415.660 947.370 1415.940 ;
        RECT 946.470 1415.040 946.750 1415.320 ;
        RECT 947.090 1415.040 947.370 1415.320 ;
        RECT 946.470 1414.420 946.750 1414.700 ;
        RECT 947.090 1414.420 947.370 1414.700 ;
        RECT 946.470 1413.800 946.750 1414.080 ;
        RECT 947.090 1413.800 947.370 1414.080 ;
        RECT 946.470 1413.180 946.750 1413.460 ;
        RECT 947.090 1413.180 947.370 1413.460 ;
        RECT 946.470 1412.560 946.750 1412.840 ;
        RECT 947.090 1412.560 947.370 1412.840 ;
        RECT 921.470 1409.280 921.750 1409.560 ;
        RECT 922.090 1409.280 922.370 1409.560 ;
        RECT 921.470 1408.660 921.750 1408.940 ;
        RECT 922.090 1408.660 922.370 1408.940 ;
        RECT 921.470 1408.040 921.750 1408.320 ;
        RECT 922.090 1408.040 922.370 1408.320 ;
        RECT 921.470 1407.420 921.750 1407.700 ;
        RECT 922.090 1407.420 922.370 1407.700 ;
        RECT 921.470 1406.800 921.750 1407.080 ;
        RECT 922.090 1406.800 922.370 1407.080 ;
        RECT 921.470 1406.180 921.750 1406.460 ;
        RECT 922.090 1406.180 922.370 1406.460 ;
        RECT 921.470 1405.560 921.750 1405.840 ;
        RECT 922.090 1405.560 922.370 1405.840 ;
        RECT 996.470 1416.280 996.750 1416.560 ;
        RECT 997.090 1416.280 997.370 1416.560 ;
        RECT 996.470 1415.660 996.750 1415.940 ;
        RECT 997.090 1415.660 997.370 1415.940 ;
        RECT 996.470 1415.040 996.750 1415.320 ;
        RECT 997.090 1415.040 997.370 1415.320 ;
        RECT 996.470 1414.420 996.750 1414.700 ;
        RECT 997.090 1414.420 997.370 1414.700 ;
        RECT 996.470 1413.800 996.750 1414.080 ;
        RECT 997.090 1413.800 997.370 1414.080 ;
        RECT 996.470 1413.180 996.750 1413.460 ;
        RECT 997.090 1413.180 997.370 1413.460 ;
        RECT 996.470 1412.560 996.750 1412.840 ;
        RECT 997.090 1412.560 997.370 1412.840 ;
        RECT 971.470 1409.280 971.750 1409.560 ;
        RECT 972.090 1409.280 972.370 1409.560 ;
        RECT 971.470 1408.660 971.750 1408.940 ;
        RECT 972.090 1408.660 972.370 1408.940 ;
        RECT 971.470 1408.040 971.750 1408.320 ;
        RECT 972.090 1408.040 972.370 1408.320 ;
        RECT 971.470 1407.420 971.750 1407.700 ;
        RECT 972.090 1407.420 972.370 1407.700 ;
        RECT 971.470 1406.800 971.750 1407.080 ;
        RECT 972.090 1406.800 972.370 1407.080 ;
        RECT 971.470 1406.180 971.750 1406.460 ;
        RECT 972.090 1406.180 972.370 1406.460 ;
        RECT 971.470 1405.560 971.750 1405.840 ;
        RECT 972.090 1405.560 972.370 1405.840 ;
        RECT 1046.470 1416.280 1046.750 1416.560 ;
        RECT 1047.090 1416.280 1047.370 1416.560 ;
        RECT 1046.470 1415.660 1046.750 1415.940 ;
        RECT 1047.090 1415.660 1047.370 1415.940 ;
        RECT 1046.470 1415.040 1046.750 1415.320 ;
        RECT 1047.090 1415.040 1047.370 1415.320 ;
        RECT 1046.470 1414.420 1046.750 1414.700 ;
        RECT 1047.090 1414.420 1047.370 1414.700 ;
        RECT 1046.470 1413.800 1046.750 1414.080 ;
        RECT 1047.090 1413.800 1047.370 1414.080 ;
        RECT 1046.470 1413.180 1046.750 1413.460 ;
        RECT 1047.090 1413.180 1047.370 1413.460 ;
        RECT 1046.470 1412.560 1046.750 1412.840 ;
        RECT 1047.090 1412.560 1047.370 1412.840 ;
        RECT 1021.470 1409.280 1021.750 1409.560 ;
        RECT 1022.090 1409.280 1022.370 1409.560 ;
        RECT 1021.470 1408.660 1021.750 1408.940 ;
        RECT 1022.090 1408.660 1022.370 1408.940 ;
        RECT 1021.470 1408.040 1021.750 1408.320 ;
        RECT 1022.090 1408.040 1022.370 1408.320 ;
        RECT 1021.470 1407.420 1021.750 1407.700 ;
        RECT 1022.090 1407.420 1022.370 1407.700 ;
        RECT 1021.470 1406.800 1021.750 1407.080 ;
        RECT 1022.090 1406.800 1022.370 1407.080 ;
        RECT 1021.470 1406.180 1021.750 1406.460 ;
        RECT 1022.090 1406.180 1022.370 1406.460 ;
        RECT 1021.470 1405.560 1021.750 1405.840 ;
        RECT 1022.090 1405.560 1022.370 1405.840 ;
        RECT 1096.470 1416.280 1096.750 1416.560 ;
        RECT 1097.090 1416.280 1097.370 1416.560 ;
        RECT 1096.470 1415.660 1096.750 1415.940 ;
        RECT 1097.090 1415.660 1097.370 1415.940 ;
        RECT 1096.470 1415.040 1096.750 1415.320 ;
        RECT 1097.090 1415.040 1097.370 1415.320 ;
        RECT 1096.470 1414.420 1096.750 1414.700 ;
        RECT 1097.090 1414.420 1097.370 1414.700 ;
        RECT 1096.470 1413.800 1096.750 1414.080 ;
        RECT 1097.090 1413.800 1097.370 1414.080 ;
        RECT 1096.470 1413.180 1096.750 1413.460 ;
        RECT 1097.090 1413.180 1097.370 1413.460 ;
        RECT 1096.470 1412.560 1096.750 1412.840 ;
        RECT 1097.090 1412.560 1097.370 1412.840 ;
        RECT 1071.470 1409.280 1071.750 1409.560 ;
        RECT 1072.090 1409.280 1072.370 1409.560 ;
        RECT 1071.470 1408.660 1071.750 1408.940 ;
        RECT 1072.090 1408.660 1072.370 1408.940 ;
        RECT 1071.470 1408.040 1071.750 1408.320 ;
        RECT 1072.090 1408.040 1072.370 1408.320 ;
        RECT 1071.470 1407.420 1071.750 1407.700 ;
        RECT 1072.090 1407.420 1072.370 1407.700 ;
        RECT 1071.470 1406.800 1071.750 1407.080 ;
        RECT 1072.090 1406.800 1072.370 1407.080 ;
        RECT 1071.470 1406.180 1071.750 1406.460 ;
        RECT 1072.090 1406.180 1072.370 1406.460 ;
        RECT 1071.470 1405.560 1071.750 1405.840 ;
        RECT 1072.090 1405.560 1072.370 1405.840 ;
        RECT 1146.470 1416.280 1146.750 1416.560 ;
        RECT 1147.090 1416.280 1147.370 1416.560 ;
        RECT 1146.470 1415.660 1146.750 1415.940 ;
        RECT 1147.090 1415.660 1147.370 1415.940 ;
        RECT 1146.470 1415.040 1146.750 1415.320 ;
        RECT 1147.090 1415.040 1147.370 1415.320 ;
        RECT 1146.470 1414.420 1146.750 1414.700 ;
        RECT 1147.090 1414.420 1147.370 1414.700 ;
        RECT 1146.470 1413.800 1146.750 1414.080 ;
        RECT 1147.090 1413.800 1147.370 1414.080 ;
        RECT 1146.470 1413.180 1146.750 1413.460 ;
        RECT 1147.090 1413.180 1147.370 1413.460 ;
        RECT 1146.470 1412.560 1146.750 1412.840 ;
        RECT 1147.090 1412.560 1147.370 1412.840 ;
        RECT 1121.470 1409.280 1121.750 1409.560 ;
        RECT 1122.090 1409.280 1122.370 1409.560 ;
        RECT 1121.470 1408.660 1121.750 1408.940 ;
        RECT 1122.090 1408.660 1122.370 1408.940 ;
        RECT 1121.470 1408.040 1121.750 1408.320 ;
        RECT 1122.090 1408.040 1122.370 1408.320 ;
        RECT 1121.470 1407.420 1121.750 1407.700 ;
        RECT 1122.090 1407.420 1122.370 1407.700 ;
        RECT 1121.470 1406.800 1121.750 1407.080 ;
        RECT 1122.090 1406.800 1122.370 1407.080 ;
        RECT 1121.470 1406.180 1121.750 1406.460 ;
        RECT 1122.090 1406.180 1122.370 1406.460 ;
        RECT 1121.470 1405.560 1121.750 1405.840 ;
        RECT 1122.090 1405.560 1122.370 1405.840 ;
        RECT 1196.470 1416.280 1196.750 1416.560 ;
        RECT 1197.090 1416.280 1197.370 1416.560 ;
        RECT 1196.470 1415.660 1196.750 1415.940 ;
        RECT 1197.090 1415.660 1197.370 1415.940 ;
        RECT 1196.470 1415.040 1196.750 1415.320 ;
        RECT 1197.090 1415.040 1197.370 1415.320 ;
        RECT 1196.470 1414.420 1196.750 1414.700 ;
        RECT 1197.090 1414.420 1197.370 1414.700 ;
        RECT 1196.470 1413.800 1196.750 1414.080 ;
        RECT 1197.090 1413.800 1197.370 1414.080 ;
        RECT 1196.470 1413.180 1196.750 1413.460 ;
        RECT 1197.090 1413.180 1197.370 1413.460 ;
        RECT 1196.470 1412.560 1196.750 1412.840 ;
        RECT 1197.090 1412.560 1197.370 1412.840 ;
        RECT 1171.470 1409.280 1171.750 1409.560 ;
        RECT 1172.090 1409.280 1172.370 1409.560 ;
        RECT 1171.470 1408.660 1171.750 1408.940 ;
        RECT 1172.090 1408.660 1172.370 1408.940 ;
        RECT 1171.470 1408.040 1171.750 1408.320 ;
        RECT 1172.090 1408.040 1172.370 1408.320 ;
        RECT 1171.470 1407.420 1171.750 1407.700 ;
        RECT 1172.090 1407.420 1172.370 1407.700 ;
        RECT 1171.470 1406.800 1171.750 1407.080 ;
        RECT 1172.090 1406.800 1172.370 1407.080 ;
        RECT 1171.470 1406.180 1171.750 1406.460 ;
        RECT 1172.090 1406.180 1172.370 1406.460 ;
        RECT 1171.470 1405.560 1171.750 1405.840 ;
        RECT 1172.090 1405.560 1172.370 1405.840 ;
        RECT 1246.470 1416.280 1246.750 1416.560 ;
        RECT 1247.090 1416.280 1247.370 1416.560 ;
        RECT 1246.470 1415.660 1246.750 1415.940 ;
        RECT 1247.090 1415.660 1247.370 1415.940 ;
        RECT 1246.470 1415.040 1246.750 1415.320 ;
        RECT 1247.090 1415.040 1247.370 1415.320 ;
        RECT 1246.470 1414.420 1246.750 1414.700 ;
        RECT 1247.090 1414.420 1247.370 1414.700 ;
        RECT 1246.470 1413.800 1246.750 1414.080 ;
        RECT 1247.090 1413.800 1247.370 1414.080 ;
        RECT 1246.470 1413.180 1246.750 1413.460 ;
        RECT 1247.090 1413.180 1247.370 1413.460 ;
        RECT 1246.470 1412.560 1246.750 1412.840 ;
        RECT 1247.090 1412.560 1247.370 1412.840 ;
        RECT 1221.470 1409.280 1221.750 1409.560 ;
        RECT 1222.090 1409.280 1222.370 1409.560 ;
        RECT 1221.470 1408.660 1221.750 1408.940 ;
        RECT 1222.090 1408.660 1222.370 1408.940 ;
        RECT 1221.470 1408.040 1221.750 1408.320 ;
        RECT 1222.090 1408.040 1222.370 1408.320 ;
        RECT 1221.470 1407.420 1221.750 1407.700 ;
        RECT 1222.090 1407.420 1222.370 1407.700 ;
        RECT 1221.470 1406.800 1221.750 1407.080 ;
        RECT 1222.090 1406.800 1222.370 1407.080 ;
        RECT 1221.470 1406.180 1221.750 1406.460 ;
        RECT 1222.090 1406.180 1222.370 1406.460 ;
        RECT 1221.470 1405.560 1221.750 1405.840 ;
        RECT 1222.090 1405.560 1222.370 1405.840 ;
        RECT 1296.470 1416.280 1296.750 1416.560 ;
        RECT 1297.090 1416.280 1297.370 1416.560 ;
        RECT 1296.470 1415.660 1296.750 1415.940 ;
        RECT 1297.090 1415.660 1297.370 1415.940 ;
        RECT 1296.470 1415.040 1296.750 1415.320 ;
        RECT 1297.090 1415.040 1297.370 1415.320 ;
        RECT 1296.470 1414.420 1296.750 1414.700 ;
        RECT 1297.090 1414.420 1297.370 1414.700 ;
        RECT 1296.470 1413.800 1296.750 1414.080 ;
        RECT 1297.090 1413.800 1297.370 1414.080 ;
        RECT 1296.470 1413.180 1296.750 1413.460 ;
        RECT 1297.090 1413.180 1297.370 1413.460 ;
        RECT 1296.470 1412.560 1296.750 1412.840 ;
        RECT 1297.090 1412.560 1297.370 1412.840 ;
        RECT 1271.470 1409.280 1271.750 1409.560 ;
        RECT 1272.090 1409.280 1272.370 1409.560 ;
        RECT 1271.470 1408.660 1271.750 1408.940 ;
        RECT 1272.090 1408.660 1272.370 1408.940 ;
        RECT 1271.470 1408.040 1271.750 1408.320 ;
        RECT 1272.090 1408.040 1272.370 1408.320 ;
        RECT 1271.470 1407.420 1271.750 1407.700 ;
        RECT 1272.090 1407.420 1272.370 1407.700 ;
        RECT 1271.470 1406.800 1271.750 1407.080 ;
        RECT 1272.090 1406.800 1272.370 1407.080 ;
        RECT 1271.470 1406.180 1271.750 1406.460 ;
        RECT 1272.090 1406.180 1272.370 1406.460 ;
        RECT 1271.470 1405.560 1271.750 1405.840 ;
        RECT 1272.090 1405.560 1272.370 1405.840 ;
        RECT 1346.470 1416.280 1346.750 1416.560 ;
        RECT 1347.090 1416.280 1347.370 1416.560 ;
        RECT 1346.470 1415.660 1346.750 1415.940 ;
        RECT 1347.090 1415.660 1347.370 1415.940 ;
        RECT 1346.470 1415.040 1346.750 1415.320 ;
        RECT 1347.090 1415.040 1347.370 1415.320 ;
        RECT 1346.470 1414.420 1346.750 1414.700 ;
        RECT 1347.090 1414.420 1347.370 1414.700 ;
        RECT 1346.470 1413.800 1346.750 1414.080 ;
        RECT 1347.090 1413.800 1347.370 1414.080 ;
        RECT 1346.470 1413.180 1346.750 1413.460 ;
        RECT 1347.090 1413.180 1347.370 1413.460 ;
        RECT 1346.470 1412.560 1346.750 1412.840 ;
        RECT 1347.090 1412.560 1347.370 1412.840 ;
        RECT 1321.470 1409.280 1321.750 1409.560 ;
        RECT 1322.090 1409.280 1322.370 1409.560 ;
        RECT 1321.470 1408.660 1321.750 1408.940 ;
        RECT 1322.090 1408.660 1322.370 1408.940 ;
        RECT 1321.470 1408.040 1321.750 1408.320 ;
        RECT 1322.090 1408.040 1322.370 1408.320 ;
        RECT 1321.470 1407.420 1321.750 1407.700 ;
        RECT 1322.090 1407.420 1322.370 1407.700 ;
        RECT 1321.470 1406.800 1321.750 1407.080 ;
        RECT 1322.090 1406.800 1322.370 1407.080 ;
        RECT 1321.470 1406.180 1321.750 1406.460 ;
        RECT 1322.090 1406.180 1322.370 1406.460 ;
        RECT 1321.470 1405.560 1321.750 1405.840 ;
        RECT 1322.090 1405.560 1322.370 1405.840 ;
        RECT 1396.470 1416.280 1396.750 1416.560 ;
        RECT 1397.090 1416.280 1397.370 1416.560 ;
        RECT 1396.470 1415.660 1396.750 1415.940 ;
        RECT 1397.090 1415.660 1397.370 1415.940 ;
        RECT 1396.470 1415.040 1396.750 1415.320 ;
        RECT 1397.090 1415.040 1397.370 1415.320 ;
        RECT 1396.470 1414.420 1396.750 1414.700 ;
        RECT 1397.090 1414.420 1397.370 1414.700 ;
        RECT 1396.470 1413.800 1396.750 1414.080 ;
        RECT 1397.090 1413.800 1397.370 1414.080 ;
        RECT 1396.470 1413.180 1396.750 1413.460 ;
        RECT 1397.090 1413.180 1397.370 1413.460 ;
        RECT 1396.470 1412.560 1396.750 1412.840 ;
        RECT 1397.090 1412.560 1397.370 1412.840 ;
        RECT 1371.470 1409.280 1371.750 1409.560 ;
        RECT 1372.090 1409.280 1372.370 1409.560 ;
        RECT 1371.470 1408.660 1371.750 1408.940 ;
        RECT 1372.090 1408.660 1372.370 1408.940 ;
        RECT 1371.470 1408.040 1371.750 1408.320 ;
        RECT 1372.090 1408.040 1372.370 1408.320 ;
        RECT 1371.470 1407.420 1371.750 1407.700 ;
        RECT 1372.090 1407.420 1372.370 1407.700 ;
        RECT 1371.470 1406.800 1371.750 1407.080 ;
        RECT 1372.090 1406.800 1372.370 1407.080 ;
        RECT 1371.470 1406.180 1371.750 1406.460 ;
        RECT 1372.090 1406.180 1372.370 1406.460 ;
        RECT 1371.470 1405.560 1371.750 1405.840 ;
        RECT 1372.090 1405.560 1372.370 1405.840 ;
        RECT 1446.470 1416.280 1446.750 1416.560 ;
        RECT 1447.090 1416.280 1447.370 1416.560 ;
        RECT 1446.470 1415.660 1446.750 1415.940 ;
        RECT 1447.090 1415.660 1447.370 1415.940 ;
        RECT 1446.470 1415.040 1446.750 1415.320 ;
        RECT 1447.090 1415.040 1447.370 1415.320 ;
        RECT 1446.470 1414.420 1446.750 1414.700 ;
        RECT 1447.090 1414.420 1447.370 1414.700 ;
        RECT 1446.470 1413.800 1446.750 1414.080 ;
        RECT 1447.090 1413.800 1447.370 1414.080 ;
        RECT 1446.470 1413.180 1446.750 1413.460 ;
        RECT 1447.090 1413.180 1447.370 1413.460 ;
        RECT 1446.470 1412.560 1446.750 1412.840 ;
        RECT 1447.090 1412.560 1447.370 1412.840 ;
        RECT 1421.470 1409.280 1421.750 1409.560 ;
        RECT 1422.090 1409.280 1422.370 1409.560 ;
        RECT 1421.470 1408.660 1421.750 1408.940 ;
        RECT 1422.090 1408.660 1422.370 1408.940 ;
        RECT 1421.470 1408.040 1421.750 1408.320 ;
        RECT 1422.090 1408.040 1422.370 1408.320 ;
        RECT 1421.470 1407.420 1421.750 1407.700 ;
        RECT 1422.090 1407.420 1422.370 1407.700 ;
        RECT 1421.470 1406.800 1421.750 1407.080 ;
        RECT 1422.090 1406.800 1422.370 1407.080 ;
        RECT 1421.470 1406.180 1421.750 1406.460 ;
        RECT 1422.090 1406.180 1422.370 1406.460 ;
        RECT 1421.470 1405.560 1421.750 1405.840 ;
        RECT 1422.090 1405.560 1422.370 1405.840 ;
        RECT 1496.470 1416.280 1496.750 1416.560 ;
        RECT 1497.090 1416.280 1497.370 1416.560 ;
        RECT 1496.470 1415.660 1496.750 1415.940 ;
        RECT 1497.090 1415.660 1497.370 1415.940 ;
        RECT 1496.470 1415.040 1496.750 1415.320 ;
        RECT 1497.090 1415.040 1497.370 1415.320 ;
        RECT 1496.470 1414.420 1496.750 1414.700 ;
        RECT 1497.090 1414.420 1497.370 1414.700 ;
        RECT 1496.470 1413.800 1496.750 1414.080 ;
        RECT 1497.090 1413.800 1497.370 1414.080 ;
        RECT 1496.470 1413.180 1496.750 1413.460 ;
        RECT 1497.090 1413.180 1497.370 1413.460 ;
        RECT 1496.470 1412.560 1496.750 1412.840 ;
        RECT 1497.090 1412.560 1497.370 1412.840 ;
        RECT 1471.470 1409.280 1471.750 1409.560 ;
        RECT 1472.090 1409.280 1472.370 1409.560 ;
        RECT 1471.470 1408.660 1471.750 1408.940 ;
        RECT 1472.090 1408.660 1472.370 1408.940 ;
        RECT 1471.470 1408.040 1471.750 1408.320 ;
        RECT 1472.090 1408.040 1472.370 1408.320 ;
        RECT 1471.470 1407.420 1471.750 1407.700 ;
        RECT 1472.090 1407.420 1472.370 1407.700 ;
        RECT 1471.470 1406.800 1471.750 1407.080 ;
        RECT 1472.090 1406.800 1472.370 1407.080 ;
        RECT 1471.470 1406.180 1471.750 1406.460 ;
        RECT 1472.090 1406.180 1472.370 1406.460 ;
        RECT 1471.470 1405.560 1471.750 1405.840 ;
        RECT 1472.090 1405.560 1472.370 1405.840 ;
        RECT 1546.470 1416.280 1546.750 1416.560 ;
        RECT 1547.090 1416.280 1547.370 1416.560 ;
        RECT 1546.470 1415.660 1546.750 1415.940 ;
        RECT 1547.090 1415.660 1547.370 1415.940 ;
        RECT 1546.470 1415.040 1546.750 1415.320 ;
        RECT 1547.090 1415.040 1547.370 1415.320 ;
        RECT 1546.470 1414.420 1546.750 1414.700 ;
        RECT 1547.090 1414.420 1547.370 1414.700 ;
        RECT 1546.470 1413.800 1546.750 1414.080 ;
        RECT 1547.090 1413.800 1547.370 1414.080 ;
        RECT 1546.470 1413.180 1546.750 1413.460 ;
        RECT 1547.090 1413.180 1547.370 1413.460 ;
        RECT 1546.470 1412.560 1546.750 1412.840 ;
        RECT 1547.090 1412.560 1547.370 1412.840 ;
        RECT 1521.470 1409.280 1521.750 1409.560 ;
        RECT 1522.090 1409.280 1522.370 1409.560 ;
        RECT 1521.470 1408.660 1521.750 1408.940 ;
        RECT 1522.090 1408.660 1522.370 1408.940 ;
        RECT 1521.470 1408.040 1521.750 1408.320 ;
        RECT 1522.090 1408.040 1522.370 1408.320 ;
        RECT 1521.470 1407.420 1521.750 1407.700 ;
        RECT 1522.090 1407.420 1522.370 1407.700 ;
        RECT 1521.470 1406.800 1521.750 1407.080 ;
        RECT 1522.090 1406.800 1522.370 1407.080 ;
        RECT 1521.470 1406.180 1521.750 1406.460 ;
        RECT 1522.090 1406.180 1522.370 1406.460 ;
        RECT 1521.470 1405.560 1521.750 1405.840 ;
        RECT 1522.090 1405.560 1522.370 1405.840 ;
        RECT 1596.470 1416.280 1596.750 1416.560 ;
        RECT 1597.090 1416.280 1597.370 1416.560 ;
        RECT 1596.470 1415.660 1596.750 1415.940 ;
        RECT 1597.090 1415.660 1597.370 1415.940 ;
        RECT 1596.470 1415.040 1596.750 1415.320 ;
        RECT 1597.090 1415.040 1597.370 1415.320 ;
        RECT 1596.470 1414.420 1596.750 1414.700 ;
        RECT 1597.090 1414.420 1597.370 1414.700 ;
        RECT 1596.470 1413.800 1596.750 1414.080 ;
        RECT 1597.090 1413.800 1597.370 1414.080 ;
        RECT 1596.470 1413.180 1596.750 1413.460 ;
        RECT 1597.090 1413.180 1597.370 1413.460 ;
        RECT 1596.470 1412.560 1596.750 1412.840 ;
        RECT 1597.090 1412.560 1597.370 1412.840 ;
        RECT 1571.470 1409.280 1571.750 1409.560 ;
        RECT 1572.090 1409.280 1572.370 1409.560 ;
        RECT 1571.470 1408.660 1571.750 1408.940 ;
        RECT 1572.090 1408.660 1572.370 1408.940 ;
        RECT 1571.470 1408.040 1571.750 1408.320 ;
        RECT 1572.090 1408.040 1572.370 1408.320 ;
        RECT 1571.470 1407.420 1571.750 1407.700 ;
        RECT 1572.090 1407.420 1572.370 1407.700 ;
        RECT 1571.470 1406.800 1571.750 1407.080 ;
        RECT 1572.090 1406.800 1572.370 1407.080 ;
        RECT 1571.470 1406.180 1571.750 1406.460 ;
        RECT 1572.090 1406.180 1572.370 1406.460 ;
        RECT 1571.470 1405.560 1571.750 1405.840 ;
        RECT 1572.090 1405.560 1572.370 1405.840 ;
        RECT 1646.470 1416.280 1646.750 1416.560 ;
        RECT 1647.090 1416.280 1647.370 1416.560 ;
        RECT 1646.470 1415.660 1646.750 1415.940 ;
        RECT 1647.090 1415.660 1647.370 1415.940 ;
        RECT 1646.470 1415.040 1646.750 1415.320 ;
        RECT 1647.090 1415.040 1647.370 1415.320 ;
        RECT 1646.470 1414.420 1646.750 1414.700 ;
        RECT 1647.090 1414.420 1647.370 1414.700 ;
        RECT 1646.470 1413.800 1646.750 1414.080 ;
        RECT 1647.090 1413.800 1647.370 1414.080 ;
        RECT 1646.470 1413.180 1646.750 1413.460 ;
        RECT 1647.090 1413.180 1647.370 1413.460 ;
        RECT 1646.470 1412.560 1646.750 1412.840 ;
        RECT 1647.090 1412.560 1647.370 1412.840 ;
        RECT 1621.470 1409.280 1621.750 1409.560 ;
        RECT 1622.090 1409.280 1622.370 1409.560 ;
        RECT 1621.470 1408.660 1621.750 1408.940 ;
        RECT 1622.090 1408.660 1622.370 1408.940 ;
        RECT 1621.470 1408.040 1621.750 1408.320 ;
        RECT 1622.090 1408.040 1622.370 1408.320 ;
        RECT 1621.470 1407.420 1621.750 1407.700 ;
        RECT 1622.090 1407.420 1622.370 1407.700 ;
        RECT 1621.470 1406.800 1621.750 1407.080 ;
        RECT 1622.090 1406.800 1622.370 1407.080 ;
        RECT 1621.470 1406.180 1621.750 1406.460 ;
        RECT 1622.090 1406.180 1622.370 1406.460 ;
        RECT 1621.470 1405.560 1621.750 1405.840 ;
        RECT 1622.090 1405.560 1622.370 1405.840 ;
        RECT 1696.470 1416.280 1696.750 1416.560 ;
        RECT 1697.090 1416.280 1697.370 1416.560 ;
        RECT 1696.470 1415.660 1696.750 1415.940 ;
        RECT 1697.090 1415.660 1697.370 1415.940 ;
        RECT 1696.470 1415.040 1696.750 1415.320 ;
        RECT 1697.090 1415.040 1697.370 1415.320 ;
        RECT 1696.470 1414.420 1696.750 1414.700 ;
        RECT 1697.090 1414.420 1697.370 1414.700 ;
        RECT 1696.470 1413.800 1696.750 1414.080 ;
        RECT 1697.090 1413.800 1697.370 1414.080 ;
        RECT 1696.470 1413.180 1696.750 1413.460 ;
        RECT 1697.090 1413.180 1697.370 1413.460 ;
        RECT 1696.470 1412.560 1696.750 1412.840 ;
        RECT 1697.090 1412.560 1697.370 1412.840 ;
        RECT 1671.470 1409.280 1671.750 1409.560 ;
        RECT 1672.090 1409.280 1672.370 1409.560 ;
        RECT 1671.470 1408.660 1671.750 1408.940 ;
        RECT 1672.090 1408.660 1672.370 1408.940 ;
        RECT 1671.470 1408.040 1671.750 1408.320 ;
        RECT 1672.090 1408.040 1672.370 1408.320 ;
        RECT 1671.470 1407.420 1671.750 1407.700 ;
        RECT 1672.090 1407.420 1672.370 1407.700 ;
        RECT 1671.470 1406.800 1671.750 1407.080 ;
        RECT 1672.090 1406.800 1672.370 1407.080 ;
        RECT 1671.470 1406.180 1671.750 1406.460 ;
        RECT 1672.090 1406.180 1672.370 1406.460 ;
        RECT 1671.470 1405.560 1671.750 1405.840 ;
        RECT 1672.090 1405.560 1672.370 1405.840 ;
        RECT 1746.470 1416.280 1746.750 1416.560 ;
        RECT 1747.090 1416.280 1747.370 1416.560 ;
        RECT 1746.470 1415.660 1746.750 1415.940 ;
        RECT 1747.090 1415.660 1747.370 1415.940 ;
        RECT 1746.470 1415.040 1746.750 1415.320 ;
        RECT 1747.090 1415.040 1747.370 1415.320 ;
        RECT 1746.470 1414.420 1746.750 1414.700 ;
        RECT 1747.090 1414.420 1747.370 1414.700 ;
        RECT 1746.470 1413.800 1746.750 1414.080 ;
        RECT 1747.090 1413.800 1747.370 1414.080 ;
        RECT 1746.470 1413.180 1746.750 1413.460 ;
        RECT 1747.090 1413.180 1747.370 1413.460 ;
        RECT 1746.470 1412.560 1746.750 1412.840 ;
        RECT 1747.090 1412.560 1747.370 1412.840 ;
        RECT 1721.470 1409.280 1721.750 1409.560 ;
        RECT 1722.090 1409.280 1722.370 1409.560 ;
        RECT 1721.470 1408.660 1721.750 1408.940 ;
        RECT 1722.090 1408.660 1722.370 1408.940 ;
        RECT 1721.470 1408.040 1721.750 1408.320 ;
        RECT 1722.090 1408.040 1722.370 1408.320 ;
        RECT 1721.470 1407.420 1721.750 1407.700 ;
        RECT 1722.090 1407.420 1722.370 1407.700 ;
        RECT 1721.470 1406.800 1721.750 1407.080 ;
        RECT 1722.090 1406.800 1722.370 1407.080 ;
        RECT 1721.470 1406.180 1721.750 1406.460 ;
        RECT 1722.090 1406.180 1722.370 1406.460 ;
        RECT 1721.470 1405.560 1721.750 1405.840 ;
        RECT 1722.090 1405.560 1722.370 1405.840 ;
        RECT 1796.470 1416.280 1796.750 1416.560 ;
        RECT 1797.090 1416.280 1797.370 1416.560 ;
        RECT 1796.470 1415.660 1796.750 1415.940 ;
        RECT 1797.090 1415.660 1797.370 1415.940 ;
        RECT 1796.470 1415.040 1796.750 1415.320 ;
        RECT 1797.090 1415.040 1797.370 1415.320 ;
        RECT 1796.470 1414.420 1796.750 1414.700 ;
        RECT 1797.090 1414.420 1797.370 1414.700 ;
        RECT 1796.470 1413.800 1796.750 1414.080 ;
        RECT 1797.090 1413.800 1797.370 1414.080 ;
        RECT 1796.470 1413.180 1796.750 1413.460 ;
        RECT 1797.090 1413.180 1797.370 1413.460 ;
        RECT 1796.470 1412.560 1796.750 1412.840 ;
        RECT 1797.090 1412.560 1797.370 1412.840 ;
        RECT 1771.470 1409.280 1771.750 1409.560 ;
        RECT 1772.090 1409.280 1772.370 1409.560 ;
        RECT 1771.470 1408.660 1771.750 1408.940 ;
        RECT 1772.090 1408.660 1772.370 1408.940 ;
        RECT 1771.470 1408.040 1771.750 1408.320 ;
        RECT 1772.090 1408.040 1772.370 1408.320 ;
        RECT 1771.470 1407.420 1771.750 1407.700 ;
        RECT 1772.090 1407.420 1772.370 1407.700 ;
        RECT 1771.470 1406.800 1771.750 1407.080 ;
        RECT 1772.090 1406.800 1772.370 1407.080 ;
        RECT 1771.470 1406.180 1771.750 1406.460 ;
        RECT 1772.090 1406.180 1772.370 1406.460 ;
        RECT 1771.470 1405.560 1771.750 1405.840 ;
        RECT 1772.090 1405.560 1772.370 1405.840 ;
        RECT 1846.470 1416.280 1846.750 1416.560 ;
        RECT 1847.090 1416.280 1847.370 1416.560 ;
        RECT 1846.470 1415.660 1846.750 1415.940 ;
        RECT 1847.090 1415.660 1847.370 1415.940 ;
        RECT 1846.470 1415.040 1846.750 1415.320 ;
        RECT 1847.090 1415.040 1847.370 1415.320 ;
        RECT 1846.470 1414.420 1846.750 1414.700 ;
        RECT 1847.090 1414.420 1847.370 1414.700 ;
        RECT 1846.470 1413.800 1846.750 1414.080 ;
        RECT 1847.090 1413.800 1847.370 1414.080 ;
        RECT 1846.470 1413.180 1846.750 1413.460 ;
        RECT 1847.090 1413.180 1847.370 1413.460 ;
        RECT 1846.470 1412.560 1846.750 1412.840 ;
        RECT 1847.090 1412.560 1847.370 1412.840 ;
        RECT 1821.470 1409.280 1821.750 1409.560 ;
        RECT 1822.090 1409.280 1822.370 1409.560 ;
        RECT 1821.470 1408.660 1821.750 1408.940 ;
        RECT 1822.090 1408.660 1822.370 1408.940 ;
        RECT 1821.470 1408.040 1821.750 1408.320 ;
        RECT 1822.090 1408.040 1822.370 1408.320 ;
        RECT 1821.470 1407.420 1821.750 1407.700 ;
        RECT 1822.090 1407.420 1822.370 1407.700 ;
        RECT 1821.470 1406.800 1821.750 1407.080 ;
        RECT 1822.090 1406.800 1822.370 1407.080 ;
        RECT 1821.470 1406.180 1821.750 1406.460 ;
        RECT 1822.090 1406.180 1822.370 1406.460 ;
        RECT 1821.470 1405.560 1821.750 1405.840 ;
        RECT 1822.090 1405.560 1822.370 1405.840 ;
        RECT 1896.470 1416.280 1896.750 1416.560 ;
        RECT 1897.090 1416.280 1897.370 1416.560 ;
        RECT 1896.470 1415.660 1896.750 1415.940 ;
        RECT 1897.090 1415.660 1897.370 1415.940 ;
        RECT 1896.470 1415.040 1896.750 1415.320 ;
        RECT 1897.090 1415.040 1897.370 1415.320 ;
        RECT 1896.470 1414.420 1896.750 1414.700 ;
        RECT 1897.090 1414.420 1897.370 1414.700 ;
        RECT 1896.470 1413.800 1896.750 1414.080 ;
        RECT 1897.090 1413.800 1897.370 1414.080 ;
        RECT 1896.470 1413.180 1896.750 1413.460 ;
        RECT 1897.090 1413.180 1897.370 1413.460 ;
        RECT 1896.470 1412.560 1896.750 1412.840 ;
        RECT 1897.090 1412.560 1897.370 1412.840 ;
        RECT 1871.470 1409.280 1871.750 1409.560 ;
        RECT 1872.090 1409.280 1872.370 1409.560 ;
        RECT 1871.470 1408.660 1871.750 1408.940 ;
        RECT 1872.090 1408.660 1872.370 1408.940 ;
        RECT 1871.470 1408.040 1871.750 1408.320 ;
        RECT 1872.090 1408.040 1872.370 1408.320 ;
        RECT 1871.470 1407.420 1871.750 1407.700 ;
        RECT 1872.090 1407.420 1872.370 1407.700 ;
        RECT 1871.470 1406.800 1871.750 1407.080 ;
        RECT 1872.090 1406.800 1872.370 1407.080 ;
        RECT 1871.470 1406.180 1871.750 1406.460 ;
        RECT 1872.090 1406.180 1872.370 1406.460 ;
        RECT 1871.470 1405.560 1871.750 1405.840 ;
        RECT 1872.090 1405.560 1872.370 1405.840 ;
        RECT 1946.470 1416.280 1946.750 1416.560 ;
        RECT 1947.090 1416.280 1947.370 1416.560 ;
        RECT 1946.470 1415.660 1946.750 1415.940 ;
        RECT 1947.090 1415.660 1947.370 1415.940 ;
        RECT 1946.470 1415.040 1946.750 1415.320 ;
        RECT 1947.090 1415.040 1947.370 1415.320 ;
        RECT 1946.470 1414.420 1946.750 1414.700 ;
        RECT 1947.090 1414.420 1947.370 1414.700 ;
        RECT 1946.470 1413.800 1946.750 1414.080 ;
        RECT 1947.090 1413.800 1947.370 1414.080 ;
        RECT 1946.470 1413.180 1946.750 1413.460 ;
        RECT 1947.090 1413.180 1947.370 1413.460 ;
        RECT 1946.470 1412.560 1946.750 1412.840 ;
        RECT 1947.090 1412.560 1947.370 1412.840 ;
        RECT 1921.470 1409.280 1921.750 1409.560 ;
        RECT 1922.090 1409.280 1922.370 1409.560 ;
        RECT 1921.470 1408.660 1921.750 1408.940 ;
        RECT 1922.090 1408.660 1922.370 1408.940 ;
        RECT 1921.470 1408.040 1921.750 1408.320 ;
        RECT 1922.090 1408.040 1922.370 1408.320 ;
        RECT 1921.470 1407.420 1921.750 1407.700 ;
        RECT 1922.090 1407.420 1922.370 1407.700 ;
        RECT 1921.470 1406.800 1921.750 1407.080 ;
        RECT 1922.090 1406.800 1922.370 1407.080 ;
        RECT 1921.470 1406.180 1921.750 1406.460 ;
        RECT 1922.090 1406.180 1922.370 1406.460 ;
        RECT 1921.470 1405.560 1921.750 1405.840 ;
        RECT 1922.090 1405.560 1922.370 1405.840 ;
        RECT 1996.470 1416.280 1996.750 1416.560 ;
        RECT 1997.090 1416.280 1997.370 1416.560 ;
        RECT 1996.470 1415.660 1996.750 1415.940 ;
        RECT 1997.090 1415.660 1997.370 1415.940 ;
        RECT 1996.470 1415.040 1996.750 1415.320 ;
        RECT 1997.090 1415.040 1997.370 1415.320 ;
        RECT 1996.470 1414.420 1996.750 1414.700 ;
        RECT 1997.090 1414.420 1997.370 1414.700 ;
        RECT 1996.470 1413.800 1996.750 1414.080 ;
        RECT 1997.090 1413.800 1997.370 1414.080 ;
        RECT 1996.470 1413.180 1996.750 1413.460 ;
        RECT 1997.090 1413.180 1997.370 1413.460 ;
        RECT 1996.470 1412.560 1996.750 1412.840 ;
        RECT 1997.090 1412.560 1997.370 1412.840 ;
        RECT 1971.470 1409.280 1971.750 1409.560 ;
        RECT 1972.090 1409.280 1972.370 1409.560 ;
        RECT 1971.470 1408.660 1971.750 1408.940 ;
        RECT 1972.090 1408.660 1972.370 1408.940 ;
        RECT 1971.470 1408.040 1971.750 1408.320 ;
        RECT 1972.090 1408.040 1972.370 1408.320 ;
        RECT 1971.470 1407.420 1971.750 1407.700 ;
        RECT 1972.090 1407.420 1972.370 1407.700 ;
        RECT 1971.470 1406.800 1971.750 1407.080 ;
        RECT 1972.090 1406.800 1972.370 1407.080 ;
        RECT 1971.470 1406.180 1971.750 1406.460 ;
        RECT 1972.090 1406.180 1972.370 1406.460 ;
        RECT 1971.470 1405.560 1971.750 1405.840 ;
        RECT 1972.090 1405.560 1972.370 1405.840 ;
        RECT 2046.470 1416.280 2046.750 1416.560 ;
        RECT 2047.090 1416.280 2047.370 1416.560 ;
        RECT 2046.470 1415.660 2046.750 1415.940 ;
        RECT 2047.090 1415.660 2047.370 1415.940 ;
        RECT 2046.470 1415.040 2046.750 1415.320 ;
        RECT 2047.090 1415.040 2047.370 1415.320 ;
        RECT 2046.470 1414.420 2046.750 1414.700 ;
        RECT 2047.090 1414.420 2047.370 1414.700 ;
        RECT 2046.470 1413.800 2046.750 1414.080 ;
        RECT 2047.090 1413.800 2047.370 1414.080 ;
        RECT 2046.470 1413.180 2046.750 1413.460 ;
        RECT 2047.090 1413.180 2047.370 1413.460 ;
        RECT 2046.470 1412.560 2046.750 1412.840 ;
        RECT 2047.090 1412.560 2047.370 1412.840 ;
        RECT 2021.470 1409.280 2021.750 1409.560 ;
        RECT 2022.090 1409.280 2022.370 1409.560 ;
        RECT 2021.470 1408.660 2021.750 1408.940 ;
        RECT 2022.090 1408.660 2022.370 1408.940 ;
        RECT 2021.470 1408.040 2021.750 1408.320 ;
        RECT 2022.090 1408.040 2022.370 1408.320 ;
        RECT 2021.470 1407.420 2021.750 1407.700 ;
        RECT 2022.090 1407.420 2022.370 1407.700 ;
        RECT 2021.470 1406.800 2021.750 1407.080 ;
        RECT 2022.090 1406.800 2022.370 1407.080 ;
        RECT 2021.470 1406.180 2021.750 1406.460 ;
        RECT 2022.090 1406.180 2022.370 1406.460 ;
        RECT 2021.470 1405.560 2021.750 1405.840 ;
        RECT 2022.090 1405.560 2022.370 1405.840 ;
        RECT 2096.470 1416.280 2096.750 1416.560 ;
        RECT 2097.090 1416.280 2097.370 1416.560 ;
        RECT 2096.470 1415.660 2096.750 1415.940 ;
        RECT 2097.090 1415.660 2097.370 1415.940 ;
        RECT 2096.470 1415.040 2096.750 1415.320 ;
        RECT 2097.090 1415.040 2097.370 1415.320 ;
        RECT 2096.470 1414.420 2096.750 1414.700 ;
        RECT 2097.090 1414.420 2097.370 1414.700 ;
        RECT 2096.470 1413.800 2096.750 1414.080 ;
        RECT 2097.090 1413.800 2097.370 1414.080 ;
        RECT 2096.470 1413.180 2096.750 1413.460 ;
        RECT 2097.090 1413.180 2097.370 1413.460 ;
        RECT 2096.470 1412.560 2096.750 1412.840 ;
        RECT 2097.090 1412.560 2097.370 1412.840 ;
        RECT 2071.470 1409.280 2071.750 1409.560 ;
        RECT 2072.090 1409.280 2072.370 1409.560 ;
        RECT 2071.470 1408.660 2071.750 1408.940 ;
        RECT 2072.090 1408.660 2072.370 1408.940 ;
        RECT 2071.470 1408.040 2071.750 1408.320 ;
        RECT 2072.090 1408.040 2072.370 1408.320 ;
        RECT 2071.470 1407.420 2071.750 1407.700 ;
        RECT 2072.090 1407.420 2072.370 1407.700 ;
        RECT 2071.470 1406.800 2071.750 1407.080 ;
        RECT 2072.090 1406.800 2072.370 1407.080 ;
        RECT 2071.470 1406.180 2071.750 1406.460 ;
        RECT 2072.090 1406.180 2072.370 1406.460 ;
        RECT 2071.470 1405.560 2071.750 1405.840 ;
        RECT 2072.090 1405.560 2072.370 1405.840 ;
        RECT 2146.470 1416.280 2146.750 1416.560 ;
        RECT 2147.090 1416.280 2147.370 1416.560 ;
        RECT 2146.470 1415.660 2146.750 1415.940 ;
        RECT 2147.090 1415.660 2147.370 1415.940 ;
        RECT 2146.470 1415.040 2146.750 1415.320 ;
        RECT 2147.090 1415.040 2147.370 1415.320 ;
        RECT 2146.470 1414.420 2146.750 1414.700 ;
        RECT 2147.090 1414.420 2147.370 1414.700 ;
        RECT 2146.470 1413.800 2146.750 1414.080 ;
        RECT 2147.090 1413.800 2147.370 1414.080 ;
        RECT 2146.470 1413.180 2146.750 1413.460 ;
        RECT 2147.090 1413.180 2147.370 1413.460 ;
        RECT 2146.470 1412.560 2146.750 1412.840 ;
        RECT 2147.090 1412.560 2147.370 1412.840 ;
        RECT 2121.470 1409.280 2121.750 1409.560 ;
        RECT 2122.090 1409.280 2122.370 1409.560 ;
        RECT 2121.470 1408.660 2121.750 1408.940 ;
        RECT 2122.090 1408.660 2122.370 1408.940 ;
        RECT 2121.470 1408.040 2121.750 1408.320 ;
        RECT 2122.090 1408.040 2122.370 1408.320 ;
        RECT 2121.470 1407.420 2121.750 1407.700 ;
        RECT 2122.090 1407.420 2122.370 1407.700 ;
        RECT 2121.470 1406.800 2121.750 1407.080 ;
        RECT 2122.090 1406.800 2122.370 1407.080 ;
        RECT 2121.470 1406.180 2121.750 1406.460 ;
        RECT 2122.090 1406.180 2122.370 1406.460 ;
        RECT 2121.470 1405.560 2121.750 1405.840 ;
        RECT 2122.090 1405.560 2122.370 1405.840 ;
        RECT 2196.470 1416.280 2196.750 1416.560 ;
        RECT 2197.090 1416.280 2197.370 1416.560 ;
        RECT 2196.470 1415.660 2196.750 1415.940 ;
        RECT 2197.090 1415.660 2197.370 1415.940 ;
        RECT 2196.470 1415.040 2196.750 1415.320 ;
        RECT 2197.090 1415.040 2197.370 1415.320 ;
        RECT 2196.470 1414.420 2196.750 1414.700 ;
        RECT 2197.090 1414.420 2197.370 1414.700 ;
        RECT 2196.470 1413.800 2196.750 1414.080 ;
        RECT 2197.090 1413.800 2197.370 1414.080 ;
        RECT 2196.470 1413.180 2196.750 1413.460 ;
        RECT 2197.090 1413.180 2197.370 1413.460 ;
        RECT 2196.470 1412.560 2196.750 1412.840 ;
        RECT 2197.090 1412.560 2197.370 1412.840 ;
        RECT 2171.470 1409.280 2171.750 1409.560 ;
        RECT 2172.090 1409.280 2172.370 1409.560 ;
        RECT 2171.470 1408.660 2171.750 1408.940 ;
        RECT 2172.090 1408.660 2172.370 1408.940 ;
        RECT 2171.470 1408.040 2171.750 1408.320 ;
        RECT 2172.090 1408.040 2172.370 1408.320 ;
        RECT 2171.470 1407.420 2171.750 1407.700 ;
        RECT 2172.090 1407.420 2172.370 1407.700 ;
        RECT 2171.470 1406.800 2171.750 1407.080 ;
        RECT 2172.090 1406.800 2172.370 1407.080 ;
        RECT 2171.470 1406.180 2171.750 1406.460 ;
        RECT 2172.090 1406.180 2172.370 1406.460 ;
        RECT 2171.470 1405.560 2171.750 1405.840 ;
        RECT 2172.090 1405.560 2172.370 1405.840 ;
        RECT 2246.470 1416.280 2246.750 1416.560 ;
        RECT 2247.090 1416.280 2247.370 1416.560 ;
        RECT 2246.470 1415.660 2246.750 1415.940 ;
        RECT 2247.090 1415.660 2247.370 1415.940 ;
        RECT 2246.470 1415.040 2246.750 1415.320 ;
        RECT 2247.090 1415.040 2247.370 1415.320 ;
        RECT 2246.470 1414.420 2246.750 1414.700 ;
        RECT 2247.090 1414.420 2247.370 1414.700 ;
        RECT 2246.470 1413.800 2246.750 1414.080 ;
        RECT 2247.090 1413.800 2247.370 1414.080 ;
        RECT 2246.470 1413.180 2246.750 1413.460 ;
        RECT 2247.090 1413.180 2247.370 1413.460 ;
        RECT 2246.470 1412.560 2246.750 1412.840 ;
        RECT 2247.090 1412.560 2247.370 1412.840 ;
        RECT 2221.470 1409.280 2221.750 1409.560 ;
        RECT 2222.090 1409.280 2222.370 1409.560 ;
        RECT 2221.470 1408.660 2221.750 1408.940 ;
        RECT 2222.090 1408.660 2222.370 1408.940 ;
        RECT 2221.470 1408.040 2221.750 1408.320 ;
        RECT 2222.090 1408.040 2222.370 1408.320 ;
        RECT 2221.470 1407.420 2221.750 1407.700 ;
        RECT 2222.090 1407.420 2222.370 1407.700 ;
        RECT 2221.470 1406.800 2221.750 1407.080 ;
        RECT 2222.090 1406.800 2222.370 1407.080 ;
        RECT 2221.470 1406.180 2221.750 1406.460 ;
        RECT 2222.090 1406.180 2222.370 1406.460 ;
        RECT 2221.470 1405.560 2221.750 1405.840 ;
        RECT 2222.090 1405.560 2222.370 1405.840 ;
        RECT 2296.470 1416.280 2296.750 1416.560 ;
        RECT 2297.090 1416.280 2297.370 1416.560 ;
        RECT 2296.470 1415.660 2296.750 1415.940 ;
        RECT 2297.090 1415.660 2297.370 1415.940 ;
        RECT 2296.470 1415.040 2296.750 1415.320 ;
        RECT 2297.090 1415.040 2297.370 1415.320 ;
        RECT 2296.470 1414.420 2296.750 1414.700 ;
        RECT 2297.090 1414.420 2297.370 1414.700 ;
        RECT 2296.470 1413.800 2296.750 1414.080 ;
        RECT 2297.090 1413.800 2297.370 1414.080 ;
        RECT 2296.470 1413.180 2296.750 1413.460 ;
        RECT 2297.090 1413.180 2297.370 1413.460 ;
        RECT 2296.470 1412.560 2296.750 1412.840 ;
        RECT 2297.090 1412.560 2297.370 1412.840 ;
        RECT 2271.470 1409.280 2271.750 1409.560 ;
        RECT 2272.090 1409.280 2272.370 1409.560 ;
        RECT 2271.470 1408.660 2271.750 1408.940 ;
        RECT 2272.090 1408.660 2272.370 1408.940 ;
        RECT 2271.470 1408.040 2271.750 1408.320 ;
        RECT 2272.090 1408.040 2272.370 1408.320 ;
        RECT 2271.470 1407.420 2271.750 1407.700 ;
        RECT 2272.090 1407.420 2272.370 1407.700 ;
        RECT 2271.470 1406.800 2271.750 1407.080 ;
        RECT 2272.090 1406.800 2272.370 1407.080 ;
        RECT 2271.470 1406.180 2271.750 1406.460 ;
        RECT 2272.090 1406.180 2272.370 1406.460 ;
        RECT 2271.470 1405.560 2271.750 1405.840 ;
        RECT 2272.090 1405.560 2272.370 1405.840 ;
        RECT 2346.470 1416.280 2346.750 1416.560 ;
        RECT 2347.090 1416.280 2347.370 1416.560 ;
        RECT 2346.470 1415.660 2346.750 1415.940 ;
        RECT 2347.090 1415.660 2347.370 1415.940 ;
        RECT 2346.470 1415.040 2346.750 1415.320 ;
        RECT 2347.090 1415.040 2347.370 1415.320 ;
        RECT 2346.470 1414.420 2346.750 1414.700 ;
        RECT 2347.090 1414.420 2347.370 1414.700 ;
        RECT 2346.470 1413.800 2346.750 1414.080 ;
        RECT 2347.090 1413.800 2347.370 1414.080 ;
        RECT 2346.470 1413.180 2346.750 1413.460 ;
        RECT 2347.090 1413.180 2347.370 1413.460 ;
        RECT 2346.470 1412.560 2346.750 1412.840 ;
        RECT 2347.090 1412.560 2347.370 1412.840 ;
        RECT 2321.470 1409.280 2321.750 1409.560 ;
        RECT 2322.090 1409.280 2322.370 1409.560 ;
        RECT 2321.470 1408.660 2321.750 1408.940 ;
        RECT 2322.090 1408.660 2322.370 1408.940 ;
        RECT 2321.470 1408.040 2321.750 1408.320 ;
        RECT 2322.090 1408.040 2322.370 1408.320 ;
        RECT 2321.470 1407.420 2321.750 1407.700 ;
        RECT 2322.090 1407.420 2322.370 1407.700 ;
        RECT 2321.470 1406.800 2321.750 1407.080 ;
        RECT 2322.090 1406.800 2322.370 1407.080 ;
        RECT 2321.470 1406.180 2321.750 1406.460 ;
        RECT 2322.090 1406.180 2322.370 1406.460 ;
        RECT 2321.470 1405.560 2321.750 1405.840 ;
        RECT 2322.090 1405.560 2322.370 1405.840 ;
        RECT 2396.470 1416.280 2396.750 1416.560 ;
        RECT 2397.090 1416.280 2397.370 1416.560 ;
        RECT 2396.470 1415.660 2396.750 1415.940 ;
        RECT 2397.090 1415.660 2397.370 1415.940 ;
        RECT 2396.470 1415.040 2396.750 1415.320 ;
        RECT 2397.090 1415.040 2397.370 1415.320 ;
        RECT 2396.470 1414.420 2396.750 1414.700 ;
        RECT 2397.090 1414.420 2397.370 1414.700 ;
        RECT 2396.470 1413.800 2396.750 1414.080 ;
        RECT 2397.090 1413.800 2397.370 1414.080 ;
        RECT 2396.470 1413.180 2396.750 1413.460 ;
        RECT 2397.090 1413.180 2397.370 1413.460 ;
        RECT 2396.470 1412.560 2396.750 1412.840 ;
        RECT 2397.090 1412.560 2397.370 1412.840 ;
        RECT 2371.470 1409.280 2371.750 1409.560 ;
        RECT 2372.090 1409.280 2372.370 1409.560 ;
        RECT 2371.470 1408.660 2371.750 1408.940 ;
        RECT 2372.090 1408.660 2372.370 1408.940 ;
        RECT 2371.470 1408.040 2371.750 1408.320 ;
        RECT 2372.090 1408.040 2372.370 1408.320 ;
        RECT 2371.470 1407.420 2371.750 1407.700 ;
        RECT 2372.090 1407.420 2372.370 1407.700 ;
        RECT 2371.470 1406.800 2371.750 1407.080 ;
        RECT 2372.090 1406.800 2372.370 1407.080 ;
        RECT 2371.470 1406.180 2371.750 1406.460 ;
        RECT 2372.090 1406.180 2372.370 1406.460 ;
        RECT 2371.470 1405.560 2371.750 1405.840 ;
        RECT 2372.090 1405.560 2372.370 1405.840 ;
        RECT 2446.470 1416.280 2446.750 1416.560 ;
        RECT 2447.090 1416.280 2447.370 1416.560 ;
        RECT 2446.470 1415.660 2446.750 1415.940 ;
        RECT 2447.090 1415.660 2447.370 1415.940 ;
        RECT 2446.470 1415.040 2446.750 1415.320 ;
        RECT 2447.090 1415.040 2447.370 1415.320 ;
        RECT 2446.470 1414.420 2446.750 1414.700 ;
        RECT 2447.090 1414.420 2447.370 1414.700 ;
        RECT 2446.470 1413.800 2446.750 1414.080 ;
        RECT 2447.090 1413.800 2447.370 1414.080 ;
        RECT 2446.470 1413.180 2446.750 1413.460 ;
        RECT 2447.090 1413.180 2447.370 1413.460 ;
        RECT 2446.470 1412.560 2446.750 1412.840 ;
        RECT 2447.090 1412.560 2447.370 1412.840 ;
        RECT 2421.470 1409.280 2421.750 1409.560 ;
        RECT 2422.090 1409.280 2422.370 1409.560 ;
        RECT 2421.470 1408.660 2421.750 1408.940 ;
        RECT 2422.090 1408.660 2422.370 1408.940 ;
        RECT 2421.470 1408.040 2421.750 1408.320 ;
        RECT 2422.090 1408.040 2422.370 1408.320 ;
        RECT 2421.470 1407.420 2421.750 1407.700 ;
        RECT 2422.090 1407.420 2422.370 1407.700 ;
        RECT 2421.470 1406.800 2421.750 1407.080 ;
        RECT 2422.090 1406.800 2422.370 1407.080 ;
        RECT 2421.470 1406.180 2421.750 1406.460 ;
        RECT 2422.090 1406.180 2422.370 1406.460 ;
        RECT 2421.470 1405.560 2421.750 1405.840 ;
        RECT 2422.090 1405.560 2422.370 1405.840 ;
        RECT 2496.470 1416.280 2496.750 1416.560 ;
        RECT 2497.090 1416.280 2497.370 1416.560 ;
        RECT 2496.470 1415.660 2496.750 1415.940 ;
        RECT 2497.090 1415.660 2497.370 1415.940 ;
        RECT 2496.470 1415.040 2496.750 1415.320 ;
        RECT 2497.090 1415.040 2497.370 1415.320 ;
        RECT 2496.470 1414.420 2496.750 1414.700 ;
        RECT 2497.090 1414.420 2497.370 1414.700 ;
        RECT 2496.470 1413.800 2496.750 1414.080 ;
        RECT 2497.090 1413.800 2497.370 1414.080 ;
        RECT 2496.470 1413.180 2496.750 1413.460 ;
        RECT 2497.090 1413.180 2497.370 1413.460 ;
        RECT 2496.470 1412.560 2496.750 1412.840 ;
        RECT 2497.090 1412.560 2497.370 1412.840 ;
        RECT 2471.470 1409.280 2471.750 1409.560 ;
        RECT 2472.090 1409.280 2472.370 1409.560 ;
        RECT 2471.470 1408.660 2471.750 1408.940 ;
        RECT 2472.090 1408.660 2472.370 1408.940 ;
        RECT 2471.470 1408.040 2471.750 1408.320 ;
        RECT 2472.090 1408.040 2472.370 1408.320 ;
        RECT 2471.470 1407.420 2471.750 1407.700 ;
        RECT 2472.090 1407.420 2472.370 1407.700 ;
        RECT 2471.470 1406.800 2471.750 1407.080 ;
        RECT 2472.090 1406.800 2472.370 1407.080 ;
        RECT 2471.470 1406.180 2471.750 1406.460 ;
        RECT 2472.090 1406.180 2472.370 1406.460 ;
        RECT 2471.470 1405.560 2471.750 1405.840 ;
        RECT 2472.090 1405.560 2472.370 1405.840 ;
        RECT 2546.470 1416.280 2546.750 1416.560 ;
        RECT 2547.090 1416.280 2547.370 1416.560 ;
        RECT 2546.470 1415.660 2546.750 1415.940 ;
        RECT 2547.090 1415.660 2547.370 1415.940 ;
        RECT 2546.470 1415.040 2546.750 1415.320 ;
        RECT 2547.090 1415.040 2547.370 1415.320 ;
        RECT 2546.470 1414.420 2546.750 1414.700 ;
        RECT 2547.090 1414.420 2547.370 1414.700 ;
        RECT 2546.470 1413.800 2546.750 1414.080 ;
        RECT 2547.090 1413.800 2547.370 1414.080 ;
        RECT 2546.470 1413.180 2546.750 1413.460 ;
        RECT 2547.090 1413.180 2547.370 1413.460 ;
        RECT 2546.470 1412.560 2546.750 1412.840 ;
        RECT 2547.090 1412.560 2547.370 1412.840 ;
        RECT 2521.470 1409.280 2521.750 1409.560 ;
        RECT 2522.090 1409.280 2522.370 1409.560 ;
        RECT 2521.470 1408.660 2521.750 1408.940 ;
        RECT 2522.090 1408.660 2522.370 1408.940 ;
        RECT 2521.470 1408.040 2521.750 1408.320 ;
        RECT 2522.090 1408.040 2522.370 1408.320 ;
        RECT 2521.470 1407.420 2521.750 1407.700 ;
        RECT 2522.090 1407.420 2522.370 1407.700 ;
        RECT 2521.470 1406.800 2521.750 1407.080 ;
        RECT 2522.090 1406.800 2522.370 1407.080 ;
        RECT 2521.470 1406.180 2521.750 1406.460 ;
        RECT 2522.090 1406.180 2522.370 1406.460 ;
        RECT 2521.470 1405.560 2521.750 1405.840 ;
        RECT 2522.090 1405.560 2522.370 1405.840 ;
        RECT 2596.470 1416.280 2596.750 1416.560 ;
        RECT 2597.090 1416.280 2597.370 1416.560 ;
        RECT 2596.470 1415.660 2596.750 1415.940 ;
        RECT 2597.090 1415.660 2597.370 1415.940 ;
        RECT 2596.470 1415.040 2596.750 1415.320 ;
        RECT 2597.090 1415.040 2597.370 1415.320 ;
        RECT 2596.470 1414.420 2596.750 1414.700 ;
        RECT 2597.090 1414.420 2597.370 1414.700 ;
        RECT 2596.470 1413.800 2596.750 1414.080 ;
        RECT 2597.090 1413.800 2597.370 1414.080 ;
        RECT 2596.470 1413.180 2596.750 1413.460 ;
        RECT 2597.090 1413.180 2597.370 1413.460 ;
        RECT 2596.470 1412.560 2596.750 1412.840 ;
        RECT 2597.090 1412.560 2597.370 1412.840 ;
        RECT 2571.470 1409.280 2571.750 1409.560 ;
        RECT 2572.090 1409.280 2572.370 1409.560 ;
        RECT 2571.470 1408.660 2571.750 1408.940 ;
        RECT 2572.090 1408.660 2572.370 1408.940 ;
        RECT 2571.470 1408.040 2571.750 1408.320 ;
        RECT 2572.090 1408.040 2572.370 1408.320 ;
        RECT 2571.470 1407.420 2571.750 1407.700 ;
        RECT 2572.090 1407.420 2572.370 1407.700 ;
        RECT 2571.470 1406.800 2571.750 1407.080 ;
        RECT 2572.090 1406.800 2572.370 1407.080 ;
        RECT 2571.470 1406.180 2571.750 1406.460 ;
        RECT 2572.090 1406.180 2572.370 1406.460 ;
        RECT 2571.470 1405.560 2571.750 1405.840 ;
        RECT 2572.090 1405.560 2572.370 1405.840 ;
        RECT 2646.470 1416.280 2646.750 1416.560 ;
        RECT 2647.090 1416.280 2647.370 1416.560 ;
        RECT 2646.470 1415.660 2646.750 1415.940 ;
        RECT 2647.090 1415.660 2647.370 1415.940 ;
        RECT 2646.470 1415.040 2646.750 1415.320 ;
        RECT 2647.090 1415.040 2647.370 1415.320 ;
        RECT 2646.470 1414.420 2646.750 1414.700 ;
        RECT 2647.090 1414.420 2647.370 1414.700 ;
        RECT 2646.470 1413.800 2646.750 1414.080 ;
        RECT 2647.090 1413.800 2647.370 1414.080 ;
        RECT 2646.470 1413.180 2646.750 1413.460 ;
        RECT 2647.090 1413.180 2647.370 1413.460 ;
        RECT 2646.470 1412.560 2646.750 1412.840 ;
        RECT 2647.090 1412.560 2647.370 1412.840 ;
        RECT 2621.470 1409.280 2621.750 1409.560 ;
        RECT 2622.090 1409.280 2622.370 1409.560 ;
        RECT 2621.470 1408.660 2621.750 1408.940 ;
        RECT 2622.090 1408.660 2622.370 1408.940 ;
        RECT 2621.470 1408.040 2621.750 1408.320 ;
        RECT 2622.090 1408.040 2622.370 1408.320 ;
        RECT 2621.470 1407.420 2621.750 1407.700 ;
        RECT 2622.090 1407.420 2622.370 1407.700 ;
        RECT 2621.470 1406.800 2621.750 1407.080 ;
        RECT 2622.090 1406.800 2622.370 1407.080 ;
        RECT 2621.470 1406.180 2621.750 1406.460 ;
        RECT 2622.090 1406.180 2622.370 1406.460 ;
        RECT 2621.470 1405.560 2621.750 1405.840 ;
        RECT 2622.090 1405.560 2622.370 1405.840 ;
        RECT 2696.470 1416.280 2696.750 1416.560 ;
        RECT 2697.090 1416.280 2697.370 1416.560 ;
        RECT 2696.470 1415.660 2696.750 1415.940 ;
        RECT 2697.090 1415.660 2697.370 1415.940 ;
        RECT 2696.470 1415.040 2696.750 1415.320 ;
        RECT 2697.090 1415.040 2697.370 1415.320 ;
        RECT 2696.470 1414.420 2696.750 1414.700 ;
        RECT 2697.090 1414.420 2697.370 1414.700 ;
        RECT 2696.470 1413.800 2696.750 1414.080 ;
        RECT 2697.090 1413.800 2697.370 1414.080 ;
        RECT 2696.470 1413.180 2696.750 1413.460 ;
        RECT 2697.090 1413.180 2697.370 1413.460 ;
        RECT 2696.470 1412.560 2696.750 1412.840 ;
        RECT 2697.090 1412.560 2697.370 1412.840 ;
        RECT 2671.470 1409.280 2671.750 1409.560 ;
        RECT 2672.090 1409.280 2672.370 1409.560 ;
        RECT 2671.470 1408.660 2671.750 1408.940 ;
        RECT 2672.090 1408.660 2672.370 1408.940 ;
        RECT 2671.470 1408.040 2671.750 1408.320 ;
        RECT 2672.090 1408.040 2672.370 1408.320 ;
        RECT 2671.470 1407.420 2671.750 1407.700 ;
        RECT 2672.090 1407.420 2672.370 1407.700 ;
        RECT 2671.470 1406.800 2671.750 1407.080 ;
        RECT 2672.090 1406.800 2672.370 1407.080 ;
        RECT 2671.470 1406.180 2671.750 1406.460 ;
        RECT 2672.090 1406.180 2672.370 1406.460 ;
        RECT 2671.470 1405.560 2671.750 1405.840 ;
        RECT 2672.090 1405.560 2672.370 1405.840 ;
        RECT 2746.470 1416.280 2746.750 1416.560 ;
        RECT 2747.090 1416.280 2747.370 1416.560 ;
        RECT 2746.470 1415.660 2746.750 1415.940 ;
        RECT 2747.090 1415.660 2747.370 1415.940 ;
        RECT 2746.470 1415.040 2746.750 1415.320 ;
        RECT 2747.090 1415.040 2747.370 1415.320 ;
        RECT 2746.470 1414.420 2746.750 1414.700 ;
        RECT 2747.090 1414.420 2747.370 1414.700 ;
        RECT 2746.470 1413.800 2746.750 1414.080 ;
        RECT 2747.090 1413.800 2747.370 1414.080 ;
        RECT 2746.470 1413.180 2746.750 1413.460 ;
        RECT 2747.090 1413.180 2747.370 1413.460 ;
        RECT 2746.470 1412.560 2746.750 1412.840 ;
        RECT 2747.090 1412.560 2747.370 1412.840 ;
        RECT 2721.470 1409.280 2721.750 1409.560 ;
        RECT 2722.090 1409.280 2722.370 1409.560 ;
        RECT 2721.470 1408.660 2721.750 1408.940 ;
        RECT 2722.090 1408.660 2722.370 1408.940 ;
        RECT 2721.470 1408.040 2721.750 1408.320 ;
        RECT 2722.090 1408.040 2722.370 1408.320 ;
        RECT 2721.470 1407.420 2721.750 1407.700 ;
        RECT 2722.090 1407.420 2722.370 1407.700 ;
        RECT 2721.470 1406.800 2721.750 1407.080 ;
        RECT 2722.090 1406.800 2722.370 1407.080 ;
        RECT 2721.470 1406.180 2721.750 1406.460 ;
        RECT 2722.090 1406.180 2722.370 1406.460 ;
        RECT 2721.470 1405.560 2721.750 1405.840 ;
        RECT 2722.090 1405.560 2722.370 1405.840 ;
        RECT 2954.850 1416.580 2955.130 1416.860 ;
        RECT 2955.470 1416.580 2955.750 1416.860 ;
        RECT 2956.090 1416.580 2956.370 1416.860 ;
        RECT 2956.710 1416.580 2956.990 1416.860 ;
        RECT 2957.330 1416.580 2957.610 1416.860 ;
        RECT 2957.950 1416.580 2958.230 1416.860 ;
        RECT 2958.570 1416.580 2958.850 1416.860 ;
        RECT 2954.850 1415.960 2955.130 1416.240 ;
        RECT 2955.470 1415.960 2955.750 1416.240 ;
        RECT 2956.090 1415.960 2956.370 1416.240 ;
        RECT 2956.710 1415.960 2956.990 1416.240 ;
        RECT 2957.330 1415.960 2957.610 1416.240 ;
        RECT 2957.950 1415.960 2958.230 1416.240 ;
        RECT 2958.570 1415.960 2958.850 1416.240 ;
        RECT 2954.850 1415.340 2955.130 1415.620 ;
        RECT 2955.470 1415.340 2955.750 1415.620 ;
        RECT 2956.090 1415.340 2956.370 1415.620 ;
        RECT 2956.710 1415.340 2956.990 1415.620 ;
        RECT 2957.330 1415.340 2957.610 1415.620 ;
        RECT 2957.950 1415.340 2958.230 1415.620 ;
        RECT 2958.570 1415.340 2958.850 1415.620 ;
        RECT 2954.850 1414.720 2955.130 1415.000 ;
        RECT 2955.470 1414.720 2955.750 1415.000 ;
        RECT 2956.090 1414.720 2956.370 1415.000 ;
        RECT 2956.710 1414.720 2956.990 1415.000 ;
        RECT 2957.330 1414.720 2957.610 1415.000 ;
        RECT 2957.950 1414.720 2958.230 1415.000 ;
        RECT 2958.570 1414.720 2958.850 1415.000 ;
        RECT 2954.850 1414.100 2955.130 1414.380 ;
        RECT 2955.470 1414.100 2955.750 1414.380 ;
        RECT 2956.090 1414.100 2956.370 1414.380 ;
        RECT 2956.710 1414.100 2956.990 1414.380 ;
        RECT 2957.330 1414.100 2957.610 1414.380 ;
        RECT 2957.950 1414.100 2958.230 1414.380 ;
        RECT 2958.570 1414.100 2958.850 1414.380 ;
        RECT 2954.850 1413.480 2955.130 1413.760 ;
        RECT 2955.470 1413.480 2955.750 1413.760 ;
        RECT 2956.090 1413.480 2956.370 1413.760 ;
        RECT 2956.710 1413.480 2956.990 1413.760 ;
        RECT 2957.330 1413.480 2957.610 1413.760 ;
        RECT 2957.950 1413.480 2958.230 1413.760 ;
        RECT 2958.570 1413.480 2958.850 1413.760 ;
        RECT 2954.850 1412.860 2955.130 1413.140 ;
        RECT 2955.470 1412.860 2955.750 1413.140 ;
        RECT 2956.090 1412.860 2956.370 1413.140 ;
        RECT 2956.710 1412.860 2956.990 1413.140 ;
        RECT 2957.330 1412.860 2957.610 1413.140 ;
        RECT 2957.950 1412.860 2958.230 1413.140 ;
        RECT 2958.570 1412.860 2958.850 1413.140 ;
        RECT 2771.470 1409.280 2771.750 1409.560 ;
        RECT 2772.090 1409.280 2772.370 1409.560 ;
        RECT 2771.470 1408.660 2771.750 1408.940 ;
        RECT 2772.090 1408.660 2772.370 1408.940 ;
        RECT 2771.470 1408.040 2771.750 1408.320 ;
        RECT 2772.090 1408.040 2772.370 1408.320 ;
        RECT 2771.470 1407.420 2771.750 1407.700 ;
        RECT 2772.090 1407.420 2772.370 1407.700 ;
        RECT 2771.470 1406.800 2771.750 1407.080 ;
        RECT 2772.090 1406.800 2772.370 1407.080 ;
        RECT 2771.470 1406.180 2771.750 1406.460 ;
        RECT 2772.090 1406.180 2772.370 1406.460 ;
        RECT 2771.470 1405.560 2771.750 1405.840 ;
        RECT 2772.090 1405.560 2772.370 1405.840 ;
        RECT 396.500 1367.830 396.780 1368.110 ;
        RECT 398.000 1367.830 398.280 1368.110 ;
        RECT 399.500 1367.830 399.780 1368.110 ;
        RECT 396.500 1332.830 396.780 1333.110 ;
        RECT 398.000 1332.830 398.280 1333.110 ;
        RECT 399.500 1332.830 399.780 1333.110 ;
        RECT 396.500 1297.830 396.780 1298.110 ;
        RECT 398.000 1297.830 398.280 1298.110 ;
        RECT 399.500 1297.830 399.780 1298.110 ;
        RECT 395.740 1276.580 396.020 1276.860 ;
        RECT 396.360 1276.580 396.640 1276.860 ;
        RECT 396.980 1276.580 397.260 1276.860 ;
        RECT 397.600 1276.580 397.880 1276.860 ;
        RECT 398.220 1276.580 398.500 1276.860 ;
        RECT 398.840 1276.580 399.120 1276.860 ;
        RECT 399.460 1276.580 399.740 1276.860 ;
        RECT 395.740 1275.960 396.020 1276.240 ;
        RECT 396.360 1275.960 396.640 1276.240 ;
        RECT 396.980 1275.960 397.260 1276.240 ;
        RECT 397.600 1275.960 397.880 1276.240 ;
        RECT 398.220 1275.960 398.500 1276.240 ;
        RECT 398.840 1275.960 399.120 1276.240 ;
        RECT 399.460 1275.960 399.740 1276.240 ;
        RECT 396.420 1244.960 396.700 1245.240 ;
        RECT 397.920 1244.960 398.200 1245.240 ;
        RECT 399.420 1244.960 399.700 1245.240 ;
        RECT 396.500 1162.830 396.780 1163.110 ;
        RECT 398.000 1162.830 398.280 1163.110 ;
        RECT 399.500 1162.830 399.780 1163.110 ;
        RECT 395.740 1146.580 396.020 1146.860 ;
        RECT 396.360 1146.580 396.640 1146.860 ;
        RECT 396.980 1146.580 397.260 1146.860 ;
        RECT 397.600 1146.580 397.880 1146.860 ;
        RECT 398.220 1146.580 398.500 1146.860 ;
        RECT 398.840 1146.580 399.120 1146.860 ;
        RECT 399.460 1146.580 399.740 1146.860 ;
        RECT 395.740 1145.960 396.020 1146.240 ;
        RECT 396.360 1145.960 396.640 1146.240 ;
        RECT 396.980 1145.960 397.260 1146.240 ;
        RECT 397.600 1145.960 397.880 1146.240 ;
        RECT 398.220 1145.960 398.500 1146.240 ;
        RECT 398.840 1145.960 399.120 1146.240 ;
        RECT 399.460 1145.960 399.740 1146.240 ;
        RECT 396.500 1127.830 396.780 1128.110 ;
        RECT 398.000 1127.830 398.280 1128.110 ;
        RECT 399.500 1127.830 399.780 1128.110 ;
        RECT 396.500 1092.830 396.780 1093.110 ;
        RECT 398.000 1092.830 398.280 1093.110 ;
        RECT 399.500 1092.830 399.780 1093.110 ;
        RECT 396.420 1039.960 396.700 1040.240 ;
        RECT 397.920 1039.960 398.200 1040.240 ;
        RECT 399.420 1039.960 399.700 1040.240 ;
        RECT 395.740 1016.580 396.020 1016.860 ;
        RECT 396.360 1016.580 396.640 1016.860 ;
        RECT 396.980 1016.580 397.260 1016.860 ;
        RECT 397.600 1016.580 397.880 1016.860 ;
        RECT 398.220 1016.580 398.500 1016.860 ;
        RECT 398.840 1016.580 399.120 1016.860 ;
        RECT 399.460 1016.580 399.740 1016.860 ;
        RECT 395.740 1015.960 396.020 1016.240 ;
        RECT 396.360 1015.960 396.640 1016.240 ;
        RECT 396.980 1015.960 397.260 1016.240 ;
        RECT 397.600 1015.960 397.880 1016.240 ;
        RECT 398.220 1015.960 398.500 1016.240 ;
        RECT 398.840 1015.960 399.120 1016.240 ;
        RECT 399.460 1015.960 399.740 1016.240 ;
        RECT 396.500 957.830 396.780 958.110 ;
        RECT 398.000 957.830 398.280 958.110 ;
        RECT 399.500 957.830 399.780 958.110 ;
        RECT 396.500 922.830 396.780 923.110 ;
        RECT 398.000 922.830 398.280 923.110 ;
        RECT 399.500 922.830 399.780 923.110 ;
        RECT 396.500 887.830 396.780 888.110 ;
        RECT 398.000 887.830 398.280 888.110 ;
        RECT 399.500 887.830 399.780 888.110 ;
        RECT 395.740 886.580 396.020 886.860 ;
        RECT 396.360 886.580 396.640 886.860 ;
        RECT 396.980 886.580 397.260 886.860 ;
        RECT 397.600 886.580 397.880 886.860 ;
        RECT 398.220 886.580 398.500 886.860 ;
        RECT 398.840 886.580 399.120 886.860 ;
        RECT 399.460 886.580 399.740 886.860 ;
        RECT 395.740 885.960 396.020 886.240 ;
        RECT 396.360 885.960 396.640 886.240 ;
        RECT 396.980 885.960 397.260 886.240 ;
        RECT 397.600 885.960 397.880 886.240 ;
        RECT 398.220 885.960 398.500 886.240 ;
        RECT 398.840 885.960 399.120 886.240 ;
        RECT 399.460 885.960 399.740 886.240 ;
        RECT 395.740 756.580 396.020 756.860 ;
        RECT 396.360 756.580 396.640 756.860 ;
        RECT 396.980 756.580 397.260 756.860 ;
        RECT 397.600 756.580 397.880 756.860 ;
        RECT 398.220 756.580 398.500 756.860 ;
        RECT 398.840 756.580 399.120 756.860 ;
        RECT 399.460 756.580 399.740 756.860 ;
        RECT 395.740 755.960 396.020 756.240 ;
        RECT 396.360 755.960 396.640 756.240 ;
        RECT 396.980 755.960 397.260 756.240 ;
        RECT 397.600 755.960 397.880 756.240 ;
        RECT 398.220 755.960 398.500 756.240 ;
        RECT 398.840 755.960 399.120 756.240 ;
        RECT 399.460 755.960 399.740 756.240 ;
        RECT 395.740 626.580 396.020 626.860 ;
        RECT 396.360 626.580 396.640 626.860 ;
        RECT 396.980 626.580 397.260 626.860 ;
        RECT 397.600 626.580 397.880 626.860 ;
        RECT 398.220 626.580 398.500 626.860 ;
        RECT 398.840 626.580 399.120 626.860 ;
        RECT 399.460 626.580 399.740 626.860 ;
        RECT 395.740 625.960 396.020 626.240 ;
        RECT 396.360 625.960 396.640 626.240 ;
        RECT 396.980 625.960 397.260 626.240 ;
        RECT 397.600 625.960 397.880 626.240 ;
        RECT 398.220 625.960 398.500 626.240 ;
        RECT 398.840 625.960 399.120 626.240 ;
        RECT 399.460 625.960 399.740 626.240 ;
        RECT 395.740 496.580 396.020 496.860 ;
        RECT 396.360 496.580 396.640 496.860 ;
        RECT 396.980 496.580 397.260 496.860 ;
        RECT 397.600 496.580 397.880 496.860 ;
        RECT 398.220 496.580 398.500 496.860 ;
        RECT 398.840 496.580 399.120 496.860 ;
        RECT 399.460 496.580 399.740 496.860 ;
        RECT 395.740 495.960 396.020 496.240 ;
        RECT 396.360 495.960 396.640 496.240 ;
        RECT 396.980 495.960 397.260 496.240 ;
        RECT 397.600 495.960 397.880 496.240 ;
        RECT 398.220 495.960 398.500 496.240 ;
        RECT 398.840 495.960 399.120 496.240 ;
        RECT 399.460 495.960 399.740 496.240 ;
        RECT 2954.850 1276.580 2955.130 1276.860 ;
        RECT 2955.470 1276.580 2955.750 1276.860 ;
        RECT 2956.090 1276.580 2956.370 1276.860 ;
        RECT 2956.710 1276.580 2956.990 1276.860 ;
        RECT 2957.330 1276.580 2957.610 1276.860 ;
        RECT 2957.950 1276.580 2958.230 1276.860 ;
        RECT 2958.570 1276.580 2958.850 1276.860 ;
        RECT 2954.850 1275.960 2955.130 1276.240 ;
        RECT 2955.470 1275.960 2955.750 1276.240 ;
        RECT 2956.090 1275.960 2956.370 1276.240 ;
        RECT 2956.710 1275.960 2956.990 1276.240 ;
        RECT 2957.330 1275.960 2957.610 1276.240 ;
        RECT 2957.950 1275.960 2958.230 1276.240 ;
        RECT 2958.570 1275.960 2958.850 1276.240 ;
        RECT 2954.850 1146.580 2955.130 1146.860 ;
        RECT 2955.470 1146.580 2955.750 1146.860 ;
        RECT 2956.090 1146.580 2956.370 1146.860 ;
        RECT 2956.710 1146.580 2956.990 1146.860 ;
        RECT 2957.330 1146.580 2957.610 1146.860 ;
        RECT 2957.950 1146.580 2958.230 1146.860 ;
        RECT 2958.570 1146.580 2958.850 1146.860 ;
        RECT 2954.850 1145.960 2955.130 1146.240 ;
        RECT 2955.470 1145.960 2955.750 1146.240 ;
        RECT 2956.090 1145.960 2956.370 1146.240 ;
        RECT 2956.710 1145.960 2956.990 1146.240 ;
        RECT 2957.330 1145.960 2957.610 1146.240 ;
        RECT 2957.950 1145.960 2958.230 1146.240 ;
        RECT 2958.570 1145.960 2958.850 1146.240 ;
        RECT 2954.850 1016.580 2955.130 1016.860 ;
        RECT 2955.470 1016.580 2955.750 1016.860 ;
        RECT 2956.090 1016.580 2956.370 1016.860 ;
        RECT 2956.710 1016.580 2956.990 1016.860 ;
        RECT 2957.330 1016.580 2957.610 1016.860 ;
        RECT 2957.950 1016.580 2958.230 1016.860 ;
        RECT 2958.570 1016.580 2958.850 1016.860 ;
        RECT 2954.850 1015.960 2955.130 1016.240 ;
        RECT 2955.470 1015.960 2955.750 1016.240 ;
        RECT 2956.090 1015.960 2956.370 1016.240 ;
        RECT 2956.710 1015.960 2956.990 1016.240 ;
        RECT 2957.330 1015.960 2957.610 1016.240 ;
        RECT 2957.950 1015.960 2958.230 1016.240 ;
        RECT 2958.570 1015.960 2958.850 1016.240 ;
        RECT 2954.850 886.580 2955.130 886.860 ;
        RECT 2955.470 886.580 2955.750 886.860 ;
        RECT 2956.090 886.580 2956.370 886.860 ;
        RECT 2956.710 886.580 2956.990 886.860 ;
        RECT 2957.330 886.580 2957.610 886.860 ;
        RECT 2957.950 886.580 2958.230 886.860 ;
        RECT 2958.570 886.580 2958.850 886.860 ;
        RECT 2954.850 885.960 2955.130 886.240 ;
        RECT 2955.470 885.960 2955.750 886.240 ;
        RECT 2956.090 885.960 2956.370 886.240 ;
        RECT 2956.710 885.960 2956.990 886.240 ;
        RECT 2957.330 885.960 2957.610 886.240 ;
        RECT 2957.950 885.960 2958.230 886.240 ;
        RECT 2958.570 885.960 2958.850 886.240 ;
        RECT 2954.850 756.580 2955.130 756.860 ;
        RECT 2955.470 756.580 2955.750 756.860 ;
        RECT 2956.090 756.580 2956.370 756.860 ;
        RECT 2956.710 756.580 2956.990 756.860 ;
        RECT 2957.330 756.580 2957.610 756.860 ;
        RECT 2957.950 756.580 2958.230 756.860 ;
        RECT 2958.570 756.580 2958.850 756.860 ;
        RECT 2954.850 755.960 2955.130 756.240 ;
        RECT 2955.470 755.960 2955.750 756.240 ;
        RECT 2956.090 755.960 2956.370 756.240 ;
        RECT 2956.710 755.960 2956.990 756.240 ;
        RECT 2957.330 755.960 2957.610 756.240 ;
        RECT 2957.950 755.960 2958.230 756.240 ;
        RECT 2958.570 755.960 2958.850 756.240 ;
        RECT 2954.850 626.580 2955.130 626.860 ;
        RECT 2955.470 626.580 2955.750 626.860 ;
        RECT 2956.090 626.580 2956.370 626.860 ;
        RECT 2956.710 626.580 2956.990 626.860 ;
        RECT 2957.330 626.580 2957.610 626.860 ;
        RECT 2957.950 626.580 2958.230 626.860 ;
        RECT 2958.570 626.580 2958.850 626.860 ;
        RECT 2954.850 625.960 2955.130 626.240 ;
        RECT 2955.470 625.960 2955.750 626.240 ;
        RECT 2956.090 625.960 2956.370 626.240 ;
        RECT 2956.710 625.960 2956.990 626.240 ;
        RECT 2957.330 625.960 2957.610 626.240 ;
        RECT 2957.950 625.960 2958.230 626.240 ;
        RECT 2958.570 625.960 2958.850 626.240 ;
        RECT 2954.795 600.405 2955.075 600.685 ;
        RECT 2956.295 600.405 2956.575 600.685 ;
        RECT 2957.795 600.405 2958.075 600.685 ;
        RECT 2954.795 584.865 2955.075 585.145 ;
        RECT 2956.295 584.865 2956.575 585.145 ;
        RECT 2957.795 584.865 2958.075 585.145 ;
        RECT 2954.795 569.325 2955.075 569.605 ;
        RECT 2956.295 569.325 2956.575 569.605 ;
        RECT 2957.795 569.325 2958.075 569.605 ;
        RECT 2954.850 496.580 2955.130 496.860 ;
        RECT 2955.470 496.580 2955.750 496.860 ;
        RECT 2956.090 496.580 2956.370 496.860 ;
        RECT 2956.710 496.580 2956.990 496.860 ;
        RECT 2957.330 496.580 2957.610 496.860 ;
        RECT 2957.950 496.580 2958.230 496.860 ;
        RECT 2958.570 496.580 2958.850 496.860 ;
        RECT 2954.850 495.960 2955.130 496.240 ;
        RECT 2955.470 495.960 2955.750 496.240 ;
        RECT 2956.090 495.960 2956.370 496.240 ;
        RECT 2956.710 495.960 2956.990 496.240 ;
        RECT 2957.330 495.960 2957.610 496.240 ;
        RECT 2957.950 495.960 2958.230 496.240 ;
        RECT 2958.570 495.960 2958.850 496.240 ;
        RECT 396.040 399.760 396.320 400.040 ;
        RECT 396.660 399.760 396.940 400.040 ;
        RECT 397.280 399.760 397.560 400.040 ;
        RECT 397.900 399.760 398.180 400.040 ;
        RECT 398.520 399.760 398.800 400.040 ;
        RECT 399.140 399.760 399.420 400.040 ;
        RECT 399.760 399.760 400.040 400.040 ;
        RECT 396.040 399.140 396.320 399.420 ;
        RECT 396.660 399.140 396.940 399.420 ;
        RECT 397.280 399.140 397.560 399.420 ;
        RECT 397.900 399.140 398.180 399.420 ;
        RECT 398.520 399.140 398.800 399.420 ;
        RECT 399.140 399.140 399.420 399.420 ;
        RECT 399.760 399.140 400.040 399.420 ;
        RECT 396.040 398.520 396.320 398.800 ;
        RECT 396.660 398.520 396.940 398.800 ;
        RECT 397.280 398.520 397.560 398.800 ;
        RECT 397.900 398.520 398.180 398.800 ;
        RECT 398.520 398.520 398.800 398.800 ;
        RECT 399.140 398.520 399.420 398.800 ;
        RECT 399.760 398.520 400.040 398.800 ;
        RECT 396.040 397.900 396.320 398.180 ;
        RECT 396.660 397.900 396.940 398.180 ;
        RECT 397.280 397.900 397.560 398.180 ;
        RECT 397.900 397.900 398.180 398.180 ;
        RECT 398.520 397.900 398.800 398.180 ;
        RECT 399.140 397.900 399.420 398.180 ;
        RECT 399.760 397.900 400.040 398.180 ;
        RECT 396.040 397.280 396.320 397.560 ;
        RECT 396.660 397.280 396.940 397.560 ;
        RECT 397.280 397.280 397.560 397.560 ;
        RECT 397.900 397.280 398.180 397.560 ;
        RECT 398.520 397.280 398.800 397.560 ;
        RECT 399.140 397.280 399.420 397.560 ;
        RECT 399.760 397.280 400.040 397.560 ;
        RECT 396.040 396.660 396.320 396.940 ;
        RECT 396.660 396.660 396.940 396.940 ;
        RECT 397.280 396.660 397.560 396.940 ;
        RECT 397.900 396.660 398.180 396.940 ;
        RECT 398.520 396.660 398.800 396.940 ;
        RECT 399.140 396.660 399.420 396.940 ;
        RECT 399.760 396.660 400.040 396.940 ;
        RECT 396.040 396.040 396.320 396.320 ;
        RECT 396.660 396.040 396.940 396.320 ;
        RECT 397.280 396.040 397.560 396.320 ;
        RECT 397.900 396.040 398.180 396.320 ;
        RECT 398.520 396.040 398.800 396.320 ;
        RECT 399.140 396.040 399.420 396.320 ;
        RECT 399.760 396.040 400.040 396.320 ;
        RECT 389.040 392.760 389.320 393.040 ;
        RECT 389.660 392.760 389.940 393.040 ;
        RECT 390.280 392.760 390.560 393.040 ;
        RECT 390.900 392.760 391.180 393.040 ;
        RECT 391.520 392.760 391.800 393.040 ;
        RECT 392.140 392.760 392.420 393.040 ;
        RECT 392.760 392.760 393.040 393.040 ;
        RECT 389.040 392.140 389.320 392.420 ;
        RECT 389.660 392.140 389.940 392.420 ;
        RECT 390.280 392.140 390.560 392.420 ;
        RECT 390.900 392.140 391.180 392.420 ;
        RECT 391.520 392.140 391.800 392.420 ;
        RECT 392.140 392.140 392.420 392.420 ;
        RECT 392.760 392.140 393.040 392.420 ;
        RECT 389.040 391.520 389.320 391.800 ;
        RECT 389.660 391.520 389.940 391.800 ;
        RECT 390.280 391.520 390.560 391.800 ;
        RECT 390.900 391.520 391.180 391.800 ;
        RECT 391.520 391.520 391.800 391.800 ;
        RECT 392.140 391.520 392.420 391.800 ;
        RECT 392.760 391.520 393.040 391.800 ;
        RECT 389.040 390.900 389.320 391.180 ;
        RECT 389.660 390.900 389.940 391.180 ;
        RECT 390.280 390.900 390.560 391.180 ;
        RECT 390.900 390.900 391.180 391.180 ;
        RECT 391.520 390.900 391.800 391.180 ;
        RECT 392.140 390.900 392.420 391.180 ;
        RECT 392.760 390.900 393.040 391.180 ;
        RECT 389.040 390.280 389.320 390.560 ;
        RECT 389.660 390.280 389.940 390.560 ;
        RECT 390.280 390.280 390.560 390.560 ;
        RECT 390.900 390.280 391.180 390.560 ;
        RECT 391.520 390.280 391.800 390.560 ;
        RECT 392.140 390.280 392.420 390.560 ;
        RECT 392.760 390.280 393.040 390.560 ;
        RECT 389.040 389.660 389.320 389.940 ;
        RECT 389.660 389.660 389.940 389.940 ;
        RECT 390.280 389.660 390.560 389.940 ;
        RECT 390.900 389.660 391.180 389.940 ;
        RECT 391.520 389.660 391.800 389.940 ;
        RECT 392.140 389.660 392.420 389.940 ;
        RECT 392.760 389.660 393.040 389.940 ;
        RECT 389.040 389.040 389.320 389.320 ;
        RECT 389.660 389.040 389.940 389.320 ;
        RECT 390.280 389.040 390.560 389.320 ;
        RECT 390.900 389.040 391.180 389.320 ;
        RECT 391.520 389.040 391.800 389.320 ;
        RECT 392.140 389.040 392.420 389.320 ;
        RECT 392.760 389.040 393.040 389.320 ;
        RECT 496.470 399.760 496.750 400.040 ;
        RECT 497.090 399.760 497.370 400.040 ;
        RECT 496.470 399.140 496.750 399.420 ;
        RECT 497.090 399.140 497.370 399.420 ;
        RECT 496.470 398.520 496.750 398.800 ;
        RECT 497.090 398.520 497.370 398.800 ;
        RECT 496.470 397.900 496.750 398.180 ;
        RECT 497.090 397.900 497.370 398.180 ;
        RECT 496.470 397.280 496.750 397.560 ;
        RECT 497.090 397.280 497.370 397.560 ;
        RECT 496.470 396.660 496.750 396.940 ;
        RECT 497.090 396.660 497.370 396.940 ;
        RECT 496.470 396.040 496.750 396.320 ;
        RECT 497.090 396.040 497.370 396.320 ;
        RECT 471.470 392.760 471.750 393.040 ;
        RECT 472.090 392.760 472.370 393.040 ;
        RECT 471.470 392.140 471.750 392.420 ;
        RECT 472.090 392.140 472.370 392.420 ;
        RECT 471.470 391.520 471.750 391.800 ;
        RECT 472.090 391.520 472.370 391.800 ;
        RECT 471.470 390.900 471.750 391.180 ;
        RECT 472.090 390.900 472.370 391.180 ;
        RECT 471.470 390.280 471.750 390.560 ;
        RECT 472.090 390.280 472.370 390.560 ;
        RECT 471.470 389.660 471.750 389.940 ;
        RECT 472.090 389.660 472.370 389.940 ;
        RECT 471.470 389.040 471.750 389.320 ;
        RECT 472.090 389.040 472.370 389.320 ;
        RECT 521.470 392.760 521.750 393.040 ;
        RECT 522.090 392.760 522.370 393.040 ;
        RECT 521.470 392.140 521.750 392.420 ;
        RECT 522.090 392.140 522.370 392.420 ;
        RECT 521.470 391.520 521.750 391.800 ;
        RECT 522.090 391.520 522.370 391.800 ;
        RECT 521.470 390.900 521.750 391.180 ;
        RECT 522.090 390.900 522.370 391.180 ;
        RECT 521.470 390.280 521.750 390.560 ;
        RECT 522.090 390.280 522.370 390.560 ;
        RECT 521.470 389.660 521.750 389.940 ;
        RECT 522.090 389.660 522.370 389.940 ;
        RECT 521.470 389.040 521.750 389.320 ;
        RECT 522.090 389.040 522.370 389.320 ;
        RECT 536.650 399.760 536.930 400.040 ;
        RECT 537.270 399.760 537.550 400.040 ;
        RECT 537.890 399.760 538.170 400.040 ;
        RECT 538.510 399.760 538.790 400.040 ;
        RECT 539.130 399.760 539.410 400.040 ;
        RECT 539.750 399.760 540.030 400.040 ;
        RECT 540.370 399.760 540.650 400.040 ;
        RECT 540.990 399.760 541.270 400.040 ;
        RECT 541.610 399.760 541.890 400.040 ;
        RECT 542.230 399.760 542.510 400.040 ;
        RECT 542.850 399.760 543.130 400.040 ;
        RECT 543.470 399.760 543.750 400.040 ;
        RECT 544.090 399.760 544.370 400.040 ;
        RECT 544.710 399.760 544.990 400.040 ;
        RECT 545.330 399.760 545.610 400.040 ;
        RECT 536.650 399.140 536.930 399.420 ;
        RECT 537.270 399.140 537.550 399.420 ;
        RECT 537.890 399.140 538.170 399.420 ;
        RECT 538.510 399.140 538.790 399.420 ;
        RECT 539.130 399.140 539.410 399.420 ;
        RECT 539.750 399.140 540.030 399.420 ;
        RECT 540.370 399.140 540.650 399.420 ;
        RECT 540.990 399.140 541.270 399.420 ;
        RECT 541.610 399.140 541.890 399.420 ;
        RECT 542.230 399.140 542.510 399.420 ;
        RECT 542.850 399.140 543.130 399.420 ;
        RECT 543.470 399.140 543.750 399.420 ;
        RECT 544.090 399.140 544.370 399.420 ;
        RECT 544.710 399.140 544.990 399.420 ;
        RECT 545.330 399.140 545.610 399.420 ;
        RECT 536.650 398.520 536.930 398.800 ;
        RECT 537.270 398.520 537.550 398.800 ;
        RECT 537.890 398.520 538.170 398.800 ;
        RECT 538.510 398.520 538.790 398.800 ;
        RECT 539.130 398.520 539.410 398.800 ;
        RECT 539.750 398.520 540.030 398.800 ;
        RECT 540.370 398.520 540.650 398.800 ;
        RECT 540.990 398.520 541.270 398.800 ;
        RECT 541.610 398.520 541.890 398.800 ;
        RECT 542.230 398.520 542.510 398.800 ;
        RECT 542.850 398.520 543.130 398.800 ;
        RECT 543.470 398.520 543.750 398.800 ;
        RECT 544.090 398.520 544.370 398.800 ;
        RECT 544.710 398.520 544.990 398.800 ;
        RECT 545.330 398.520 545.610 398.800 ;
        RECT 536.650 397.900 536.930 398.180 ;
        RECT 537.270 397.900 537.550 398.180 ;
        RECT 537.890 397.900 538.170 398.180 ;
        RECT 538.510 397.900 538.790 398.180 ;
        RECT 539.130 397.900 539.410 398.180 ;
        RECT 539.750 397.900 540.030 398.180 ;
        RECT 540.370 397.900 540.650 398.180 ;
        RECT 540.990 397.900 541.270 398.180 ;
        RECT 541.610 397.900 541.890 398.180 ;
        RECT 542.230 397.900 542.510 398.180 ;
        RECT 542.850 397.900 543.130 398.180 ;
        RECT 543.470 397.900 543.750 398.180 ;
        RECT 544.090 397.900 544.370 398.180 ;
        RECT 544.710 397.900 544.990 398.180 ;
        RECT 545.330 397.900 545.610 398.180 ;
        RECT 536.650 397.280 536.930 397.560 ;
        RECT 537.270 397.280 537.550 397.560 ;
        RECT 537.890 397.280 538.170 397.560 ;
        RECT 538.510 397.280 538.790 397.560 ;
        RECT 539.130 397.280 539.410 397.560 ;
        RECT 539.750 397.280 540.030 397.560 ;
        RECT 540.370 397.280 540.650 397.560 ;
        RECT 540.990 397.280 541.270 397.560 ;
        RECT 541.610 397.280 541.890 397.560 ;
        RECT 542.230 397.280 542.510 397.560 ;
        RECT 542.850 397.280 543.130 397.560 ;
        RECT 543.470 397.280 543.750 397.560 ;
        RECT 544.090 397.280 544.370 397.560 ;
        RECT 544.710 397.280 544.990 397.560 ;
        RECT 545.330 397.280 545.610 397.560 ;
        RECT 536.650 396.660 536.930 396.940 ;
        RECT 537.270 396.660 537.550 396.940 ;
        RECT 537.890 396.660 538.170 396.940 ;
        RECT 538.510 396.660 538.790 396.940 ;
        RECT 539.130 396.660 539.410 396.940 ;
        RECT 539.750 396.660 540.030 396.940 ;
        RECT 540.370 396.660 540.650 396.940 ;
        RECT 540.990 396.660 541.270 396.940 ;
        RECT 541.610 396.660 541.890 396.940 ;
        RECT 542.230 396.660 542.510 396.940 ;
        RECT 542.850 396.660 543.130 396.940 ;
        RECT 543.470 396.660 543.750 396.940 ;
        RECT 544.090 396.660 544.370 396.940 ;
        RECT 544.710 396.660 544.990 396.940 ;
        RECT 545.330 396.660 545.610 396.940 ;
        RECT 536.650 396.040 536.930 396.320 ;
        RECT 537.270 396.040 537.550 396.320 ;
        RECT 537.890 396.040 538.170 396.320 ;
        RECT 538.510 396.040 538.790 396.320 ;
        RECT 539.130 396.040 539.410 396.320 ;
        RECT 539.750 396.040 540.030 396.320 ;
        RECT 540.370 396.040 540.650 396.320 ;
        RECT 540.990 396.040 541.270 396.320 ;
        RECT 541.610 396.040 541.890 396.320 ;
        RECT 542.230 396.040 542.510 396.320 ;
        RECT 542.850 396.040 543.130 396.320 ;
        RECT 543.470 396.040 543.750 396.320 ;
        RECT 544.090 396.040 544.370 396.320 ;
        RECT 544.710 396.040 544.990 396.320 ;
        RECT 545.330 396.040 545.610 396.320 ;
        RECT 549.050 399.760 549.330 400.040 ;
        RECT 549.670 399.760 549.950 400.040 ;
        RECT 550.290 399.760 550.570 400.040 ;
        RECT 550.910 399.760 551.190 400.040 ;
        RECT 551.530 399.760 551.810 400.040 ;
        RECT 552.150 399.760 552.430 400.040 ;
        RECT 552.770 399.760 553.050 400.040 ;
        RECT 553.390 399.760 553.670 400.040 ;
        RECT 554.010 399.760 554.290 400.040 ;
        RECT 554.630 399.760 554.910 400.040 ;
        RECT 555.250 399.760 555.530 400.040 ;
        RECT 555.870 399.760 556.150 400.040 ;
        RECT 556.490 399.760 556.770 400.040 ;
        RECT 557.110 399.760 557.390 400.040 ;
        RECT 557.730 399.760 558.010 400.040 ;
        RECT 558.350 399.760 558.630 400.040 ;
        RECT 549.050 399.140 549.330 399.420 ;
        RECT 549.670 399.140 549.950 399.420 ;
        RECT 550.290 399.140 550.570 399.420 ;
        RECT 550.910 399.140 551.190 399.420 ;
        RECT 551.530 399.140 551.810 399.420 ;
        RECT 552.150 399.140 552.430 399.420 ;
        RECT 552.770 399.140 553.050 399.420 ;
        RECT 553.390 399.140 553.670 399.420 ;
        RECT 554.010 399.140 554.290 399.420 ;
        RECT 554.630 399.140 554.910 399.420 ;
        RECT 555.250 399.140 555.530 399.420 ;
        RECT 555.870 399.140 556.150 399.420 ;
        RECT 556.490 399.140 556.770 399.420 ;
        RECT 557.110 399.140 557.390 399.420 ;
        RECT 557.730 399.140 558.010 399.420 ;
        RECT 558.350 399.140 558.630 399.420 ;
        RECT 549.050 398.520 549.330 398.800 ;
        RECT 549.670 398.520 549.950 398.800 ;
        RECT 550.290 398.520 550.570 398.800 ;
        RECT 550.910 398.520 551.190 398.800 ;
        RECT 551.530 398.520 551.810 398.800 ;
        RECT 552.150 398.520 552.430 398.800 ;
        RECT 552.770 398.520 553.050 398.800 ;
        RECT 553.390 398.520 553.670 398.800 ;
        RECT 554.010 398.520 554.290 398.800 ;
        RECT 554.630 398.520 554.910 398.800 ;
        RECT 555.250 398.520 555.530 398.800 ;
        RECT 555.870 398.520 556.150 398.800 ;
        RECT 556.490 398.520 556.770 398.800 ;
        RECT 557.110 398.520 557.390 398.800 ;
        RECT 557.730 398.520 558.010 398.800 ;
        RECT 558.350 398.520 558.630 398.800 ;
        RECT 549.050 397.900 549.330 398.180 ;
        RECT 549.670 397.900 549.950 398.180 ;
        RECT 550.290 397.900 550.570 398.180 ;
        RECT 550.910 397.900 551.190 398.180 ;
        RECT 551.530 397.900 551.810 398.180 ;
        RECT 552.150 397.900 552.430 398.180 ;
        RECT 552.770 397.900 553.050 398.180 ;
        RECT 553.390 397.900 553.670 398.180 ;
        RECT 554.010 397.900 554.290 398.180 ;
        RECT 554.630 397.900 554.910 398.180 ;
        RECT 555.250 397.900 555.530 398.180 ;
        RECT 555.870 397.900 556.150 398.180 ;
        RECT 556.490 397.900 556.770 398.180 ;
        RECT 557.110 397.900 557.390 398.180 ;
        RECT 557.730 397.900 558.010 398.180 ;
        RECT 558.350 397.900 558.630 398.180 ;
        RECT 549.050 397.280 549.330 397.560 ;
        RECT 549.670 397.280 549.950 397.560 ;
        RECT 550.290 397.280 550.570 397.560 ;
        RECT 550.910 397.280 551.190 397.560 ;
        RECT 551.530 397.280 551.810 397.560 ;
        RECT 552.150 397.280 552.430 397.560 ;
        RECT 552.770 397.280 553.050 397.560 ;
        RECT 553.390 397.280 553.670 397.560 ;
        RECT 554.010 397.280 554.290 397.560 ;
        RECT 554.630 397.280 554.910 397.560 ;
        RECT 555.250 397.280 555.530 397.560 ;
        RECT 555.870 397.280 556.150 397.560 ;
        RECT 556.490 397.280 556.770 397.560 ;
        RECT 557.110 397.280 557.390 397.560 ;
        RECT 557.730 397.280 558.010 397.560 ;
        RECT 558.350 397.280 558.630 397.560 ;
        RECT 549.050 396.660 549.330 396.940 ;
        RECT 549.670 396.660 549.950 396.940 ;
        RECT 550.290 396.660 550.570 396.940 ;
        RECT 550.910 396.660 551.190 396.940 ;
        RECT 551.530 396.660 551.810 396.940 ;
        RECT 552.150 396.660 552.430 396.940 ;
        RECT 552.770 396.660 553.050 396.940 ;
        RECT 553.390 396.660 553.670 396.940 ;
        RECT 554.010 396.660 554.290 396.940 ;
        RECT 554.630 396.660 554.910 396.940 ;
        RECT 555.250 396.660 555.530 396.940 ;
        RECT 555.870 396.660 556.150 396.940 ;
        RECT 556.490 396.660 556.770 396.940 ;
        RECT 557.110 396.660 557.390 396.940 ;
        RECT 557.730 396.660 558.010 396.940 ;
        RECT 558.350 396.660 558.630 396.940 ;
        RECT 549.050 396.040 549.330 396.320 ;
        RECT 549.670 396.040 549.950 396.320 ;
        RECT 550.290 396.040 550.570 396.320 ;
        RECT 550.910 396.040 551.190 396.320 ;
        RECT 551.530 396.040 551.810 396.320 ;
        RECT 552.150 396.040 552.430 396.320 ;
        RECT 552.770 396.040 553.050 396.320 ;
        RECT 553.390 396.040 553.670 396.320 ;
        RECT 554.010 396.040 554.290 396.320 ;
        RECT 554.630 396.040 554.910 396.320 ;
        RECT 555.250 396.040 555.530 396.320 ;
        RECT 555.870 396.040 556.150 396.320 ;
        RECT 556.490 396.040 556.770 396.320 ;
        RECT 557.110 396.040 557.390 396.320 ;
        RECT 557.730 396.040 558.010 396.320 ;
        RECT 558.350 396.040 558.630 396.320 ;
        RECT 560.900 399.760 561.180 400.040 ;
        RECT 561.520 399.760 561.800 400.040 ;
        RECT 562.140 399.760 562.420 400.040 ;
        RECT 562.760 399.760 563.040 400.040 ;
        RECT 563.380 399.760 563.660 400.040 ;
        RECT 564.000 399.760 564.280 400.040 ;
        RECT 564.620 399.760 564.900 400.040 ;
        RECT 565.240 399.760 565.520 400.040 ;
        RECT 565.860 399.760 566.140 400.040 ;
        RECT 566.480 399.760 566.760 400.040 ;
        RECT 567.100 399.760 567.380 400.040 ;
        RECT 567.720 399.760 568.000 400.040 ;
        RECT 568.340 399.760 568.620 400.040 ;
        RECT 568.960 399.760 569.240 400.040 ;
        RECT 569.580 399.760 569.860 400.040 ;
        RECT 570.200 399.760 570.480 400.040 ;
        RECT 560.900 399.140 561.180 399.420 ;
        RECT 561.520 399.140 561.800 399.420 ;
        RECT 562.140 399.140 562.420 399.420 ;
        RECT 562.760 399.140 563.040 399.420 ;
        RECT 563.380 399.140 563.660 399.420 ;
        RECT 564.000 399.140 564.280 399.420 ;
        RECT 564.620 399.140 564.900 399.420 ;
        RECT 565.240 399.140 565.520 399.420 ;
        RECT 565.860 399.140 566.140 399.420 ;
        RECT 566.480 399.140 566.760 399.420 ;
        RECT 567.100 399.140 567.380 399.420 ;
        RECT 567.720 399.140 568.000 399.420 ;
        RECT 568.340 399.140 568.620 399.420 ;
        RECT 568.960 399.140 569.240 399.420 ;
        RECT 569.580 399.140 569.860 399.420 ;
        RECT 570.200 399.140 570.480 399.420 ;
        RECT 560.900 398.520 561.180 398.800 ;
        RECT 561.520 398.520 561.800 398.800 ;
        RECT 562.140 398.520 562.420 398.800 ;
        RECT 562.760 398.520 563.040 398.800 ;
        RECT 563.380 398.520 563.660 398.800 ;
        RECT 564.000 398.520 564.280 398.800 ;
        RECT 564.620 398.520 564.900 398.800 ;
        RECT 565.240 398.520 565.520 398.800 ;
        RECT 565.860 398.520 566.140 398.800 ;
        RECT 566.480 398.520 566.760 398.800 ;
        RECT 567.100 398.520 567.380 398.800 ;
        RECT 567.720 398.520 568.000 398.800 ;
        RECT 568.340 398.520 568.620 398.800 ;
        RECT 568.960 398.520 569.240 398.800 ;
        RECT 569.580 398.520 569.860 398.800 ;
        RECT 570.200 398.520 570.480 398.800 ;
        RECT 560.900 397.900 561.180 398.180 ;
        RECT 561.520 397.900 561.800 398.180 ;
        RECT 562.140 397.900 562.420 398.180 ;
        RECT 562.760 397.900 563.040 398.180 ;
        RECT 563.380 397.900 563.660 398.180 ;
        RECT 564.000 397.900 564.280 398.180 ;
        RECT 564.620 397.900 564.900 398.180 ;
        RECT 565.240 397.900 565.520 398.180 ;
        RECT 565.860 397.900 566.140 398.180 ;
        RECT 566.480 397.900 566.760 398.180 ;
        RECT 567.100 397.900 567.380 398.180 ;
        RECT 567.720 397.900 568.000 398.180 ;
        RECT 568.340 397.900 568.620 398.180 ;
        RECT 568.960 397.900 569.240 398.180 ;
        RECT 569.580 397.900 569.860 398.180 ;
        RECT 570.200 397.900 570.480 398.180 ;
        RECT 560.900 397.280 561.180 397.560 ;
        RECT 561.520 397.280 561.800 397.560 ;
        RECT 562.140 397.280 562.420 397.560 ;
        RECT 562.760 397.280 563.040 397.560 ;
        RECT 563.380 397.280 563.660 397.560 ;
        RECT 564.000 397.280 564.280 397.560 ;
        RECT 564.620 397.280 564.900 397.560 ;
        RECT 565.240 397.280 565.520 397.560 ;
        RECT 565.860 397.280 566.140 397.560 ;
        RECT 566.480 397.280 566.760 397.560 ;
        RECT 567.100 397.280 567.380 397.560 ;
        RECT 567.720 397.280 568.000 397.560 ;
        RECT 568.340 397.280 568.620 397.560 ;
        RECT 568.960 397.280 569.240 397.560 ;
        RECT 569.580 397.280 569.860 397.560 ;
        RECT 570.200 397.280 570.480 397.560 ;
        RECT 560.900 396.660 561.180 396.940 ;
        RECT 561.520 396.660 561.800 396.940 ;
        RECT 562.140 396.660 562.420 396.940 ;
        RECT 562.760 396.660 563.040 396.940 ;
        RECT 563.380 396.660 563.660 396.940 ;
        RECT 564.000 396.660 564.280 396.940 ;
        RECT 564.620 396.660 564.900 396.940 ;
        RECT 565.240 396.660 565.520 396.940 ;
        RECT 565.860 396.660 566.140 396.940 ;
        RECT 566.480 396.660 566.760 396.940 ;
        RECT 567.100 396.660 567.380 396.940 ;
        RECT 567.720 396.660 568.000 396.940 ;
        RECT 568.340 396.660 568.620 396.940 ;
        RECT 568.960 396.660 569.240 396.940 ;
        RECT 569.580 396.660 569.860 396.940 ;
        RECT 570.200 396.660 570.480 396.940 ;
        RECT 560.900 396.040 561.180 396.320 ;
        RECT 561.520 396.040 561.800 396.320 ;
        RECT 562.140 396.040 562.420 396.320 ;
        RECT 562.760 396.040 563.040 396.320 ;
        RECT 563.380 396.040 563.660 396.320 ;
        RECT 564.000 396.040 564.280 396.320 ;
        RECT 564.620 396.040 564.900 396.320 ;
        RECT 565.240 396.040 565.520 396.320 ;
        RECT 565.860 396.040 566.140 396.320 ;
        RECT 566.480 396.040 566.760 396.320 ;
        RECT 567.100 396.040 567.380 396.320 ;
        RECT 567.720 396.040 568.000 396.320 ;
        RECT 568.340 396.040 568.620 396.320 ;
        RECT 568.960 396.040 569.240 396.320 ;
        RECT 569.580 396.040 569.860 396.320 ;
        RECT 570.200 396.040 570.480 396.320 ;
        RECT 574.430 399.760 574.710 400.040 ;
        RECT 575.050 399.760 575.330 400.040 ;
        RECT 575.670 399.760 575.950 400.040 ;
        RECT 576.290 399.760 576.570 400.040 ;
        RECT 576.910 399.760 577.190 400.040 ;
        RECT 577.530 399.760 577.810 400.040 ;
        RECT 578.150 399.760 578.430 400.040 ;
        RECT 578.770 399.760 579.050 400.040 ;
        RECT 579.390 399.760 579.670 400.040 ;
        RECT 580.010 399.760 580.290 400.040 ;
        RECT 580.630 399.760 580.910 400.040 ;
        RECT 581.250 399.760 581.530 400.040 ;
        RECT 581.870 399.760 582.150 400.040 ;
        RECT 582.490 399.760 582.770 400.040 ;
        RECT 583.110 399.760 583.390 400.040 ;
        RECT 583.730 399.760 584.010 400.040 ;
        RECT 574.430 399.140 574.710 399.420 ;
        RECT 575.050 399.140 575.330 399.420 ;
        RECT 575.670 399.140 575.950 399.420 ;
        RECT 576.290 399.140 576.570 399.420 ;
        RECT 576.910 399.140 577.190 399.420 ;
        RECT 577.530 399.140 577.810 399.420 ;
        RECT 578.150 399.140 578.430 399.420 ;
        RECT 578.770 399.140 579.050 399.420 ;
        RECT 579.390 399.140 579.670 399.420 ;
        RECT 580.010 399.140 580.290 399.420 ;
        RECT 580.630 399.140 580.910 399.420 ;
        RECT 581.250 399.140 581.530 399.420 ;
        RECT 581.870 399.140 582.150 399.420 ;
        RECT 582.490 399.140 582.770 399.420 ;
        RECT 583.110 399.140 583.390 399.420 ;
        RECT 583.730 399.140 584.010 399.420 ;
        RECT 574.430 398.520 574.710 398.800 ;
        RECT 575.050 398.520 575.330 398.800 ;
        RECT 575.670 398.520 575.950 398.800 ;
        RECT 576.290 398.520 576.570 398.800 ;
        RECT 576.910 398.520 577.190 398.800 ;
        RECT 577.530 398.520 577.810 398.800 ;
        RECT 578.150 398.520 578.430 398.800 ;
        RECT 578.770 398.520 579.050 398.800 ;
        RECT 579.390 398.520 579.670 398.800 ;
        RECT 580.010 398.520 580.290 398.800 ;
        RECT 580.630 398.520 580.910 398.800 ;
        RECT 581.250 398.520 581.530 398.800 ;
        RECT 581.870 398.520 582.150 398.800 ;
        RECT 582.490 398.520 582.770 398.800 ;
        RECT 583.110 398.520 583.390 398.800 ;
        RECT 583.730 398.520 584.010 398.800 ;
        RECT 574.430 397.900 574.710 398.180 ;
        RECT 575.050 397.900 575.330 398.180 ;
        RECT 575.670 397.900 575.950 398.180 ;
        RECT 576.290 397.900 576.570 398.180 ;
        RECT 576.910 397.900 577.190 398.180 ;
        RECT 577.530 397.900 577.810 398.180 ;
        RECT 578.150 397.900 578.430 398.180 ;
        RECT 578.770 397.900 579.050 398.180 ;
        RECT 579.390 397.900 579.670 398.180 ;
        RECT 580.010 397.900 580.290 398.180 ;
        RECT 580.630 397.900 580.910 398.180 ;
        RECT 581.250 397.900 581.530 398.180 ;
        RECT 581.870 397.900 582.150 398.180 ;
        RECT 582.490 397.900 582.770 398.180 ;
        RECT 583.110 397.900 583.390 398.180 ;
        RECT 583.730 397.900 584.010 398.180 ;
        RECT 574.430 397.280 574.710 397.560 ;
        RECT 575.050 397.280 575.330 397.560 ;
        RECT 575.670 397.280 575.950 397.560 ;
        RECT 576.290 397.280 576.570 397.560 ;
        RECT 576.910 397.280 577.190 397.560 ;
        RECT 577.530 397.280 577.810 397.560 ;
        RECT 578.150 397.280 578.430 397.560 ;
        RECT 578.770 397.280 579.050 397.560 ;
        RECT 579.390 397.280 579.670 397.560 ;
        RECT 580.010 397.280 580.290 397.560 ;
        RECT 580.630 397.280 580.910 397.560 ;
        RECT 581.250 397.280 581.530 397.560 ;
        RECT 581.870 397.280 582.150 397.560 ;
        RECT 582.490 397.280 582.770 397.560 ;
        RECT 583.110 397.280 583.390 397.560 ;
        RECT 583.730 397.280 584.010 397.560 ;
        RECT 574.430 396.660 574.710 396.940 ;
        RECT 575.050 396.660 575.330 396.940 ;
        RECT 575.670 396.660 575.950 396.940 ;
        RECT 576.290 396.660 576.570 396.940 ;
        RECT 576.910 396.660 577.190 396.940 ;
        RECT 577.530 396.660 577.810 396.940 ;
        RECT 578.150 396.660 578.430 396.940 ;
        RECT 578.770 396.660 579.050 396.940 ;
        RECT 579.390 396.660 579.670 396.940 ;
        RECT 580.010 396.660 580.290 396.940 ;
        RECT 580.630 396.660 580.910 396.940 ;
        RECT 581.250 396.660 581.530 396.940 ;
        RECT 581.870 396.660 582.150 396.940 ;
        RECT 582.490 396.660 582.770 396.940 ;
        RECT 583.110 396.660 583.390 396.940 ;
        RECT 583.730 396.660 584.010 396.940 ;
        RECT 574.430 396.040 574.710 396.320 ;
        RECT 575.050 396.040 575.330 396.320 ;
        RECT 575.670 396.040 575.950 396.320 ;
        RECT 576.290 396.040 576.570 396.320 ;
        RECT 576.910 396.040 577.190 396.320 ;
        RECT 577.530 396.040 577.810 396.320 ;
        RECT 578.150 396.040 578.430 396.320 ;
        RECT 578.770 396.040 579.050 396.320 ;
        RECT 579.390 396.040 579.670 396.320 ;
        RECT 580.010 396.040 580.290 396.320 ;
        RECT 580.630 396.040 580.910 396.320 ;
        RECT 581.250 396.040 581.530 396.320 ;
        RECT 581.870 396.040 582.150 396.320 ;
        RECT 582.490 396.040 582.770 396.320 ;
        RECT 583.110 396.040 583.390 396.320 ;
        RECT 583.730 396.040 584.010 396.320 ;
        RECT 586.280 399.760 586.560 400.040 ;
        RECT 586.900 399.760 587.180 400.040 ;
        RECT 587.520 399.760 587.800 400.040 ;
        RECT 588.140 399.760 588.420 400.040 ;
        RECT 588.760 399.760 589.040 400.040 ;
        RECT 589.380 399.760 589.660 400.040 ;
        RECT 590.000 399.760 590.280 400.040 ;
        RECT 590.620 399.760 590.900 400.040 ;
        RECT 591.240 399.760 591.520 400.040 ;
        RECT 591.860 399.760 592.140 400.040 ;
        RECT 592.480 399.760 592.760 400.040 ;
        RECT 593.100 399.760 593.380 400.040 ;
        RECT 593.720 399.760 594.000 400.040 ;
        RECT 594.340 399.760 594.620 400.040 ;
        RECT 594.960 399.760 595.240 400.040 ;
        RECT 595.580 399.760 595.860 400.040 ;
        RECT 586.280 399.140 586.560 399.420 ;
        RECT 586.900 399.140 587.180 399.420 ;
        RECT 587.520 399.140 587.800 399.420 ;
        RECT 588.140 399.140 588.420 399.420 ;
        RECT 588.760 399.140 589.040 399.420 ;
        RECT 589.380 399.140 589.660 399.420 ;
        RECT 590.000 399.140 590.280 399.420 ;
        RECT 590.620 399.140 590.900 399.420 ;
        RECT 591.240 399.140 591.520 399.420 ;
        RECT 591.860 399.140 592.140 399.420 ;
        RECT 592.480 399.140 592.760 399.420 ;
        RECT 593.100 399.140 593.380 399.420 ;
        RECT 593.720 399.140 594.000 399.420 ;
        RECT 594.340 399.140 594.620 399.420 ;
        RECT 594.960 399.140 595.240 399.420 ;
        RECT 595.580 399.140 595.860 399.420 ;
        RECT 586.280 398.520 586.560 398.800 ;
        RECT 586.900 398.520 587.180 398.800 ;
        RECT 587.520 398.520 587.800 398.800 ;
        RECT 588.140 398.520 588.420 398.800 ;
        RECT 588.760 398.520 589.040 398.800 ;
        RECT 589.380 398.520 589.660 398.800 ;
        RECT 590.000 398.520 590.280 398.800 ;
        RECT 590.620 398.520 590.900 398.800 ;
        RECT 591.240 398.520 591.520 398.800 ;
        RECT 591.860 398.520 592.140 398.800 ;
        RECT 592.480 398.520 592.760 398.800 ;
        RECT 593.100 398.520 593.380 398.800 ;
        RECT 593.720 398.520 594.000 398.800 ;
        RECT 594.340 398.520 594.620 398.800 ;
        RECT 594.960 398.520 595.240 398.800 ;
        RECT 595.580 398.520 595.860 398.800 ;
        RECT 586.280 397.900 586.560 398.180 ;
        RECT 586.900 397.900 587.180 398.180 ;
        RECT 587.520 397.900 587.800 398.180 ;
        RECT 588.140 397.900 588.420 398.180 ;
        RECT 588.760 397.900 589.040 398.180 ;
        RECT 589.380 397.900 589.660 398.180 ;
        RECT 590.000 397.900 590.280 398.180 ;
        RECT 590.620 397.900 590.900 398.180 ;
        RECT 591.240 397.900 591.520 398.180 ;
        RECT 591.860 397.900 592.140 398.180 ;
        RECT 592.480 397.900 592.760 398.180 ;
        RECT 593.100 397.900 593.380 398.180 ;
        RECT 593.720 397.900 594.000 398.180 ;
        RECT 594.340 397.900 594.620 398.180 ;
        RECT 594.960 397.900 595.240 398.180 ;
        RECT 595.580 397.900 595.860 398.180 ;
        RECT 586.280 397.280 586.560 397.560 ;
        RECT 586.900 397.280 587.180 397.560 ;
        RECT 587.520 397.280 587.800 397.560 ;
        RECT 588.140 397.280 588.420 397.560 ;
        RECT 588.760 397.280 589.040 397.560 ;
        RECT 589.380 397.280 589.660 397.560 ;
        RECT 590.000 397.280 590.280 397.560 ;
        RECT 590.620 397.280 590.900 397.560 ;
        RECT 591.240 397.280 591.520 397.560 ;
        RECT 591.860 397.280 592.140 397.560 ;
        RECT 592.480 397.280 592.760 397.560 ;
        RECT 593.100 397.280 593.380 397.560 ;
        RECT 593.720 397.280 594.000 397.560 ;
        RECT 594.340 397.280 594.620 397.560 ;
        RECT 594.960 397.280 595.240 397.560 ;
        RECT 595.580 397.280 595.860 397.560 ;
        RECT 586.280 396.660 586.560 396.940 ;
        RECT 586.900 396.660 587.180 396.940 ;
        RECT 587.520 396.660 587.800 396.940 ;
        RECT 588.140 396.660 588.420 396.940 ;
        RECT 588.760 396.660 589.040 396.940 ;
        RECT 589.380 396.660 589.660 396.940 ;
        RECT 590.000 396.660 590.280 396.940 ;
        RECT 590.620 396.660 590.900 396.940 ;
        RECT 591.240 396.660 591.520 396.940 ;
        RECT 591.860 396.660 592.140 396.940 ;
        RECT 592.480 396.660 592.760 396.940 ;
        RECT 593.100 396.660 593.380 396.940 ;
        RECT 593.720 396.660 594.000 396.940 ;
        RECT 594.340 396.660 594.620 396.940 ;
        RECT 594.960 396.660 595.240 396.940 ;
        RECT 595.580 396.660 595.860 396.940 ;
        RECT 586.280 396.040 586.560 396.320 ;
        RECT 586.900 396.040 587.180 396.320 ;
        RECT 587.520 396.040 587.800 396.320 ;
        RECT 588.140 396.040 588.420 396.320 ;
        RECT 588.760 396.040 589.040 396.320 ;
        RECT 589.380 396.040 589.660 396.320 ;
        RECT 590.000 396.040 590.280 396.320 ;
        RECT 590.620 396.040 590.900 396.320 ;
        RECT 591.240 396.040 591.520 396.320 ;
        RECT 591.860 396.040 592.140 396.320 ;
        RECT 592.480 396.040 592.760 396.320 ;
        RECT 593.100 396.040 593.380 396.320 ;
        RECT 593.720 396.040 594.000 396.320 ;
        RECT 594.340 396.040 594.620 396.320 ;
        RECT 594.960 396.040 595.240 396.320 ;
        RECT 595.580 396.040 595.860 396.320 ;
        RECT 599.300 399.760 599.580 400.040 ;
        RECT 599.920 399.760 600.200 400.040 ;
        RECT 600.540 399.760 600.820 400.040 ;
        RECT 601.160 399.760 601.440 400.040 ;
        RECT 601.780 399.760 602.060 400.040 ;
        RECT 602.400 399.760 602.680 400.040 ;
        RECT 603.020 399.760 603.300 400.040 ;
        RECT 603.640 399.760 603.920 400.040 ;
        RECT 604.260 399.760 604.540 400.040 ;
        RECT 604.880 399.760 605.160 400.040 ;
        RECT 605.500 399.760 605.780 400.040 ;
        RECT 606.120 399.760 606.400 400.040 ;
        RECT 606.740 399.760 607.020 400.040 ;
        RECT 607.360 399.760 607.640 400.040 ;
        RECT 607.980 399.760 608.260 400.040 ;
        RECT 599.300 399.140 599.580 399.420 ;
        RECT 599.920 399.140 600.200 399.420 ;
        RECT 600.540 399.140 600.820 399.420 ;
        RECT 601.160 399.140 601.440 399.420 ;
        RECT 601.780 399.140 602.060 399.420 ;
        RECT 602.400 399.140 602.680 399.420 ;
        RECT 603.020 399.140 603.300 399.420 ;
        RECT 603.640 399.140 603.920 399.420 ;
        RECT 604.260 399.140 604.540 399.420 ;
        RECT 604.880 399.140 605.160 399.420 ;
        RECT 605.500 399.140 605.780 399.420 ;
        RECT 606.120 399.140 606.400 399.420 ;
        RECT 606.740 399.140 607.020 399.420 ;
        RECT 607.360 399.140 607.640 399.420 ;
        RECT 607.980 399.140 608.260 399.420 ;
        RECT 599.300 398.520 599.580 398.800 ;
        RECT 599.920 398.520 600.200 398.800 ;
        RECT 600.540 398.520 600.820 398.800 ;
        RECT 601.160 398.520 601.440 398.800 ;
        RECT 601.780 398.520 602.060 398.800 ;
        RECT 602.400 398.520 602.680 398.800 ;
        RECT 603.020 398.520 603.300 398.800 ;
        RECT 603.640 398.520 603.920 398.800 ;
        RECT 604.260 398.520 604.540 398.800 ;
        RECT 604.880 398.520 605.160 398.800 ;
        RECT 605.500 398.520 605.780 398.800 ;
        RECT 606.120 398.520 606.400 398.800 ;
        RECT 606.740 398.520 607.020 398.800 ;
        RECT 607.360 398.520 607.640 398.800 ;
        RECT 607.980 398.520 608.260 398.800 ;
        RECT 599.300 397.900 599.580 398.180 ;
        RECT 599.920 397.900 600.200 398.180 ;
        RECT 600.540 397.900 600.820 398.180 ;
        RECT 601.160 397.900 601.440 398.180 ;
        RECT 601.780 397.900 602.060 398.180 ;
        RECT 602.400 397.900 602.680 398.180 ;
        RECT 603.020 397.900 603.300 398.180 ;
        RECT 603.640 397.900 603.920 398.180 ;
        RECT 604.260 397.900 604.540 398.180 ;
        RECT 604.880 397.900 605.160 398.180 ;
        RECT 605.500 397.900 605.780 398.180 ;
        RECT 606.120 397.900 606.400 398.180 ;
        RECT 606.740 397.900 607.020 398.180 ;
        RECT 607.360 397.900 607.640 398.180 ;
        RECT 607.980 397.900 608.260 398.180 ;
        RECT 599.300 397.280 599.580 397.560 ;
        RECT 599.920 397.280 600.200 397.560 ;
        RECT 600.540 397.280 600.820 397.560 ;
        RECT 601.160 397.280 601.440 397.560 ;
        RECT 601.780 397.280 602.060 397.560 ;
        RECT 602.400 397.280 602.680 397.560 ;
        RECT 603.020 397.280 603.300 397.560 ;
        RECT 603.640 397.280 603.920 397.560 ;
        RECT 604.260 397.280 604.540 397.560 ;
        RECT 604.880 397.280 605.160 397.560 ;
        RECT 605.500 397.280 605.780 397.560 ;
        RECT 606.120 397.280 606.400 397.560 ;
        RECT 606.740 397.280 607.020 397.560 ;
        RECT 607.360 397.280 607.640 397.560 ;
        RECT 607.980 397.280 608.260 397.560 ;
        RECT 599.300 396.660 599.580 396.940 ;
        RECT 599.920 396.660 600.200 396.940 ;
        RECT 600.540 396.660 600.820 396.940 ;
        RECT 601.160 396.660 601.440 396.940 ;
        RECT 601.780 396.660 602.060 396.940 ;
        RECT 602.400 396.660 602.680 396.940 ;
        RECT 603.020 396.660 603.300 396.940 ;
        RECT 603.640 396.660 603.920 396.940 ;
        RECT 604.260 396.660 604.540 396.940 ;
        RECT 604.880 396.660 605.160 396.940 ;
        RECT 605.500 396.660 605.780 396.940 ;
        RECT 606.120 396.660 606.400 396.940 ;
        RECT 606.740 396.660 607.020 396.940 ;
        RECT 607.360 396.660 607.640 396.940 ;
        RECT 607.980 396.660 608.260 396.940 ;
        RECT 599.300 396.040 599.580 396.320 ;
        RECT 599.920 396.040 600.200 396.320 ;
        RECT 600.540 396.040 600.820 396.320 ;
        RECT 601.160 396.040 601.440 396.320 ;
        RECT 601.780 396.040 602.060 396.320 ;
        RECT 602.400 396.040 602.680 396.320 ;
        RECT 603.020 396.040 603.300 396.320 ;
        RECT 603.640 396.040 603.920 396.320 ;
        RECT 604.260 396.040 604.540 396.320 ;
        RECT 604.880 396.040 605.160 396.320 ;
        RECT 605.500 396.040 605.780 396.320 ;
        RECT 606.120 396.040 606.400 396.320 ;
        RECT 606.740 396.040 607.020 396.320 ;
        RECT 607.360 396.040 607.640 396.320 ;
        RECT 607.980 396.040 608.260 396.320 ;
        RECT 646.470 399.760 646.750 400.040 ;
        RECT 647.090 399.760 647.370 400.040 ;
        RECT 646.470 399.140 646.750 399.420 ;
        RECT 647.090 399.140 647.370 399.420 ;
        RECT 646.470 398.520 646.750 398.800 ;
        RECT 647.090 398.520 647.370 398.800 ;
        RECT 646.470 397.900 646.750 398.180 ;
        RECT 647.090 397.900 647.370 398.180 ;
        RECT 646.470 397.280 646.750 397.560 ;
        RECT 647.090 397.280 647.370 397.560 ;
        RECT 646.470 396.660 646.750 396.940 ;
        RECT 647.090 396.660 647.370 396.940 ;
        RECT 646.470 396.040 646.750 396.320 ;
        RECT 647.090 396.040 647.370 396.320 ;
        RECT 621.470 392.760 621.750 393.040 ;
        RECT 622.090 392.760 622.370 393.040 ;
        RECT 621.470 392.140 621.750 392.420 ;
        RECT 622.090 392.140 622.370 392.420 ;
        RECT 621.470 391.520 621.750 391.800 ;
        RECT 622.090 391.520 622.370 391.800 ;
        RECT 621.470 390.900 621.750 391.180 ;
        RECT 622.090 390.900 622.370 391.180 ;
        RECT 621.470 390.280 621.750 390.560 ;
        RECT 622.090 390.280 622.370 390.560 ;
        RECT 621.470 389.660 621.750 389.940 ;
        RECT 622.090 389.660 622.370 389.940 ;
        RECT 621.470 389.040 621.750 389.320 ;
        RECT 622.090 389.040 622.370 389.320 ;
        RECT 696.470 399.760 696.750 400.040 ;
        RECT 697.090 399.760 697.370 400.040 ;
        RECT 696.470 399.140 696.750 399.420 ;
        RECT 697.090 399.140 697.370 399.420 ;
        RECT 696.470 398.520 696.750 398.800 ;
        RECT 697.090 398.520 697.370 398.800 ;
        RECT 696.470 397.900 696.750 398.180 ;
        RECT 697.090 397.900 697.370 398.180 ;
        RECT 696.470 397.280 696.750 397.560 ;
        RECT 697.090 397.280 697.370 397.560 ;
        RECT 696.470 396.660 696.750 396.940 ;
        RECT 697.090 396.660 697.370 396.940 ;
        RECT 696.470 396.040 696.750 396.320 ;
        RECT 697.090 396.040 697.370 396.320 ;
        RECT 671.470 392.760 671.750 393.040 ;
        RECT 672.090 392.760 672.370 393.040 ;
        RECT 671.470 392.140 671.750 392.420 ;
        RECT 672.090 392.140 672.370 392.420 ;
        RECT 671.470 391.520 671.750 391.800 ;
        RECT 672.090 391.520 672.370 391.800 ;
        RECT 671.470 390.900 671.750 391.180 ;
        RECT 672.090 390.900 672.370 391.180 ;
        RECT 671.470 390.280 671.750 390.560 ;
        RECT 672.090 390.280 672.370 390.560 ;
        RECT 671.470 389.660 671.750 389.940 ;
        RECT 672.090 389.660 672.370 389.940 ;
        RECT 671.470 389.040 671.750 389.320 ;
        RECT 672.090 389.040 672.370 389.320 ;
        RECT 746.470 399.760 746.750 400.040 ;
        RECT 747.090 399.760 747.370 400.040 ;
        RECT 746.470 399.140 746.750 399.420 ;
        RECT 747.090 399.140 747.370 399.420 ;
        RECT 746.470 398.520 746.750 398.800 ;
        RECT 747.090 398.520 747.370 398.800 ;
        RECT 746.470 397.900 746.750 398.180 ;
        RECT 747.090 397.900 747.370 398.180 ;
        RECT 746.470 397.280 746.750 397.560 ;
        RECT 747.090 397.280 747.370 397.560 ;
        RECT 746.470 396.660 746.750 396.940 ;
        RECT 747.090 396.660 747.370 396.940 ;
        RECT 746.470 396.040 746.750 396.320 ;
        RECT 747.090 396.040 747.370 396.320 ;
        RECT 721.470 392.760 721.750 393.040 ;
        RECT 722.090 392.760 722.370 393.040 ;
        RECT 721.470 392.140 721.750 392.420 ;
        RECT 722.090 392.140 722.370 392.420 ;
        RECT 721.470 391.520 721.750 391.800 ;
        RECT 722.090 391.520 722.370 391.800 ;
        RECT 721.470 390.900 721.750 391.180 ;
        RECT 722.090 390.900 722.370 391.180 ;
        RECT 721.470 390.280 721.750 390.560 ;
        RECT 722.090 390.280 722.370 390.560 ;
        RECT 721.470 389.660 721.750 389.940 ;
        RECT 722.090 389.660 722.370 389.940 ;
        RECT 721.470 389.040 721.750 389.320 ;
        RECT 722.090 389.040 722.370 389.320 ;
        RECT 796.470 399.760 796.750 400.040 ;
        RECT 797.090 399.760 797.370 400.040 ;
        RECT 796.470 399.140 796.750 399.420 ;
        RECT 797.090 399.140 797.370 399.420 ;
        RECT 796.470 398.520 796.750 398.800 ;
        RECT 797.090 398.520 797.370 398.800 ;
        RECT 796.470 397.900 796.750 398.180 ;
        RECT 797.090 397.900 797.370 398.180 ;
        RECT 796.470 397.280 796.750 397.560 ;
        RECT 797.090 397.280 797.370 397.560 ;
        RECT 796.470 396.660 796.750 396.940 ;
        RECT 797.090 396.660 797.370 396.940 ;
        RECT 796.470 396.040 796.750 396.320 ;
        RECT 797.090 396.040 797.370 396.320 ;
        RECT 771.470 392.760 771.750 393.040 ;
        RECT 772.090 392.760 772.370 393.040 ;
        RECT 771.470 392.140 771.750 392.420 ;
        RECT 772.090 392.140 772.370 392.420 ;
        RECT 771.470 391.520 771.750 391.800 ;
        RECT 772.090 391.520 772.370 391.800 ;
        RECT 771.470 390.900 771.750 391.180 ;
        RECT 772.090 390.900 772.370 391.180 ;
        RECT 771.470 390.280 771.750 390.560 ;
        RECT 772.090 390.280 772.370 390.560 ;
        RECT 771.470 389.660 771.750 389.940 ;
        RECT 772.090 389.660 772.370 389.940 ;
        RECT 771.470 389.040 771.750 389.320 ;
        RECT 772.090 389.040 772.370 389.320 ;
        RECT 846.470 399.760 846.750 400.040 ;
        RECT 847.090 399.760 847.370 400.040 ;
        RECT 846.470 399.140 846.750 399.420 ;
        RECT 847.090 399.140 847.370 399.420 ;
        RECT 846.470 398.520 846.750 398.800 ;
        RECT 847.090 398.520 847.370 398.800 ;
        RECT 846.470 397.900 846.750 398.180 ;
        RECT 847.090 397.900 847.370 398.180 ;
        RECT 846.470 397.280 846.750 397.560 ;
        RECT 847.090 397.280 847.370 397.560 ;
        RECT 846.470 396.660 846.750 396.940 ;
        RECT 847.090 396.660 847.370 396.940 ;
        RECT 846.470 396.040 846.750 396.320 ;
        RECT 847.090 396.040 847.370 396.320 ;
        RECT 821.470 392.760 821.750 393.040 ;
        RECT 822.090 392.760 822.370 393.040 ;
        RECT 821.470 392.140 821.750 392.420 ;
        RECT 822.090 392.140 822.370 392.420 ;
        RECT 821.470 391.520 821.750 391.800 ;
        RECT 822.090 391.520 822.370 391.800 ;
        RECT 821.470 390.900 821.750 391.180 ;
        RECT 822.090 390.900 822.370 391.180 ;
        RECT 821.470 390.280 821.750 390.560 ;
        RECT 822.090 390.280 822.370 390.560 ;
        RECT 821.470 389.660 821.750 389.940 ;
        RECT 822.090 389.660 822.370 389.940 ;
        RECT 821.470 389.040 821.750 389.320 ;
        RECT 822.090 389.040 822.370 389.320 ;
        RECT 896.470 399.760 896.750 400.040 ;
        RECT 897.090 399.760 897.370 400.040 ;
        RECT 896.470 399.140 896.750 399.420 ;
        RECT 897.090 399.140 897.370 399.420 ;
        RECT 896.470 398.520 896.750 398.800 ;
        RECT 897.090 398.520 897.370 398.800 ;
        RECT 896.470 397.900 896.750 398.180 ;
        RECT 897.090 397.900 897.370 398.180 ;
        RECT 896.470 397.280 896.750 397.560 ;
        RECT 897.090 397.280 897.370 397.560 ;
        RECT 896.470 396.660 896.750 396.940 ;
        RECT 897.090 396.660 897.370 396.940 ;
        RECT 896.470 396.040 896.750 396.320 ;
        RECT 897.090 396.040 897.370 396.320 ;
        RECT 871.470 392.760 871.750 393.040 ;
        RECT 872.090 392.760 872.370 393.040 ;
        RECT 871.470 392.140 871.750 392.420 ;
        RECT 872.090 392.140 872.370 392.420 ;
        RECT 871.470 391.520 871.750 391.800 ;
        RECT 872.090 391.520 872.370 391.800 ;
        RECT 871.470 390.900 871.750 391.180 ;
        RECT 872.090 390.900 872.370 391.180 ;
        RECT 871.470 390.280 871.750 390.560 ;
        RECT 872.090 390.280 872.370 390.560 ;
        RECT 871.470 389.660 871.750 389.940 ;
        RECT 872.090 389.660 872.370 389.940 ;
        RECT 871.470 389.040 871.750 389.320 ;
        RECT 872.090 389.040 872.370 389.320 ;
        RECT 946.470 399.760 946.750 400.040 ;
        RECT 947.090 399.760 947.370 400.040 ;
        RECT 946.470 399.140 946.750 399.420 ;
        RECT 947.090 399.140 947.370 399.420 ;
        RECT 946.470 398.520 946.750 398.800 ;
        RECT 947.090 398.520 947.370 398.800 ;
        RECT 946.470 397.900 946.750 398.180 ;
        RECT 947.090 397.900 947.370 398.180 ;
        RECT 946.470 397.280 946.750 397.560 ;
        RECT 947.090 397.280 947.370 397.560 ;
        RECT 946.470 396.660 946.750 396.940 ;
        RECT 947.090 396.660 947.370 396.940 ;
        RECT 946.470 396.040 946.750 396.320 ;
        RECT 947.090 396.040 947.370 396.320 ;
        RECT 921.470 392.760 921.750 393.040 ;
        RECT 922.090 392.760 922.370 393.040 ;
        RECT 921.470 392.140 921.750 392.420 ;
        RECT 922.090 392.140 922.370 392.420 ;
        RECT 921.470 391.520 921.750 391.800 ;
        RECT 922.090 391.520 922.370 391.800 ;
        RECT 921.470 390.900 921.750 391.180 ;
        RECT 922.090 390.900 922.370 391.180 ;
        RECT 921.470 390.280 921.750 390.560 ;
        RECT 922.090 390.280 922.370 390.560 ;
        RECT 921.470 389.660 921.750 389.940 ;
        RECT 922.090 389.660 922.370 389.940 ;
        RECT 921.470 389.040 921.750 389.320 ;
        RECT 922.090 389.040 922.370 389.320 ;
        RECT 996.470 399.760 996.750 400.040 ;
        RECT 997.090 399.760 997.370 400.040 ;
        RECT 996.470 399.140 996.750 399.420 ;
        RECT 997.090 399.140 997.370 399.420 ;
        RECT 996.470 398.520 996.750 398.800 ;
        RECT 997.090 398.520 997.370 398.800 ;
        RECT 996.470 397.900 996.750 398.180 ;
        RECT 997.090 397.900 997.370 398.180 ;
        RECT 996.470 397.280 996.750 397.560 ;
        RECT 997.090 397.280 997.370 397.560 ;
        RECT 996.470 396.660 996.750 396.940 ;
        RECT 997.090 396.660 997.370 396.940 ;
        RECT 996.470 396.040 996.750 396.320 ;
        RECT 997.090 396.040 997.370 396.320 ;
        RECT 971.470 392.760 971.750 393.040 ;
        RECT 972.090 392.760 972.370 393.040 ;
        RECT 971.470 392.140 971.750 392.420 ;
        RECT 972.090 392.140 972.370 392.420 ;
        RECT 971.470 391.520 971.750 391.800 ;
        RECT 972.090 391.520 972.370 391.800 ;
        RECT 971.470 390.900 971.750 391.180 ;
        RECT 972.090 390.900 972.370 391.180 ;
        RECT 971.470 390.280 971.750 390.560 ;
        RECT 972.090 390.280 972.370 390.560 ;
        RECT 971.470 389.660 971.750 389.940 ;
        RECT 972.090 389.660 972.370 389.940 ;
        RECT 971.470 389.040 971.750 389.320 ;
        RECT 972.090 389.040 972.370 389.320 ;
        RECT 1046.470 399.760 1046.750 400.040 ;
        RECT 1047.090 399.760 1047.370 400.040 ;
        RECT 1046.470 399.140 1046.750 399.420 ;
        RECT 1047.090 399.140 1047.370 399.420 ;
        RECT 1046.470 398.520 1046.750 398.800 ;
        RECT 1047.090 398.520 1047.370 398.800 ;
        RECT 1046.470 397.900 1046.750 398.180 ;
        RECT 1047.090 397.900 1047.370 398.180 ;
        RECT 1046.470 397.280 1046.750 397.560 ;
        RECT 1047.090 397.280 1047.370 397.560 ;
        RECT 1046.470 396.660 1046.750 396.940 ;
        RECT 1047.090 396.660 1047.370 396.940 ;
        RECT 1046.470 396.040 1046.750 396.320 ;
        RECT 1047.090 396.040 1047.370 396.320 ;
        RECT 1021.470 392.760 1021.750 393.040 ;
        RECT 1022.090 392.760 1022.370 393.040 ;
        RECT 1021.470 392.140 1021.750 392.420 ;
        RECT 1022.090 392.140 1022.370 392.420 ;
        RECT 1021.470 391.520 1021.750 391.800 ;
        RECT 1022.090 391.520 1022.370 391.800 ;
        RECT 1021.470 390.900 1021.750 391.180 ;
        RECT 1022.090 390.900 1022.370 391.180 ;
        RECT 1021.470 390.280 1021.750 390.560 ;
        RECT 1022.090 390.280 1022.370 390.560 ;
        RECT 1021.470 389.660 1021.750 389.940 ;
        RECT 1022.090 389.660 1022.370 389.940 ;
        RECT 1021.470 389.040 1021.750 389.320 ;
        RECT 1022.090 389.040 1022.370 389.320 ;
        RECT 1096.470 399.760 1096.750 400.040 ;
        RECT 1097.090 399.760 1097.370 400.040 ;
        RECT 1096.470 399.140 1096.750 399.420 ;
        RECT 1097.090 399.140 1097.370 399.420 ;
        RECT 1096.470 398.520 1096.750 398.800 ;
        RECT 1097.090 398.520 1097.370 398.800 ;
        RECT 1096.470 397.900 1096.750 398.180 ;
        RECT 1097.090 397.900 1097.370 398.180 ;
        RECT 1096.470 397.280 1096.750 397.560 ;
        RECT 1097.090 397.280 1097.370 397.560 ;
        RECT 1096.470 396.660 1096.750 396.940 ;
        RECT 1097.090 396.660 1097.370 396.940 ;
        RECT 1096.470 396.040 1096.750 396.320 ;
        RECT 1097.090 396.040 1097.370 396.320 ;
        RECT 1071.470 392.760 1071.750 393.040 ;
        RECT 1072.090 392.760 1072.370 393.040 ;
        RECT 1071.470 392.140 1071.750 392.420 ;
        RECT 1072.090 392.140 1072.370 392.420 ;
        RECT 1071.470 391.520 1071.750 391.800 ;
        RECT 1072.090 391.520 1072.370 391.800 ;
        RECT 1071.470 390.900 1071.750 391.180 ;
        RECT 1072.090 390.900 1072.370 391.180 ;
        RECT 1071.470 390.280 1071.750 390.560 ;
        RECT 1072.090 390.280 1072.370 390.560 ;
        RECT 1071.470 389.660 1071.750 389.940 ;
        RECT 1072.090 389.660 1072.370 389.940 ;
        RECT 1071.470 389.040 1071.750 389.320 ;
        RECT 1072.090 389.040 1072.370 389.320 ;
        RECT 1146.470 399.760 1146.750 400.040 ;
        RECT 1147.090 399.760 1147.370 400.040 ;
        RECT 1146.470 399.140 1146.750 399.420 ;
        RECT 1147.090 399.140 1147.370 399.420 ;
        RECT 1146.470 398.520 1146.750 398.800 ;
        RECT 1147.090 398.520 1147.370 398.800 ;
        RECT 1146.470 397.900 1146.750 398.180 ;
        RECT 1147.090 397.900 1147.370 398.180 ;
        RECT 1146.470 397.280 1146.750 397.560 ;
        RECT 1147.090 397.280 1147.370 397.560 ;
        RECT 1146.470 396.660 1146.750 396.940 ;
        RECT 1147.090 396.660 1147.370 396.940 ;
        RECT 1146.470 396.040 1146.750 396.320 ;
        RECT 1147.090 396.040 1147.370 396.320 ;
        RECT 1121.470 392.760 1121.750 393.040 ;
        RECT 1122.090 392.760 1122.370 393.040 ;
        RECT 1121.470 392.140 1121.750 392.420 ;
        RECT 1122.090 392.140 1122.370 392.420 ;
        RECT 1121.470 391.520 1121.750 391.800 ;
        RECT 1122.090 391.520 1122.370 391.800 ;
        RECT 1121.470 390.900 1121.750 391.180 ;
        RECT 1122.090 390.900 1122.370 391.180 ;
        RECT 1121.470 390.280 1121.750 390.560 ;
        RECT 1122.090 390.280 1122.370 390.560 ;
        RECT 1121.470 389.660 1121.750 389.940 ;
        RECT 1122.090 389.660 1122.370 389.940 ;
        RECT 1121.470 389.040 1121.750 389.320 ;
        RECT 1122.090 389.040 1122.370 389.320 ;
        RECT 1196.470 399.760 1196.750 400.040 ;
        RECT 1197.090 399.760 1197.370 400.040 ;
        RECT 1196.470 399.140 1196.750 399.420 ;
        RECT 1197.090 399.140 1197.370 399.420 ;
        RECT 1196.470 398.520 1196.750 398.800 ;
        RECT 1197.090 398.520 1197.370 398.800 ;
        RECT 1196.470 397.900 1196.750 398.180 ;
        RECT 1197.090 397.900 1197.370 398.180 ;
        RECT 1196.470 397.280 1196.750 397.560 ;
        RECT 1197.090 397.280 1197.370 397.560 ;
        RECT 1196.470 396.660 1196.750 396.940 ;
        RECT 1197.090 396.660 1197.370 396.940 ;
        RECT 1196.470 396.040 1196.750 396.320 ;
        RECT 1197.090 396.040 1197.370 396.320 ;
        RECT 1171.470 392.760 1171.750 393.040 ;
        RECT 1172.090 392.760 1172.370 393.040 ;
        RECT 1171.470 392.140 1171.750 392.420 ;
        RECT 1172.090 392.140 1172.370 392.420 ;
        RECT 1171.470 391.520 1171.750 391.800 ;
        RECT 1172.090 391.520 1172.370 391.800 ;
        RECT 1171.470 390.900 1171.750 391.180 ;
        RECT 1172.090 390.900 1172.370 391.180 ;
        RECT 1171.470 390.280 1171.750 390.560 ;
        RECT 1172.090 390.280 1172.370 390.560 ;
        RECT 1171.470 389.660 1171.750 389.940 ;
        RECT 1172.090 389.660 1172.370 389.940 ;
        RECT 1171.470 389.040 1171.750 389.320 ;
        RECT 1172.090 389.040 1172.370 389.320 ;
        RECT 1246.470 399.760 1246.750 400.040 ;
        RECT 1247.090 399.760 1247.370 400.040 ;
        RECT 1246.470 399.140 1246.750 399.420 ;
        RECT 1247.090 399.140 1247.370 399.420 ;
        RECT 1246.470 398.520 1246.750 398.800 ;
        RECT 1247.090 398.520 1247.370 398.800 ;
        RECT 1246.470 397.900 1246.750 398.180 ;
        RECT 1247.090 397.900 1247.370 398.180 ;
        RECT 1246.470 397.280 1246.750 397.560 ;
        RECT 1247.090 397.280 1247.370 397.560 ;
        RECT 1246.470 396.660 1246.750 396.940 ;
        RECT 1247.090 396.660 1247.370 396.940 ;
        RECT 1246.470 396.040 1246.750 396.320 ;
        RECT 1247.090 396.040 1247.370 396.320 ;
        RECT 1221.470 392.760 1221.750 393.040 ;
        RECT 1222.090 392.760 1222.370 393.040 ;
        RECT 1221.470 392.140 1221.750 392.420 ;
        RECT 1222.090 392.140 1222.370 392.420 ;
        RECT 1221.470 391.520 1221.750 391.800 ;
        RECT 1222.090 391.520 1222.370 391.800 ;
        RECT 1221.470 390.900 1221.750 391.180 ;
        RECT 1222.090 390.900 1222.370 391.180 ;
        RECT 1221.470 390.280 1221.750 390.560 ;
        RECT 1222.090 390.280 1222.370 390.560 ;
        RECT 1221.470 389.660 1221.750 389.940 ;
        RECT 1222.090 389.660 1222.370 389.940 ;
        RECT 1221.470 389.040 1221.750 389.320 ;
        RECT 1222.090 389.040 1222.370 389.320 ;
        RECT 1296.470 399.760 1296.750 400.040 ;
        RECT 1297.090 399.760 1297.370 400.040 ;
        RECT 1296.470 399.140 1296.750 399.420 ;
        RECT 1297.090 399.140 1297.370 399.420 ;
        RECT 1296.470 398.520 1296.750 398.800 ;
        RECT 1297.090 398.520 1297.370 398.800 ;
        RECT 1296.470 397.900 1296.750 398.180 ;
        RECT 1297.090 397.900 1297.370 398.180 ;
        RECT 1296.470 397.280 1296.750 397.560 ;
        RECT 1297.090 397.280 1297.370 397.560 ;
        RECT 1296.470 396.660 1296.750 396.940 ;
        RECT 1297.090 396.660 1297.370 396.940 ;
        RECT 1296.470 396.040 1296.750 396.320 ;
        RECT 1297.090 396.040 1297.370 396.320 ;
        RECT 1271.470 392.760 1271.750 393.040 ;
        RECT 1272.090 392.760 1272.370 393.040 ;
        RECT 1271.470 392.140 1271.750 392.420 ;
        RECT 1272.090 392.140 1272.370 392.420 ;
        RECT 1271.470 391.520 1271.750 391.800 ;
        RECT 1272.090 391.520 1272.370 391.800 ;
        RECT 1271.470 390.900 1271.750 391.180 ;
        RECT 1272.090 390.900 1272.370 391.180 ;
        RECT 1271.470 390.280 1271.750 390.560 ;
        RECT 1272.090 390.280 1272.370 390.560 ;
        RECT 1271.470 389.660 1271.750 389.940 ;
        RECT 1272.090 389.660 1272.370 389.940 ;
        RECT 1271.470 389.040 1271.750 389.320 ;
        RECT 1272.090 389.040 1272.370 389.320 ;
        RECT 1346.470 399.760 1346.750 400.040 ;
        RECT 1347.090 399.760 1347.370 400.040 ;
        RECT 1346.470 399.140 1346.750 399.420 ;
        RECT 1347.090 399.140 1347.370 399.420 ;
        RECT 1346.470 398.520 1346.750 398.800 ;
        RECT 1347.090 398.520 1347.370 398.800 ;
        RECT 1346.470 397.900 1346.750 398.180 ;
        RECT 1347.090 397.900 1347.370 398.180 ;
        RECT 1346.470 397.280 1346.750 397.560 ;
        RECT 1347.090 397.280 1347.370 397.560 ;
        RECT 1346.470 396.660 1346.750 396.940 ;
        RECT 1347.090 396.660 1347.370 396.940 ;
        RECT 1346.470 396.040 1346.750 396.320 ;
        RECT 1347.090 396.040 1347.370 396.320 ;
        RECT 1361.650 399.760 1361.930 400.040 ;
        RECT 1362.270 399.760 1362.550 400.040 ;
        RECT 1362.890 399.760 1363.170 400.040 ;
        RECT 1363.510 399.760 1363.790 400.040 ;
        RECT 1364.130 399.760 1364.410 400.040 ;
        RECT 1364.750 399.760 1365.030 400.040 ;
        RECT 1365.370 399.760 1365.650 400.040 ;
        RECT 1365.990 399.760 1366.270 400.040 ;
        RECT 1366.610 399.760 1366.890 400.040 ;
        RECT 1367.230 399.760 1367.510 400.040 ;
        RECT 1367.850 399.760 1368.130 400.040 ;
        RECT 1368.470 399.760 1368.750 400.040 ;
        RECT 1369.090 399.760 1369.370 400.040 ;
        RECT 1369.710 399.760 1369.990 400.040 ;
        RECT 1370.330 399.760 1370.610 400.040 ;
        RECT 1361.650 399.140 1361.930 399.420 ;
        RECT 1362.270 399.140 1362.550 399.420 ;
        RECT 1362.890 399.140 1363.170 399.420 ;
        RECT 1363.510 399.140 1363.790 399.420 ;
        RECT 1364.130 399.140 1364.410 399.420 ;
        RECT 1364.750 399.140 1365.030 399.420 ;
        RECT 1365.370 399.140 1365.650 399.420 ;
        RECT 1365.990 399.140 1366.270 399.420 ;
        RECT 1366.610 399.140 1366.890 399.420 ;
        RECT 1367.230 399.140 1367.510 399.420 ;
        RECT 1367.850 399.140 1368.130 399.420 ;
        RECT 1368.470 399.140 1368.750 399.420 ;
        RECT 1369.090 399.140 1369.370 399.420 ;
        RECT 1369.710 399.140 1369.990 399.420 ;
        RECT 1370.330 399.140 1370.610 399.420 ;
        RECT 1361.650 398.520 1361.930 398.800 ;
        RECT 1362.270 398.520 1362.550 398.800 ;
        RECT 1362.890 398.520 1363.170 398.800 ;
        RECT 1363.510 398.520 1363.790 398.800 ;
        RECT 1364.130 398.520 1364.410 398.800 ;
        RECT 1364.750 398.520 1365.030 398.800 ;
        RECT 1365.370 398.520 1365.650 398.800 ;
        RECT 1365.990 398.520 1366.270 398.800 ;
        RECT 1366.610 398.520 1366.890 398.800 ;
        RECT 1367.230 398.520 1367.510 398.800 ;
        RECT 1367.850 398.520 1368.130 398.800 ;
        RECT 1368.470 398.520 1368.750 398.800 ;
        RECT 1369.090 398.520 1369.370 398.800 ;
        RECT 1369.710 398.520 1369.990 398.800 ;
        RECT 1370.330 398.520 1370.610 398.800 ;
        RECT 1361.650 397.900 1361.930 398.180 ;
        RECT 1362.270 397.900 1362.550 398.180 ;
        RECT 1362.890 397.900 1363.170 398.180 ;
        RECT 1363.510 397.900 1363.790 398.180 ;
        RECT 1364.130 397.900 1364.410 398.180 ;
        RECT 1364.750 397.900 1365.030 398.180 ;
        RECT 1365.370 397.900 1365.650 398.180 ;
        RECT 1365.990 397.900 1366.270 398.180 ;
        RECT 1366.610 397.900 1366.890 398.180 ;
        RECT 1367.230 397.900 1367.510 398.180 ;
        RECT 1367.850 397.900 1368.130 398.180 ;
        RECT 1368.470 397.900 1368.750 398.180 ;
        RECT 1369.090 397.900 1369.370 398.180 ;
        RECT 1369.710 397.900 1369.990 398.180 ;
        RECT 1370.330 397.900 1370.610 398.180 ;
        RECT 1361.650 397.280 1361.930 397.560 ;
        RECT 1362.270 397.280 1362.550 397.560 ;
        RECT 1362.890 397.280 1363.170 397.560 ;
        RECT 1363.510 397.280 1363.790 397.560 ;
        RECT 1364.130 397.280 1364.410 397.560 ;
        RECT 1364.750 397.280 1365.030 397.560 ;
        RECT 1365.370 397.280 1365.650 397.560 ;
        RECT 1365.990 397.280 1366.270 397.560 ;
        RECT 1366.610 397.280 1366.890 397.560 ;
        RECT 1367.230 397.280 1367.510 397.560 ;
        RECT 1367.850 397.280 1368.130 397.560 ;
        RECT 1368.470 397.280 1368.750 397.560 ;
        RECT 1369.090 397.280 1369.370 397.560 ;
        RECT 1369.710 397.280 1369.990 397.560 ;
        RECT 1370.330 397.280 1370.610 397.560 ;
        RECT 1361.650 396.660 1361.930 396.940 ;
        RECT 1362.270 396.660 1362.550 396.940 ;
        RECT 1362.890 396.660 1363.170 396.940 ;
        RECT 1363.510 396.660 1363.790 396.940 ;
        RECT 1364.130 396.660 1364.410 396.940 ;
        RECT 1364.750 396.660 1365.030 396.940 ;
        RECT 1365.370 396.660 1365.650 396.940 ;
        RECT 1365.990 396.660 1366.270 396.940 ;
        RECT 1366.610 396.660 1366.890 396.940 ;
        RECT 1367.230 396.660 1367.510 396.940 ;
        RECT 1367.850 396.660 1368.130 396.940 ;
        RECT 1368.470 396.660 1368.750 396.940 ;
        RECT 1369.090 396.660 1369.370 396.940 ;
        RECT 1369.710 396.660 1369.990 396.940 ;
        RECT 1370.330 396.660 1370.610 396.940 ;
        RECT 1361.650 396.040 1361.930 396.320 ;
        RECT 1362.270 396.040 1362.550 396.320 ;
        RECT 1362.890 396.040 1363.170 396.320 ;
        RECT 1363.510 396.040 1363.790 396.320 ;
        RECT 1364.130 396.040 1364.410 396.320 ;
        RECT 1364.750 396.040 1365.030 396.320 ;
        RECT 1365.370 396.040 1365.650 396.320 ;
        RECT 1365.990 396.040 1366.270 396.320 ;
        RECT 1366.610 396.040 1366.890 396.320 ;
        RECT 1367.230 396.040 1367.510 396.320 ;
        RECT 1367.850 396.040 1368.130 396.320 ;
        RECT 1368.470 396.040 1368.750 396.320 ;
        RECT 1369.090 396.040 1369.370 396.320 ;
        RECT 1369.710 396.040 1369.990 396.320 ;
        RECT 1370.330 396.040 1370.610 396.320 ;
        RECT 1321.470 392.760 1321.750 393.040 ;
        RECT 1322.090 392.760 1322.370 393.040 ;
        RECT 1321.470 392.140 1321.750 392.420 ;
        RECT 1322.090 392.140 1322.370 392.420 ;
        RECT 1321.470 391.520 1321.750 391.800 ;
        RECT 1322.090 391.520 1322.370 391.800 ;
        RECT 1321.470 390.900 1321.750 391.180 ;
        RECT 1322.090 390.900 1322.370 391.180 ;
        RECT 1321.470 390.280 1321.750 390.560 ;
        RECT 1322.090 390.280 1322.370 390.560 ;
        RECT 1321.470 389.660 1321.750 389.940 ;
        RECT 1322.090 389.660 1322.370 389.940 ;
        RECT 1321.470 389.040 1321.750 389.320 ;
        RECT 1322.090 389.040 1322.370 389.320 ;
        RECT 1374.050 399.760 1374.330 400.040 ;
        RECT 1374.670 399.760 1374.950 400.040 ;
        RECT 1375.290 399.760 1375.570 400.040 ;
        RECT 1375.910 399.760 1376.190 400.040 ;
        RECT 1376.530 399.760 1376.810 400.040 ;
        RECT 1377.150 399.760 1377.430 400.040 ;
        RECT 1377.770 399.760 1378.050 400.040 ;
        RECT 1378.390 399.760 1378.670 400.040 ;
        RECT 1379.010 399.760 1379.290 400.040 ;
        RECT 1379.630 399.760 1379.910 400.040 ;
        RECT 1380.250 399.760 1380.530 400.040 ;
        RECT 1380.870 399.760 1381.150 400.040 ;
        RECT 1381.490 399.760 1381.770 400.040 ;
        RECT 1382.110 399.760 1382.390 400.040 ;
        RECT 1382.730 399.760 1383.010 400.040 ;
        RECT 1383.350 399.760 1383.630 400.040 ;
        RECT 1374.050 399.140 1374.330 399.420 ;
        RECT 1374.670 399.140 1374.950 399.420 ;
        RECT 1375.290 399.140 1375.570 399.420 ;
        RECT 1375.910 399.140 1376.190 399.420 ;
        RECT 1376.530 399.140 1376.810 399.420 ;
        RECT 1377.150 399.140 1377.430 399.420 ;
        RECT 1377.770 399.140 1378.050 399.420 ;
        RECT 1378.390 399.140 1378.670 399.420 ;
        RECT 1379.010 399.140 1379.290 399.420 ;
        RECT 1379.630 399.140 1379.910 399.420 ;
        RECT 1380.250 399.140 1380.530 399.420 ;
        RECT 1380.870 399.140 1381.150 399.420 ;
        RECT 1381.490 399.140 1381.770 399.420 ;
        RECT 1382.110 399.140 1382.390 399.420 ;
        RECT 1382.730 399.140 1383.010 399.420 ;
        RECT 1383.350 399.140 1383.630 399.420 ;
        RECT 1374.050 398.520 1374.330 398.800 ;
        RECT 1374.670 398.520 1374.950 398.800 ;
        RECT 1375.290 398.520 1375.570 398.800 ;
        RECT 1375.910 398.520 1376.190 398.800 ;
        RECT 1376.530 398.520 1376.810 398.800 ;
        RECT 1377.150 398.520 1377.430 398.800 ;
        RECT 1377.770 398.520 1378.050 398.800 ;
        RECT 1378.390 398.520 1378.670 398.800 ;
        RECT 1379.010 398.520 1379.290 398.800 ;
        RECT 1379.630 398.520 1379.910 398.800 ;
        RECT 1380.250 398.520 1380.530 398.800 ;
        RECT 1380.870 398.520 1381.150 398.800 ;
        RECT 1381.490 398.520 1381.770 398.800 ;
        RECT 1382.110 398.520 1382.390 398.800 ;
        RECT 1382.730 398.520 1383.010 398.800 ;
        RECT 1383.350 398.520 1383.630 398.800 ;
        RECT 1374.050 397.900 1374.330 398.180 ;
        RECT 1374.670 397.900 1374.950 398.180 ;
        RECT 1375.290 397.900 1375.570 398.180 ;
        RECT 1375.910 397.900 1376.190 398.180 ;
        RECT 1376.530 397.900 1376.810 398.180 ;
        RECT 1377.150 397.900 1377.430 398.180 ;
        RECT 1377.770 397.900 1378.050 398.180 ;
        RECT 1378.390 397.900 1378.670 398.180 ;
        RECT 1379.010 397.900 1379.290 398.180 ;
        RECT 1379.630 397.900 1379.910 398.180 ;
        RECT 1380.250 397.900 1380.530 398.180 ;
        RECT 1380.870 397.900 1381.150 398.180 ;
        RECT 1381.490 397.900 1381.770 398.180 ;
        RECT 1382.110 397.900 1382.390 398.180 ;
        RECT 1382.730 397.900 1383.010 398.180 ;
        RECT 1383.350 397.900 1383.630 398.180 ;
        RECT 1374.050 397.280 1374.330 397.560 ;
        RECT 1374.670 397.280 1374.950 397.560 ;
        RECT 1375.290 397.280 1375.570 397.560 ;
        RECT 1375.910 397.280 1376.190 397.560 ;
        RECT 1376.530 397.280 1376.810 397.560 ;
        RECT 1377.150 397.280 1377.430 397.560 ;
        RECT 1377.770 397.280 1378.050 397.560 ;
        RECT 1378.390 397.280 1378.670 397.560 ;
        RECT 1379.010 397.280 1379.290 397.560 ;
        RECT 1379.630 397.280 1379.910 397.560 ;
        RECT 1380.250 397.280 1380.530 397.560 ;
        RECT 1380.870 397.280 1381.150 397.560 ;
        RECT 1381.490 397.280 1381.770 397.560 ;
        RECT 1382.110 397.280 1382.390 397.560 ;
        RECT 1382.730 397.280 1383.010 397.560 ;
        RECT 1383.350 397.280 1383.630 397.560 ;
        RECT 1374.050 396.660 1374.330 396.940 ;
        RECT 1374.670 396.660 1374.950 396.940 ;
        RECT 1375.290 396.660 1375.570 396.940 ;
        RECT 1375.910 396.660 1376.190 396.940 ;
        RECT 1376.530 396.660 1376.810 396.940 ;
        RECT 1377.150 396.660 1377.430 396.940 ;
        RECT 1377.770 396.660 1378.050 396.940 ;
        RECT 1378.390 396.660 1378.670 396.940 ;
        RECT 1379.010 396.660 1379.290 396.940 ;
        RECT 1379.630 396.660 1379.910 396.940 ;
        RECT 1380.250 396.660 1380.530 396.940 ;
        RECT 1380.870 396.660 1381.150 396.940 ;
        RECT 1381.490 396.660 1381.770 396.940 ;
        RECT 1382.110 396.660 1382.390 396.940 ;
        RECT 1382.730 396.660 1383.010 396.940 ;
        RECT 1383.350 396.660 1383.630 396.940 ;
        RECT 1374.050 396.040 1374.330 396.320 ;
        RECT 1374.670 396.040 1374.950 396.320 ;
        RECT 1375.290 396.040 1375.570 396.320 ;
        RECT 1375.910 396.040 1376.190 396.320 ;
        RECT 1376.530 396.040 1376.810 396.320 ;
        RECT 1377.150 396.040 1377.430 396.320 ;
        RECT 1377.770 396.040 1378.050 396.320 ;
        RECT 1378.390 396.040 1378.670 396.320 ;
        RECT 1379.010 396.040 1379.290 396.320 ;
        RECT 1379.630 396.040 1379.910 396.320 ;
        RECT 1380.250 396.040 1380.530 396.320 ;
        RECT 1380.870 396.040 1381.150 396.320 ;
        RECT 1381.490 396.040 1381.770 396.320 ;
        RECT 1382.110 396.040 1382.390 396.320 ;
        RECT 1382.730 396.040 1383.010 396.320 ;
        RECT 1383.350 396.040 1383.630 396.320 ;
        RECT 1385.900 399.760 1386.180 400.040 ;
        RECT 1386.520 399.760 1386.800 400.040 ;
        RECT 1387.140 399.760 1387.420 400.040 ;
        RECT 1387.760 399.760 1388.040 400.040 ;
        RECT 1388.380 399.760 1388.660 400.040 ;
        RECT 1389.000 399.760 1389.280 400.040 ;
        RECT 1389.620 399.760 1389.900 400.040 ;
        RECT 1390.240 399.760 1390.520 400.040 ;
        RECT 1390.860 399.760 1391.140 400.040 ;
        RECT 1391.480 399.760 1391.760 400.040 ;
        RECT 1392.100 399.760 1392.380 400.040 ;
        RECT 1392.720 399.760 1393.000 400.040 ;
        RECT 1393.340 399.760 1393.620 400.040 ;
        RECT 1393.960 399.760 1394.240 400.040 ;
        RECT 1394.580 399.760 1394.860 400.040 ;
        RECT 1395.200 399.760 1395.480 400.040 ;
        RECT 1385.900 399.140 1386.180 399.420 ;
        RECT 1386.520 399.140 1386.800 399.420 ;
        RECT 1387.140 399.140 1387.420 399.420 ;
        RECT 1387.760 399.140 1388.040 399.420 ;
        RECT 1388.380 399.140 1388.660 399.420 ;
        RECT 1389.000 399.140 1389.280 399.420 ;
        RECT 1389.620 399.140 1389.900 399.420 ;
        RECT 1390.240 399.140 1390.520 399.420 ;
        RECT 1390.860 399.140 1391.140 399.420 ;
        RECT 1391.480 399.140 1391.760 399.420 ;
        RECT 1392.100 399.140 1392.380 399.420 ;
        RECT 1392.720 399.140 1393.000 399.420 ;
        RECT 1393.340 399.140 1393.620 399.420 ;
        RECT 1393.960 399.140 1394.240 399.420 ;
        RECT 1394.580 399.140 1394.860 399.420 ;
        RECT 1395.200 399.140 1395.480 399.420 ;
        RECT 1385.900 398.520 1386.180 398.800 ;
        RECT 1386.520 398.520 1386.800 398.800 ;
        RECT 1387.140 398.520 1387.420 398.800 ;
        RECT 1387.760 398.520 1388.040 398.800 ;
        RECT 1388.380 398.520 1388.660 398.800 ;
        RECT 1389.000 398.520 1389.280 398.800 ;
        RECT 1389.620 398.520 1389.900 398.800 ;
        RECT 1390.240 398.520 1390.520 398.800 ;
        RECT 1390.860 398.520 1391.140 398.800 ;
        RECT 1391.480 398.520 1391.760 398.800 ;
        RECT 1392.100 398.520 1392.380 398.800 ;
        RECT 1392.720 398.520 1393.000 398.800 ;
        RECT 1393.340 398.520 1393.620 398.800 ;
        RECT 1393.960 398.520 1394.240 398.800 ;
        RECT 1394.580 398.520 1394.860 398.800 ;
        RECT 1395.200 398.520 1395.480 398.800 ;
        RECT 1385.900 397.900 1386.180 398.180 ;
        RECT 1386.520 397.900 1386.800 398.180 ;
        RECT 1387.140 397.900 1387.420 398.180 ;
        RECT 1387.760 397.900 1388.040 398.180 ;
        RECT 1388.380 397.900 1388.660 398.180 ;
        RECT 1389.000 397.900 1389.280 398.180 ;
        RECT 1389.620 397.900 1389.900 398.180 ;
        RECT 1390.240 397.900 1390.520 398.180 ;
        RECT 1390.860 397.900 1391.140 398.180 ;
        RECT 1391.480 397.900 1391.760 398.180 ;
        RECT 1392.100 397.900 1392.380 398.180 ;
        RECT 1392.720 397.900 1393.000 398.180 ;
        RECT 1393.340 397.900 1393.620 398.180 ;
        RECT 1393.960 397.900 1394.240 398.180 ;
        RECT 1394.580 397.900 1394.860 398.180 ;
        RECT 1395.200 397.900 1395.480 398.180 ;
        RECT 1385.900 397.280 1386.180 397.560 ;
        RECT 1386.520 397.280 1386.800 397.560 ;
        RECT 1387.140 397.280 1387.420 397.560 ;
        RECT 1387.760 397.280 1388.040 397.560 ;
        RECT 1388.380 397.280 1388.660 397.560 ;
        RECT 1389.000 397.280 1389.280 397.560 ;
        RECT 1389.620 397.280 1389.900 397.560 ;
        RECT 1390.240 397.280 1390.520 397.560 ;
        RECT 1390.860 397.280 1391.140 397.560 ;
        RECT 1391.480 397.280 1391.760 397.560 ;
        RECT 1392.100 397.280 1392.380 397.560 ;
        RECT 1392.720 397.280 1393.000 397.560 ;
        RECT 1393.340 397.280 1393.620 397.560 ;
        RECT 1393.960 397.280 1394.240 397.560 ;
        RECT 1394.580 397.280 1394.860 397.560 ;
        RECT 1395.200 397.280 1395.480 397.560 ;
        RECT 1385.900 396.660 1386.180 396.940 ;
        RECT 1386.520 396.660 1386.800 396.940 ;
        RECT 1387.140 396.660 1387.420 396.940 ;
        RECT 1387.760 396.660 1388.040 396.940 ;
        RECT 1388.380 396.660 1388.660 396.940 ;
        RECT 1389.000 396.660 1389.280 396.940 ;
        RECT 1389.620 396.660 1389.900 396.940 ;
        RECT 1390.240 396.660 1390.520 396.940 ;
        RECT 1390.860 396.660 1391.140 396.940 ;
        RECT 1391.480 396.660 1391.760 396.940 ;
        RECT 1392.100 396.660 1392.380 396.940 ;
        RECT 1392.720 396.660 1393.000 396.940 ;
        RECT 1393.340 396.660 1393.620 396.940 ;
        RECT 1393.960 396.660 1394.240 396.940 ;
        RECT 1394.580 396.660 1394.860 396.940 ;
        RECT 1395.200 396.660 1395.480 396.940 ;
        RECT 1385.900 396.040 1386.180 396.320 ;
        RECT 1386.520 396.040 1386.800 396.320 ;
        RECT 1387.140 396.040 1387.420 396.320 ;
        RECT 1387.760 396.040 1388.040 396.320 ;
        RECT 1388.380 396.040 1388.660 396.320 ;
        RECT 1389.000 396.040 1389.280 396.320 ;
        RECT 1389.620 396.040 1389.900 396.320 ;
        RECT 1390.240 396.040 1390.520 396.320 ;
        RECT 1390.860 396.040 1391.140 396.320 ;
        RECT 1391.480 396.040 1391.760 396.320 ;
        RECT 1392.100 396.040 1392.380 396.320 ;
        RECT 1392.720 396.040 1393.000 396.320 ;
        RECT 1393.340 396.040 1393.620 396.320 ;
        RECT 1393.960 396.040 1394.240 396.320 ;
        RECT 1394.580 396.040 1394.860 396.320 ;
        RECT 1395.200 396.040 1395.480 396.320 ;
        RECT 1399.430 399.760 1399.710 400.040 ;
        RECT 1400.050 399.760 1400.330 400.040 ;
        RECT 1400.670 399.760 1400.950 400.040 ;
        RECT 1401.290 399.760 1401.570 400.040 ;
        RECT 1401.910 399.760 1402.190 400.040 ;
        RECT 1402.530 399.760 1402.810 400.040 ;
        RECT 1403.150 399.760 1403.430 400.040 ;
        RECT 1403.770 399.760 1404.050 400.040 ;
        RECT 1404.390 399.760 1404.670 400.040 ;
        RECT 1405.010 399.760 1405.290 400.040 ;
        RECT 1405.630 399.760 1405.910 400.040 ;
        RECT 1406.250 399.760 1406.530 400.040 ;
        RECT 1406.870 399.760 1407.150 400.040 ;
        RECT 1407.490 399.760 1407.770 400.040 ;
        RECT 1408.110 399.760 1408.390 400.040 ;
        RECT 1408.730 399.760 1409.010 400.040 ;
        RECT 1399.430 399.140 1399.710 399.420 ;
        RECT 1400.050 399.140 1400.330 399.420 ;
        RECT 1400.670 399.140 1400.950 399.420 ;
        RECT 1401.290 399.140 1401.570 399.420 ;
        RECT 1401.910 399.140 1402.190 399.420 ;
        RECT 1402.530 399.140 1402.810 399.420 ;
        RECT 1403.150 399.140 1403.430 399.420 ;
        RECT 1403.770 399.140 1404.050 399.420 ;
        RECT 1404.390 399.140 1404.670 399.420 ;
        RECT 1405.010 399.140 1405.290 399.420 ;
        RECT 1405.630 399.140 1405.910 399.420 ;
        RECT 1406.250 399.140 1406.530 399.420 ;
        RECT 1406.870 399.140 1407.150 399.420 ;
        RECT 1407.490 399.140 1407.770 399.420 ;
        RECT 1408.110 399.140 1408.390 399.420 ;
        RECT 1408.730 399.140 1409.010 399.420 ;
        RECT 1399.430 398.520 1399.710 398.800 ;
        RECT 1400.050 398.520 1400.330 398.800 ;
        RECT 1400.670 398.520 1400.950 398.800 ;
        RECT 1401.290 398.520 1401.570 398.800 ;
        RECT 1401.910 398.520 1402.190 398.800 ;
        RECT 1402.530 398.520 1402.810 398.800 ;
        RECT 1403.150 398.520 1403.430 398.800 ;
        RECT 1403.770 398.520 1404.050 398.800 ;
        RECT 1404.390 398.520 1404.670 398.800 ;
        RECT 1405.010 398.520 1405.290 398.800 ;
        RECT 1405.630 398.520 1405.910 398.800 ;
        RECT 1406.250 398.520 1406.530 398.800 ;
        RECT 1406.870 398.520 1407.150 398.800 ;
        RECT 1407.490 398.520 1407.770 398.800 ;
        RECT 1408.110 398.520 1408.390 398.800 ;
        RECT 1408.730 398.520 1409.010 398.800 ;
        RECT 1399.430 397.900 1399.710 398.180 ;
        RECT 1400.050 397.900 1400.330 398.180 ;
        RECT 1400.670 397.900 1400.950 398.180 ;
        RECT 1401.290 397.900 1401.570 398.180 ;
        RECT 1401.910 397.900 1402.190 398.180 ;
        RECT 1402.530 397.900 1402.810 398.180 ;
        RECT 1403.150 397.900 1403.430 398.180 ;
        RECT 1403.770 397.900 1404.050 398.180 ;
        RECT 1404.390 397.900 1404.670 398.180 ;
        RECT 1405.010 397.900 1405.290 398.180 ;
        RECT 1405.630 397.900 1405.910 398.180 ;
        RECT 1406.250 397.900 1406.530 398.180 ;
        RECT 1406.870 397.900 1407.150 398.180 ;
        RECT 1407.490 397.900 1407.770 398.180 ;
        RECT 1408.110 397.900 1408.390 398.180 ;
        RECT 1408.730 397.900 1409.010 398.180 ;
        RECT 1399.430 397.280 1399.710 397.560 ;
        RECT 1400.050 397.280 1400.330 397.560 ;
        RECT 1400.670 397.280 1400.950 397.560 ;
        RECT 1401.290 397.280 1401.570 397.560 ;
        RECT 1401.910 397.280 1402.190 397.560 ;
        RECT 1402.530 397.280 1402.810 397.560 ;
        RECT 1403.150 397.280 1403.430 397.560 ;
        RECT 1403.770 397.280 1404.050 397.560 ;
        RECT 1404.390 397.280 1404.670 397.560 ;
        RECT 1405.010 397.280 1405.290 397.560 ;
        RECT 1405.630 397.280 1405.910 397.560 ;
        RECT 1406.250 397.280 1406.530 397.560 ;
        RECT 1406.870 397.280 1407.150 397.560 ;
        RECT 1407.490 397.280 1407.770 397.560 ;
        RECT 1408.110 397.280 1408.390 397.560 ;
        RECT 1408.730 397.280 1409.010 397.560 ;
        RECT 1399.430 396.660 1399.710 396.940 ;
        RECT 1400.050 396.660 1400.330 396.940 ;
        RECT 1400.670 396.660 1400.950 396.940 ;
        RECT 1401.290 396.660 1401.570 396.940 ;
        RECT 1401.910 396.660 1402.190 396.940 ;
        RECT 1402.530 396.660 1402.810 396.940 ;
        RECT 1403.150 396.660 1403.430 396.940 ;
        RECT 1403.770 396.660 1404.050 396.940 ;
        RECT 1404.390 396.660 1404.670 396.940 ;
        RECT 1405.010 396.660 1405.290 396.940 ;
        RECT 1405.630 396.660 1405.910 396.940 ;
        RECT 1406.250 396.660 1406.530 396.940 ;
        RECT 1406.870 396.660 1407.150 396.940 ;
        RECT 1407.490 396.660 1407.770 396.940 ;
        RECT 1408.110 396.660 1408.390 396.940 ;
        RECT 1408.730 396.660 1409.010 396.940 ;
        RECT 1399.430 396.040 1399.710 396.320 ;
        RECT 1400.050 396.040 1400.330 396.320 ;
        RECT 1400.670 396.040 1400.950 396.320 ;
        RECT 1401.290 396.040 1401.570 396.320 ;
        RECT 1401.910 396.040 1402.190 396.320 ;
        RECT 1402.530 396.040 1402.810 396.320 ;
        RECT 1403.150 396.040 1403.430 396.320 ;
        RECT 1403.770 396.040 1404.050 396.320 ;
        RECT 1404.390 396.040 1404.670 396.320 ;
        RECT 1405.010 396.040 1405.290 396.320 ;
        RECT 1405.630 396.040 1405.910 396.320 ;
        RECT 1406.250 396.040 1406.530 396.320 ;
        RECT 1406.870 396.040 1407.150 396.320 ;
        RECT 1407.490 396.040 1407.770 396.320 ;
        RECT 1408.110 396.040 1408.390 396.320 ;
        RECT 1408.730 396.040 1409.010 396.320 ;
        RECT 1411.280 399.760 1411.560 400.040 ;
        RECT 1411.900 399.760 1412.180 400.040 ;
        RECT 1412.520 399.760 1412.800 400.040 ;
        RECT 1413.140 399.760 1413.420 400.040 ;
        RECT 1413.760 399.760 1414.040 400.040 ;
        RECT 1414.380 399.760 1414.660 400.040 ;
        RECT 1415.000 399.760 1415.280 400.040 ;
        RECT 1415.620 399.760 1415.900 400.040 ;
        RECT 1416.240 399.760 1416.520 400.040 ;
        RECT 1416.860 399.760 1417.140 400.040 ;
        RECT 1417.480 399.760 1417.760 400.040 ;
        RECT 1418.100 399.760 1418.380 400.040 ;
        RECT 1418.720 399.760 1419.000 400.040 ;
        RECT 1419.340 399.760 1419.620 400.040 ;
        RECT 1419.960 399.760 1420.240 400.040 ;
        RECT 1420.580 399.760 1420.860 400.040 ;
        RECT 1411.280 399.140 1411.560 399.420 ;
        RECT 1411.900 399.140 1412.180 399.420 ;
        RECT 1412.520 399.140 1412.800 399.420 ;
        RECT 1413.140 399.140 1413.420 399.420 ;
        RECT 1413.760 399.140 1414.040 399.420 ;
        RECT 1414.380 399.140 1414.660 399.420 ;
        RECT 1415.000 399.140 1415.280 399.420 ;
        RECT 1415.620 399.140 1415.900 399.420 ;
        RECT 1416.240 399.140 1416.520 399.420 ;
        RECT 1416.860 399.140 1417.140 399.420 ;
        RECT 1417.480 399.140 1417.760 399.420 ;
        RECT 1418.100 399.140 1418.380 399.420 ;
        RECT 1418.720 399.140 1419.000 399.420 ;
        RECT 1419.340 399.140 1419.620 399.420 ;
        RECT 1419.960 399.140 1420.240 399.420 ;
        RECT 1420.580 399.140 1420.860 399.420 ;
        RECT 1411.280 398.520 1411.560 398.800 ;
        RECT 1411.900 398.520 1412.180 398.800 ;
        RECT 1412.520 398.520 1412.800 398.800 ;
        RECT 1413.140 398.520 1413.420 398.800 ;
        RECT 1413.760 398.520 1414.040 398.800 ;
        RECT 1414.380 398.520 1414.660 398.800 ;
        RECT 1415.000 398.520 1415.280 398.800 ;
        RECT 1415.620 398.520 1415.900 398.800 ;
        RECT 1416.240 398.520 1416.520 398.800 ;
        RECT 1416.860 398.520 1417.140 398.800 ;
        RECT 1417.480 398.520 1417.760 398.800 ;
        RECT 1418.100 398.520 1418.380 398.800 ;
        RECT 1418.720 398.520 1419.000 398.800 ;
        RECT 1419.340 398.520 1419.620 398.800 ;
        RECT 1419.960 398.520 1420.240 398.800 ;
        RECT 1420.580 398.520 1420.860 398.800 ;
        RECT 1411.280 397.900 1411.560 398.180 ;
        RECT 1411.900 397.900 1412.180 398.180 ;
        RECT 1412.520 397.900 1412.800 398.180 ;
        RECT 1413.140 397.900 1413.420 398.180 ;
        RECT 1413.760 397.900 1414.040 398.180 ;
        RECT 1414.380 397.900 1414.660 398.180 ;
        RECT 1415.000 397.900 1415.280 398.180 ;
        RECT 1415.620 397.900 1415.900 398.180 ;
        RECT 1416.240 397.900 1416.520 398.180 ;
        RECT 1416.860 397.900 1417.140 398.180 ;
        RECT 1417.480 397.900 1417.760 398.180 ;
        RECT 1418.100 397.900 1418.380 398.180 ;
        RECT 1418.720 397.900 1419.000 398.180 ;
        RECT 1419.340 397.900 1419.620 398.180 ;
        RECT 1419.960 397.900 1420.240 398.180 ;
        RECT 1420.580 397.900 1420.860 398.180 ;
        RECT 1411.280 397.280 1411.560 397.560 ;
        RECT 1411.900 397.280 1412.180 397.560 ;
        RECT 1412.520 397.280 1412.800 397.560 ;
        RECT 1413.140 397.280 1413.420 397.560 ;
        RECT 1413.760 397.280 1414.040 397.560 ;
        RECT 1414.380 397.280 1414.660 397.560 ;
        RECT 1415.000 397.280 1415.280 397.560 ;
        RECT 1415.620 397.280 1415.900 397.560 ;
        RECT 1416.240 397.280 1416.520 397.560 ;
        RECT 1416.860 397.280 1417.140 397.560 ;
        RECT 1417.480 397.280 1417.760 397.560 ;
        RECT 1418.100 397.280 1418.380 397.560 ;
        RECT 1418.720 397.280 1419.000 397.560 ;
        RECT 1419.340 397.280 1419.620 397.560 ;
        RECT 1419.960 397.280 1420.240 397.560 ;
        RECT 1420.580 397.280 1420.860 397.560 ;
        RECT 1411.280 396.660 1411.560 396.940 ;
        RECT 1411.900 396.660 1412.180 396.940 ;
        RECT 1412.520 396.660 1412.800 396.940 ;
        RECT 1413.140 396.660 1413.420 396.940 ;
        RECT 1413.760 396.660 1414.040 396.940 ;
        RECT 1414.380 396.660 1414.660 396.940 ;
        RECT 1415.000 396.660 1415.280 396.940 ;
        RECT 1415.620 396.660 1415.900 396.940 ;
        RECT 1416.240 396.660 1416.520 396.940 ;
        RECT 1416.860 396.660 1417.140 396.940 ;
        RECT 1417.480 396.660 1417.760 396.940 ;
        RECT 1418.100 396.660 1418.380 396.940 ;
        RECT 1418.720 396.660 1419.000 396.940 ;
        RECT 1419.340 396.660 1419.620 396.940 ;
        RECT 1419.960 396.660 1420.240 396.940 ;
        RECT 1420.580 396.660 1420.860 396.940 ;
        RECT 1411.280 396.040 1411.560 396.320 ;
        RECT 1411.900 396.040 1412.180 396.320 ;
        RECT 1412.520 396.040 1412.800 396.320 ;
        RECT 1413.140 396.040 1413.420 396.320 ;
        RECT 1413.760 396.040 1414.040 396.320 ;
        RECT 1414.380 396.040 1414.660 396.320 ;
        RECT 1415.000 396.040 1415.280 396.320 ;
        RECT 1415.620 396.040 1415.900 396.320 ;
        RECT 1416.240 396.040 1416.520 396.320 ;
        RECT 1416.860 396.040 1417.140 396.320 ;
        RECT 1417.480 396.040 1417.760 396.320 ;
        RECT 1418.100 396.040 1418.380 396.320 ;
        RECT 1418.720 396.040 1419.000 396.320 ;
        RECT 1419.340 396.040 1419.620 396.320 ;
        RECT 1419.960 396.040 1420.240 396.320 ;
        RECT 1420.580 396.040 1420.860 396.320 ;
        RECT 1424.300 399.760 1424.580 400.040 ;
        RECT 1424.920 399.760 1425.200 400.040 ;
        RECT 1425.540 399.760 1425.820 400.040 ;
        RECT 1426.160 399.760 1426.440 400.040 ;
        RECT 1426.780 399.760 1427.060 400.040 ;
        RECT 1427.400 399.760 1427.680 400.040 ;
        RECT 1428.020 399.760 1428.300 400.040 ;
        RECT 1428.640 399.760 1428.920 400.040 ;
        RECT 1429.260 399.760 1429.540 400.040 ;
        RECT 1429.880 399.760 1430.160 400.040 ;
        RECT 1430.500 399.760 1430.780 400.040 ;
        RECT 1431.120 399.760 1431.400 400.040 ;
        RECT 1431.740 399.760 1432.020 400.040 ;
        RECT 1432.360 399.760 1432.640 400.040 ;
        RECT 1432.980 399.760 1433.260 400.040 ;
        RECT 1424.300 399.140 1424.580 399.420 ;
        RECT 1424.920 399.140 1425.200 399.420 ;
        RECT 1425.540 399.140 1425.820 399.420 ;
        RECT 1426.160 399.140 1426.440 399.420 ;
        RECT 1426.780 399.140 1427.060 399.420 ;
        RECT 1427.400 399.140 1427.680 399.420 ;
        RECT 1428.020 399.140 1428.300 399.420 ;
        RECT 1428.640 399.140 1428.920 399.420 ;
        RECT 1429.260 399.140 1429.540 399.420 ;
        RECT 1429.880 399.140 1430.160 399.420 ;
        RECT 1430.500 399.140 1430.780 399.420 ;
        RECT 1431.120 399.140 1431.400 399.420 ;
        RECT 1431.740 399.140 1432.020 399.420 ;
        RECT 1432.360 399.140 1432.640 399.420 ;
        RECT 1432.980 399.140 1433.260 399.420 ;
        RECT 1424.300 398.520 1424.580 398.800 ;
        RECT 1424.920 398.520 1425.200 398.800 ;
        RECT 1425.540 398.520 1425.820 398.800 ;
        RECT 1426.160 398.520 1426.440 398.800 ;
        RECT 1426.780 398.520 1427.060 398.800 ;
        RECT 1427.400 398.520 1427.680 398.800 ;
        RECT 1428.020 398.520 1428.300 398.800 ;
        RECT 1428.640 398.520 1428.920 398.800 ;
        RECT 1429.260 398.520 1429.540 398.800 ;
        RECT 1429.880 398.520 1430.160 398.800 ;
        RECT 1430.500 398.520 1430.780 398.800 ;
        RECT 1431.120 398.520 1431.400 398.800 ;
        RECT 1431.740 398.520 1432.020 398.800 ;
        RECT 1432.360 398.520 1432.640 398.800 ;
        RECT 1432.980 398.520 1433.260 398.800 ;
        RECT 1424.300 397.900 1424.580 398.180 ;
        RECT 1424.920 397.900 1425.200 398.180 ;
        RECT 1425.540 397.900 1425.820 398.180 ;
        RECT 1426.160 397.900 1426.440 398.180 ;
        RECT 1426.780 397.900 1427.060 398.180 ;
        RECT 1427.400 397.900 1427.680 398.180 ;
        RECT 1428.020 397.900 1428.300 398.180 ;
        RECT 1428.640 397.900 1428.920 398.180 ;
        RECT 1429.260 397.900 1429.540 398.180 ;
        RECT 1429.880 397.900 1430.160 398.180 ;
        RECT 1430.500 397.900 1430.780 398.180 ;
        RECT 1431.120 397.900 1431.400 398.180 ;
        RECT 1431.740 397.900 1432.020 398.180 ;
        RECT 1432.360 397.900 1432.640 398.180 ;
        RECT 1432.980 397.900 1433.260 398.180 ;
        RECT 1424.300 397.280 1424.580 397.560 ;
        RECT 1424.920 397.280 1425.200 397.560 ;
        RECT 1425.540 397.280 1425.820 397.560 ;
        RECT 1426.160 397.280 1426.440 397.560 ;
        RECT 1426.780 397.280 1427.060 397.560 ;
        RECT 1427.400 397.280 1427.680 397.560 ;
        RECT 1428.020 397.280 1428.300 397.560 ;
        RECT 1428.640 397.280 1428.920 397.560 ;
        RECT 1429.260 397.280 1429.540 397.560 ;
        RECT 1429.880 397.280 1430.160 397.560 ;
        RECT 1430.500 397.280 1430.780 397.560 ;
        RECT 1431.120 397.280 1431.400 397.560 ;
        RECT 1431.740 397.280 1432.020 397.560 ;
        RECT 1432.360 397.280 1432.640 397.560 ;
        RECT 1432.980 397.280 1433.260 397.560 ;
        RECT 1424.300 396.660 1424.580 396.940 ;
        RECT 1424.920 396.660 1425.200 396.940 ;
        RECT 1425.540 396.660 1425.820 396.940 ;
        RECT 1426.160 396.660 1426.440 396.940 ;
        RECT 1426.780 396.660 1427.060 396.940 ;
        RECT 1427.400 396.660 1427.680 396.940 ;
        RECT 1428.020 396.660 1428.300 396.940 ;
        RECT 1428.640 396.660 1428.920 396.940 ;
        RECT 1429.260 396.660 1429.540 396.940 ;
        RECT 1429.880 396.660 1430.160 396.940 ;
        RECT 1430.500 396.660 1430.780 396.940 ;
        RECT 1431.120 396.660 1431.400 396.940 ;
        RECT 1431.740 396.660 1432.020 396.940 ;
        RECT 1432.360 396.660 1432.640 396.940 ;
        RECT 1432.980 396.660 1433.260 396.940 ;
        RECT 1424.300 396.040 1424.580 396.320 ;
        RECT 1424.920 396.040 1425.200 396.320 ;
        RECT 1425.540 396.040 1425.820 396.320 ;
        RECT 1426.160 396.040 1426.440 396.320 ;
        RECT 1426.780 396.040 1427.060 396.320 ;
        RECT 1427.400 396.040 1427.680 396.320 ;
        RECT 1428.020 396.040 1428.300 396.320 ;
        RECT 1428.640 396.040 1428.920 396.320 ;
        RECT 1429.260 396.040 1429.540 396.320 ;
        RECT 1429.880 396.040 1430.160 396.320 ;
        RECT 1430.500 396.040 1430.780 396.320 ;
        RECT 1431.120 396.040 1431.400 396.320 ;
        RECT 1431.740 396.040 1432.020 396.320 ;
        RECT 1432.360 396.040 1432.640 396.320 ;
        RECT 1432.980 396.040 1433.260 396.320 ;
        RECT 1446.470 399.760 1446.750 400.040 ;
        RECT 1447.090 399.760 1447.370 400.040 ;
        RECT 1446.470 399.140 1446.750 399.420 ;
        RECT 1447.090 399.140 1447.370 399.420 ;
        RECT 1446.470 398.520 1446.750 398.800 ;
        RECT 1447.090 398.520 1447.370 398.800 ;
        RECT 1446.470 397.900 1446.750 398.180 ;
        RECT 1447.090 397.900 1447.370 398.180 ;
        RECT 1446.470 397.280 1446.750 397.560 ;
        RECT 1447.090 397.280 1447.370 397.560 ;
        RECT 1446.470 396.660 1446.750 396.940 ;
        RECT 1447.090 396.660 1447.370 396.940 ;
        RECT 1446.470 396.040 1446.750 396.320 ;
        RECT 1447.090 396.040 1447.370 396.320 ;
        RECT 1496.470 399.760 1496.750 400.040 ;
        RECT 1497.090 399.760 1497.370 400.040 ;
        RECT 1496.470 399.140 1496.750 399.420 ;
        RECT 1497.090 399.140 1497.370 399.420 ;
        RECT 1496.470 398.520 1496.750 398.800 ;
        RECT 1497.090 398.520 1497.370 398.800 ;
        RECT 1496.470 397.900 1496.750 398.180 ;
        RECT 1497.090 397.900 1497.370 398.180 ;
        RECT 1496.470 397.280 1496.750 397.560 ;
        RECT 1497.090 397.280 1497.370 397.560 ;
        RECT 1496.470 396.660 1496.750 396.940 ;
        RECT 1497.090 396.660 1497.370 396.940 ;
        RECT 1496.470 396.040 1496.750 396.320 ;
        RECT 1497.090 396.040 1497.370 396.320 ;
        RECT 1471.470 392.760 1471.750 393.040 ;
        RECT 1472.090 392.760 1472.370 393.040 ;
        RECT 1471.470 392.140 1471.750 392.420 ;
        RECT 1472.090 392.140 1472.370 392.420 ;
        RECT 1471.470 391.520 1471.750 391.800 ;
        RECT 1472.090 391.520 1472.370 391.800 ;
        RECT 1471.470 390.900 1471.750 391.180 ;
        RECT 1472.090 390.900 1472.370 391.180 ;
        RECT 1471.470 390.280 1471.750 390.560 ;
        RECT 1472.090 390.280 1472.370 390.560 ;
        RECT 1471.470 389.660 1471.750 389.940 ;
        RECT 1472.090 389.660 1472.370 389.940 ;
        RECT 1471.470 389.040 1471.750 389.320 ;
        RECT 1472.090 389.040 1472.370 389.320 ;
        RECT 1546.470 399.760 1546.750 400.040 ;
        RECT 1547.090 399.760 1547.370 400.040 ;
        RECT 1546.470 399.140 1546.750 399.420 ;
        RECT 1547.090 399.140 1547.370 399.420 ;
        RECT 1546.470 398.520 1546.750 398.800 ;
        RECT 1547.090 398.520 1547.370 398.800 ;
        RECT 1546.470 397.900 1546.750 398.180 ;
        RECT 1547.090 397.900 1547.370 398.180 ;
        RECT 1546.470 397.280 1546.750 397.560 ;
        RECT 1547.090 397.280 1547.370 397.560 ;
        RECT 1546.470 396.660 1546.750 396.940 ;
        RECT 1547.090 396.660 1547.370 396.940 ;
        RECT 1546.470 396.040 1546.750 396.320 ;
        RECT 1547.090 396.040 1547.370 396.320 ;
        RECT 1521.470 392.760 1521.750 393.040 ;
        RECT 1522.090 392.760 1522.370 393.040 ;
        RECT 1521.470 392.140 1521.750 392.420 ;
        RECT 1522.090 392.140 1522.370 392.420 ;
        RECT 1521.470 391.520 1521.750 391.800 ;
        RECT 1522.090 391.520 1522.370 391.800 ;
        RECT 1521.470 390.900 1521.750 391.180 ;
        RECT 1522.090 390.900 1522.370 391.180 ;
        RECT 1521.470 390.280 1521.750 390.560 ;
        RECT 1522.090 390.280 1522.370 390.560 ;
        RECT 1521.470 389.660 1521.750 389.940 ;
        RECT 1522.090 389.660 1522.370 389.940 ;
        RECT 1521.470 389.040 1521.750 389.320 ;
        RECT 1522.090 389.040 1522.370 389.320 ;
        RECT 1596.470 399.760 1596.750 400.040 ;
        RECT 1597.090 399.760 1597.370 400.040 ;
        RECT 1596.470 399.140 1596.750 399.420 ;
        RECT 1597.090 399.140 1597.370 399.420 ;
        RECT 1596.470 398.520 1596.750 398.800 ;
        RECT 1597.090 398.520 1597.370 398.800 ;
        RECT 1596.470 397.900 1596.750 398.180 ;
        RECT 1597.090 397.900 1597.370 398.180 ;
        RECT 1596.470 397.280 1596.750 397.560 ;
        RECT 1597.090 397.280 1597.370 397.560 ;
        RECT 1596.470 396.660 1596.750 396.940 ;
        RECT 1597.090 396.660 1597.370 396.940 ;
        RECT 1596.470 396.040 1596.750 396.320 ;
        RECT 1597.090 396.040 1597.370 396.320 ;
        RECT 1571.470 392.760 1571.750 393.040 ;
        RECT 1572.090 392.760 1572.370 393.040 ;
        RECT 1571.470 392.140 1571.750 392.420 ;
        RECT 1572.090 392.140 1572.370 392.420 ;
        RECT 1571.470 391.520 1571.750 391.800 ;
        RECT 1572.090 391.520 1572.370 391.800 ;
        RECT 1571.470 390.900 1571.750 391.180 ;
        RECT 1572.090 390.900 1572.370 391.180 ;
        RECT 1571.470 390.280 1571.750 390.560 ;
        RECT 1572.090 390.280 1572.370 390.560 ;
        RECT 1571.470 389.660 1571.750 389.940 ;
        RECT 1572.090 389.660 1572.370 389.940 ;
        RECT 1571.470 389.040 1571.750 389.320 ;
        RECT 1572.090 389.040 1572.370 389.320 ;
        RECT 1646.470 399.760 1646.750 400.040 ;
        RECT 1647.090 399.760 1647.370 400.040 ;
        RECT 1646.470 399.140 1646.750 399.420 ;
        RECT 1647.090 399.140 1647.370 399.420 ;
        RECT 1646.470 398.520 1646.750 398.800 ;
        RECT 1647.090 398.520 1647.370 398.800 ;
        RECT 1646.470 397.900 1646.750 398.180 ;
        RECT 1647.090 397.900 1647.370 398.180 ;
        RECT 1646.470 397.280 1646.750 397.560 ;
        RECT 1647.090 397.280 1647.370 397.560 ;
        RECT 1646.470 396.660 1646.750 396.940 ;
        RECT 1647.090 396.660 1647.370 396.940 ;
        RECT 1646.470 396.040 1646.750 396.320 ;
        RECT 1647.090 396.040 1647.370 396.320 ;
        RECT 1621.470 392.760 1621.750 393.040 ;
        RECT 1622.090 392.760 1622.370 393.040 ;
        RECT 1621.470 392.140 1621.750 392.420 ;
        RECT 1622.090 392.140 1622.370 392.420 ;
        RECT 1621.470 391.520 1621.750 391.800 ;
        RECT 1622.090 391.520 1622.370 391.800 ;
        RECT 1621.470 390.900 1621.750 391.180 ;
        RECT 1622.090 390.900 1622.370 391.180 ;
        RECT 1621.470 390.280 1621.750 390.560 ;
        RECT 1622.090 390.280 1622.370 390.560 ;
        RECT 1621.470 389.660 1621.750 389.940 ;
        RECT 1622.090 389.660 1622.370 389.940 ;
        RECT 1621.470 389.040 1621.750 389.320 ;
        RECT 1622.090 389.040 1622.370 389.320 ;
        RECT 1696.470 399.760 1696.750 400.040 ;
        RECT 1697.090 399.760 1697.370 400.040 ;
        RECT 1696.470 399.140 1696.750 399.420 ;
        RECT 1697.090 399.140 1697.370 399.420 ;
        RECT 1696.470 398.520 1696.750 398.800 ;
        RECT 1697.090 398.520 1697.370 398.800 ;
        RECT 1696.470 397.900 1696.750 398.180 ;
        RECT 1697.090 397.900 1697.370 398.180 ;
        RECT 1696.470 397.280 1696.750 397.560 ;
        RECT 1697.090 397.280 1697.370 397.560 ;
        RECT 1696.470 396.660 1696.750 396.940 ;
        RECT 1697.090 396.660 1697.370 396.940 ;
        RECT 1696.470 396.040 1696.750 396.320 ;
        RECT 1697.090 396.040 1697.370 396.320 ;
        RECT 1671.470 392.760 1671.750 393.040 ;
        RECT 1672.090 392.760 1672.370 393.040 ;
        RECT 1671.470 392.140 1671.750 392.420 ;
        RECT 1672.090 392.140 1672.370 392.420 ;
        RECT 1671.470 391.520 1671.750 391.800 ;
        RECT 1672.090 391.520 1672.370 391.800 ;
        RECT 1671.470 390.900 1671.750 391.180 ;
        RECT 1672.090 390.900 1672.370 391.180 ;
        RECT 1671.470 390.280 1671.750 390.560 ;
        RECT 1672.090 390.280 1672.370 390.560 ;
        RECT 1671.470 389.660 1671.750 389.940 ;
        RECT 1672.090 389.660 1672.370 389.940 ;
        RECT 1671.470 389.040 1671.750 389.320 ;
        RECT 1672.090 389.040 1672.370 389.320 ;
        RECT 1746.470 399.760 1746.750 400.040 ;
        RECT 1747.090 399.760 1747.370 400.040 ;
        RECT 1746.470 399.140 1746.750 399.420 ;
        RECT 1747.090 399.140 1747.370 399.420 ;
        RECT 1746.470 398.520 1746.750 398.800 ;
        RECT 1747.090 398.520 1747.370 398.800 ;
        RECT 1746.470 397.900 1746.750 398.180 ;
        RECT 1747.090 397.900 1747.370 398.180 ;
        RECT 1746.470 397.280 1746.750 397.560 ;
        RECT 1747.090 397.280 1747.370 397.560 ;
        RECT 1746.470 396.660 1746.750 396.940 ;
        RECT 1747.090 396.660 1747.370 396.940 ;
        RECT 1746.470 396.040 1746.750 396.320 ;
        RECT 1747.090 396.040 1747.370 396.320 ;
        RECT 1721.470 392.760 1721.750 393.040 ;
        RECT 1722.090 392.760 1722.370 393.040 ;
        RECT 1721.470 392.140 1721.750 392.420 ;
        RECT 1722.090 392.140 1722.370 392.420 ;
        RECT 1721.470 391.520 1721.750 391.800 ;
        RECT 1722.090 391.520 1722.370 391.800 ;
        RECT 1721.470 390.900 1721.750 391.180 ;
        RECT 1722.090 390.900 1722.370 391.180 ;
        RECT 1721.470 390.280 1721.750 390.560 ;
        RECT 1722.090 390.280 1722.370 390.560 ;
        RECT 1721.470 389.660 1721.750 389.940 ;
        RECT 1722.090 389.660 1722.370 389.940 ;
        RECT 1721.470 389.040 1721.750 389.320 ;
        RECT 1722.090 389.040 1722.370 389.320 ;
        RECT 1796.470 399.760 1796.750 400.040 ;
        RECT 1797.090 399.760 1797.370 400.040 ;
        RECT 1796.470 399.140 1796.750 399.420 ;
        RECT 1797.090 399.140 1797.370 399.420 ;
        RECT 1796.470 398.520 1796.750 398.800 ;
        RECT 1797.090 398.520 1797.370 398.800 ;
        RECT 1796.470 397.900 1796.750 398.180 ;
        RECT 1797.090 397.900 1797.370 398.180 ;
        RECT 1796.470 397.280 1796.750 397.560 ;
        RECT 1797.090 397.280 1797.370 397.560 ;
        RECT 1796.470 396.660 1796.750 396.940 ;
        RECT 1797.090 396.660 1797.370 396.940 ;
        RECT 1796.470 396.040 1796.750 396.320 ;
        RECT 1797.090 396.040 1797.370 396.320 ;
        RECT 1771.470 392.760 1771.750 393.040 ;
        RECT 1772.090 392.760 1772.370 393.040 ;
        RECT 1771.470 392.140 1771.750 392.420 ;
        RECT 1772.090 392.140 1772.370 392.420 ;
        RECT 1771.470 391.520 1771.750 391.800 ;
        RECT 1772.090 391.520 1772.370 391.800 ;
        RECT 1771.470 390.900 1771.750 391.180 ;
        RECT 1772.090 390.900 1772.370 391.180 ;
        RECT 1771.470 390.280 1771.750 390.560 ;
        RECT 1772.090 390.280 1772.370 390.560 ;
        RECT 1771.470 389.660 1771.750 389.940 ;
        RECT 1772.090 389.660 1772.370 389.940 ;
        RECT 1771.470 389.040 1771.750 389.320 ;
        RECT 1772.090 389.040 1772.370 389.320 ;
        RECT 1846.470 399.760 1846.750 400.040 ;
        RECT 1847.090 399.760 1847.370 400.040 ;
        RECT 1846.470 399.140 1846.750 399.420 ;
        RECT 1847.090 399.140 1847.370 399.420 ;
        RECT 1846.470 398.520 1846.750 398.800 ;
        RECT 1847.090 398.520 1847.370 398.800 ;
        RECT 1846.470 397.900 1846.750 398.180 ;
        RECT 1847.090 397.900 1847.370 398.180 ;
        RECT 1846.470 397.280 1846.750 397.560 ;
        RECT 1847.090 397.280 1847.370 397.560 ;
        RECT 1846.470 396.660 1846.750 396.940 ;
        RECT 1847.090 396.660 1847.370 396.940 ;
        RECT 1846.470 396.040 1846.750 396.320 ;
        RECT 1847.090 396.040 1847.370 396.320 ;
        RECT 1821.470 392.760 1821.750 393.040 ;
        RECT 1822.090 392.760 1822.370 393.040 ;
        RECT 1821.470 392.140 1821.750 392.420 ;
        RECT 1822.090 392.140 1822.370 392.420 ;
        RECT 1821.470 391.520 1821.750 391.800 ;
        RECT 1822.090 391.520 1822.370 391.800 ;
        RECT 1821.470 390.900 1821.750 391.180 ;
        RECT 1822.090 390.900 1822.370 391.180 ;
        RECT 1821.470 390.280 1821.750 390.560 ;
        RECT 1822.090 390.280 1822.370 390.560 ;
        RECT 1821.470 389.660 1821.750 389.940 ;
        RECT 1822.090 389.660 1822.370 389.940 ;
        RECT 1821.470 389.040 1821.750 389.320 ;
        RECT 1822.090 389.040 1822.370 389.320 ;
        RECT 1896.470 399.760 1896.750 400.040 ;
        RECT 1897.090 399.760 1897.370 400.040 ;
        RECT 1896.470 399.140 1896.750 399.420 ;
        RECT 1897.090 399.140 1897.370 399.420 ;
        RECT 1896.470 398.520 1896.750 398.800 ;
        RECT 1897.090 398.520 1897.370 398.800 ;
        RECT 1896.470 397.900 1896.750 398.180 ;
        RECT 1897.090 397.900 1897.370 398.180 ;
        RECT 1896.470 397.280 1896.750 397.560 ;
        RECT 1897.090 397.280 1897.370 397.560 ;
        RECT 1896.470 396.660 1896.750 396.940 ;
        RECT 1897.090 396.660 1897.370 396.940 ;
        RECT 1896.470 396.040 1896.750 396.320 ;
        RECT 1897.090 396.040 1897.370 396.320 ;
        RECT 1871.470 392.760 1871.750 393.040 ;
        RECT 1872.090 392.760 1872.370 393.040 ;
        RECT 1871.470 392.140 1871.750 392.420 ;
        RECT 1872.090 392.140 1872.370 392.420 ;
        RECT 1871.470 391.520 1871.750 391.800 ;
        RECT 1872.090 391.520 1872.370 391.800 ;
        RECT 1871.470 390.900 1871.750 391.180 ;
        RECT 1872.090 390.900 1872.370 391.180 ;
        RECT 1871.470 390.280 1871.750 390.560 ;
        RECT 1872.090 390.280 1872.370 390.560 ;
        RECT 1871.470 389.660 1871.750 389.940 ;
        RECT 1872.090 389.660 1872.370 389.940 ;
        RECT 1871.470 389.040 1871.750 389.320 ;
        RECT 1872.090 389.040 1872.370 389.320 ;
        RECT 1946.470 399.760 1946.750 400.040 ;
        RECT 1947.090 399.760 1947.370 400.040 ;
        RECT 1946.470 399.140 1946.750 399.420 ;
        RECT 1947.090 399.140 1947.370 399.420 ;
        RECT 1946.470 398.520 1946.750 398.800 ;
        RECT 1947.090 398.520 1947.370 398.800 ;
        RECT 1946.470 397.900 1946.750 398.180 ;
        RECT 1947.090 397.900 1947.370 398.180 ;
        RECT 1946.470 397.280 1946.750 397.560 ;
        RECT 1947.090 397.280 1947.370 397.560 ;
        RECT 1946.470 396.660 1946.750 396.940 ;
        RECT 1947.090 396.660 1947.370 396.940 ;
        RECT 1946.470 396.040 1946.750 396.320 ;
        RECT 1947.090 396.040 1947.370 396.320 ;
        RECT 1921.470 392.760 1921.750 393.040 ;
        RECT 1922.090 392.760 1922.370 393.040 ;
        RECT 1921.470 392.140 1921.750 392.420 ;
        RECT 1922.090 392.140 1922.370 392.420 ;
        RECT 1921.470 391.520 1921.750 391.800 ;
        RECT 1922.090 391.520 1922.370 391.800 ;
        RECT 1921.470 390.900 1921.750 391.180 ;
        RECT 1922.090 390.900 1922.370 391.180 ;
        RECT 1921.470 390.280 1921.750 390.560 ;
        RECT 1922.090 390.280 1922.370 390.560 ;
        RECT 1921.470 389.660 1921.750 389.940 ;
        RECT 1922.090 389.660 1922.370 389.940 ;
        RECT 1921.470 389.040 1921.750 389.320 ;
        RECT 1922.090 389.040 1922.370 389.320 ;
        RECT 1996.470 399.760 1996.750 400.040 ;
        RECT 1997.090 399.760 1997.370 400.040 ;
        RECT 1996.470 399.140 1996.750 399.420 ;
        RECT 1997.090 399.140 1997.370 399.420 ;
        RECT 1996.470 398.520 1996.750 398.800 ;
        RECT 1997.090 398.520 1997.370 398.800 ;
        RECT 1996.470 397.900 1996.750 398.180 ;
        RECT 1997.090 397.900 1997.370 398.180 ;
        RECT 1996.470 397.280 1996.750 397.560 ;
        RECT 1997.090 397.280 1997.370 397.560 ;
        RECT 1996.470 396.660 1996.750 396.940 ;
        RECT 1997.090 396.660 1997.370 396.940 ;
        RECT 1996.470 396.040 1996.750 396.320 ;
        RECT 1997.090 396.040 1997.370 396.320 ;
        RECT 1971.470 392.760 1971.750 393.040 ;
        RECT 1972.090 392.760 1972.370 393.040 ;
        RECT 1971.470 392.140 1971.750 392.420 ;
        RECT 1972.090 392.140 1972.370 392.420 ;
        RECT 1971.470 391.520 1971.750 391.800 ;
        RECT 1972.090 391.520 1972.370 391.800 ;
        RECT 1971.470 390.900 1971.750 391.180 ;
        RECT 1972.090 390.900 1972.370 391.180 ;
        RECT 1971.470 390.280 1971.750 390.560 ;
        RECT 1972.090 390.280 1972.370 390.560 ;
        RECT 1971.470 389.660 1971.750 389.940 ;
        RECT 1972.090 389.660 1972.370 389.940 ;
        RECT 1971.470 389.040 1971.750 389.320 ;
        RECT 1972.090 389.040 1972.370 389.320 ;
        RECT 2046.470 399.760 2046.750 400.040 ;
        RECT 2047.090 399.760 2047.370 400.040 ;
        RECT 2046.470 399.140 2046.750 399.420 ;
        RECT 2047.090 399.140 2047.370 399.420 ;
        RECT 2046.470 398.520 2046.750 398.800 ;
        RECT 2047.090 398.520 2047.370 398.800 ;
        RECT 2046.470 397.900 2046.750 398.180 ;
        RECT 2047.090 397.900 2047.370 398.180 ;
        RECT 2046.470 397.280 2046.750 397.560 ;
        RECT 2047.090 397.280 2047.370 397.560 ;
        RECT 2046.470 396.660 2046.750 396.940 ;
        RECT 2047.090 396.660 2047.370 396.940 ;
        RECT 2046.470 396.040 2046.750 396.320 ;
        RECT 2047.090 396.040 2047.370 396.320 ;
        RECT 2021.470 392.760 2021.750 393.040 ;
        RECT 2022.090 392.760 2022.370 393.040 ;
        RECT 2021.470 392.140 2021.750 392.420 ;
        RECT 2022.090 392.140 2022.370 392.420 ;
        RECT 2021.470 391.520 2021.750 391.800 ;
        RECT 2022.090 391.520 2022.370 391.800 ;
        RECT 2021.470 390.900 2021.750 391.180 ;
        RECT 2022.090 390.900 2022.370 391.180 ;
        RECT 2021.470 390.280 2021.750 390.560 ;
        RECT 2022.090 390.280 2022.370 390.560 ;
        RECT 2021.470 389.660 2021.750 389.940 ;
        RECT 2022.090 389.660 2022.370 389.940 ;
        RECT 2021.470 389.040 2021.750 389.320 ;
        RECT 2022.090 389.040 2022.370 389.320 ;
        RECT 2096.470 399.760 2096.750 400.040 ;
        RECT 2097.090 399.760 2097.370 400.040 ;
        RECT 2096.470 399.140 2096.750 399.420 ;
        RECT 2097.090 399.140 2097.370 399.420 ;
        RECT 2096.470 398.520 2096.750 398.800 ;
        RECT 2097.090 398.520 2097.370 398.800 ;
        RECT 2096.470 397.900 2096.750 398.180 ;
        RECT 2097.090 397.900 2097.370 398.180 ;
        RECT 2096.470 397.280 2096.750 397.560 ;
        RECT 2097.090 397.280 2097.370 397.560 ;
        RECT 2096.470 396.660 2096.750 396.940 ;
        RECT 2097.090 396.660 2097.370 396.940 ;
        RECT 2096.470 396.040 2096.750 396.320 ;
        RECT 2097.090 396.040 2097.370 396.320 ;
        RECT 2071.470 392.760 2071.750 393.040 ;
        RECT 2072.090 392.760 2072.370 393.040 ;
        RECT 2071.470 392.140 2071.750 392.420 ;
        RECT 2072.090 392.140 2072.370 392.420 ;
        RECT 2071.470 391.520 2071.750 391.800 ;
        RECT 2072.090 391.520 2072.370 391.800 ;
        RECT 2071.470 390.900 2071.750 391.180 ;
        RECT 2072.090 390.900 2072.370 391.180 ;
        RECT 2071.470 390.280 2071.750 390.560 ;
        RECT 2072.090 390.280 2072.370 390.560 ;
        RECT 2071.470 389.660 2071.750 389.940 ;
        RECT 2072.090 389.660 2072.370 389.940 ;
        RECT 2071.470 389.040 2071.750 389.320 ;
        RECT 2072.090 389.040 2072.370 389.320 ;
        RECT 2146.470 399.760 2146.750 400.040 ;
        RECT 2147.090 399.760 2147.370 400.040 ;
        RECT 2146.470 399.140 2146.750 399.420 ;
        RECT 2147.090 399.140 2147.370 399.420 ;
        RECT 2146.470 398.520 2146.750 398.800 ;
        RECT 2147.090 398.520 2147.370 398.800 ;
        RECT 2146.470 397.900 2146.750 398.180 ;
        RECT 2147.090 397.900 2147.370 398.180 ;
        RECT 2146.470 397.280 2146.750 397.560 ;
        RECT 2147.090 397.280 2147.370 397.560 ;
        RECT 2146.470 396.660 2146.750 396.940 ;
        RECT 2147.090 396.660 2147.370 396.940 ;
        RECT 2146.470 396.040 2146.750 396.320 ;
        RECT 2147.090 396.040 2147.370 396.320 ;
        RECT 2121.470 392.760 2121.750 393.040 ;
        RECT 2122.090 392.760 2122.370 393.040 ;
        RECT 2121.470 392.140 2121.750 392.420 ;
        RECT 2122.090 392.140 2122.370 392.420 ;
        RECT 2121.470 391.520 2121.750 391.800 ;
        RECT 2122.090 391.520 2122.370 391.800 ;
        RECT 2121.470 390.900 2121.750 391.180 ;
        RECT 2122.090 390.900 2122.370 391.180 ;
        RECT 2121.470 390.280 2121.750 390.560 ;
        RECT 2122.090 390.280 2122.370 390.560 ;
        RECT 2121.470 389.660 2121.750 389.940 ;
        RECT 2122.090 389.660 2122.370 389.940 ;
        RECT 2121.470 389.040 2121.750 389.320 ;
        RECT 2122.090 389.040 2122.370 389.320 ;
        RECT 2196.470 399.760 2196.750 400.040 ;
        RECT 2197.090 399.760 2197.370 400.040 ;
        RECT 2196.470 399.140 2196.750 399.420 ;
        RECT 2197.090 399.140 2197.370 399.420 ;
        RECT 2196.470 398.520 2196.750 398.800 ;
        RECT 2197.090 398.520 2197.370 398.800 ;
        RECT 2196.470 397.900 2196.750 398.180 ;
        RECT 2197.090 397.900 2197.370 398.180 ;
        RECT 2196.470 397.280 2196.750 397.560 ;
        RECT 2197.090 397.280 2197.370 397.560 ;
        RECT 2196.470 396.660 2196.750 396.940 ;
        RECT 2197.090 396.660 2197.370 396.940 ;
        RECT 2196.470 396.040 2196.750 396.320 ;
        RECT 2197.090 396.040 2197.370 396.320 ;
        RECT 2171.470 392.760 2171.750 393.040 ;
        RECT 2172.090 392.760 2172.370 393.040 ;
        RECT 2171.470 392.140 2171.750 392.420 ;
        RECT 2172.090 392.140 2172.370 392.420 ;
        RECT 2171.470 391.520 2171.750 391.800 ;
        RECT 2172.090 391.520 2172.370 391.800 ;
        RECT 2171.470 390.900 2171.750 391.180 ;
        RECT 2172.090 390.900 2172.370 391.180 ;
        RECT 2171.470 390.280 2171.750 390.560 ;
        RECT 2172.090 390.280 2172.370 390.560 ;
        RECT 2171.470 389.660 2171.750 389.940 ;
        RECT 2172.090 389.660 2172.370 389.940 ;
        RECT 2171.470 389.040 2171.750 389.320 ;
        RECT 2172.090 389.040 2172.370 389.320 ;
        RECT 2246.470 399.760 2246.750 400.040 ;
        RECT 2247.090 399.760 2247.370 400.040 ;
        RECT 2246.470 399.140 2246.750 399.420 ;
        RECT 2247.090 399.140 2247.370 399.420 ;
        RECT 2246.470 398.520 2246.750 398.800 ;
        RECT 2247.090 398.520 2247.370 398.800 ;
        RECT 2246.470 397.900 2246.750 398.180 ;
        RECT 2247.090 397.900 2247.370 398.180 ;
        RECT 2246.470 397.280 2246.750 397.560 ;
        RECT 2247.090 397.280 2247.370 397.560 ;
        RECT 2246.470 396.660 2246.750 396.940 ;
        RECT 2247.090 396.660 2247.370 396.940 ;
        RECT 2246.470 396.040 2246.750 396.320 ;
        RECT 2247.090 396.040 2247.370 396.320 ;
        RECT 2221.470 392.760 2221.750 393.040 ;
        RECT 2222.090 392.760 2222.370 393.040 ;
        RECT 2221.470 392.140 2221.750 392.420 ;
        RECT 2222.090 392.140 2222.370 392.420 ;
        RECT 2221.470 391.520 2221.750 391.800 ;
        RECT 2222.090 391.520 2222.370 391.800 ;
        RECT 2221.470 390.900 2221.750 391.180 ;
        RECT 2222.090 390.900 2222.370 391.180 ;
        RECT 2221.470 390.280 2221.750 390.560 ;
        RECT 2222.090 390.280 2222.370 390.560 ;
        RECT 2221.470 389.660 2221.750 389.940 ;
        RECT 2222.090 389.660 2222.370 389.940 ;
        RECT 2221.470 389.040 2221.750 389.320 ;
        RECT 2222.090 389.040 2222.370 389.320 ;
        RECT 2296.470 399.760 2296.750 400.040 ;
        RECT 2297.090 399.760 2297.370 400.040 ;
        RECT 2296.470 399.140 2296.750 399.420 ;
        RECT 2297.090 399.140 2297.370 399.420 ;
        RECT 2296.470 398.520 2296.750 398.800 ;
        RECT 2297.090 398.520 2297.370 398.800 ;
        RECT 2296.470 397.900 2296.750 398.180 ;
        RECT 2297.090 397.900 2297.370 398.180 ;
        RECT 2296.470 397.280 2296.750 397.560 ;
        RECT 2297.090 397.280 2297.370 397.560 ;
        RECT 2296.470 396.660 2296.750 396.940 ;
        RECT 2297.090 396.660 2297.370 396.940 ;
        RECT 2296.470 396.040 2296.750 396.320 ;
        RECT 2297.090 396.040 2297.370 396.320 ;
        RECT 2271.470 392.760 2271.750 393.040 ;
        RECT 2272.090 392.760 2272.370 393.040 ;
        RECT 2271.470 392.140 2271.750 392.420 ;
        RECT 2272.090 392.140 2272.370 392.420 ;
        RECT 2271.470 391.520 2271.750 391.800 ;
        RECT 2272.090 391.520 2272.370 391.800 ;
        RECT 2271.470 390.900 2271.750 391.180 ;
        RECT 2272.090 390.900 2272.370 391.180 ;
        RECT 2271.470 390.280 2271.750 390.560 ;
        RECT 2272.090 390.280 2272.370 390.560 ;
        RECT 2271.470 389.660 2271.750 389.940 ;
        RECT 2272.090 389.660 2272.370 389.940 ;
        RECT 2271.470 389.040 2271.750 389.320 ;
        RECT 2272.090 389.040 2272.370 389.320 ;
        RECT 2346.470 399.760 2346.750 400.040 ;
        RECT 2347.090 399.760 2347.370 400.040 ;
        RECT 2346.470 399.140 2346.750 399.420 ;
        RECT 2347.090 399.140 2347.370 399.420 ;
        RECT 2346.470 398.520 2346.750 398.800 ;
        RECT 2347.090 398.520 2347.370 398.800 ;
        RECT 2346.470 397.900 2346.750 398.180 ;
        RECT 2347.090 397.900 2347.370 398.180 ;
        RECT 2346.470 397.280 2346.750 397.560 ;
        RECT 2347.090 397.280 2347.370 397.560 ;
        RECT 2346.470 396.660 2346.750 396.940 ;
        RECT 2347.090 396.660 2347.370 396.940 ;
        RECT 2346.470 396.040 2346.750 396.320 ;
        RECT 2347.090 396.040 2347.370 396.320 ;
        RECT 2321.470 392.760 2321.750 393.040 ;
        RECT 2322.090 392.760 2322.370 393.040 ;
        RECT 2321.470 392.140 2321.750 392.420 ;
        RECT 2322.090 392.140 2322.370 392.420 ;
        RECT 2321.470 391.520 2321.750 391.800 ;
        RECT 2322.090 391.520 2322.370 391.800 ;
        RECT 2321.470 390.900 2321.750 391.180 ;
        RECT 2322.090 390.900 2322.370 391.180 ;
        RECT 2321.470 390.280 2321.750 390.560 ;
        RECT 2322.090 390.280 2322.370 390.560 ;
        RECT 2321.470 389.660 2321.750 389.940 ;
        RECT 2322.090 389.660 2322.370 389.940 ;
        RECT 2321.470 389.040 2321.750 389.320 ;
        RECT 2322.090 389.040 2322.370 389.320 ;
        RECT 2396.470 399.760 2396.750 400.040 ;
        RECT 2397.090 399.760 2397.370 400.040 ;
        RECT 2396.470 399.140 2396.750 399.420 ;
        RECT 2397.090 399.140 2397.370 399.420 ;
        RECT 2396.470 398.520 2396.750 398.800 ;
        RECT 2397.090 398.520 2397.370 398.800 ;
        RECT 2396.470 397.900 2396.750 398.180 ;
        RECT 2397.090 397.900 2397.370 398.180 ;
        RECT 2396.470 397.280 2396.750 397.560 ;
        RECT 2397.090 397.280 2397.370 397.560 ;
        RECT 2396.470 396.660 2396.750 396.940 ;
        RECT 2397.090 396.660 2397.370 396.940 ;
        RECT 2396.470 396.040 2396.750 396.320 ;
        RECT 2397.090 396.040 2397.370 396.320 ;
        RECT 2371.470 392.760 2371.750 393.040 ;
        RECT 2372.090 392.760 2372.370 393.040 ;
        RECT 2371.470 392.140 2371.750 392.420 ;
        RECT 2372.090 392.140 2372.370 392.420 ;
        RECT 2371.470 391.520 2371.750 391.800 ;
        RECT 2372.090 391.520 2372.370 391.800 ;
        RECT 2371.470 390.900 2371.750 391.180 ;
        RECT 2372.090 390.900 2372.370 391.180 ;
        RECT 2371.470 390.280 2371.750 390.560 ;
        RECT 2372.090 390.280 2372.370 390.560 ;
        RECT 2371.470 389.660 2371.750 389.940 ;
        RECT 2372.090 389.660 2372.370 389.940 ;
        RECT 2371.470 389.040 2371.750 389.320 ;
        RECT 2372.090 389.040 2372.370 389.320 ;
        RECT 2446.470 399.760 2446.750 400.040 ;
        RECT 2447.090 399.760 2447.370 400.040 ;
        RECT 2446.470 399.140 2446.750 399.420 ;
        RECT 2447.090 399.140 2447.370 399.420 ;
        RECT 2446.470 398.520 2446.750 398.800 ;
        RECT 2447.090 398.520 2447.370 398.800 ;
        RECT 2446.470 397.900 2446.750 398.180 ;
        RECT 2447.090 397.900 2447.370 398.180 ;
        RECT 2446.470 397.280 2446.750 397.560 ;
        RECT 2447.090 397.280 2447.370 397.560 ;
        RECT 2446.470 396.660 2446.750 396.940 ;
        RECT 2447.090 396.660 2447.370 396.940 ;
        RECT 2446.470 396.040 2446.750 396.320 ;
        RECT 2447.090 396.040 2447.370 396.320 ;
        RECT 2421.470 392.760 2421.750 393.040 ;
        RECT 2422.090 392.760 2422.370 393.040 ;
        RECT 2421.470 392.140 2421.750 392.420 ;
        RECT 2422.090 392.140 2422.370 392.420 ;
        RECT 2421.470 391.520 2421.750 391.800 ;
        RECT 2422.090 391.520 2422.370 391.800 ;
        RECT 2421.470 390.900 2421.750 391.180 ;
        RECT 2422.090 390.900 2422.370 391.180 ;
        RECT 2421.470 390.280 2421.750 390.560 ;
        RECT 2422.090 390.280 2422.370 390.560 ;
        RECT 2421.470 389.660 2421.750 389.940 ;
        RECT 2422.090 389.660 2422.370 389.940 ;
        RECT 2421.470 389.040 2421.750 389.320 ;
        RECT 2422.090 389.040 2422.370 389.320 ;
        RECT 2496.470 399.760 2496.750 400.040 ;
        RECT 2497.090 399.760 2497.370 400.040 ;
        RECT 2496.470 399.140 2496.750 399.420 ;
        RECT 2497.090 399.140 2497.370 399.420 ;
        RECT 2496.470 398.520 2496.750 398.800 ;
        RECT 2497.090 398.520 2497.370 398.800 ;
        RECT 2496.470 397.900 2496.750 398.180 ;
        RECT 2497.090 397.900 2497.370 398.180 ;
        RECT 2496.470 397.280 2496.750 397.560 ;
        RECT 2497.090 397.280 2497.370 397.560 ;
        RECT 2496.470 396.660 2496.750 396.940 ;
        RECT 2497.090 396.660 2497.370 396.940 ;
        RECT 2496.470 396.040 2496.750 396.320 ;
        RECT 2497.090 396.040 2497.370 396.320 ;
        RECT 2471.470 392.760 2471.750 393.040 ;
        RECT 2472.090 392.760 2472.370 393.040 ;
        RECT 2471.470 392.140 2471.750 392.420 ;
        RECT 2472.090 392.140 2472.370 392.420 ;
        RECT 2471.470 391.520 2471.750 391.800 ;
        RECT 2472.090 391.520 2472.370 391.800 ;
        RECT 2471.470 390.900 2471.750 391.180 ;
        RECT 2472.090 390.900 2472.370 391.180 ;
        RECT 2471.470 390.280 2471.750 390.560 ;
        RECT 2472.090 390.280 2472.370 390.560 ;
        RECT 2471.470 389.660 2471.750 389.940 ;
        RECT 2472.090 389.660 2472.370 389.940 ;
        RECT 2471.470 389.040 2471.750 389.320 ;
        RECT 2472.090 389.040 2472.370 389.320 ;
        RECT 2546.470 399.760 2546.750 400.040 ;
        RECT 2547.090 399.760 2547.370 400.040 ;
        RECT 2546.470 399.140 2546.750 399.420 ;
        RECT 2547.090 399.140 2547.370 399.420 ;
        RECT 2546.470 398.520 2546.750 398.800 ;
        RECT 2547.090 398.520 2547.370 398.800 ;
        RECT 2546.470 397.900 2546.750 398.180 ;
        RECT 2547.090 397.900 2547.370 398.180 ;
        RECT 2546.470 397.280 2546.750 397.560 ;
        RECT 2547.090 397.280 2547.370 397.560 ;
        RECT 2546.470 396.660 2546.750 396.940 ;
        RECT 2547.090 396.660 2547.370 396.940 ;
        RECT 2546.470 396.040 2546.750 396.320 ;
        RECT 2547.090 396.040 2547.370 396.320 ;
        RECT 2521.470 392.760 2521.750 393.040 ;
        RECT 2522.090 392.760 2522.370 393.040 ;
        RECT 2521.470 392.140 2521.750 392.420 ;
        RECT 2522.090 392.140 2522.370 392.420 ;
        RECT 2521.470 391.520 2521.750 391.800 ;
        RECT 2522.090 391.520 2522.370 391.800 ;
        RECT 2521.470 390.900 2521.750 391.180 ;
        RECT 2522.090 390.900 2522.370 391.180 ;
        RECT 2521.470 390.280 2521.750 390.560 ;
        RECT 2522.090 390.280 2522.370 390.560 ;
        RECT 2521.470 389.660 2521.750 389.940 ;
        RECT 2522.090 389.660 2522.370 389.940 ;
        RECT 2521.470 389.040 2521.750 389.320 ;
        RECT 2522.090 389.040 2522.370 389.320 ;
        RECT 2596.470 399.760 2596.750 400.040 ;
        RECT 2597.090 399.760 2597.370 400.040 ;
        RECT 2596.470 399.140 2596.750 399.420 ;
        RECT 2597.090 399.140 2597.370 399.420 ;
        RECT 2596.470 398.520 2596.750 398.800 ;
        RECT 2597.090 398.520 2597.370 398.800 ;
        RECT 2596.470 397.900 2596.750 398.180 ;
        RECT 2597.090 397.900 2597.370 398.180 ;
        RECT 2596.470 397.280 2596.750 397.560 ;
        RECT 2597.090 397.280 2597.370 397.560 ;
        RECT 2596.470 396.660 2596.750 396.940 ;
        RECT 2597.090 396.660 2597.370 396.940 ;
        RECT 2596.470 396.040 2596.750 396.320 ;
        RECT 2597.090 396.040 2597.370 396.320 ;
        RECT 2571.470 392.760 2571.750 393.040 ;
        RECT 2572.090 392.760 2572.370 393.040 ;
        RECT 2571.470 392.140 2571.750 392.420 ;
        RECT 2572.090 392.140 2572.370 392.420 ;
        RECT 2571.470 391.520 2571.750 391.800 ;
        RECT 2572.090 391.520 2572.370 391.800 ;
        RECT 2571.470 390.900 2571.750 391.180 ;
        RECT 2572.090 390.900 2572.370 391.180 ;
        RECT 2571.470 390.280 2571.750 390.560 ;
        RECT 2572.090 390.280 2572.370 390.560 ;
        RECT 2571.470 389.660 2571.750 389.940 ;
        RECT 2572.090 389.660 2572.370 389.940 ;
        RECT 2571.470 389.040 2571.750 389.320 ;
        RECT 2572.090 389.040 2572.370 389.320 ;
        RECT 2646.470 399.760 2646.750 400.040 ;
        RECT 2647.090 399.760 2647.370 400.040 ;
        RECT 2646.470 399.140 2646.750 399.420 ;
        RECT 2647.090 399.140 2647.370 399.420 ;
        RECT 2646.470 398.520 2646.750 398.800 ;
        RECT 2647.090 398.520 2647.370 398.800 ;
        RECT 2646.470 397.900 2646.750 398.180 ;
        RECT 2647.090 397.900 2647.370 398.180 ;
        RECT 2646.470 397.280 2646.750 397.560 ;
        RECT 2647.090 397.280 2647.370 397.560 ;
        RECT 2646.470 396.660 2646.750 396.940 ;
        RECT 2647.090 396.660 2647.370 396.940 ;
        RECT 2646.470 396.040 2646.750 396.320 ;
        RECT 2647.090 396.040 2647.370 396.320 ;
        RECT 2621.470 392.760 2621.750 393.040 ;
        RECT 2622.090 392.760 2622.370 393.040 ;
        RECT 2621.470 392.140 2621.750 392.420 ;
        RECT 2622.090 392.140 2622.370 392.420 ;
        RECT 2621.470 391.520 2621.750 391.800 ;
        RECT 2622.090 391.520 2622.370 391.800 ;
        RECT 2621.470 390.900 2621.750 391.180 ;
        RECT 2622.090 390.900 2622.370 391.180 ;
        RECT 2621.470 390.280 2621.750 390.560 ;
        RECT 2622.090 390.280 2622.370 390.560 ;
        RECT 2621.470 389.660 2621.750 389.940 ;
        RECT 2622.090 389.660 2622.370 389.940 ;
        RECT 2621.470 389.040 2621.750 389.320 ;
        RECT 2622.090 389.040 2622.370 389.320 ;
        RECT 2696.470 399.760 2696.750 400.040 ;
        RECT 2697.090 399.760 2697.370 400.040 ;
        RECT 2696.470 399.140 2696.750 399.420 ;
        RECT 2697.090 399.140 2697.370 399.420 ;
        RECT 2696.470 398.520 2696.750 398.800 ;
        RECT 2697.090 398.520 2697.370 398.800 ;
        RECT 2696.470 397.900 2696.750 398.180 ;
        RECT 2697.090 397.900 2697.370 398.180 ;
        RECT 2696.470 397.280 2696.750 397.560 ;
        RECT 2697.090 397.280 2697.370 397.560 ;
        RECT 2696.470 396.660 2696.750 396.940 ;
        RECT 2697.090 396.660 2697.370 396.940 ;
        RECT 2696.470 396.040 2696.750 396.320 ;
        RECT 2697.090 396.040 2697.370 396.320 ;
        RECT 2671.470 392.760 2671.750 393.040 ;
        RECT 2672.090 392.760 2672.370 393.040 ;
        RECT 2671.470 392.140 2671.750 392.420 ;
        RECT 2672.090 392.140 2672.370 392.420 ;
        RECT 2671.470 391.520 2671.750 391.800 ;
        RECT 2672.090 391.520 2672.370 391.800 ;
        RECT 2671.470 390.900 2671.750 391.180 ;
        RECT 2672.090 390.900 2672.370 391.180 ;
        RECT 2671.470 390.280 2671.750 390.560 ;
        RECT 2672.090 390.280 2672.370 390.560 ;
        RECT 2671.470 389.660 2671.750 389.940 ;
        RECT 2672.090 389.660 2672.370 389.940 ;
        RECT 2671.470 389.040 2671.750 389.320 ;
        RECT 2672.090 389.040 2672.370 389.320 ;
        RECT 2746.470 399.760 2746.750 400.040 ;
        RECT 2747.090 399.760 2747.370 400.040 ;
        RECT 2746.470 399.140 2746.750 399.420 ;
        RECT 2747.090 399.140 2747.370 399.420 ;
        RECT 2746.470 398.520 2746.750 398.800 ;
        RECT 2747.090 398.520 2747.370 398.800 ;
        RECT 2746.470 397.900 2746.750 398.180 ;
        RECT 2747.090 397.900 2747.370 398.180 ;
        RECT 2746.470 397.280 2746.750 397.560 ;
        RECT 2747.090 397.280 2747.370 397.560 ;
        RECT 2746.470 396.660 2746.750 396.940 ;
        RECT 2747.090 396.660 2747.370 396.940 ;
        RECT 2746.470 396.040 2746.750 396.320 ;
        RECT 2747.090 396.040 2747.370 396.320 ;
        RECT 2721.470 392.760 2721.750 393.040 ;
        RECT 2722.090 392.760 2722.370 393.040 ;
        RECT 2721.470 392.140 2721.750 392.420 ;
        RECT 2722.090 392.140 2722.370 392.420 ;
        RECT 2721.470 391.520 2721.750 391.800 ;
        RECT 2722.090 391.520 2722.370 391.800 ;
        RECT 2721.470 390.900 2721.750 391.180 ;
        RECT 2722.090 390.900 2722.370 391.180 ;
        RECT 2721.470 390.280 2721.750 390.560 ;
        RECT 2722.090 390.280 2722.370 390.560 ;
        RECT 2721.470 389.660 2721.750 389.940 ;
        RECT 2722.090 389.660 2722.370 389.940 ;
        RECT 2721.470 389.040 2721.750 389.320 ;
        RECT 2722.090 389.040 2722.370 389.320 ;
        RECT 2954.850 399.760 2955.130 400.040 ;
        RECT 2955.470 399.760 2955.750 400.040 ;
        RECT 2956.090 399.760 2956.370 400.040 ;
        RECT 2956.710 399.760 2956.990 400.040 ;
        RECT 2957.330 399.760 2957.610 400.040 ;
        RECT 2957.950 399.760 2958.230 400.040 ;
        RECT 2958.570 399.760 2958.850 400.040 ;
        RECT 2954.850 399.140 2955.130 399.420 ;
        RECT 2955.470 399.140 2955.750 399.420 ;
        RECT 2956.090 399.140 2956.370 399.420 ;
        RECT 2956.710 399.140 2956.990 399.420 ;
        RECT 2957.330 399.140 2957.610 399.420 ;
        RECT 2957.950 399.140 2958.230 399.420 ;
        RECT 2958.570 399.140 2958.850 399.420 ;
        RECT 2954.850 398.520 2955.130 398.800 ;
        RECT 2955.470 398.520 2955.750 398.800 ;
        RECT 2956.090 398.520 2956.370 398.800 ;
        RECT 2956.710 398.520 2956.990 398.800 ;
        RECT 2957.330 398.520 2957.610 398.800 ;
        RECT 2957.950 398.520 2958.230 398.800 ;
        RECT 2958.570 398.520 2958.850 398.800 ;
        RECT 2954.850 397.900 2955.130 398.180 ;
        RECT 2955.470 397.900 2955.750 398.180 ;
        RECT 2956.090 397.900 2956.370 398.180 ;
        RECT 2956.710 397.900 2956.990 398.180 ;
        RECT 2957.330 397.900 2957.610 398.180 ;
        RECT 2957.950 397.900 2958.230 398.180 ;
        RECT 2958.570 397.900 2958.850 398.180 ;
        RECT 2954.850 397.280 2955.130 397.560 ;
        RECT 2955.470 397.280 2955.750 397.560 ;
        RECT 2956.090 397.280 2956.370 397.560 ;
        RECT 2956.710 397.280 2956.990 397.560 ;
        RECT 2957.330 397.280 2957.610 397.560 ;
        RECT 2957.950 397.280 2958.230 397.560 ;
        RECT 2958.570 397.280 2958.850 397.560 ;
        RECT 2954.850 396.660 2955.130 396.940 ;
        RECT 2955.470 396.660 2955.750 396.940 ;
        RECT 2956.090 396.660 2956.370 396.940 ;
        RECT 2956.710 396.660 2956.990 396.940 ;
        RECT 2957.330 396.660 2957.610 396.940 ;
        RECT 2957.950 396.660 2958.230 396.940 ;
        RECT 2958.570 396.660 2958.850 396.940 ;
        RECT 2954.850 396.040 2955.130 396.320 ;
        RECT 2955.470 396.040 2955.750 396.320 ;
        RECT 2956.090 396.040 2956.370 396.320 ;
        RECT 2956.710 396.040 2956.990 396.320 ;
        RECT 2957.330 396.040 2957.610 396.320 ;
        RECT 2957.950 396.040 2958.230 396.320 ;
        RECT 2958.570 396.040 2958.850 396.320 ;
        RECT 2961.550 1528.350 2961.830 1528.630 ;
        RECT 2962.170 1528.350 2962.450 1528.630 ;
        RECT 2962.790 1528.350 2963.070 1528.630 ;
        RECT 2963.410 1528.350 2963.690 1528.630 ;
        RECT 2964.030 1528.350 2964.310 1528.630 ;
        RECT 2964.650 1528.350 2964.930 1528.630 ;
        RECT 2965.270 1528.350 2965.550 1528.630 ;
        RECT 2961.550 1527.730 2961.830 1528.010 ;
        RECT 2962.170 1527.730 2962.450 1528.010 ;
        RECT 2962.790 1527.730 2963.070 1528.010 ;
        RECT 2963.410 1527.730 2963.690 1528.010 ;
        RECT 2964.030 1527.730 2964.310 1528.010 ;
        RECT 2964.650 1527.730 2964.930 1528.010 ;
        RECT 2965.270 1527.730 2965.550 1528.010 ;
        RECT 2961.550 1527.110 2961.830 1527.390 ;
        RECT 2962.170 1527.110 2962.450 1527.390 ;
        RECT 2962.790 1527.110 2963.070 1527.390 ;
        RECT 2963.410 1527.110 2963.690 1527.390 ;
        RECT 2964.030 1527.110 2964.310 1527.390 ;
        RECT 2964.650 1527.110 2964.930 1527.390 ;
        RECT 2965.270 1527.110 2965.550 1527.390 ;
        RECT 2961.550 1526.490 2961.830 1526.770 ;
        RECT 2962.170 1526.490 2962.450 1526.770 ;
        RECT 2962.790 1526.490 2963.070 1526.770 ;
        RECT 2963.410 1526.490 2963.690 1526.770 ;
        RECT 2964.030 1526.490 2964.310 1526.770 ;
        RECT 2964.650 1526.490 2964.930 1526.770 ;
        RECT 2965.270 1526.490 2965.550 1526.770 ;
        RECT 2961.550 1525.870 2961.830 1526.150 ;
        RECT 2962.170 1525.870 2962.450 1526.150 ;
        RECT 2962.790 1525.870 2963.070 1526.150 ;
        RECT 2963.410 1525.870 2963.690 1526.150 ;
        RECT 2964.030 1525.870 2964.310 1526.150 ;
        RECT 2964.650 1525.870 2964.930 1526.150 ;
        RECT 2965.270 1525.870 2965.550 1526.150 ;
        RECT 2961.550 1525.250 2961.830 1525.530 ;
        RECT 2962.170 1525.250 2962.450 1525.530 ;
        RECT 2962.790 1525.250 2963.070 1525.530 ;
        RECT 2963.410 1525.250 2963.690 1525.530 ;
        RECT 2964.030 1525.250 2964.310 1525.530 ;
        RECT 2964.650 1525.250 2964.930 1525.530 ;
        RECT 2965.270 1525.250 2965.550 1525.530 ;
        RECT 2961.550 1524.630 2961.830 1524.910 ;
        RECT 2962.170 1524.630 2962.450 1524.910 ;
        RECT 2962.790 1524.630 2963.070 1524.910 ;
        RECT 2963.410 1524.630 2963.690 1524.910 ;
        RECT 2964.030 1524.630 2964.310 1524.910 ;
        RECT 2964.650 1524.630 2964.930 1524.910 ;
        RECT 2965.270 1524.630 2965.550 1524.910 ;
        RECT 3174.300 1535.650 3174.580 1535.930 ;
        RECT 3174.920 1535.650 3175.200 1535.930 ;
        RECT 3174.300 1535.030 3174.580 1535.310 ;
        RECT 3174.920 1535.030 3175.200 1535.310 ;
        RECT 3174.300 1534.410 3174.580 1534.690 ;
        RECT 3174.920 1534.410 3175.200 1534.690 ;
        RECT 3174.300 1533.790 3174.580 1534.070 ;
        RECT 3174.920 1533.790 3175.200 1534.070 ;
        RECT 3174.300 1533.170 3174.580 1533.450 ;
        RECT 3174.920 1533.170 3175.200 1533.450 ;
        RECT 3174.300 1532.550 3174.580 1532.830 ;
        RECT 3174.920 1532.550 3175.200 1532.830 ;
        RECT 3174.300 1531.930 3174.580 1532.210 ;
        RECT 3174.920 1531.930 3175.200 1532.210 ;
        RECT 3166.325 1528.650 3166.605 1528.930 ;
        RECT 3166.945 1528.650 3167.225 1528.930 ;
        RECT 3166.325 1528.030 3166.605 1528.310 ;
        RECT 3166.945 1528.030 3167.225 1528.310 ;
        RECT 3166.325 1527.410 3166.605 1527.690 ;
        RECT 3166.945 1527.410 3167.225 1527.690 ;
        RECT 3166.325 1526.790 3166.605 1527.070 ;
        RECT 3166.945 1526.790 3167.225 1527.070 ;
        RECT 3166.325 1526.170 3166.605 1526.450 ;
        RECT 3166.945 1526.170 3167.225 1526.450 ;
        RECT 3166.325 1525.550 3166.605 1525.830 ;
        RECT 3166.945 1525.550 3167.225 1525.830 ;
        RECT 3166.325 1524.930 3166.605 1525.210 ;
        RECT 3166.945 1524.930 3167.225 1525.210 ;
        RECT 3190.250 1535.650 3190.530 1535.930 ;
        RECT 3190.870 1535.650 3191.150 1535.930 ;
        RECT 3190.250 1535.030 3190.530 1535.310 ;
        RECT 3190.870 1535.030 3191.150 1535.310 ;
        RECT 3190.250 1534.410 3190.530 1534.690 ;
        RECT 3190.870 1534.410 3191.150 1534.690 ;
        RECT 3190.250 1533.790 3190.530 1534.070 ;
        RECT 3190.870 1533.790 3191.150 1534.070 ;
        RECT 3190.250 1533.170 3190.530 1533.450 ;
        RECT 3190.870 1533.170 3191.150 1533.450 ;
        RECT 3190.250 1532.550 3190.530 1532.830 ;
        RECT 3190.870 1532.550 3191.150 1532.830 ;
        RECT 3190.250 1531.930 3190.530 1532.210 ;
        RECT 3190.870 1531.930 3191.150 1532.210 ;
        RECT 3182.275 1528.650 3182.555 1528.930 ;
        RECT 3182.895 1528.650 3183.175 1528.930 ;
        RECT 3182.275 1528.030 3182.555 1528.310 ;
        RECT 3182.895 1528.030 3183.175 1528.310 ;
        RECT 3182.275 1527.410 3182.555 1527.690 ;
        RECT 3182.895 1527.410 3183.175 1527.690 ;
        RECT 3182.275 1526.790 3182.555 1527.070 ;
        RECT 3182.895 1526.790 3183.175 1527.070 ;
        RECT 3182.275 1526.170 3182.555 1526.450 ;
        RECT 3182.895 1526.170 3183.175 1526.450 ;
        RECT 3182.275 1525.550 3182.555 1525.830 ;
        RECT 3182.895 1525.550 3183.175 1525.830 ;
        RECT 3182.275 1524.930 3182.555 1525.210 ;
        RECT 3182.895 1524.930 3183.175 1525.210 ;
        RECT 3206.200 1535.650 3206.480 1535.930 ;
        RECT 3206.820 1535.650 3207.100 1535.930 ;
        RECT 3206.200 1535.030 3206.480 1535.310 ;
        RECT 3206.820 1535.030 3207.100 1535.310 ;
        RECT 3206.200 1534.410 3206.480 1534.690 ;
        RECT 3206.820 1534.410 3207.100 1534.690 ;
        RECT 3206.200 1533.790 3206.480 1534.070 ;
        RECT 3206.820 1533.790 3207.100 1534.070 ;
        RECT 3206.200 1533.170 3206.480 1533.450 ;
        RECT 3206.820 1533.170 3207.100 1533.450 ;
        RECT 3206.200 1532.550 3206.480 1532.830 ;
        RECT 3206.820 1532.550 3207.100 1532.830 ;
        RECT 3206.200 1531.930 3206.480 1532.210 ;
        RECT 3206.820 1531.930 3207.100 1532.210 ;
        RECT 3198.225 1528.650 3198.505 1528.930 ;
        RECT 3198.845 1528.650 3199.125 1528.930 ;
        RECT 3198.225 1528.030 3198.505 1528.310 ;
        RECT 3198.845 1528.030 3199.125 1528.310 ;
        RECT 3198.225 1527.410 3198.505 1527.690 ;
        RECT 3198.845 1527.410 3199.125 1527.690 ;
        RECT 3198.225 1526.790 3198.505 1527.070 ;
        RECT 3198.845 1526.790 3199.125 1527.070 ;
        RECT 3198.225 1526.170 3198.505 1526.450 ;
        RECT 3198.845 1526.170 3199.125 1526.450 ;
        RECT 3198.225 1525.550 3198.505 1525.830 ;
        RECT 3198.845 1525.550 3199.125 1525.830 ;
        RECT 3198.225 1524.930 3198.505 1525.210 ;
        RECT 3198.845 1524.930 3199.125 1525.210 ;
        RECT 3214.175 1528.650 3214.455 1528.930 ;
        RECT 3214.795 1528.650 3215.075 1528.930 ;
        RECT 3214.175 1528.030 3214.455 1528.310 ;
        RECT 3214.795 1528.030 3215.075 1528.310 ;
        RECT 3214.175 1527.410 3214.455 1527.690 ;
        RECT 3214.795 1527.410 3215.075 1527.690 ;
        RECT 3214.175 1526.790 3214.455 1527.070 ;
        RECT 3214.795 1526.790 3215.075 1527.070 ;
        RECT 3214.175 1526.170 3214.455 1526.450 ;
        RECT 3214.795 1526.170 3215.075 1526.450 ;
        RECT 3214.175 1525.550 3214.455 1525.830 ;
        RECT 3214.795 1525.550 3215.075 1525.830 ;
        RECT 3214.175 1524.930 3214.455 1525.210 ;
        RECT 3214.795 1524.930 3215.075 1525.210 ;
        RECT 3490.220 1566.890 3490.500 1567.170 ;
        RECT 3491.720 1566.890 3492.000 1567.170 ;
        RECT 3493.220 1566.890 3493.500 1567.170 ;
        RECT 3490.260 1535.650 3490.540 1535.930 ;
        RECT 3490.880 1535.650 3491.160 1535.930 ;
        RECT 3491.500 1535.650 3491.780 1535.930 ;
        RECT 3492.120 1535.650 3492.400 1535.930 ;
        RECT 3492.740 1535.650 3493.020 1535.930 ;
        RECT 3493.360 1535.650 3493.640 1535.930 ;
        RECT 3493.980 1535.650 3494.260 1535.930 ;
        RECT 3490.260 1535.030 3490.540 1535.310 ;
        RECT 3490.880 1535.030 3491.160 1535.310 ;
        RECT 3491.500 1535.030 3491.780 1535.310 ;
        RECT 3492.120 1535.030 3492.400 1535.310 ;
        RECT 3492.740 1535.030 3493.020 1535.310 ;
        RECT 3493.360 1535.030 3493.640 1535.310 ;
        RECT 3493.980 1535.030 3494.260 1535.310 ;
        RECT 3490.260 1534.410 3490.540 1534.690 ;
        RECT 3490.880 1534.410 3491.160 1534.690 ;
        RECT 3491.500 1534.410 3491.780 1534.690 ;
        RECT 3492.120 1534.410 3492.400 1534.690 ;
        RECT 3492.740 1534.410 3493.020 1534.690 ;
        RECT 3493.360 1534.410 3493.640 1534.690 ;
        RECT 3493.980 1534.410 3494.260 1534.690 ;
        RECT 3490.260 1533.790 3490.540 1534.070 ;
        RECT 3490.880 1533.790 3491.160 1534.070 ;
        RECT 3491.500 1533.790 3491.780 1534.070 ;
        RECT 3492.120 1533.790 3492.400 1534.070 ;
        RECT 3492.740 1533.790 3493.020 1534.070 ;
        RECT 3493.360 1533.790 3493.640 1534.070 ;
        RECT 3493.980 1533.790 3494.260 1534.070 ;
        RECT 3490.260 1533.170 3490.540 1533.450 ;
        RECT 3490.880 1533.170 3491.160 1533.450 ;
        RECT 3491.500 1533.170 3491.780 1533.450 ;
        RECT 3492.120 1533.170 3492.400 1533.450 ;
        RECT 3492.740 1533.170 3493.020 1533.450 ;
        RECT 3493.360 1533.170 3493.640 1533.450 ;
        RECT 3493.980 1533.170 3494.260 1533.450 ;
        RECT 3490.260 1532.550 3490.540 1532.830 ;
        RECT 3490.880 1532.550 3491.160 1532.830 ;
        RECT 3491.500 1532.550 3491.780 1532.830 ;
        RECT 3492.120 1532.550 3492.400 1532.830 ;
        RECT 3492.740 1532.550 3493.020 1532.830 ;
        RECT 3493.360 1532.550 3493.640 1532.830 ;
        RECT 3493.980 1532.550 3494.260 1532.830 ;
        RECT 3490.260 1531.930 3490.540 1532.210 ;
        RECT 3490.880 1531.930 3491.160 1532.210 ;
        RECT 3491.500 1531.930 3491.780 1532.210 ;
        RECT 3492.120 1531.930 3492.400 1532.210 ;
        RECT 3492.740 1531.930 3493.020 1532.210 ;
        RECT 3493.360 1531.930 3493.640 1532.210 ;
        RECT 3493.980 1531.930 3494.260 1532.210 ;
        RECT 2961.850 1409.580 2962.130 1409.860 ;
        RECT 2962.470 1409.580 2962.750 1409.860 ;
        RECT 2963.090 1409.580 2963.370 1409.860 ;
        RECT 2963.710 1409.580 2963.990 1409.860 ;
        RECT 2964.330 1409.580 2964.610 1409.860 ;
        RECT 2964.950 1409.580 2965.230 1409.860 ;
        RECT 2965.570 1409.580 2965.850 1409.860 ;
        RECT 2961.850 1408.960 2962.130 1409.240 ;
        RECT 2962.470 1408.960 2962.750 1409.240 ;
        RECT 2963.090 1408.960 2963.370 1409.240 ;
        RECT 2963.710 1408.960 2963.990 1409.240 ;
        RECT 2964.330 1408.960 2964.610 1409.240 ;
        RECT 2964.950 1408.960 2965.230 1409.240 ;
        RECT 2965.570 1408.960 2965.850 1409.240 ;
        RECT 2961.850 1408.340 2962.130 1408.620 ;
        RECT 2962.470 1408.340 2962.750 1408.620 ;
        RECT 2963.090 1408.340 2963.370 1408.620 ;
        RECT 2963.710 1408.340 2963.990 1408.620 ;
        RECT 2964.330 1408.340 2964.610 1408.620 ;
        RECT 2964.950 1408.340 2965.230 1408.620 ;
        RECT 2965.570 1408.340 2965.850 1408.620 ;
        RECT 2961.850 1407.720 2962.130 1408.000 ;
        RECT 2962.470 1407.720 2962.750 1408.000 ;
        RECT 2963.090 1407.720 2963.370 1408.000 ;
        RECT 2963.710 1407.720 2963.990 1408.000 ;
        RECT 2964.330 1407.720 2964.610 1408.000 ;
        RECT 2964.950 1407.720 2965.230 1408.000 ;
        RECT 2965.570 1407.720 2965.850 1408.000 ;
        RECT 2961.850 1407.100 2962.130 1407.380 ;
        RECT 2962.470 1407.100 2962.750 1407.380 ;
        RECT 2963.090 1407.100 2963.370 1407.380 ;
        RECT 2963.710 1407.100 2963.990 1407.380 ;
        RECT 2964.330 1407.100 2964.610 1407.380 ;
        RECT 2964.950 1407.100 2965.230 1407.380 ;
        RECT 2965.570 1407.100 2965.850 1407.380 ;
        RECT 2961.850 1406.480 2962.130 1406.760 ;
        RECT 2962.470 1406.480 2962.750 1406.760 ;
        RECT 2963.090 1406.480 2963.370 1406.760 ;
        RECT 2963.710 1406.480 2963.990 1406.760 ;
        RECT 2964.330 1406.480 2964.610 1406.760 ;
        RECT 2964.950 1406.480 2965.230 1406.760 ;
        RECT 2965.570 1406.480 2965.850 1406.760 ;
        RECT 2961.850 1405.860 2962.130 1406.140 ;
        RECT 2962.470 1405.860 2962.750 1406.140 ;
        RECT 2963.090 1405.860 2963.370 1406.140 ;
        RECT 2963.710 1405.860 2963.990 1406.140 ;
        RECT 2964.330 1405.860 2964.610 1406.140 ;
        RECT 2964.950 1405.860 2965.230 1406.140 ;
        RECT 2965.570 1405.860 2965.850 1406.140 ;
        RECT 2961.850 1341.580 2962.130 1341.860 ;
        RECT 2962.470 1341.580 2962.750 1341.860 ;
        RECT 2963.090 1341.580 2963.370 1341.860 ;
        RECT 2963.710 1341.580 2963.990 1341.860 ;
        RECT 2964.330 1341.580 2964.610 1341.860 ;
        RECT 2964.950 1341.580 2965.230 1341.860 ;
        RECT 2965.570 1341.580 2965.850 1341.860 ;
        RECT 2961.850 1340.960 2962.130 1341.240 ;
        RECT 2962.470 1340.960 2962.750 1341.240 ;
        RECT 2963.090 1340.960 2963.370 1341.240 ;
        RECT 2963.710 1340.960 2963.990 1341.240 ;
        RECT 2964.330 1340.960 2964.610 1341.240 ;
        RECT 2964.950 1340.960 2965.230 1341.240 ;
        RECT 2965.570 1340.960 2965.850 1341.240 ;
        RECT 2961.850 1211.580 2962.130 1211.860 ;
        RECT 2962.470 1211.580 2962.750 1211.860 ;
        RECT 2963.090 1211.580 2963.370 1211.860 ;
        RECT 2963.710 1211.580 2963.990 1211.860 ;
        RECT 2964.330 1211.580 2964.610 1211.860 ;
        RECT 2964.950 1211.580 2965.230 1211.860 ;
        RECT 2965.570 1211.580 2965.850 1211.860 ;
        RECT 2961.850 1210.960 2962.130 1211.240 ;
        RECT 2962.470 1210.960 2962.750 1211.240 ;
        RECT 2963.090 1210.960 2963.370 1211.240 ;
        RECT 2963.710 1210.960 2963.990 1211.240 ;
        RECT 2964.330 1210.960 2964.610 1211.240 ;
        RECT 2964.950 1210.960 2965.230 1211.240 ;
        RECT 2965.570 1210.960 2965.850 1211.240 ;
        RECT 2961.850 1081.580 2962.130 1081.860 ;
        RECT 2962.470 1081.580 2962.750 1081.860 ;
        RECT 2963.090 1081.580 2963.370 1081.860 ;
        RECT 2963.710 1081.580 2963.990 1081.860 ;
        RECT 2964.330 1081.580 2964.610 1081.860 ;
        RECT 2964.950 1081.580 2965.230 1081.860 ;
        RECT 2965.570 1081.580 2965.850 1081.860 ;
        RECT 2961.850 1080.960 2962.130 1081.240 ;
        RECT 2962.470 1080.960 2962.750 1081.240 ;
        RECT 2963.090 1080.960 2963.370 1081.240 ;
        RECT 2963.710 1080.960 2963.990 1081.240 ;
        RECT 2964.330 1080.960 2964.610 1081.240 ;
        RECT 2964.950 1080.960 2965.230 1081.240 ;
        RECT 2965.570 1080.960 2965.850 1081.240 ;
        RECT 2961.850 951.580 2962.130 951.860 ;
        RECT 2962.470 951.580 2962.750 951.860 ;
        RECT 2963.090 951.580 2963.370 951.860 ;
        RECT 2963.710 951.580 2963.990 951.860 ;
        RECT 2964.330 951.580 2964.610 951.860 ;
        RECT 2964.950 951.580 2965.230 951.860 ;
        RECT 2965.570 951.580 2965.850 951.860 ;
        RECT 2961.850 950.960 2962.130 951.240 ;
        RECT 2962.470 950.960 2962.750 951.240 ;
        RECT 2963.090 950.960 2963.370 951.240 ;
        RECT 2963.710 950.960 2963.990 951.240 ;
        RECT 2964.330 950.960 2964.610 951.240 ;
        RECT 2964.950 950.960 2965.230 951.240 ;
        RECT 2965.570 950.960 2965.850 951.240 ;
        RECT 2961.850 821.580 2962.130 821.860 ;
        RECT 2962.470 821.580 2962.750 821.860 ;
        RECT 2963.090 821.580 2963.370 821.860 ;
        RECT 2963.710 821.580 2963.990 821.860 ;
        RECT 2964.330 821.580 2964.610 821.860 ;
        RECT 2964.950 821.580 2965.230 821.860 ;
        RECT 2965.570 821.580 2965.850 821.860 ;
        RECT 2961.850 820.960 2962.130 821.240 ;
        RECT 2962.470 820.960 2962.750 821.240 ;
        RECT 2963.090 820.960 2963.370 821.240 ;
        RECT 2963.710 820.960 2963.990 821.240 ;
        RECT 2964.330 820.960 2964.610 821.240 ;
        RECT 2964.950 820.960 2965.230 821.240 ;
        RECT 2965.570 820.960 2965.850 821.240 ;
        RECT 2961.850 691.580 2962.130 691.860 ;
        RECT 2962.470 691.580 2962.750 691.860 ;
        RECT 2963.090 691.580 2963.370 691.860 ;
        RECT 2963.710 691.580 2963.990 691.860 ;
        RECT 2964.330 691.580 2964.610 691.860 ;
        RECT 2964.950 691.580 2965.230 691.860 ;
        RECT 2965.570 691.580 2965.850 691.860 ;
        RECT 2961.850 690.960 2962.130 691.240 ;
        RECT 2962.470 690.960 2962.750 691.240 ;
        RECT 2963.090 690.960 2963.370 691.240 ;
        RECT 2963.710 690.960 2963.990 691.240 ;
        RECT 2964.330 690.960 2964.610 691.240 ;
        RECT 2964.950 690.960 2965.230 691.240 ;
        RECT 2965.570 690.960 2965.850 691.240 ;
        RECT 2961.795 608.175 2962.075 608.455 ;
        RECT 2963.295 608.175 2963.575 608.455 ;
        RECT 2964.795 608.175 2965.075 608.455 ;
        RECT 2961.795 592.635 2962.075 592.915 ;
        RECT 2963.295 592.635 2963.575 592.915 ;
        RECT 2964.795 592.635 2965.075 592.915 ;
        RECT 2961.795 577.095 2962.075 577.375 ;
        RECT 2963.295 577.095 2963.575 577.375 ;
        RECT 2964.795 577.095 2965.075 577.375 ;
        RECT 2961.850 561.580 2962.130 561.860 ;
        RECT 2962.470 561.580 2962.750 561.860 ;
        RECT 2963.090 561.580 2963.370 561.860 ;
        RECT 2963.710 561.580 2963.990 561.860 ;
        RECT 2964.330 561.580 2964.610 561.860 ;
        RECT 2964.950 561.580 2965.230 561.860 ;
        RECT 2965.570 561.580 2965.850 561.860 ;
        RECT 2961.850 560.960 2962.130 561.240 ;
        RECT 2962.470 560.960 2962.750 561.240 ;
        RECT 2963.090 560.960 2963.370 561.240 ;
        RECT 2963.710 560.960 2963.990 561.240 ;
        RECT 2964.330 560.960 2964.610 561.240 ;
        RECT 2964.950 560.960 2965.230 561.240 ;
        RECT 2965.570 560.960 2965.850 561.240 ;
        RECT 3490.300 1449.760 3490.580 1450.040 ;
        RECT 3491.800 1449.760 3492.080 1450.040 ;
        RECT 3493.300 1449.760 3493.580 1450.040 ;
        RECT 3490.220 1419.345 3490.500 1419.625 ;
        RECT 3491.720 1419.345 3492.000 1419.625 ;
        RECT 3493.220 1419.345 3493.500 1419.625 ;
        RECT 3490.220 1386.890 3490.500 1387.170 ;
        RECT 3491.720 1386.890 3492.000 1387.170 ;
        RECT 3493.220 1386.890 3493.500 1387.170 ;
        RECT 3490.220 1351.890 3490.500 1352.170 ;
        RECT 3491.720 1351.890 3492.000 1352.170 ;
        RECT 3493.220 1351.890 3493.500 1352.170 ;
        RECT 3490.220 1316.890 3490.500 1317.170 ;
        RECT 3491.720 1316.890 3492.000 1317.170 ;
        RECT 3493.220 1316.890 3493.500 1317.170 ;
        RECT 3490.220 1266.165 3490.500 1266.445 ;
        RECT 3491.720 1266.165 3492.000 1266.445 ;
        RECT 3493.220 1266.165 3493.500 1266.445 ;
        RECT 3490.300 1234.760 3490.580 1235.040 ;
        RECT 3491.800 1234.760 3492.080 1235.040 ;
        RECT 3493.300 1234.760 3493.580 1235.040 ;
        RECT 3490.220 1171.890 3490.500 1172.170 ;
        RECT 3491.720 1171.890 3492.000 1172.170 ;
        RECT 3493.220 1171.890 3493.500 1172.170 ;
        RECT 3490.220 1136.890 3490.500 1137.170 ;
        RECT 3491.720 1136.890 3492.000 1137.170 ;
        RECT 3493.220 1136.890 3493.500 1137.170 ;
        RECT 3490.220 1112.985 3490.500 1113.265 ;
        RECT 3491.720 1112.985 3492.000 1113.265 ;
        RECT 3493.220 1112.985 3493.500 1113.265 ;
        RECT 3490.220 1101.890 3490.500 1102.170 ;
        RECT 3491.720 1101.890 3492.000 1102.170 ;
        RECT 3493.220 1101.890 3493.500 1102.170 ;
        RECT 3490.300 1019.760 3490.580 1020.040 ;
        RECT 3491.800 1019.760 3492.080 1020.040 ;
        RECT 3493.300 1019.760 3493.580 1020.040 ;
        RECT 3490.220 959.805 3490.500 960.085 ;
        RECT 3491.720 959.805 3492.000 960.085 ;
        RECT 3493.220 959.805 3493.500 960.085 ;
        RECT 3490.220 956.890 3490.500 957.170 ;
        RECT 3491.720 956.890 3492.000 957.170 ;
        RECT 3493.220 956.890 3493.500 957.170 ;
        RECT 3490.220 921.890 3490.500 922.170 ;
        RECT 3491.720 921.890 3492.000 922.170 ;
        RECT 3493.220 921.890 3493.500 922.170 ;
        RECT 3490.220 886.890 3490.500 887.170 ;
        RECT 3491.720 886.890 3492.000 887.170 ;
        RECT 3493.220 886.890 3493.500 887.170 ;
        RECT 3490.220 806.625 3490.500 806.905 ;
        RECT 3491.720 806.625 3492.000 806.905 ;
        RECT 3493.220 806.625 3493.500 806.905 ;
        RECT 3490.300 804.760 3490.580 805.040 ;
        RECT 3491.800 804.760 3492.080 805.040 ;
        RECT 3493.300 804.760 3493.580 805.040 ;
        RECT 3490.220 741.890 3490.500 742.170 ;
        RECT 3491.720 741.890 3492.000 742.170 ;
        RECT 3493.220 741.890 3493.500 742.170 ;
        RECT 3490.220 706.890 3490.500 707.170 ;
        RECT 3491.720 706.890 3492.000 707.170 ;
        RECT 3493.220 706.890 3493.500 707.170 ;
        RECT 3490.220 671.810 3490.500 672.090 ;
        RECT 3491.720 671.810 3492.000 672.090 ;
        RECT 3493.220 671.810 3493.500 672.090 ;
        RECT 3490.220 664.735 3490.500 665.015 ;
        RECT 3491.720 664.735 3492.000 665.015 ;
        RECT 3493.220 664.735 3493.500 665.015 ;
        RECT 3490.300 589.760 3490.580 590.040 ;
        RECT 3491.800 589.760 3492.080 590.040 ;
        RECT 3493.300 589.760 3493.580 590.040 ;
        RECT 3490.220 526.890 3490.500 527.170 ;
        RECT 3491.720 526.890 3492.000 527.170 ;
        RECT 3493.220 526.890 3493.500 527.170 ;
        RECT 2961.850 431.580 2962.130 431.860 ;
        RECT 2962.470 431.580 2962.750 431.860 ;
        RECT 2963.090 431.580 2963.370 431.860 ;
        RECT 2963.710 431.580 2963.990 431.860 ;
        RECT 2964.330 431.580 2964.610 431.860 ;
        RECT 2964.950 431.580 2965.230 431.860 ;
        RECT 2965.570 431.580 2965.850 431.860 ;
        RECT 2961.850 430.960 2962.130 431.240 ;
        RECT 2962.470 430.960 2962.750 431.240 ;
        RECT 2963.090 430.960 2963.370 431.240 ;
        RECT 2963.710 430.960 2963.990 431.240 ;
        RECT 2964.330 430.960 2964.610 431.240 ;
        RECT 2964.950 430.960 2965.230 431.240 ;
        RECT 2965.570 430.960 2965.850 431.240 ;
        RECT 2771.470 392.760 2771.750 393.040 ;
        RECT 2772.090 392.760 2772.370 393.040 ;
        RECT 2771.470 392.140 2771.750 392.420 ;
        RECT 2772.090 392.140 2772.370 392.420 ;
        RECT 2771.470 391.520 2771.750 391.800 ;
        RECT 2772.090 391.520 2772.370 391.800 ;
        RECT 2771.470 390.900 2771.750 391.180 ;
        RECT 2772.090 390.900 2772.370 391.180 ;
        RECT 2771.470 390.280 2771.750 390.560 ;
        RECT 2772.090 390.280 2772.370 390.560 ;
        RECT 2771.470 389.660 2771.750 389.940 ;
        RECT 2772.090 389.660 2772.370 389.940 ;
        RECT 2771.470 389.040 2771.750 389.320 ;
        RECT 2772.090 389.040 2772.370 389.320 ;
        RECT 3340.300 497.265 3340.580 497.545 ;
        RECT 3340.920 497.265 3341.200 497.545 ;
        RECT 3341.540 497.265 3341.820 497.545 ;
        RECT 3342.160 497.265 3342.440 497.545 ;
        RECT 3342.780 497.265 3343.060 497.545 ;
        RECT 3343.400 497.265 3343.680 497.545 ;
        RECT 3340.300 496.645 3340.580 496.925 ;
        RECT 3340.920 496.645 3341.200 496.925 ;
        RECT 3341.540 496.645 3341.820 496.925 ;
        RECT 3342.160 496.645 3342.440 496.925 ;
        RECT 3342.780 496.645 3343.060 496.925 ;
        RECT 3343.400 496.645 3343.680 496.925 ;
        RECT 3340.300 496.025 3340.580 496.305 ;
        RECT 3340.920 496.025 3341.200 496.305 ;
        RECT 3341.540 496.025 3341.820 496.305 ;
        RECT 3342.160 496.025 3342.440 496.305 ;
        RECT 3342.780 496.025 3343.060 496.305 ;
        RECT 3343.400 496.025 3343.680 496.305 ;
        RECT 3340.300 495.405 3340.580 495.685 ;
        RECT 3340.920 495.405 3341.200 495.685 ;
        RECT 3341.540 495.405 3341.820 495.685 ;
        RECT 3342.160 495.405 3342.440 495.685 ;
        RECT 3342.780 495.405 3343.060 495.685 ;
        RECT 3343.400 495.405 3343.680 495.685 ;
        RECT 3340.300 494.785 3340.580 495.065 ;
        RECT 3340.920 494.785 3341.200 495.065 ;
        RECT 3341.540 494.785 3341.820 495.065 ;
        RECT 3342.160 494.785 3342.440 495.065 ;
        RECT 3342.780 494.785 3343.060 495.065 ;
        RECT 3343.400 494.785 3343.680 495.065 ;
        RECT 3340.300 494.165 3340.580 494.445 ;
        RECT 3340.920 494.165 3341.200 494.445 ;
        RECT 3341.540 494.165 3341.820 494.445 ;
        RECT 3342.160 494.165 3342.440 494.445 ;
        RECT 3342.780 494.165 3343.060 494.445 ;
        RECT 3343.400 494.165 3343.680 494.445 ;
        RECT 3340.300 493.545 3340.580 493.825 ;
        RECT 3340.920 493.545 3341.200 493.825 ;
        RECT 3341.540 493.545 3341.820 493.825 ;
        RECT 3342.160 493.545 3342.440 493.825 ;
        RECT 3342.780 493.545 3343.060 493.825 ;
        RECT 3343.400 493.545 3343.680 493.825 ;
        RECT 2961.850 392.760 2962.130 393.040 ;
        RECT 2962.470 392.760 2962.750 393.040 ;
        RECT 2963.090 392.760 2963.370 393.040 ;
        RECT 2963.710 392.760 2963.990 393.040 ;
        RECT 2964.330 392.760 2964.610 393.040 ;
        RECT 2964.950 392.760 2965.230 393.040 ;
        RECT 2965.570 392.760 2965.850 393.040 ;
        RECT 2961.850 392.140 2962.130 392.420 ;
        RECT 2962.470 392.140 2962.750 392.420 ;
        RECT 2963.090 392.140 2963.370 392.420 ;
        RECT 2963.710 392.140 2963.990 392.420 ;
        RECT 2964.330 392.140 2964.610 392.420 ;
        RECT 2964.950 392.140 2965.230 392.420 ;
        RECT 2965.570 392.140 2965.850 392.420 ;
        RECT 2961.850 391.520 2962.130 391.800 ;
        RECT 2962.470 391.520 2962.750 391.800 ;
        RECT 2963.090 391.520 2963.370 391.800 ;
        RECT 2963.710 391.520 2963.990 391.800 ;
        RECT 2964.330 391.520 2964.610 391.800 ;
        RECT 2964.950 391.520 2965.230 391.800 ;
        RECT 2965.570 391.520 2965.850 391.800 ;
        RECT 2961.850 390.900 2962.130 391.180 ;
        RECT 2962.470 390.900 2962.750 391.180 ;
        RECT 2963.090 390.900 2963.370 391.180 ;
        RECT 2963.710 390.900 2963.990 391.180 ;
        RECT 2964.330 390.900 2964.610 391.180 ;
        RECT 2964.950 390.900 2965.230 391.180 ;
        RECT 2965.570 390.900 2965.850 391.180 ;
        RECT 2961.850 390.280 2962.130 390.560 ;
        RECT 2962.470 390.280 2962.750 390.560 ;
        RECT 2963.090 390.280 2963.370 390.560 ;
        RECT 2963.710 390.280 2963.990 390.560 ;
        RECT 2964.330 390.280 2964.610 390.560 ;
        RECT 2964.950 390.280 2965.230 390.560 ;
        RECT 2965.570 390.280 2965.850 390.560 ;
        RECT 2961.850 389.660 2962.130 389.940 ;
        RECT 2962.470 389.660 2962.750 389.940 ;
        RECT 2963.090 389.660 2963.370 389.940 ;
        RECT 2963.710 389.660 2963.990 389.940 ;
        RECT 2964.330 389.660 2964.610 389.940 ;
        RECT 2964.950 389.660 2965.230 389.940 ;
        RECT 2965.570 389.660 2965.850 389.940 ;
        RECT 2961.850 389.040 2962.130 389.320 ;
        RECT 2962.470 389.040 2962.750 389.320 ;
        RECT 2963.090 389.040 2963.370 389.320 ;
        RECT 2963.710 389.040 2963.990 389.320 ;
        RECT 2964.330 389.040 2964.610 389.320 ;
        RECT 2964.950 389.040 2965.230 389.320 ;
        RECT 2965.570 389.040 2965.850 389.320 ;
        RECT 3011.650 399.760 3011.930 400.040 ;
        RECT 3012.270 399.760 3012.550 400.040 ;
        RECT 3012.890 399.760 3013.170 400.040 ;
        RECT 3013.510 399.760 3013.790 400.040 ;
        RECT 3014.130 399.760 3014.410 400.040 ;
        RECT 3014.750 399.760 3015.030 400.040 ;
        RECT 3015.370 399.760 3015.650 400.040 ;
        RECT 3015.990 399.760 3016.270 400.040 ;
        RECT 3016.610 399.760 3016.890 400.040 ;
        RECT 3017.230 399.760 3017.510 400.040 ;
        RECT 3017.850 399.760 3018.130 400.040 ;
        RECT 3018.470 399.760 3018.750 400.040 ;
        RECT 3019.090 399.760 3019.370 400.040 ;
        RECT 3019.710 399.760 3019.990 400.040 ;
        RECT 3020.330 399.760 3020.610 400.040 ;
        RECT 3011.650 399.140 3011.930 399.420 ;
        RECT 3012.270 399.140 3012.550 399.420 ;
        RECT 3012.890 399.140 3013.170 399.420 ;
        RECT 3013.510 399.140 3013.790 399.420 ;
        RECT 3014.130 399.140 3014.410 399.420 ;
        RECT 3014.750 399.140 3015.030 399.420 ;
        RECT 3015.370 399.140 3015.650 399.420 ;
        RECT 3015.990 399.140 3016.270 399.420 ;
        RECT 3016.610 399.140 3016.890 399.420 ;
        RECT 3017.230 399.140 3017.510 399.420 ;
        RECT 3017.850 399.140 3018.130 399.420 ;
        RECT 3018.470 399.140 3018.750 399.420 ;
        RECT 3019.090 399.140 3019.370 399.420 ;
        RECT 3019.710 399.140 3019.990 399.420 ;
        RECT 3020.330 399.140 3020.610 399.420 ;
        RECT 3011.650 398.520 3011.930 398.800 ;
        RECT 3012.270 398.520 3012.550 398.800 ;
        RECT 3012.890 398.520 3013.170 398.800 ;
        RECT 3013.510 398.520 3013.790 398.800 ;
        RECT 3014.130 398.520 3014.410 398.800 ;
        RECT 3014.750 398.520 3015.030 398.800 ;
        RECT 3015.370 398.520 3015.650 398.800 ;
        RECT 3015.990 398.520 3016.270 398.800 ;
        RECT 3016.610 398.520 3016.890 398.800 ;
        RECT 3017.230 398.520 3017.510 398.800 ;
        RECT 3017.850 398.520 3018.130 398.800 ;
        RECT 3018.470 398.520 3018.750 398.800 ;
        RECT 3019.090 398.520 3019.370 398.800 ;
        RECT 3019.710 398.520 3019.990 398.800 ;
        RECT 3020.330 398.520 3020.610 398.800 ;
        RECT 3011.650 397.900 3011.930 398.180 ;
        RECT 3012.270 397.900 3012.550 398.180 ;
        RECT 3012.890 397.900 3013.170 398.180 ;
        RECT 3013.510 397.900 3013.790 398.180 ;
        RECT 3014.130 397.900 3014.410 398.180 ;
        RECT 3014.750 397.900 3015.030 398.180 ;
        RECT 3015.370 397.900 3015.650 398.180 ;
        RECT 3015.990 397.900 3016.270 398.180 ;
        RECT 3016.610 397.900 3016.890 398.180 ;
        RECT 3017.230 397.900 3017.510 398.180 ;
        RECT 3017.850 397.900 3018.130 398.180 ;
        RECT 3018.470 397.900 3018.750 398.180 ;
        RECT 3019.090 397.900 3019.370 398.180 ;
        RECT 3019.710 397.900 3019.990 398.180 ;
        RECT 3020.330 397.900 3020.610 398.180 ;
        RECT 3011.650 397.280 3011.930 397.560 ;
        RECT 3012.270 397.280 3012.550 397.560 ;
        RECT 3012.890 397.280 3013.170 397.560 ;
        RECT 3013.510 397.280 3013.790 397.560 ;
        RECT 3014.130 397.280 3014.410 397.560 ;
        RECT 3014.750 397.280 3015.030 397.560 ;
        RECT 3015.370 397.280 3015.650 397.560 ;
        RECT 3015.990 397.280 3016.270 397.560 ;
        RECT 3016.610 397.280 3016.890 397.560 ;
        RECT 3017.230 397.280 3017.510 397.560 ;
        RECT 3017.850 397.280 3018.130 397.560 ;
        RECT 3018.470 397.280 3018.750 397.560 ;
        RECT 3019.090 397.280 3019.370 397.560 ;
        RECT 3019.710 397.280 3019.990 397.560 ;
        RECT 3020.330 397.280 3020.610 397.560 ;
        RECT 3011.650 396.660 3011.930 396.940 ;
        RECT 3012.270 396.660 3012.550 396.940 ;
        RECT 3012.890 396.660 3013.170 396.940 ;
        RECT 3013.510 396.660 3013.790 396.940 ;
        RECT 3014.130 396.660 3014.410 396.940 ;
        RECT 3014.750 396.660 3015.030 396.940 ;
        RECT 3015.370 396.660 3015.650 396.940 ;
        RECT 3015.990 396.660 3016.270 396.940 ;
        RECT 3016.610 396.660 3016.890 396.940 ;
        RECT 3017.230 396.660 3017.510 396.940 ;
        RECT 3017.850 396.660 3018.130 396.940 ;
        RECT 3018.470 396.660 3018.750 396.940 ;
        RECT 3019.090 396.660 3019.370 396.940 ;
        RECT 3019.710 396.660 3019.990 396.940 ;
        RECT 3020.330 396.660 3020.610 396.940 ;
        RECT 3011.650 396.040 3011.930 396.320 ;
        RECT 3012.270 396.040 3012.550 396.320 ;
        RECT 3012.890 396.040 3013.170 396.320 ;
        RECT 3013.510 396.040 3013.790 396.320 ;
        RECT 3014.130 396.040 3014.410 396.320 ;
        RECT 3014.750 396.040 3015.030 396.320 ;
        RECT 3015.370 396.040 3015.650 396.320 ;
        RECT 3015.990 396.040 3016.270 396.320 ;
        RECT 3016.610 396.040 3016.890 396.320 ;
        RECT 3017.230 396.040 3017.510 396.320 ;
        RECT 3017.850 396.040 3018.130 396.320 ;
        RECT 3018.470 396.040 3018.750 396.320 ;
        RECT 3019.090 396.040 3019.370 396.320 ;
        RECT 3019.710 396.040 3019.990 396.320 ;
        RECT 3020.330 396.040 3020.610 396.320 ;
        RECT 3024.050 399.760 3024.330 400.040 ;
        RECT 3024.670 399.760 3024.950 400.040 ;
        RECT 3025.290 399.760 3025.570 400.040 ;
        RECT 3025.910 399.760 3026.190 400.040 ;
        RECT 3026.530 399.760 3026.810 400.040 ;
        RECT 3027.150 399.760 3027.430 400.040 ;
        RECT 3027.770 399.760 3028.050 400.040 ;
        RECT 3028.390 399.760 3028.670 400.040 ;
        RECT 3029.010 399.760 3029.290 400.040 ;
        RECT 3029.630 399.760 3029.910 400.040 ;
        RECT 3030.250 399.760 3030.530 400.040 ;
        RECT 3030.870 399.760 3031.150 400.040 ;
        RECT 3031.490 399.760 3031.770 400.040 ;
        RECT 3032.110 399.760 3032.390 400.040 ;
        RECT 3032.730 399.760 3033.010 400.040 ;
        RECT 3033.350 399.760 3033.630 400.040 ;
        RECT 3024.050 399.140 3024.330 399.420 ;
        RECT 3024.670 399.140 3024.950 399.420 ;
        RECT 3025.290 399.140 3025.570 399.420 ;
        RECT 3025.910 399.140 3026.190 399.420 ;
        RECT 3026.530 399.140 3026.810 399.420 ;
        RECT 3027.150 399.140 3027.430 399.420 ;
        RECT 3027.770 399.140 3028.050 399.420 ;
        RECT 3028.390 399.140 3028.670 399.420 ;
        RECT 3029.010 399.140 3029.290 399.420 ;
        RECT 3029.630 399.140 3029.910 399.420 ;
        RECT 3030.250 399.140 3030.530 399.420 ;
        RECT 3030.870 399.140 3031.150 399.420 ;
        RECT 3031.490 399.140 3031.770 399.420 ;
        RECT 3032.110 399.140 3032.390 399.420 ;
        RECT 3032.730 399.140 3033.010 399.420 ;
        RECT 3033.350 399.140 3033.630 399.420 ;
        RECT 3024.050 398.520 3024.330 398.800 ;
        RECT 3024.670 398.520 3024.950 398.800 ;
        RECT 3025.290 398.520 3025.570 398.800 ;
        RECT 3025.910 398.520 3026.190 398.800 ;
        RECT 3026.530 398.520 3026.810 398.800 ;
        RECT 3027.150 398.520 3027.430 398.800 ;
        RECT 3027.770 398.520 3028.050 398.800 ;
        RECT 3028.390 398.520 3028.670 398.800 ;
        RECT 3029.010 398.520 3029.290 398.800 ;
        RECT 3029.630 398.520 3029.910 398.800 ;
        RECT 3030.250 398.520 3030.530 398.800 ;
        RECT 3030.870 398.520 3031.150 398.800 ;
        RECT 3031.490 398.520 3031.770 398.800 ;
        RECT 3032.110 398.520 3032.390 398.800 ;
        RECT 3032.730 398.520 3033.010 398.800 ;
        RECT 3033.350 398.520 3033.630 398.800 ;
        RECT 3024.050 397.900 3024.330 398.180 ;
        RECT 3024.670 397.900 3024.950 398.180 ;
        RECT 3025.290 397.900 3025.570 398.180 ;
        RECT 3025.910 397.900 3026.190 398.180 ;
        RECT 3026.530 397.900 3026.810 398.180 ;
        RECT 3027.150 397.900 3027.430 398.180 ;
        RECT 3027.770 397.900 3028.050 398.180 ;
        RECT 3028.390 397.900 3028.670 398.180 ;
        RECT 3029.010 397.900 3029.290 398.180 ;
        RECT 3029.630 397.900 3029.910 398.180 ;
        RECT 3030.250 397.900 3030.530 398.180 ;
        RECT 3030.870 397.900 3031.150 398.180 ;
        RECT 3031.490 397.900 3031.770 398.180 ;
        RECT 3032.110 397.900 3032.390 398.180 ;
        RECT 3032.730 397.900 3033.010 398.180 ;
        RECT 3033.350 397.900 3033.630 398.180 ;
        RECT 3024.050 397.280 3024.330 397.560 ;
        RECT 3024.670 397.280 3024.950 397.560 ;
        RECT 3025.290 397.280 3025.570 397.560 ;
        RECT 3025.910 397.280 3026.190 397.560 ;
        RECT 3026.530 397.280 3026.810 397.560 ;
        RECT 3027.150 397.280 3027.430 397.560 ;
        RECT 3027.770 397.280 3028.050 397.560 ;
        RECT 3028.390 397.280 3028.670 397.560 ;
        RECT 3029.010 397.280 3029.290 397.560 ;
        RECT 3029.630 397.280 3029.910 397.560 ;
        RECT 3030.250 397.280 3030.530 397.560 ;
        RECT 3030.870 397.280 3031.150 397.560 ;
        RECT 3031.490 397.280 3031.770 397.560 ;
        RECT 3032.110 397.280 3032.390 397.560 ;
        RECT 3032.730 397.280 3033.010 397.560 ;
        RECT 3033.350 397.280 3033.630 397.560 ;
        RECT 3024.050 396.660 3024.330 396.940 ;
        RECT 3024.670 396.660 3024.950 396.940 ;
        RECT 3025.290 396.660 3025.570 396.940 ;
        RECT 3025.910 396.660 3026.190 396.940 ;
        RECT 3026.530 396.660 3026.810 396.940 ;
        RECT 3027.150 396.660 3027.430 396.940 ;
        RECT 3027.770 396.660 3028.050 396.940 ;
        RECT 3028.390 396.660 3028.670 396.940 ;
        RECT 3029.010 396.660 3029.290 396.940 ;
        RECT 3029.630 396.660 3029.910 396.940 ;
        RECT 3030.250 396.660 3030.530 396.940 ;
        RECT 3030.870 396.660 3031.150 396.940 ;
        RECT 3031.490 396.660 3031.770 396.940 ;
        RECT 3032.110 396.660 3032.390 396.940 ;
        RECT 3032.730 396.660 3033.010 396.940 ;
        RECT 3033.350 396.660 3033.630 396.940 ;
        RECT 3024.050 396.040 3024.330 396.320 ;
        RECT 3024.670 396.040 3024.950 396.320 ;
        RECT 3025.290 396.040 3025.570 396.320 ;
        RECT 3025.910 396.040 3026.190 396.320 ;
        RECT 3026.530 396.040 3026.810 396.320 ;
        RECT 3027.150 396.040 3027.430 396.320 ;
        RECT 3027.770 396.040 3028.050 396.320 ;
        RECT 3028.390 396.040 3028.670 396.320 ;
        RECT 3029.010 396.040 3029.290 396.320 ;
        RECT 3029.630 396.040 3029.910 396.320 ;
        RECT 3030.250 396.040 3030.530 396.320 ;
        RECT 3030.870 396.040 3031.150 396.320 ;
        RECT 3031.490 396.040 3031.770 396.320 ;
        RECT 3032.110 396.040 3032.390 396.320 ;
        RECT 3032.730 396.040 3033.010 396.320 ;
        RECT 3033.350 396.040 3033.630 396.320 ;
        RECT 3035.900 399.760 3036.180 400.040 ;
        RECT 3036.520 399.760 3036.800 400.040 ;
        RECT 3037.140 399.760 3037.420 400.040 ;
        RECT 3037.760 399.760 3038.040 400.040 ;
        RECT 3038.380 399.760 3038.660 400.040 ;
        RECT 3039.000 399.760 3039.280 400.040 ;
        RECT 3039.620 399.760 3039.900 400.040 ;
        RECT 3040.240 399.760 3040.520 400.040 ;
        RECT 3040.860 399.760 3041.140 400.040 ;
        RECT 3041.480 399.760 3041.760 400.040 ;
        RECT 3042.100 399.760 3042.380 400.040 ;
        RECT 3042.720 399.760 3043.000 400.040 ;
        RECT 3043.340 399.760 3043.620 400.040 ;
        RECT 3043.960 399.760 3044.240 400.040 ;
        RECT 3044.580 399.760 3044.860 400.040 ;
        RECT 3045.200 399.760 3045.480 400.040 ;
        RECT 3035.900 399.140 3036.180 399.420 ;
        RECT 3036.520 399.140 3036.800 399.420 ;
        RECT 3037.140 399.140 3037.420 399.420 ;
        RECT 3037.760 399.140 3038.040 399.420 ;
        RECT 3038.380 399.140 3038.660 399.420 ;
        RECT 3039.000 399.140 3039.280 399.420 ;
        RECT 3039.620 399.140 3039.900 399.420 ;
        RECT 3040.240 399.140 3040.520 399.420 ;
        RECT 3040.860 399.140 3041.140 399.420 ;
        RECT 3041.480 399.140 3041.760 399.420 ;
        RECT 3042.100 399.140 3042.380 399.420 ;
        RECT 3042.720 399.140 3043.000 399.420 ;
        RECT 3043.340 399.140 3043.620 399.420 ;
        RECT 3043.960 399.140 3044.240 399.420 ;
        RECT 3044.580 399.140 3044.860 399.420 ;
        RECT 3045.200 399.140 3045.480 399.420 ;
        RECT 3035.900 398.520 3036.180 398.800 ;
        RECT 3036.520 398.520 3036.800 398.800 ;
        RECT 3037.140 398.520 3037.420 398.800 ;
        RECT 3037.760 398.520 3038.040 398.800 ;
        RECT 3038.380 398.520 3038.660 398.800 ;
        RECT 3039.000 398.520 3039.280 398.800 ;
        RECT 3039.620 398.520 3039.900 398.800 ;
        RECT 3040.240 398.520 3040.520 398.800 ;
        RECT 3040.860 398.520 3041.140 398.800 ;
        RECT 3041.480 398.520 3041.760 398.800 ;
        RECT 3042.100 398.520 3042.380 398.800 ;
        RECT 3042.720 398.520 3043.000 398.800 ;
        RECT 3043.340 398.520 3043.620 398.800 ;
        RECT 3043.960 398.520 3044.240 398.800 ;
        RECT 3044.580 398.520 3044.860 398.800 ;
        RECT 3045.200 398.520 3045.480 398.800 ;
        RECT 3035.900 397.900 3036.180 398.180 ;
        RECT 3036.520 397.900 3036.800 398.180 ;
        RECT 3037.140 397.900 3037.420 398.180 ;
        RECT 3037.760 397.900 3038.040 398.180 ;
        RECT 3038.380 397.900 3038.660 398.180 ;
        RECT 3039.000 397.900 3039.280 398.180 ;
        RECT 3039.620 397.900 3039.900 398.180 ;
        RECT 3040.240 397.900 3040.520 398.180 ;
        RECT 3040.860 397.900 3041.140 398.180 ;
        RECT 3041.480 397.900 3041.760 398.180 ;
        RECT 3042.100 397.900 3042.380 398.180 ;
        RECT 3042.720 397.900 3043.000 398.180 ;
        RECT 3043.340 397.900 3043.620 398.180 ;
        RECT 3043.960 397.900 3044.240 398.180 ;
        RECT 3044.580 397.900 3044.860 398.180 ;
        RECT 3045.200 397.900 3045.480 398.180 ;
        RECT 3035.900 397.280 3036.180 397.560 ;
        RECT 3036.520 397.280 3036.800 397.560 ;
        RECT 3037.140 397.280 3037.420 397.560 ;
        RECT 3037.760 397.280 3038.040 397.560 ;
        RECT 3038.380 397.280 3038.660 397.560 ;
        RECT 3039.000 397.280 3039.280 397.560 ;
        RECT 3039.620 397.280 3039.900 397.560 ;
        RECT 3040.240 397.280 3040.520 397.560 ;
        RECT 3040.860 397.280 3041.140 397.560 ;
        RECT 3041.480 397.280 3041.760 397.560 ;
        RECT 3042.100 397.280 3042.380 397.560 ;
        RECT 3042.720 397.280 3043.000 397.560 ;
        RECT 3043.340 397.280 3043.620 397.560 ;
        RECT 3043.960 397.280 3044.240 397.560 ;
        RECT 3044.580 397.280 3044.860 397.560 ;
        RECT 3045.200 397.280 3045.480 397.560 ;
        RECT 3035.900 396.660 3036.180 396.940 ;
        RECT 3036.520 396.660 3036.800 396.940 ;
        RECT 3037.140 396.660 3037.420 396.940 ;
        RECT 3037.760 396.660 3038.040 396.940 ;
        RECT 3038.380 396.660 3038.660 396.940 ;
        RECT 3039.000 396.660 3039.280 396.940 ;
        RECT 3039.620 396.660 3039.900 396.940 ;
        RECT 3040.240 396.660 3040.520 396.940 ;
        RECT 3040.860 396.660 3041.140 396.940 ;
        RECT 3041.480 396.660 3041.760 396.940 ;
        RECT 3042.100 396.660 3042.380 396.940 ;
        RECT 3042.720 396.660 3043.000 396.940 ;
        RECT 3043.340 396.660 3043.620 396.940 ;
        RECT 3043.960 396.660 3044.240 396.940 ;
        RECT 3044.580 396.660 3044.860 396.940 ;
        RECT 3045.200 396.660 3045.480 396.940 ;
        RECT 3035.900 396.040 3036.180 396.320 ;
        RECT 3036.520 396.040 3036.800 396.320 ;
        RECT 3037.140 396.040 3037.420 396.320 ;
        RECT 3037.760 396.040 3038.040 396.320 ;
        RECT 3038.380 396.040 3038.660 396.320 ;
        RECT 3039.000 396.040 3039.280 396.320 ;
        RECT 3039.620 396.040 3039.900 396.320 ;
        RECT 3040.240 396.040 3040.520 396.320 ;
        RECT 3040.860 396.040 3041.140 396.320 ;
        RECT 3041.480 396.040 3041.760 396.320 ;
        RECT 3042.100 396.040 3042.380 396.320 ;
        RECT 3042.720 396.040 3043.000 396.320 ;
        RECT 3043.340 396.040 3043.620 396.320 ;
        RECT 3043.960 396.040 3044.240 396.320 ;
        RECT 3044.580 396.040 3044.860 396.320 ;
        RECT 3045.200 396.040 3045.480 396.320 ;
        RECT 3049.430 399.760 3049.710 400.040 ;
        RECT 3050.050 399.760 3050.330 400.040 ;
        RECT 3050.670 399.760 3050.950 400.040 ;
        RECT 3051.290 399.760 3051.570 400.040 ;
        RECT 3051.910 399.760 3052.190 400.040 ;
        RECT 3052.530 399.760 3052.810 400.040 ;
        RECT 3053.150 399.760 3053.430 400.040 ;
        RECT 3053.770 399.760 3054.050 400.040 ;
        RECT 3054.390 399.760 3054.670 400.040 ;
        RECT 3055.010 399.760 3055.290 400.040 ;
        RECT 3055.630 399.760 3055.910 400.040 ;
        RECT 3056.250 399.760 3056.530 400.040 ;
        RECT 3056.870 399.760 3057.150 400.040 ;
        RECT 3057.490 399.760 3057.770 400.040 ;
        RECT 3058.110 399.760 3058.390 400.040 ;
        RECT 3058.730 399.760 3059.010 400.040 ;
        RECT 3049.430 399.140 3049.710 399.420 ;
        RECT 3050.050 399.140 3050.330 399.420 ;
        RECT 3050.670 399.140 3050.950 399.420 ;
        RECT 3051.290 399.140 3051.570 399.420 ;
        RECT 3051.910 399.140 3052.190 399.420 ;
        RECT 3052.530 399.140 3052.810 399.420 ;
        RECT 3053.150 399.140 3053.430 399.420 ;
        RECT 3053.770 399.140 3054.050 399.420 ;
        RECT 3054.390 399.140 3054.670 399.420 ;
        RECT 3055.010 399.140 3055.290 399.420 ;
        RECT 3055.630 399.140 3055.910 399.420 ;
        RECT 3056.250 399.140 3056.530 399.420 ;
        RECT 3056.870 399.140 3057.150 399.420 ;
        RECT 3057.490 399.140 3057.770 399.420 ;
        RECT 3058.110 399.140 3058.390 399.420 ;
        RECT 3058.730 399.140 3059.010 399.420 ;
        RECT 3049.430 398.520 3049.710 398.800 ;
        RECT 3050.050 398.520 3050.330 398.800 ;
        RECT 3050.670 398.520 3050.950 398.800 ;
        RECT 3051.290 398.520 3051.570 398.800 ;
        RECT 3051.910 398.520 3052.190 398.800 ;
        RECT 3052.530 398.520 3052.810 398.800 ;
        RECT 3053.150 398.520 3053.430 398.800 ;
        RECT 3053.770 398.520 3054.050 398.800 ;
        RECT 3054.390 398.520 3054.670 398.800 ;
        RECT 3055.010 398.520 3055.290 398.800 ;
        RECT 3055.630 398.520 3055.910 398.800 ;
        RECT 3056.250 398.520 3056.530 398.800 ;
        RECT 3056.870 398.520 3057.150 398.800 ;
        RECT 3057.490 398.520 3057.770 398.800 ;
        RECT 3058.110 398.520 3058.390 398.800 ;
        RECT 3058.730 398.520 3059.010 398.800 ;
        RECT 3049.430 397.900 3049.710 398.180 ;
        RECT 3050.050 397.900 3050.330 398.180 ;
        RECT 3050.670 397.900 3050.950 398.180 ;
        RECT 3051.290 397.900 3051.570 398.180 ;
        RECT 3051.910 397.900 3052.190 398.180 ;
        RECT 3052.530 397.900 3052.810 398.180 ;
        RECT 3053.150 397.900 3053.430 398.180 ;
        RECT 3053.770 397.900 3054.050 398.180 ;
        RECT 3054.390 397.900 3054.670 398.180 ;
        RECT 3055.010 397.900 3055.290 398.180 ;
        RECT 3055.630 397.900 3055.910 398.180 ;
        RECT 3056.250 397.900 3056.530 398.180 ;
        RECT 3056.870 397.900 3057.150 398.180 ;
        RECT 3057.490 397.900 3057.770 398.180 ;
        RECT 3058.110 397.900 3058.390 398.180 ;
        RECT 3058.730 397.900 3059.010 398.180 ;
        RECT 3049.430 397.280 3049.710 397.560 ;
        RECT 3050.050 397.280 3050.330 397.560 ;
        RECT 3050.670 397.280 3050.950 397.560 ;
        RECT 3051.290 397.280 3051.570 397.560 ;
        RECT 3051.910 397.280 3052.190 397.560 ;
        RECT 3052.530 397.280 3052.810 397.560 ;
        RECT 3053.150 397.280 3053.430 397.560 ;
        RECT 3053.770 397.280 3054.050 397.560 ;
        RECT 3054.390 397.280 3054.670 397.560 ;
        RECT 3055.010 397.280 3055.290 397.560 ;
        RECT 3055.630 397.280 3055.910 397.560 ;
        RECT 3056.250 397.280 3056.530 397.560 ;
        RECT 3056.870 397.280 3057.150 397.560 ;
        RECT 3057.490 397.280 3057.770 397.560 ;
        RECT 3058.110 397.280 3058.390 397.560 ;
        RECT 3058.730 397.280 3059.010 397.560 ;
        RECT 3049.430 396.660 3049.710 396.940 ;
        RECT 3050.050 396.660 3050.330 396.940 ;
        RECT 3050.670 396.660 3050.950 396.940 ;
        RECT 3051.290 396.660 3051.570 396.940 ;
        RECT 3051.910 396.660 3052.190 396.940 ;
        RECT 3052.530 396.660 3052.810 396.940 ;
        RECT 3053.150 396.660 3053.430 396.940 ;
        RECT 3053.770 396.660 3054.050 396.940 ;
        RECT 3054.390 396.660 3054.670 396.940 ;
        RECT 3055.010 396.660 3055.290 396.940 ;
        RECT 3055.630 396.660 3055.910 396.940 ;
        RECT 3056.250 396.660 3056.530 396.940 ;
        RECT 3056.870 396.660 3057.150 396.940 ;
        RECT 3057.490 396.660 3057.770 396.940 ;
        RECT 3058.110 396.660 3058.390 396.940 ;
        RECT 3058.730 396.660 3059.010 396.940 ;
        RECT 3049.430 396.040 3049.710 396.320 ;
        RECT 3050.050 396.040 3050.330 396.320 ;
        RECT 3050.670 396.040 3050.950 396.320 ;
        RECT 3051.290 396.040 3051.570 396.320 ;
        RECT 3051.910 396.040 3052.190 396.320 ;
        RECT 3052.530 396.040 3052.810 396.320 ;
        RECT 3053.150 396.040 3053.430 396.320 ;
        RECT 3053.770 396.040 3054.050 396.320 ;
        RECT 3054.390 396.040 3054.670 396.320 ;
        RECT 3055.010 396.040 3055.290 396.320 ;
        RECT 3055.630 396.040 3055.910 396.320 ;
        RECT 3056.250 396.040 3056.530 396.320 ;
        RECT 3056.870 396.040 3057.150 396.320 ;
        RECT 3057.490 396.040 3057.770 396.320 ;
        RECT 3058.110 396.040 3058.390 396.320 ;
        RECT 3058.730 396.040 3059.010 396.320 ;
        RECT 3061.280 399.760 3061.560 400.040 ;
        RECT 3061.900 399.760 3062.180 400.040 ;
        RECT 3062.520 399.760 3062.800 400.040 ;
        RECT 3063.140 399.760 3063.420 400.040 ;
        RECT 3063.760 399.760 3064.040 400.040 ;
        RECT 3064.380 399.760 3064.660 400.040 ;
        RECT 3065.000 399.760 3065.280 400.040 ;
        RECT 3065.620 399.760 3065.900 400.040 ;
        RECT 3066.240 399.760 3066.520 400.040 ;
        RECT 3066.860 399.760 3067.140 400.040 ;
        RECT 3067.480 399.760 3067.760 400.040 ;
        RECT 3068.100 399.760 3068.380 400.040 ;
        RECT 3068.720 399.760 3069.000 400.040 ;
        RECT 3069.340 399.760 3069.620 400.040 ;
        RECT 3069.960 399.760 3070.240 400.040 ;
        RECT 3070.580 399.760 3070.860 400.040 ;
        RECT 3061.280 399.140 3061.560 399.420 ;
        RECT 3061.900 399.140 3062.180 399.420 ;
        RECT 3062.520 399.140 3062.800 399.420 ;
        RECT 3063.140 399.140 3063.420 399.420 ;
        RECT 3063.760 399.140 3064.040 399.420 ;
        RECT 3064.380 399.140 3064.660 399.420 ;
        RECT 3065.000 399.140 3065.280 399.420 ;
        RECT 3065.620 399.140 3065.900 399.420 ;
        RECT 3066.240 399.140 3066.520 399.420 ;
        RECT 3066.860 399.140 3067.140 399.420 ;
        RECT 3067.480 399.140 3067.760 399.420 ;
        RECT 3068.100 399.140 3068.380 399.420 ;
        RECT 3068.720 399.140 3069.000 399.420 ;
        RECT 3069.340 399.140 3069.620 399.420 ;
        RECT 3069.960 399.140 3070.240 399.420 ;
        RECT 3070.580 399.140 3070.860 399.420 ;
        RECT 3061.280 398.520 3061.560 398.800 ;
        RECT 3061.900 398.520 3062.180 398.800 ;
        RECT 3062.520 398.520 3062.800 398.800 ;
        RECT 3063.140 398.520 3063.420 398.800 ;
        RECT 3063.760 398.520 3064.040 398.800 ;
        RECT 3064.380 398.520 3064.660 398.800 ;
        RECT 3065.000 398.520 3065.280 398.800 ;
        RECT 3065.620 398.520 3065.900 398.800 ;
        RECT 3066.240 398.520 3066.520 398.800 ;
        RECT 3066.860 398.520 3067.140 398.800 ;
        RECT 3067.480 398.520 3067.760 398.800 ;
        RECT 3068.100 398.520 3068.380 398.800 ;
        RECT 3068.720 398.520 3069.000 398.800 ;
        RECT 3069.340 398.520 3069.620 398.800 ;
        RECT 3069.960 398.520 3070.240 398.800 ;
        RECT 3070.580 398.520 3070.860 398.800 ;
        RECT 3061.280 397.900 3061.560 398.180 ;
        RECT 3061.900 397.900 3062.180 398.180 ;
        RECT 3062.520 397.900 3062.800 398.180 ;
        RECT 3063.140 397.900 3063.420 398.180 ;
        RECT 3063.760 397.900 3064.040 398.180 ;
        RECT 3064.380 397.900 3064.660 398.180 ;
        RECT 3065.000 397.900 3065.280 398.180 ;
        RECT 3065.620 397.900 3065.900 398.180 ;
        RECT 3066.240 397.900 3066.520 398.180 ;
        RECT 3066.860 397.900 3067.140 398.180 ;
        RECT 3067.480 397.900 3067.760 398.180 ;
        RECT 3068.100 397.900 3068.380 398.180 ;
        RECT 3068.720 397.900 3069.000 398.180 ;
        RECT 3069.340 397.900 3069.620 398.180 ;
        RECT 3069.960 397.900 3070.240 398.180 ;
        RECT 3070.580 397.900 3070.860 398.180 ;
        RECT 3061.280 397.280 3061.560 397.560 ;
        RECT 3061.900 397.280 3062.180 397.560 ;
        RECT 3062.520 397.280 3062.800 397.560 ;
        RECT 3063.140 397.280 3063.420 397.560 ;
        RECT 3063.760 397.280 3064.040 397.560 ;
        RECT 3064.380 397.280 3064.660 397.560 ;
        RECT 3065.000 397.280 3065.280 397.560 ;
        RECT 3065.620 397.280 3065.900 397.560 ;
        RECT 3066.240 397.280 3066.520 397.560 ;
        RECT 3066.860 397.280 3067.140 397.560 ;
        RECT 3067.480 397.280 3067.760 397.560 ;
        RECT 3068.100 397.280 3068.380 397.560 ;
        RECT 3068.720 397.280 3069.000 397.560 ;
        RECT 3069.340 397.280 3069.620 397.560 ;
        RECT 3069.960 397.280 3070.240 397.560 ;
        RECT 3070.580 397.280 3070.860 397.560 ;
        RECT 3061.280 396.660 3061.560 396.940 ;
        RECT 3061.900 396.660 3062.180 396.940 ;
        RECT 3062.520 396.660 3062.800 396.940 ;
        RECT 3063.140 396.660 3063.420 396.940 ;
        RECT 3063.760 396.660 3064.040 396.940 ;
        RECT 3064.380 396.660 3064.660 396.940 ;
        RECT 3065.000 396.660 3065.280 396.940 ;
        RECT 3065.620 396.660 3065.900 396.940 ;
        RECT 3066.240 396.660 3066.520 396.940 ;
        RECT 3066.860 396.660 3067.140 396.940 ;
        RECT 3067.480 396.660 3067.760 396.940 ;
        RECT 3068.100 396.660 3068.380 396.940 ;
        RECT 3068.720 396.660 3069.000 396.940 ;
        RECT 3069.340 396.660 3069.620 396.940 ;
        RECT 3069.960 396.660 3070.240 396.940 ;
        RECT 3070.580 396.660 3070.860 396.940 ;
        RECT 3061.280 396.040 3061.560 396.320 ;
        RECT 3061.900 396.040 3062.180 396.320 ;
        RECT 3062.520 396.040 3062.800 396.320 ;
        RECT 3063.140 396.040 3063.420 396.320 ;
        RECT 3063.760 396.040 3064.040 396.320 ;
        RECT 3064.380 396.040 3064.660 396.320 ;
        RECT 3065.000 396.040 3065.280 396.320 ;
        RECT 3065.620 396.040 3065.900 396.320 ;
        RECT 3066.240 396.040 3066.520 396.320 ;
        RECT 3066.860 396.040 3067.140 396.320 ;
        RECT 3067.480 396.040 3067.760 396.320 ;
        RECT 3068.100 396.040 3068.380 396.320 ;
        RECT 3068.720 396.040 3069.000 396.320 ;
        RECT 3069.340 396.040 3069.620 396.320 ;
        RECT 3069.960 396.040 3070.240 396.320 ;
        RECT 3070.580 396.040 3070.860 396.320 ;
        RECT 3074.300 399.760 3074.580 400.040 ;
        RECT 3074.920 399.760 3075.200 400.040 ;
        RECT 3075.540 399.760 3075.820 400.040 ;
        RECT 3076.160 399.760 3076.440 400.040 ;
        RECT 3076.780 399.760 3077.060 400.040 ;
        RECT 3077.400 399.760 3077.680 400.040 ;
        RECT 3078.020 399.760 3078.300 400.040 ;
        RECT 3078.640 399.760 3078.920 400.040 ;
        RECT 3079.260 399.760 3079.540 400.040 ;
        RECT 3079.880 399.760 3080.160 400.040 ;
        RECT 3080.500 399.760 3080.780 400.040 ;
        RECT 3081.120 399.760 3081.400 400.040 ;
        RECT 3081.740 399.760 3082.020 400.040 ;
        RECT 3082.360 399.760 3082.640 400.040 ;
        RECT 3082.980 399.760 3083.260 400.040 ;
        RECT 3074.300 399.140 3074.580 399.420 ;
        RECT 3074.920 399.140 3075.200 399.420 ;
        RECT 3075.540 399.140 3075.820 399.420 ;
        RECT 3076.160 399.140 3076.440 399.420 ;
        RECT 3076.780 399.140 3077.060 399.420 ;
        RECT 3077.400 399.140 3077.680 399.420 ;
        RECT 3078.020 399.140 3078.300 399.420 ;
        RECT 3078.640 399.140 3078.920 399.420 ;
        RECT 3079.260 399.140 3079.540 399.420 ;
        RECT 3079.880 399.140 3080.160 399.420 ;
        RECT 3080.500 399.140 3080.780 399.420 ;
        RECT 3081.120 399.140 3081.400 399.420 ;
        RECT 3081.740 399.140 3082.020 399.420 ;
        RECT 3082.360 399.140 3082.640 399.420 ;
        RECT 3082.980 399.140 3083.260 399.420 ;
        RECT 3074.300 398.520 3074.580 398.800 ;
        RECT 3074.920 398.520 3075.200 398.800 ;
        RECT 3075.540 398.520 3075.820 398.800 ;
        RECT 3076.160 398.520 3076.440 398.800 ;
        RECT 3076.780 398.520 3077.060 398.800 ;
        RECT 3077.400 398.520 3077.680 398.800 ;
        RECT 3078.020 398.520 3078.300 398.800 ;
        RECT 3078.640 398.520 3078.920 398.800 ;
        RECT 3079.260 398.520 3079.540 398.800 ;
        RECT 3079.880 398.520 3080.160 398.800 ;
        RECT 3080.500 398.520 3080.780 398.800 ;
        RECT 3081.120 398.520 3081.400 398.800 ;
        RECT 3081.740 398.520 3082.020 398.800 ;
        RECT 3082.360 398.520 3082.640 398.800 ;
        RECT 3082.980 398.520 3083.260 398.800 ;
        RECT 3074.300 397.900 3074.580 398.180 ;
        RECT 3074.920 397.900 3075.200 398.180 ;
        RECT 3075.540 397.900 3075.820 398.180 ;
        RECT 3076.160 397.900 3076.440 398.180 ;
        RECT 3076.780 397.900 3077.060 398.180 ;
        RECT 3077.400 397.900 3077.680 398.180 ;
        RECT 3078.020 397.900 3078.300 398.180 ;
        RECT 3078.640 397.900 3078.920 398.180 ;
        RECT 3079.260 397.900 3079.540 398.180 ;
        RECT 3079.880 397.900 3080.160 398.180 ;
        RECT 3080.500 397.900 3080.780 398.180 ;
        RECT 3081.120 397.900 3081.400 398.180 ;
        RECT 3081.740 397.900 3082.020 398.180 ;
        RECT 3082.360 397.900 3082.640 398.180 ;
        RECT 3082.980 397.900 3083.260 398.180 ;
        RECT 3074.300 397.280 3074.580 397.560 ;
        RECT 3074.920 397.280 3075.200 397.560 ;
        RECT 3075.540 397.280 3075.820 397.560 ;
        RECT 3076.160 397.280 3076.440 397.560 ;
        RECT 3076.780 397.280 3077.060 397.560 ;
        RECT 3077.400 397.280 3077.680 397.560 ;
        RECT 3078.020 397.280 3078.300 397.560 ;
        RECT 3078.640 397.280 3078.920 397.560 ;
        RECT 3079.260 397.280 3079.540 397.560 ;
        RECT 3079.880 397.280 3080.160 397.560 ;
        RECT 3080.500 397.280 3080.780 397.560 ;
        RECT 3081.120 397.280 3081.400 397.560 ;
        RECT 3081.740 397.280 3082.020 397.560 ;
        RECT 3082.360 397.280 3082.640 397.560 ;
        RECT 3082.980 397.280 3083.260 397.560 ;
        RECT 3074.300 396.660 3074.580 396.940 ;
        RECT 3074.920 396.660 3075.200 396.940 ;
        RECT 3075.540 396.660 3075.820 396.940 ;
        RECT 3076.160 396.660 3076.440 396.940 ;
        RECT 3076.780 396.660 3077.060 396.940 ;
        RECT 3077.400 396.660 3077.680 396.940 ;
        RECT 3078.020 396.660 3078.300 396.940 ;
        RECT 3078.640 396.660 3078.920 396.940 ;
        RECT 3079.260 396.660 3079.540 396.940 ;
        RECT 3079.880 396.660 3080.160 396.940 ;
        RECT 3080.500 396.660 3080.780 396.940 ;
        RECT 3081.120 396.660 3081.400 396.940 ;
        RECT 3081.740 396.660 3082.020 396.940 ;
        RECT 3082.360 396.660 3082.640 396.940 ;
        RECT 3082.980 396.660 3083.260 396.940 ;
        RECT 3074.300 396.040 3074.580 396.320 ;
        RECT 3074.920 396.040 3075.200 396.320 ;
        RECT 3075.540 396.040 3075.820 396.320 ;
        RECT 3076.160 396.040 3076.440 396.320 ;
        RECT 3076.780 396.040 3077.060 396.320 ;
        RECT 3077.400 396.040 3077.680 396.320 ;
        RECT 3078.020 396.040 3078.300 396.320 ;
        RECT 3078.640 396.040 3078.920 396.320 ;
        RECT 3079.260 396.040 3079.540 396.320 ;
        RECT 3079.880 396.040 3080.160 396.320 ;
        RECT 3080.500 396.040 3080.780 396.320 ;
        RECT 3081.120 396.040 3081.400 396.320 ;
        RECT 3081.740 396.040 3082.020 396.320 ;
        RECT 3082.360 396.040 3082.640 396.320 ;
        RECT 3082.980 396.040 3083.260 396.320 ;
        RECT 3143.485 399.760 3143.765 400.040 ;
        RECT 3144.105 399.760 3144.385 400.040 ;
        RECT 3143.485 399.140 3143.765 399.420 ;
        RECT 3144.105 399.140 3144.385 399.420 ;
        RECT 3143.485 398.520 3143.765 398.800 ;
        RECT 3144.105 398.520 3144.385 398.800 ;
        RECT 3143.485 397.900 3143.765 398.180 ;
        RECT 3144.105 397.900 3144.385 398.180 ;
        RECT 3143.485 397.280 3143.765 397.560 ;
        RECT 3144.105 397.280 3144.385 397.560 ;
        RECT 3143.485 396.660 3143.765 396.940 ;
        RECT 3144.105 396.660 3144.385 396.940 ;
        RECT 3143.485 396.040 3143.765 396.320 ;
        RECT 3144.105 396.040 3144.385 396.320 ;
        RECT 3123.635 392.760 3123.915 393.040 ;
        RECT 3124.255 392.760 3124.535 393.040 ;
        RECT 3123.635 392.140 3123.915 392.420 ;
        RECT 3124.255 392.140 3124.535 392.420 ;
        RECT 3123.635 391.520 3123.915 391.800 ;
        RECT 3124.255 391.520 3124.535 391.800 ;
        RECT 3123.635 390.900 3123.915 391.180 ;
        RECT 3124.255 390.900 3124.535 391.180 ;
        RECT 3123.635 390.280 3123.915 390.560 ;
        RECT 3124.255 390.280 3124.535 390.560 ;
        RECT 3123.635 389.660 3123.915 389.940 ;
        RECT 3124.255 389.660 3124.535 389.940 ;
        RECT 3123.635 389.040 3123.915 389.320 ;
        RECT 3124.255 389.040 3124.535 389.320 ;
        RECT 3183.185 399.760 3183.465 400.040 ;
        RECT 3183.805 399.760 3184.085 400.040 ;
        RECT 3183.185 399.140 3183.465 399.420 ;
        RECT 3183.805 399.140 3184.085 399.420 ;
        RECT 3183.185 398.520 3183.465 398.800 ;
        RECT 3183.805 398.520 3184.085 398.800 ;
        RECT 3183.185 397.900 3183.465 398.180 ;
        RECT 3183.805 397.900 3184.085 398.180 ;
        RECT 3183.185 397.280 3183.465 397.560 ;
        RECT 3183.805 397.280 3184.085 397.560 ;
        RECT 3183.185 396.660 3183.465 396.940 ;
        RECT 3183.805 396.660 3184.085 396.940 ;
        RECT 3183.185 396.040 3183.465 396.320 ;
        RECT 3183.805 396.040 3184.085 396.320 ;
        RECT 3163.335 392.760 3163.615 393.040 ;
        RECT 3163.955 392.760 3164.235 393.040 ;
        RECT 3163.335 392.140 3163.615 392.420 ;
        RECT 3163.955 392.140 3164.235 392.420 ;
        RECT 3163.335 391.520 3163.615 391.800 ;
        RECT 3163.955 391.520 3164.235 391.800 ;
        RECT 3163.335 390.900 3163.615 391.180 ;
        RECT 3163.955 390.900 3164.235 391.180 ;
        RECT 3163.335 390.280 3163.615 390.560 ;
        RECT 3163.955 390.280 3164.235 390.560 ;
        RECT 3163.335 389.660 3163.615 389.940 ;
        RECT 3163.955 389.660 3164.235 389.940 ;
        RECT 3163.335 389.040 3163.615 389.320 ;
        RECT 3163.955 389.040 3164.235 389.320 ;
        RECT 3222.885 399.760 3223.165 400.040 ;
        RECT 3223.505 399.760 3223.785 400.040 ;
        RECT 3222.885 399.140 3223.165 399.420 ;
        RECT 3223.505 399.140 3223.785 399.420 ;
        RECT 3222.885 398.520 3223.165 398.800 ;
        RECT 3223.505 398.520 3223.785 398.800 ;
        RECT 3222.885 397.900 3223.165 398.180 ;
        RECT 3223.505 397.900 3223.785 398.180 ;
        RECT 3222.885 397.280 3223.165 397.560 ;
        RECT 3223.505 397.280 3223.785 397.560 ;
        RECT 3222.885 396.660 3223.165 396.940 ;
        RECT 3223.505 396.660 3223.785 396.940 ;
        RECT 3222.885 396.040 3223.165 396.320 ;
        RECT 3223.505 396.040 3223.785 396.320 ;
        RECT 3203.035 392.760 3203.315 393.040 ;
        RECT 3203.655 392.760 3203.935 393.040 ;
        RECT 3203.035 392.140 3203.315 392.420 ;
        RECT 3203.655 392.140 3203.935 392.420 ;
        RECT 3203.035 391.520 3203.315 391.800 ;
        RECT 3203.655 391.520 3203.935 391.800 ;
        RECT 3203.035 390.900 3203.315 391.180 ;
        RECT 3203.655 390.900 3203.935 391.180 ;
        RECT 3203.035 390.280 3203.315 390.560 ;
        RECT 3203.655 390.280 3203.935 390.560 ;
        RECT 3203.035 389.660 3203.315 389.940 ;
        RECT 3203.655 389.660 3203.935 389.940 ;
        RECT 3203.035 389.040 3203.315 389.320 ;
        RECT 3203.655 389.040 3203.935 389.320 ;
        RECT 3350.450 497.265 3350.730 497.545 ;
        RECT 3351.070 497.265 3351.350 497.545 ;
        RECT 3351.690 497.265 3351.970 497.545 ;
        RECT 3352.310 497.265 3352.590 497.545 ;
        RECT 3352.930 497.265 3353.210 497.545 ;
        RECT 3353.550 497.265 3353.830 497.545 ;
        RECT 3350.450 496.645 3350.730 496.925 ;
        RECT 3351.070 496.645 3351.350 496.925 ;
        RECT 3351.690 496.645 3351.970 496.925 ;
        RECT 3352.310 496.645 3352.590 496.925 ;
        RECT 3352.930 496.645 3353.210 496.925 ;
        RECT 3353.550 496.645 3353.830 496.925 ;
        RECT 3350.450 496.025 3350.730 496.305 ;
        RECT 3351.070 496.025 3351.350 496.305 ;
        RECT 3351.690 496.025 3351.970 496.305 ;
        RECT 3352.310 496.025 3352.590 496.305 ;
        RECT 3352.930 496.025 3353.210 496.305 ;
        RECT 3353.550 496.025 3353.830 496.305 ;
        RECT 3350.450 495.405 3350.730 495.685 ;
        RECT 3351.070 495.405 3351.350 495.685 ;
        RECT 3351.690 495.405 3351.970 495.685 ;
        RECT 3352.310 495.405 3352.590 495.685 ;
        RECT 3352.930 495.405 3353.210 495.685 ;
        RECT 3353.550 495.405 3353.830 495.685 ;
        RECT 3350.450 494.785 3350.730 495.065 ;
        RECT 3351.070 494.785 3351.350 495.065 ;
        RECT 3351.690 494.785 3351.970 495.065 ;
        RECT 3352.310 494.785 3352.590 495.065 ;
        RECT 3352.930 494.785 3353.210 495.065 ;
        RECT 3353.550 494.785 3353.830 495.065 ;
        RECT 3350.450 494.165 3350.730 494.445 ;
        RECT 3351.070 494.165 3351.350 494.445 ;
        RECT 3351.690 494.165 3351.970 494.445 ;
        RECT 3352.310 494.165 3352.590 494.445 ;
        RECT 3352.930 494.165 3353.210 494.445 ;
        RECT 3353.550 494.165 3353.830 494.445 ;
        RECT 3350.450 493.545 3350.730 493.825 ;
        RECT 3351.070 493.545 3351.350 493.825 ;
        RECT 3351.690 493.545 3351.970 493.825 ;
        RECT 3352.310 493.545 3352.590 493.825 ;
        RECT 3352.930 493.545 3353.210 493.825 ;
        RECT 3353.550 493.545 3353.830 493.825 ;
        RECT 3350.450 399.760 3350.730 400.040 ;
        RECT 3351.070 399.760 3351.350 400.040 ;
        RECT 3351.690 399.760 3351.970 400.040 ;
        RECT 3352.310 399.760 3352.590 400.040 ;
        RECT 3352.930 399.760 3353.210 400.040 ;
        RECT 3353.550 399.760 3353.830 400.040 ;
        RECT 3350.450 399.140 3350.730 399.420 ;
        RECT 3351.070 399.140 3351.350 399.420 ;
        RECT 3351.690 399.140 3351.970 399.420 ;
        RECT 3352.310 399.140 3352.590 399.420 ;
        RECT 3352.930 399.140 3353.210 399.420 ;
        RECT 3353.550 399.140 3353.830 399.420 ;
        RECT 3350.450 398.520 3350.730 398.800 ;
        RECT 3351.070 398.520 3351.350 398.800 ;
        RECT 3351.690 398.520 3351.970 398.800 ;
        RECT 3352.310 398.520 3352.590 398.800 ;
        RECT 3352.930 398.520 3353.210 398.800 ;
        RECT 3353.550 398.520 3353.830 398.800 ;
        RECT 3350.450 397.900 3350.730 398.180 ;
        RECT 3351.070 397.900 3351.350 398.180 ;
        RECT 3351.690 397.900 3351.970 398.180 ;
        RECT 3352.310 397.900 3352.590 398.180 ;
        RECT 3352.930 397.900 3353.210 398.180 ;
        RECT 3353.550 397.900 3353.830 398.180 ;
        RECT 3350.450 397.280 3350.730 397.560 ;
        RECT 3351.070 397.280 3351.350 397.560 ;
        RECT 3351.690 397.280 3351.970 397.560 ;
        RECT 3352.310 397.280 3352.590 397.560 ;
        RECT 3352.930 397.280 3353.210 397.560 ;
        RECT 3353.550 397.280 3353.830 397.560 ;
        RECT 3350.450 396.660 3350.730 396.940 ;
        RECT 3351.070 396.660 3351.350 396.940 ;
        RECT 3351.690 396.660 3351.970 396.940 ;
        RECT 3352.310 396.660 3352.590 396.940 ;
        RECT 3352.930 396.660 3353.210 396.940 ;
        RECT 3353.550 396.660 3353.830 396.940 ;
        RECT 3350.450 396.040 3350.730 396.320 ;
        RECT 3351.070 396.040 3351.350 396.320 ;
        RECT 3351.690 396.040 3351.970 396.320 ;
        RECT 3352.310 396.040 3352.590 396.320 ;
        RECT 3352.930 396.040 3353.210 396.320 ;
        RECT 3353.550 396.040 3353.830 396.320 ;
        RECT 3490.220 491.890 3490.500 492.170 ;
        RECT 3491.720 491.890 3492.000 492.170 ;
        RECT 3493.220 491.890 3493.500 492.170 ;
        RECT 3490.220 456.890 3490.500 457.170 ;
        RECT 3491.720 456.890 3492.000 457.170 ;
        RECT 3493.220 456.890 3493.500 457.170 ;
        RECT 3490.260 399.760 3490.540 400.040 ;
        RECT 3490.880 399.760 3491.160 400.040 ;
        RECT 3491.500 399.760 3491.780 400.040 ;
        RECT 3492.120 399.760 3492.400 400.040 ;
        RECT 3492.740 399.760 3493.020 400.040 ;
        RECT 3493.360 399.760 3493.640 400.040 ;
        RECT 3493.980 399.760 3494.260 400.040 ;
        RECT 3490.260 399.140 3490.540 399.420 ;
        RECT 3490.880 399.140 3491.160 399.420 ;
        RECT 3491.500 399.140 3491.780 399.420 ;
        RECT 3492.120 399.140 3492.400 399.420 ;
        RECT 3492.740 399.140 3493.020 399.420 ;
        RECT 3493.360 399.140 3493.640 399.420 ;
        RECT 3493.980 399.140 3494.260 399.420 ;
        RECT 3490.260 398.520 3490.540 398.800 ;
        RECT 3490.880 398.520 3491.160 398.800 ;
        RECT 3491.500 398.520 3491.780 398.800 ;
        RECT 3492.120 398.520 3492.400 398.800 ;
        RECT 3492.740 398.520 3493.020 398.800 ;
        RECT 3493.360 398.520 3493.640 398.800 ;
        RECT 3493.980 398.520 3494.260 398.800 ;
        RECT 3490.260 397.900 3490.540 398.180 ;
        RECT 3490.880 397.900 3491.160 398.180 ;
        RECT 3491.500 397.900 3491.780 398.180 ;
        RECT 3492.120 397.900 3492.400 398.180 ;
        RECT 3492.740 397.900 3493.020 398.180 ;
        RECT 3493.360 397.900 3493.640 398.180 ;
        RECT 3493.980 397.900 3494.260 398.180 ;
        RECT 3490.260 397.280 3490.540 397.560 ;
        RECT 3490.880 397.280 3491.160 397.560 ;
        RECT 3491.500 397.280 3491.780 397.560 ;
        RECT 3492.120 397.280 3492.400 397.560 ;
        RECT 3492.740 397.280 3493.020 397.560 ;
        RECT 3493.360 397.280 3493.640 397.560 ;
        RECT 3493.980 397.280 3494.260 397.560 ;
        RECT 3490.260 396.660 3490.540 396.940 ;
        RECT 3490.880 396.660 3491.160 396.940 ;
        RECT 3491.500 396.660 3491.780 396.940 ;
        RECT 3492.120 396.660 3492.400 396.940 ;
        RECT 3492.740 396.660 3493.020 396.940 ;
        RECT 3493.360 396.660 3493.640 396.940 ;
        RECT 3493.980 396.660 3494.260 396.940 ;
        RECT 3490.260 396.040 3490.540 396.320 ;
        RECT 3490.880 396.040 3491.160 396.320 ;
        RECT 3491.500 396.040 3491.780 396.320 ;
        RECT 3492.120 396.040 3492.400 396.320 ;
        RECT 3492.740 396.040 3493.020 396.320 ;
        RECT 3493.360 396.040 3493.640 396.320 ;
        RECT 3493.980 396.040 3494.260 396.320 ;
        RECT 3242.735 392.760 3243.015 393.040 ;
        RECT 3243.355 392.760 3243.635 393.040 ;
        RECT 3242.735 392.140 3243.015 392.420 ;
        RECT 3243.355 392.140 3243.635 392.420 ;
        RECT 3242.735 391.520 3243.015 391.800 ;
        RECT 3243.355 391.520 3243.635 391.800 ;
        RECT 3242.735 390.900 3243.015 391.180 ;
        RECT 3243.355 390.900 3243.635 391.180 ;
        RECT 3242.735 390.280 3243.015 390.560 ;
        RECT 3243.355 390.280 3243.635 390.560 ;
        RECT 3242.735 389.660 3243.015 389.940 ;
        RECT 3243.355 389.660 3243.635 389.940 ;
        RECT 3242.735 389.040 3243.015 389.320 ;
        RECT 3243.355 389.040 3243.635 389.320 ;
        RECT 3286.650 392.760 3286.930 393.040 ;
        RECT 3287.270 392.760 3287.550 393.040 ;
        RECT 3287.890 392.760 3288.170 393.040 ;
        RECT 3288.510 392.760 3288.790 393.040 ;
        RECT 3289.130 392.760 3289.410 393.040 ;
        RECT 3289.750 392.760 3290.030 393.040 ;
        RECT 3290.370 392.760 3290.650 393.040 ;
        RECT 3290.990 392.760 3291.270 393.040 ;
        RECT 3291.610 392.760 3291.890 393.040 ;
        RECT 3292.230 392.760 3292.510 393.040 ;
        RECT 3292.850 392.760 3293.130 393.040 ;
        RECT 3293.470 392.760 3293.750 393.040 ;
        RECT 3294.090 392.760 3294.370 393.040 ;
        RECT 3294.710 392.760 3294.990 393.040 ;
        RECT 3295.330 392.760 3295.610 393.040 ;
        RECT 3286.650 392.140 3286.930 392.420 ;
        RECT 3287.270 392.140 3287.550 392.420 ;
        RECT 3287.890 392.140 3288.170 392.420 ;
        RECT 3288.510 392.140 3288.790 392.420 ;
        RECT 3289.130 392.140 3289.410 392.420 ;
        RECT 3289.750 392.140 3290.030 392.420 ;
        RECT 3290.370 392.140 3290.650 392.420 ;
        RECT 3290.990 392.140 3291.270 392.420 ;
        RECT 3291.610 392.140 3291.890 392.420 ;
        RECT 3292.230 392.140 3292.510 392.420 ;
        RECT 3292.850 392.140 3293.130 392.420 ;
        RECT 3293.470 392.140 3293.750 392.420 ;
        RECT 3294.090 392.140 3294.370 392.420 ;
        RECT 3294.710 392.140 3294.990 392.420 ;
        RECT 3295.330 392.140 3295.610 392.420 ;
        RECT 3286.650 391.520 3286.930 391.800 ;
        RECT 3287.270 391.520 3287.550 391.800 ;
        RECT 3287.890 391.520 3288.170 391.800 ;
        RECT 3288.510 391.520 3288.790 391.800 ;
        RECT 3289.130 391.520 3289.410 391.800 ;
        RECT 3289.750 391.520 3290.030 391.800 ;
        RECT 3290.370 391.520 3290.650 391.800 ;
        RECT 3290.990 391.520 3291.270 391.800 ;
        RECT 3291.610 391.520 3291.890 391.800 ;
        RECT 3292.230 391.520 3292.510 391.800 ;
        RECT 3292.850 391.520 3293.130 391.800 ;
        RECT 3293.470 391.520 3293.750 391.800 ;
        RECT 3294.090 391.520 3294.370 391.800 ;
        RECT 3294.710 391.520 3294.990 391.800 ;
        RECT 3295.330 391.520 3295.610 391.800 ;
        RECT 3286.650 390.900 3286.930 391.180 ;
        RECT 3287.270 390.900 3287.550 391.180 ;
        RECT 3287.890 390.900 3288.170 391.180 ;
        RECT 3288.510 390.900 3288.790 391.180 ;
        RECT 3289.130 390.900 3289.410 391.180 ;
        RECT 3289.750 390.900 3290.030 391.180 ;
        RECT 3290.370 390.900 3290.650 391.180 ;
        RECT 3290.990 390.900 3291.270 391.180 ;
        RECT 3291.610 390.900 3291.890 391.180 ;
        RECT 3292.230 390.900 3292.510 391.180 ;
        RECT 3292.850 390.900 3293.130 391.180 ;
        RECT 3293.470 390.900 3293.750 391.180 ;
        RECT 3294.090 390.900 3294.370 391.180 ;
        RECT 3294.710 390.900 3294.990 391.180 ;
        RECT 3295.330 390.900 3295.610 391.180 ;
        RECT 3286.650 390.280 3286.930 390.560 ;
        RECT 3287.270 390.280 3287.550 390.560 ;
        RECT 3287.890 390.280 3288.170 390.560 ;
        RECT 3288.510 390.280 3288.790 390.560 ;
        RECT 3289.130 390.280 3289.410 390.560 ;
        RECT 3289.750 390.280 3290.030 390.560 ;
        RECT 3290.370 390.280 3290.650 390.560 ;
        RECT 3290.990 390.280 3291.270 390.560 ;
        RECT 3291.610 390.280 3291.890 390.560 ;
        RECT 3292.230 390.280 3292.510 390.560 ;
        RECT 3292.850 390.280 3293.130 390.560 ;
        RECT 3293.470 390.280 3293.750 390.560 ;
        RECT 3294.090 390.280 3294.370 390.560 ;
        RECT 3294.710 390.280 3294.990 390.560 ;
        RECT 3295.330 390.280 3295.610 390.560 ;
        RECT 3286.650 389.660 3286.930 389.940 ;
        RECT 3287.270 389.660 3287.550 389.940 ;
        RECT 3287.890 389.660 3288.170 389.940 ;
        RECT 3288.510 389.660 3288.790 389.940 ;
        RECT 3289.130 389.660 3289.410 389.940 ;
        RECT 3289.750 389.660 3290.030 389.940 ;
        RECT 3290.370 389.660 3290.650 389.940 ;
        RECT 3290.990 389.660 3291.270 389.940 ;
        RECT 3291.610 389.660 3291.890 389.940 ;
        RECT 3292.230 389.660 3292.510 389.940 ;
        RECT 3292.850 389.660 3293.130 389.940 ;
        RECT 3293.470 389.660 3293.750 389.940 ;
        RECT 3294.090 389.660 3294.370 389.940 ;
        RECT 3294.710 389.660 3294.990 389.940 ;
        RECT 3295.330 389.660 3295.610 389.940 ;
        RECT 3286.650 389.040 3286.930 389.320 ;
        RECT 3287.270 389.040 3287.550 389.320 ;
        RECT 3287.890 389.040 3288.170 389.320 ;
        RECT 3288.510 389.040 3288.790 389.320 ;
        RECT 3289.130 389.040 3289.410 389.320 ;
        RECT 3289.750 389.040 3290.030 389.320 ;
        RECT 3290.370 389.040 3290.650 389.320 ;
        RECT 3290.990 389.040 3291.270 389.320 ;
        RECT 3291.610 389.040 3291.890 389.320 ;
        RECT 3292.230 389.040 3292.510 389.320 ;
        RECT 3292.850 389.040 3293.130 389.320 ;
        RECT 3293.470 389.040 3293.750 389.320 ;
        RECT 3294.090 389.040 3294.370 389.320 ;
        RECT 3294.710 389.040 3294.990 389.320 ;
        RECT 3295.330 389.040 3295.610 389.320 ;
        RECT 3299.050 392.760 3299.330 393.040 ;
        RECT 3299.670 392.760 3299.950 393.040 ;
        RECT 3300.290 392.760 3300.570 393.040 ;
        RECT 3300.910 392.760 3301.190 393.040 ;
        RECT 3301.530 392.760 3301.810 393.040 ;
        RECT 3302.150 392.760 3302.430 393.040 ;
        RECT 3302.770 392.760 3303.050 393.040 ;
        RECT 3303.390 392.760 3303.670 393.040 ;
        RECT 3304.010 392.760 3304.290 393.040 ;
        RECT 3304.630 392.760 3304.910 393.040 ;
        RECT 3305.250 392.760 3305.530 393.040 ;
        RECT 3305.870 392.760 3306.150 393.040 ;
        RECT 3306.490 392.760 3306.770 393.040 ;
        RECT 3307.110 392.760 3307.390 393.040 ;
        RECT 3307.730 392.760 3308.010 393.040 ;
        RECT 3308.350 392.760 3308.630 393.040 ;
        RECT 3299.050 392.140 3299.330 392.420 ;
        RECT 3299.670 392.140 3299.950 392.420 ;
        RECT 3300.290 392.140 3300.570 392.420 ;
        RECT 3300.910 392.140 3301.190 392.420 ;
        RECT 3301.530 392.140 3301.810 392.420 ;
        RECT 3302.150 392.140 3302.430 392.420 ;
        RECT 3302.770 392.140 3303.050 392.420 ;
        RECT 3303.390 392.140 3303.670 392.420 ;
        RECT 3304.010 392.140 3304.290 392.420 ;
        RECT 3304.630 392.140 3304.910 392.420 ;
        RECT 3305.250 392.140 3305.530 392.420 ;
        RECT 3305.870 392.140 3306.150 392.420 ;
        RECT 3306.490 392.140 3306.770 392.420 ;
        RECT 3307.110 392.140 3307.390 392.420 ;
        RECT 3307.730 392.140 3308.010 392.420 ;
        RECT 3308.350 392.140 3308.630 392.420 ;
        RECT 3299.050 391.520 3299.330 391.800 ;
        RECT 3299.670 391.520 3299.950 391.800 ;
        RECT 3300.290 391.520 3300.570 391.800 ;
        RECT 3300.910 391.520 3301.190 391.800 ;
        RECT 3301.530 391.520 3301.810 391.800 ;
        RECT 3302.150 391.520 3302.430 391.800 ;
        RECT 3302.770 391.520 3303.050 391.800 ;
        RECT 3303.390 391.520 3303.670 391.800 ;
        RECT 3304.010 391.520 3304.290 391.800 ;
        RECT 3304.630 391.520 3304.910 391.800 ;
        RECT 3305.250 391.520 3305.530 391.800 ;
        RECT 3305.870 391.520 3306.150 391.800 ;
        RECT 3306.490 391.520 3306.770 391.800 ;
        RECT 3307.110 391.520 3307.390 391.800 ;
        RECT 3307.730 391.520 3308.010 391.800 ;
        RECT 3308.350 391.520 3308.630 391.800 ;
        RECT 3299.050 390.900 3299.330 391.180 ;
        RECT 3299.670 390.900 3299.950 391.180 ;
        RECT 3300.290 390.900 3300.570 391.180 ;
        RECT 3300.910 390.900 3301.190 391.180 ;
        RECT 3301.530 390.900 3301.810 391.180 ;
        RECT 3302.150 390.900 3302.430 391.180 ;
        RECT 3302.770 390.900 3303.050 391.180 ;
        RECT 3303.390 390.900 3303.670 391.180 ;
        RECT 3304.010 390.900 3304.290 391.180 ;
        RECT 3304.630 390.900 3304.910 391.180 ;
        RECT 3305.250 390.900 3305.530 391.180 ;
        RECT 3305.870 390.900 3306.150 391.180 ;
        RECT 3306.490 390.900 3306.770 391.180 ;
        RECT 3307.110 390.900 3307.390 391.180 ;
        RECT 3307.730 390.900 3308.010 391.180 ;
        RECT 3308.350 390.900 3308.630 391.180 ;
        RECT 3299.050 390.280 3299.330 390.560 ;
        RECT 3299.670 390.280 3299.950 390.560 ;
        RECT 3300.290 390.280 3300.570 390.560 ;
        RECT 3300.910 390.280 3301.190 390.560 ;
        RECT 3301.530 390.280 3301.810 390.560 ;
        RECT 3302.150 390.280 3302.430 390.560 ;
        RECT 3302.770 390.280 3303.050 390.560 ;
        RECT 3303.390 390.280 3303.670 390.560 ;
        RECT 3304.010 390.280 3304.290 390.560 ;
        RECT 3304.630 390.280 3304.910 390.560 ;
        RECT 3305.250 390.280 3305.530 390.560 ;
        RECT 3305.870 390.280 3306.150 390.560 ;
        RECT 3306.490 390.280 3306.770 390.560 ;
        RECT 3307.110 390.280 3307.390 390.560 ;
        RECT 3307.730 390.280 3308.010 390.560 ;
        RECT 3308.350 390.280 3308.630 390.560 ;
        RECT 3299.050 389.660 3299.330 389.940 ;
        RECT 3299.670 389.660 3299.950 389.940 ;
        RECT 3300.290 389.660 3300.570 389.940 ;
        RECT 3300.910 389.660 3301.190 389.940 ;
        RECT 3301.530 389.660 3301.810 389.940 ;
        RECT 3302.150 389.660 3302.430 389.940 ;
        RECT 3302.770 389.660 3303.050 389.940 ;
        RECT 3303.390 389.660 3303.670 389.940 ;
        RECT 3304.010 389.660 3304.290 389.940 ;
        RECT 3304.630 389.660 3304.910 389.940 ;
        RECT 3305.250 389.660 3305.530 389.940 ;
        RECT 3305.870 389.660 3306.150 389.940 ;
        RECT 3306.490 389.660 3306.770 389.940 ;
        RECT 3307.110 389.660 3307.390 389.940 ;
        RECT 3307.730 389.660 3308.010 389.940 ;
        RECT 3308.350 389.660 3308.630 389.940 ;
        RECT 3299.050 389.040 3299.330 389.320 ;
        RECT 3299.670 389.040 3299.950 389.320 ;
        RECT 3300.290 389.040 3300.570 389.320 ;
        RECT 3300.910 389.040 3301.190 389.320 ;
        RECT 3301.530 389.040 3301.810 389.320 ;
        RECT 3302.150 389.040 3302.430 389.320 ;
        RECT 3302.770 389.040 3303.050 389.320 ;
        RECT 3303.390 389.040 3303.670 389.320 ;
        RECT 3304.010 389.040 3304.290 389.320 ;
        RECT 3304.630 389.040 3304.910 389.320 ;
        RECT 3305.250 389.040 3305.530 389.320 ;
        RECT 3305.870 389.040 3306.150 389.320 ;
        RECT 3306.490 389.040 3306.770 389.320 ;
        RECT 3307.110 389.040 3307.390 389.320 ;
        RECT 3307.730 389.040 3308.010 389.320 ;
        RECT 3308.350 389.040 3308.630 389.320 ;
        RECT 3310.900 392.760 3311.180 393.040 ;
        RECT 3311.520 392.760 3311.800 393.040 ;
        RECT 3312.140 392.760 3312.420 393.040 ;
        RECT 3312.760 392.760 3313.040 393.040 ;
        RECT 3313.380 392.760 3313.660 393.040 ;
        RECT 3314.000 392.760 3314.280 393.040 ;
        RECT 3314.620 392.760 3314.900 393.040 ;
        RECT 3315.240 392.760 3315.520 393.040 ;
        RECT 3315.860 392.760 3316.140 393.040 ;
        RECT 3316.480 392.760 3316.760 393.040 ;
        RECT 3317.100 392.760 3317.380 393.040 ;
        RECT 3317.720 392.760 3318.000 393.040 ;
        RECT 3318.340 392.760 3318.620 393.040 ;
        RECT 3318.960 392.760 3319.240 393.040 ;
        RECT 3319.580 392.760 3319.860 393.040 ;
        RECT 3320.200 392.760 3320.480 393.040 ;
        RECT 3310.900 392.140 3311.180 392.420 ;
        RECT 3311.520 392.140 3311.800 392.420 ;
        RECT 3312.140 392.140 3312.420 392.420 ;
        RECT 3312.760 392.140 3313.040 392.420 ;
        RECT 3313.380 392.140 3313.660 392.420 ;
        RECT 3314.000 392.140 3314.280 392.420 ;
        RECT 3314.620 392.140 3314.900 392.420 ;
        RECT 3315.240 392.140 3315.520 392.420 ;
        RECT 3315.860 392.140 3316.140 392.420 ;
        RECT 3316.480 392.140 3316.760 392.420 ;
        RECT 3317.100 392.140 3317.380 392.420 ;
        RECT 3317.720 392.140 3318.000 392.420 ;
        RECT 3318.340 392.140 3318.620 392.420 ;
        RECT 3318.960 392.140 3319.240 392.420 ;
        RECT 3319.580 392.140 3319.860 392.420 ;
        RECT 3320.200 392.140 3320.480 392.420 ;
        RECT 3310.900 391.520 3311.180 391.800 ;
        RECT 3311.520 391.520 3311.800 391.800 ;
        RECT 3312.140 391.520 3312.420 391.800 ;
        RECT 3312.760 391.520 3313.040 391.800 ;
        RECT 3313.380 391.520 3313.660 391.800 ;
        RECT 3314.000 391.520 3314.280 391.800 ;
        RECT 3314.620 391.520 3314.900 391.800 ;
        RECT 3315.240 391.520 3315.520 391.800 ;
        RECT 3315.860 391.520 3316.140 391.800 ;
        RECT 3316.480 391.520 3316.760 391.800 ;
        RECT 3317.100 391.520 3317.380 391.800 ;
        RECT 3317.720 391.520 3318.000 391.800 ;
        RECT 3318.340 391.520 3318.620 391.800 ;
        RECT 3318.960 391.520 3319.240 391.800 ;
        RECT 3319.580 391.520 3319.860 391.800 ;
        RECT 3320.200 391.520 3320.480 391.800 ;
        RECT 3310.900 390.900 3311.180 391.180 ;
        RECT 3311.520 390.900 3311.800 391.180 ;
        RECT 3312.140 390.900 3312.420 391.180 ;
        RECT 3312.760 390.900 3313.040 391.180 ;
        RECT 3313.380 390.900 3313.660 391.180 ;
        RECT 3314.000 390.900 3314.280 391.180 ;
        RECT 3314.620 390.900 3314.900 391.180 ;
        RECT 3315.240 390.900 3315.520 391.180 ;
        RECT 3315.860 390.900 3316.140 391.180 ;
        RECT 3316.480 390.900 3316.760 391.180 ;
        RECT 3317.100 390.900 3317.380 391.180 ;
        RECT 3317.720 390.900 3318.000 391.180 ;
        RECT 3318.340 390.900 3318.620 391.180 ;
        RECT 3318.960 390.900 3319.240 391.180 ;
        RECT 3319.580 390.900 3319.860 391.180 ;
        RECT 3320.200 390.900 3320.480 391.180 ;
        RECT 3310.900 390.280 3311.180 390.560 ;
        RECT 3311.520 390.280 3311.800 390.560 ;
        RECT 3312.140 390.280 3312.420 390.560 ;
        RECT 3312.760 390.280 3313.040 390.560 ;
        RECT 3313.380 390.280 3313.660 390.560 ;
        RECT 3314.000 390.280 3314.280 390.560 ;
        RECT 3314.620 390.280 3314.900 390.560 ;
        RECT 3315.240 390.280 3315.520 390.560 ;
        RECT 3315.860 390.280 3316.140 390.560 ;
        RECT 3316.480 390.280 3316.760 390.560 ;
        RECT 3317.100 390.280 3317.380 390.560 ;
        RECT 3317.720 390.280 3318.000 390.560 ;
        RECT 3318.340 390.280 3318.620 390.560 ;
        RECT 3318.960 390.280 3319.240 390.560 ;
        RECT 3319.580 390.280 3319.860 390.560 ;
        RECT 3320.200 390.280 3320.480 390.560 ;
        RECT 3310.900 389.660 3311.180 389.940 ;
        RECT 3311.520 389.660 3311.800 389.940 ;
        RECT 3312.140 389.660 3312.420 389.940 ;
        RECT 3312.760 389.660 3313.040 389.940 ;
        RECT 3313.380 389.660 3313.660 389.940 ;
        RECT 3314.000 389.660 3314.280 389.940 ;
        RECT 3314.620 389.660 3314.900 389.940 ;
        RECT 3315.240 389.660 3315.520 389.940 ;
        RECT 3315.860 389.660 3316.140 389.940 ;
        RECT 3316.480 389.660 3316.760 389.940 ;
        RECT 3317.100 389.660 3317.380 389.940 ;
        RECT 3317.720 389.660 3318.000 389.940 ;
        RECT 3318.340 389.660 3318.620 389.940 ;
        RECT 3318.960 389.660 3319.240 389.940 ;
        RECT 3319.580 389.660 3319.860 389.940 ;
        RECT 3320.200 389.660 3320.480 389.940 ;
        RECT 3310.900 389.040 3311.180 389.320 ;
        RECT 3311.520 389.040 3311.800 389.320 ;
        RECT 3312.140 389.040 3312.420 389.320 ;
        RECT 3312.760 389.040 3313.040 389.320 ;
        RECT 3313.380 389.040 3313.660 389.320 ;
        RECT 3314.000 389.040 3314.280 389.320 ;
        RECT 3314.620 389.040 3314.900 389.320 ;
        RECT 3315.240 389.040 3315.520 389.320 ;
        RECT 3315.860 389.040 3316.140 389.320 ;
        RECT 3316.480 389.040 3316.760 389.320 ;
        RECT 3317.100 389.040 3317.380 389.320 ;
        RECT 3317.720 389.040 3318.000 389.320 ;
        RECT 3318.340 389.040 3318.620 389.320 ;
        RECT 3318.960 389.040 3319.240 389.320 ;
        RECT 3319.580 389.040 3319.860 389.320 ;
        RECT 3320.200 389.040 3320.480 389.320 ;
        RECT 3324.430 392.760 3324.710 393.040 ;
        RECT 3325.050 392.760 3325.330 393.040 ;
        RECT 3325.670 392.760 3325.950 393.040 ;
        RECT 3326.290 392.760 3326.570 393.040 ;
        RECT 3326.910 392.760 3327.190 393.040 ;
        RECT 3327.530 392.760 3327.810 393.040 ;
        RECT 3328.150 392.760 3328.430 393.040 ;
        RECT 3328.770 392.760 3329.050 393.040 ;
        RECT 3329.390 392.760 3329.670 393.040 ;
        RECT 3330.010 392.760 3330.290 393.040 ;
        RECT 3330.630 392.760 3330.910 393.040 ;
        RECT 3331.250 392.760 3331.530 393.040 ;
        RECT 3331.870 392.760 3332.150 393.040 ;
        RECT 3332.490 392.760 3332.770 393.040 ;
        RECT 3333.110 392.760 3333.390 393.040 ;
        RECT 3333.730 392.760 3334.010 393.040 ;
        RECT 3324.430 392.140 3324.710 392.420 ;
        RECT 3325.050 392.140 3325.330 392.420 ;
        RECT 3325.670 392.140 3325.950 392.420 ;
        RECT 3326.290 392.140 3326.570 392.420 ;
        RECT 3326.910 392.140 3327.190 392.420 ;
        RECT 3327.530 392.140 3327.810 392.420 ;
        RECT 3328.150 392.140 3328.430 392.420 ;
        RECT 3328.770 392.140 3329.050 392.420 ;
        RECT 3329.390 392.140 3329.670 392.420 ;
        RECT 3330.010 392.140 3330.290 392.420 ;
        RECT 3330.630 392.140 3330.910 392.420 ;
        RECT 3331.250 392.140 3331.530 392.420 ;
        RECT 3331.870 392.140 3332.150 392.420 ;
        RECT 3332.490 392.140 3332.770 392.420 ;
        RECT 3333.110 392.140 3333.390 392.420 ;
        RECT 3333.730 392.140 3334.010 392.420 ;
        RECT 3324.430 391.520 3324.710 391.800 ;
        RECT 3325.050 391.520 3325.330 391.800 ;
        RECT 3325.670 391.520 3325.950 391.800 ;
        RECT 3326.290 391.520 3326.570 391.800 ;
        RECT 3326.910 391.520 3327.190 391.800 ;
        RECT 3327.530 391.520 3327.810 391.800 ;
        RECT 3328.150 391.520 3328.430 391.800 ;
        RECT 3328.770 391.520 3329.050 391.800 ;
        RECT 3329.390 391.520 3329.670 391.800 ;
        RECT 3330.010 391.520 3330.290 391.800 ;
        RECT 3330.630 391.520 3330.910 391.800 ;
        RECT 3331.250 391.520 3331.530 391.800 ;
        RECT 3331.870 391.520 3332.150 391.800 ;
        RECT 3332.490 391.520 3332.770 391.800 ;
        RECT 3333.110 391.520 3333.390 391.800 ;
        RECT 3333.730 391.520 3334.010 391.800 ;
        RECT 3324.430 390.900 3324.710 391.180 ;
        RECT 3325.050 390.900 3325.330 391.180 ;
        RECT 3325.670 390.900 3325.950 391.180 ;
        RECT 3326.290 390.900 3326.570 391.180 ;
        RECT 3326.910 390.900 3327.190 391.180 ;
        RECT 3327.530 390.900 3327.810 391.180 ;
        RECT 3328.150 390.900 3328.430 391.180 ;
        RECT 3328.770 390.900 3329.050 391.180 ;
        RECT 3329.390 390.900 3329.670 391.180 ;
        RECT 3330.010 390.900 3330.290 391.180 ;
        RECT 3330.630 390.900 3330.910 391.180 ;
        RECT 3331.250 390.900 3331.530 391.180 ;
        RECT 3331.870 390.900 3332.150 391.180 ;
        RECT 3332.490 390.900 3332.770 391.180 ;
        RECT 3333.110 390.900 3333.390 391.180 ;
        RECT 3333.730 390.900 3334.010 391.180 ;
        RECT 3324.430 390.280 3324.710 390.560 ;
        RECT 3325.050 390.280 3325.330 390.560 ;
        RECT 3325.670 390.280 3325.950 390.560 ;
        RECT 3326.290 390.280 3326.570 390.560 ;
        RECT 3326.910 390.280 3327.190 390.560 ;
        RECT 3327.530 390.280 3327.810 390.560 ;
        RECT 3328.150 390.280 3328.430 390.560 ;
        RECT 3328.770 390.280 3329.050 390.560 ;
        RECT 3329.390 390.280 3329.670 390.560 ;
        RECT 3330.010 390.280 3330.290 390.560 ;
        RECT 3330.630 390.280 3330.910 390.560 ;
        RECT 3331.250 390.280 3331.530 390.560 ;
        RECT 3331.870 390.280 3332.150 390.560 ;
        RECT 3332.490 390.280 3332.770 390.560 ;
        RECT 3333.110 390.280 3333.390 390.560 ;
        RECT 3333.730 390.280 3334.010 390.560 ;
        RECT 3324.430 389.660 3324.710 389.940 ;
        RECT 3325.050 389.660 3325.330 389.940 ;
        RECT 3325.670 389.660 3325.950 389.940 ;
        RECT 3326.290 389.660 3326.570 389.940 ;
        RECT 3326.910 389.660 3327.190 389.940 ;
        RECT 3327.530 389.660 3327.810 389.940 ;
        RECT 3328.150 389.660 3328.430 389.940 ;
        RECT 3328.770 389.660 3329.050 389.940 ;
        RECT 3329.390 389.660 3329.670 389.940 ;
        RECT 3330.010 389.660 3330.290 389.940 ;
        RECT 3330.630 389.660 3330.910 389.940 ;
        RECT 3331.250 389.660 3331.530 389.940 ;
        RECT 3331.870 389.660 3332.150 389.940 ;
        RECT 3332.490 389.660 3332.770 389.940 ;
        RECT 3333.110 389.660 3333.390 389.940 ;
        RECT 3333.730 389.660 3334.010 389.940 ;
        RECT 3324.430 389.040 3324.710 389.320 ;
        RECT 3325.050 389.040 3325.330 389.320 ;
        RECT 3325.670 389.040 3325.950 389.320 ;
        RECT 3326.290 389.040 3326.570 389.320 ;
        RECT 3326.910 389.040 3327.190 389.320 ;
        RECT 3327.530 389.040 3327.810 389.320 ;
        RECT 3328.150 389.040 3328.430 389.320 ;
        RECT 3328.770 389.040 3329.050 389.320 ;
        RECT 3329.390 389.040 3329.670 389.320 ;
        RECT 3330.010 389.040 3330.290 389.320 ;
        RECT 3330.630 389.040 3330.910 389.320 ;
        RECT 3331.250 389.040 3331.530 389.320 ;
        RECT 3331.870 389.040 3332.150 389.320 ;
        RECT 3332.490 389.040 3332.770 389.320 ;
        RECT 3333.110 389.040 3333.390 389.320 ;
        RECT 3333.730 389.040 3334.010 389.320 ;
        RECT 3336.280 392.760 3336.560 393.040 ;
        RECT 3336.900 392.760 3337.180 393.040 ;
        RECT 3337.520 392.760 3337.800 393.040 ;
        RECT 3338.140 392.760 3338.420 393.040 ;
        RECT 3338.760 392.760 3339.040 393.040 ;
        RECT 3339.380 392.760 3339.660 393.040 ;
        RECT 3340.000 392.760 3340.280 393.040 ;
        RECT 3340.620 392.760 3340.900 393.040 ;
        RECT 3341.240 392.760 3341.520 393.040 ;
        RECT 3341.860 392.760 3342.140 393.040 ;
        RECT 3342.480 392.760 3342.760 393.040 ;
        RECT 3343.100 392.760 3343.380 393.040 ;
        RECT 3343.720 392.760 3344.000 393.040 ;
        RECT 3344.340 392.760 3344.620 393.040 ;
        RECT 3344.960 392.760 3345.240 393.040 ;
        RECT 3345.580 392.760 3345.860 393.040 ;
        RECT 3336.280 392.140 3336.560 392.420 ;
        RECT 3336.900 392.140 3337.180 392.420 ;
        RECT 3337.520 392.140 3337.800 392.420 ;
        RECT 3338.140 392.140 3338.420 392.420 ;
        RECT 3338.760 392.140 3339.040 392.420 ;
        RECT 3339.380 392.140 3339.660 392.420 ;
        RECT 3340.000 392.140 3340.280 392.420 ;
        RECT 3340.620 392.140 3340.900 392.420 ;
        RECT 3341.240 392.140 3341.520 392.420 ;
        RECT 3341.860 392.140 3342.140 392.420 ;
        RECT 3342.480 392.140 3342.760 392.420 ;
        RECT 3343.100 392.140 3343.380 392.420 ;
        RECT 3343.720 392.140 3344.000 392.420 ;
        RECT 3344.340 392.140 3344.620 392.420 ;
        RECT 3344.960 392.140 3345.240 392.420 ;
        RECT 3345.580 392.140 3345.860 392.420 ;
        RECT 3336.280 391.520 3336.560 391.800 ;
        RECT 3336.900 391.520 3337.180 391.800 ;
        RECT 3337.520 391.520 3337.800 391.800 ;
        RECT 3338.140 391.520 3338.420 391.800 ;
        RECT 3338.760 391.520 3339.040 391.800 ;
        RECT 3339.380 391.520 3339.660 391.800 ;
        RECT 3340.000 391.520 3340.280 391.800 ;
        RECT 3340.620 391.520 3340.900 391.800 ;
        RECT 3341.240 391.520 3341.520 391.800 ;
        RECT 3341.860 391.520 3342.140 391.800 ;
        RECT 3342.480 391.520 3342.760 391.800 ;
        RECT 3343.100 391.520 3343.380 391.800 ;
        RECT 3343.720 391.520 3344.000 391.800 ;
        RECT 3344.340 391.520 3344.620 391.800 ;
        RECT 3344.960 391.520 3345.240 391.800 ;
        RECT 3345.580 391.520 3345.860 391.800 ;
        RECT 3336.280 390.900 3336.560 391.180 ;
        RECT 3336.900 390.900 3337.180 391.180 ;
        RECT 3337.520 390.900 3337.800 391.180 ;
        RECT 3338.140 390.900 3338.420 391.180 ;
        RECT 3338.760 390.900 3339.040 391.180 ;
        RECT 3339.380 390.900 3339.660 391.180 ;
        RECT 3340.000 390.900 3340.280 391.180 ;
        RECT 3340.620 390.900 3340.900 391.180 ;
        RECT 3341.240 390.900 3341.520 391.180 ;
        RECT 3341.860 390.900 3342.140 391.180 ;
        RECT 3342.480 390.900 3342.760 391.180 ;
        RECT 3343.100 390.900 3343.380 391.180 ;
        RECT 3343.720 390.900 3344.000 391.180 ;
        RECT 3344.340 390.900 3344.620 391.180 ;
        RECT 3344.960 390.900 3345.240 391.180 ;
        RECT 3345.580 390.900 3345.860 391.180 ;
        RECT 3336.280 390.280 3336.560 390.560 ;
        RECT 3336.900 390.280 3337.180 390.560 ;
        RECT 3337.520 390.280 3337.800 390.560 ;
        RECT 3338.140 390.280 3338.420 390.560 ;
        RECT 3338.760 390.280 3339.040 390.560 ;
        RECT 3339.380 390.280 3339.660 390.560 ;
        RECT 3340.000 390.280 3340.280 390.560 ;
        RECT 3340.620 390.280 3340.900 390.560 ;
        RECT 3341.240 390.280 3341.520 390.560 ;
        RECT 3341.860 390.280 3342.140 390.560 ;
        RECT 3342.480 390.280 3342.760 390.560 ;
        RECT 3343.100 390.280 3343.380 390.560 ;
        RECT 3343.720 390.280 3344.000 390.560 ;
        RECT 3344.340 390.280 3344.620 390.560 ;
        RECT 3344.960 390.280 3345.240 390.560 ;
        RECT 3345.580 390.280 3345.860 390.560 ;
        RECT 3336.280 389.660 3336.560 389.940 ;
        RECT 3336.900 389.660 3337.180 389.940 ;
        RECT 3337.520 389.660 3337.800 389.940 ;
        RECT 3338.140 389.660 3338.420 389.940 ;
        RECT 3338.760 389.660 3339.040 389.940 ;
        RECT 3339.380 389.660 3339.660 389.940 ;
        RECT 3340.000 389.660 3340.280 389.940 ;
        RECT 3340.620 389.660 3340.900 389.940 ;
        RECT 3341.240 389.660 3341.520 389.940 ;
        RECT 3341.860 389.660 3342.140 389.940 ;
        RECT 3342.480 389.660 3342.760 389.940 ;
        RECT 3343.100 389.660 3343.380 389.940 ;
        RECT 3343.720 389.660 3344.000 389.940 ;
        RECT 3344.340 389.660 3344.620 389.940 ;
        RECT 3344.960 389.660 3345.240 389.940 ;
        RECT 3345.580 389.660 3345.860 389.940 ;
        RECT 3336.280 389.040 3336.560 389.320 ;
        RECT 3336.900 389.040 3337.180 389.320 ;
        RECT 3337.520 389.040 3337.800 389.320 ;
        RECT 3338.140 389.040 3338.420 389.320 ;
        RECT 3338.760 389.040 3339.040 389.320 ;
        RECT 3339.380 389.040 3339.660 389.320 ;
        RECT 3340.000 389.040 3340.280 389.320 ;
        RECT 3340.620 389.040 3340.900 389.320 ;
        RECT 3341.240 389.040 3341.520 389.320 ;
        RECT 3341.860 389.040 3342.140 389.320 ;
        RECT 3342.480 389.040 3342.760 389.320 ;
        RECT 3343.100 389.040 3343.380 389.320 ;
        RECT 3343.720 389.040 3344.000 389.320 ;
        RECT 3344.340 389.040 3344.620 389.320 ;
        RECT 3344.960 389.040 3345.240 389.320 ;
        RECT 3345.580 389.040 3345.860 389.320 ;
        RECT 3349.300 392.760 3349.580 393.040 ;
        RECT 3349.920 392.760 3350.200 393.040 ;
        RECT 3350.540 392.760 3350.820 393.040 ;
        RECT 3351.160 392.760 3351.440 393.040 ;
        RECT 3351.780 392.760 3352.060 393.040 ;
        RECT 3352.400 392.760 3352.680 393.040 ;
        RECT 3353.020 392.760 3353.300 393.040 ;
        RECT 3353.640 392.760 3353.920 393.040 ;
        RECT 3354.260 392.760 3354.540 393.040 ;
        RECT 3354.880 392.760 3355.160 393.040 ;
        RECT 3355.500 392.760 3355.780 393.040 ;
        RECT 3356.120 392.760 3356.400 393.040 ;
        RECT 3356.740 392.760 3357.020 393.040 ;
        RECT 3357.360 392.760 3357.640 393.040 ;
        RECT 3357.980 392.760 3358.260 393.040 ;
        RECT 3349.300 392.140 3349.580 392.420 ;
        RECT 3349.920 392.140 3350.200 392.420 ;
        RECT 3350.540 392.140 3350.820 392.420 ;
        RECT 3351.160 392.140 3351.440 392.420 ;
        RECT 3351.780 392.140 3352.060 392.420 ;
        RECT 3352.400 392.140 3352.680 392.420 ;
        RECT 3353.020 392.140 3353.300 392.420 ;
        RECT 3353.640 392.140 3353.920 392.420 ;
        RECT 3354.260 392.140 3354.540 392.420 ;
        RECT 3354.880 392.140 3355.160 392.420 ;
        RECT 3355.500 392.140 3355.780 392.420 ;
        RECT 3356.120 392.140 3356.400 392.420 ;
        RECT 3356.740 392.140 3357.020 392.420 ;
        RECT 3357.360 392.140 3357.640 392.420 ;
        RECT 3357.980 392.140 3358.260 392.420 ;
        RECT 3349.300 391.520 3349.580 391.800 ;
        RECT 3349.920 391.520 3350.200 391.800 ;
        RECT 3350.540 391.520 3350.820 391.800 ;
        RECT 3351.160 391.520 3351.440 391.800 ;
        RECT 3351.780 391.520 3352.060 391.800 ;
        RECT 3352.400 391.520 3352.680 391.800 ;
        RECT 3353.020 391.520 3353.300 391.800 ;
        RECT 3353.640 391.520 3353.920 391.800 ;
        RECT 3354.260 391.520 3354.540 391.800 ;
        RECT 3354.880 391.520 3355.160 391.800 ;
        RECT 3355.500 391.520 3355.780 391.800 ;
        RECT 3356.120 391.520 3356.400 391.800 ;
        RECT 3356.740 391.520 3357.020 391.800 ;
        RECT 3357.360 391.520 3357.640 391.800 ;
        RECT 3357.980 391.520 3358.260 391.800 ;
        RECT 3349.300 390.900 3349.580 391.180 ;
        RECT 3349.920 390.900 3350.200 391.180 ;
        RECT 3350.540 390.900 3350.820 391.180 ;
        RECT 3351.160 390.900 3351.440 391.180 ;
        RECT 3351.780 390.900 3352.060 391.180 ;
        RECT 3352.400 390.900 3352.680 391.180 ;
        RECT 3353.020 390.900 3353.300 391.180 ;
        RECT 3353.640 390.900 3353.920 391.180 ;
        RECT 3354.260 390.900 3354.540 391.180 ;
        RECT 3354.880 390.900 3355.160 391.180 ;
        RECT 3355.500 390.900 3355.780 391.180 ;
        RECT 3356.120 390.900 3356.400 391.180 ;
        RECT 3356.740 390.900 3357.020 391.180 ;
        RECT 3357.360 390.900 3357.640 391.180 ;
        RECT 3357.980 390.900 3358.260 391.180 ;
        RECT 3349.300 390.280 3349.580 390.560 ;
        RECT 3349.920 390.280 3350.200 390.560 ;
        RECT 3350.540 390.280 3350.820 390.560 ;
        RECT 3351.160 390.280 3351.440 390.560 ;
        RECT 3351.780 390.280 3352.060 390.560 ;
        RECT 3352.400 390.280 3352.680 390.560 ;
        RECT 3353.020 390.280 3353.300 390.560 ;
        RECT 3353.640 390.280 3353.920 390.560 ;
        RECT 3354.260 390.280 3354.540 390.560 ;
        RECT 3354.880 390.280 3355.160 390.560 ;
        RECT 3355.500 390.280 3355.780 390.560 ;
        RECT 3356.120 390.280 3356.400 390.560 ;
        RECT 3356.740 390.280 3357.020 390.560 ;
        RECT 3357.360 390.280 3357.640 390.560 ;
        RECT 3357.980 390.280 3358.260 390.560 ;
        RECT 3349.300 389.660 3349.580 389.940 ;
        RECT 3349.920 389.660 3350.200 389.940 ;
        RECT 3350.540 389.660 3350.820 389.940 ;
        RECT 3351.160 389.660 3351.440 389.940 ;
        RECT 3351.780 389.660 3352.060 389.940 ;
        RECT 3352.400 389.660 3352.680 389.940 ;
        RECT 3353.020 389.660 3353.300 389.940 ;
        RECT 3353.640 389.660 3353.920 389.940 ;
        RECT 3354.260 389.660 3354.540 389.940 ;
        RECT 3354.880 389.660 3355.160 389.940 ;
        RECT 3355.500 389.660 3355.780 389.940 ;
        RECT 3356.120 389.660 3356.400 389.940 ;
        RECT 3356.740 389.660 3357.020 389.940 ;
        RECT 3357.360 389.660 3357.640 389.940 ;
        RECT 3357.980 389.660 3358.260 389.940 ;
        RECT 3349.300 389.040 3349.580 389.320 ;
        RECT 3349.920 389.040 3350.200 389.320 ;
        RECT 3350.540 389.040 3350.820 389.320 ;
        RECT 3351.160 389.040 3351.440 389.320 ;
        RECT 3351.780 389.040 3352.060 389.320 ;
        RECT 3352.400 389.040 3352.680 389.320 ;
        RECT 3353.020 389.040 3353.300 389.320 ;
        RECT 3353.640 389.040 3353.920 389.320 ;
        RECT 3354.260 389.040 3354.540 389.320 ;
        RECT 3354.880 389.040 3355.160 389.320 ;
        RECT 3355.500 389.040 3355.780 389.320 ;
        RECT 3356.120 389.040 3356.400 389.320 ;
        RECT 3356.740 389.040 3357.020 389.320 ;
        RECT 3357.360 389.040 3357.640 389.320 ;
        RECT 3357.980 389.040 3358.260 389.320 ;
        RECT 3497.220 4629.490 3497.500 4629.770 ;
        RECT 3498.720 4629.490 3499.000 4629.770 ;
        RECT 3500.220 4629.490 3500.500 4629.770 ;
        RECT 3497.220 4594.490 3497.500 4594.770 ;
        RECT 3498.720 4594.490 3499.000 4594.770 ;
        RECT 3500.220 4594.490 3500.500 4594.770 ;
        RECT 3497.720 4571.865 3498.000 4572.145 ;
        RECT 3499.220 4571.865 3499.500 4572.145 ;
        RECT 3500.720 4571.865 3501.000 4572.145 ;
        RECT 3497.720 4570.865 3498.000 4571.145 ;
        RECT 3499.220 4570.865 3499.500 4571.145 ;
        RECT 3500.720 4570.865 3501.000 4571.145 ;
        RECT 3497.220 4559.490 3497.500 4559.770 ;
        RECT 3498.720 4559.490 3499.000 4559.770 ;
        RECT 3500.220 4559.490 3500.500 4559.770 ;
        RECT 3497.485 4461.835 3497.765 4462.115 ;
        RECT 3498.985 4461.835 3499.265 4462.115 ;
        RECT 3500.485 4461.835 3500.765 4462.115 ;
        RECT 3496.960 4417.980 3497.240 4418.260 ;
        RECT 3497.580 4417.980 3497.860 4418.260 ;
        RECT 3498.200 4417.980 3498.480 4418.260 ;
        RECT 3498.820 4417.980 3499.100 4418.260 ;
        RECT 3499.440 4417.980 3499.720 4418.260 ;
        RECT 3500.060 4417.980 3500.340 4418.260 ;
        RECT 3500.680 4417.980 3500.960 4418.260 ;
        RECT 3496.960 4417.360 3497.240 4417.640 ;
        RECT 3497.580 4417.360 3497.860 4417.640 ;
        RECT 3498.200 4417.360 3498.480 4417.640 ;
        RECT 3498.820 4417.360 3499.100 4417.640 ;
        RECT 3499.440 4417.360 3499.720 4417.640 ;
        RECT 3500.060 4417.360 3500.340 4417.640 ;
        RECT 3500.680 4417.360 3500.960 4417.640 ;
        RECT 3496.960 4416.740 3497.240 4417.020 ;
        RECT 3497.580 4416.740 3497.860 4417.020 ;
        RECT 3498.200 4416.740 3498.480 4417.020 ;
        RECT 3498.820 4416.740 3499.100 4417.020 ;
        RECT 3499.440 4416.740 3499.720 4417.020 ;
        RECT 3500.060 4416.740 3500.340 4417.020 ;
        RECT 3500.680 4416.740 3500.960 4417.020 ;
        RECT 3496.960 4416.120 3497.240 4416.400 ;
        RECT 3497.580 4416.120 3497.860 4416.400 ;
        RECT 3498.200 4416.120 3498.480 4416.400 ;
        RECT 3498.820 4416.120 3499.100 4416.400 ;
        RECT 3499.440 4416.120 3499.720 4416.400 ;
        RECT 3500.060 4416.120 3500.340 4416.400 ;
        RECT 3500.680 4416.120 3500.960 4416.400 ;
        RECT 3496.960 4415.500 3497.240 4415.780 ;
        RECT 3497.580 4415.500 3497.860 4415.780 ;
        RECT 3498.200 4415.500 3498.480 4415.780 ;
        RECT 3498.820 4415.500 3499.100 4415.780 ;
        RECT 3499.440 4415.500 3499.720 4415.780 ;
        RECT 3500.060 4415.500 3500.340 4415.780 ;
        RECT 3500.680 4415.500 3500.960 4415.780 ;
        RECT 3496.960 4414.880 3497.240 4415.160 ;
        RECT 3497.580 4414.880 3497.860 4415.160 ;
        RECT 3498.200 4414.880 3498.480 4415.160 ;
        RECT 3498.820 4414.880 3499.100 4415.160 ;
        RECT 3499.440 4414.880 3499.720 4415.160 ;
        RECT 3500.060 4414.880 3500.340 4415.160 ;
        RECT 3500.680 4414.880 3500.960 4415.160 ;
        RECT 3496.960 4414.260 3497.240 4414.540 ;
        RECT 3497.580 4414.260 3497.860 4414.540 ;
        RECT 3498.200 4414.260 3498.480 4414.540 ;
        RECT 3498.820 4414.260 3499.100 4414.540 ;
        RECT 3499.440 4414.260 3499.720 4414.540 ;
        RECT 3500.060 4414.260 3500.340 4414.540 ;
        RECT 3500.680 4414.260 3500.960 4414.540 ;
        RECT 3496.960 4413.640 3497.240 4413.920 ;
        RECT 3497.580 4413.640 3497.860 4413.920 ;
        RECT 3498.200 4413.640 3498.480 4413.920 ;
        RECT 3498.820 4413.640 3499.100 4413.920 ;
        RECT 3499.440 4413.640 3499.720 4413.920 ;
        RECT 3500.060 4413.640 3500.340 4413.920 ;
        RECT 3500.680 4413.640 3500.960 4413.920 ;
        RECT 3496.960 4413.020 3497.240 4413.300 ;
        RECT 3497.580 4413.020 3497.860 4413.300 ;
        RECT 3498.200 4413.020 3498.480 4413.300 ;
        RECT 3498.820 4413.020 3499.100 4413.300 ;
        RECT 3499.440 4413.020 3499.720 4413.300 ;
        RECT 3500.060 4413.020 3500.340 4413.300 ;
        RECT 3500.680 4413.020 3500.960 4413.300 ;
        RECT 3496.960 4412.400 3497.240 4412.680 ;
        RECT 3497.580 4412.400 3497.860 4412.680 ;
        RECT 3498.200 4412.400 3498.480 4412.680 ;
        RECT 3498.820 4412.400 3499.100 4412.680 ;
        RECT 3499.440 4412.400 3499.720 4412.680 ;
        RECT 3500.060 4412.400 3500.340 4412.680 ;
        RECT 3500.680 4412.400 3500.960 4412.680 ;
        RECT 3496.960 4411.780 3497.240 4412.060 ;
        RECT 3497.580 4411.780 3497.860 4412.060 ;
        RECT 3498.200 4411.780 3498.480 4412.060 ;
        RECT 3498.820 4411.780 3499.100 4412.060 ;
        RECT 3499.440 4411.780 3499.720 4412.060 ;
        RECT 3500.060 4411.780 3500.340 4412.060 ;
        RECT 3500.680 4411.780 3500.960 4412.060 ;
        RECT 3496.960 4411.160 3497.240 4411.440 ;
        RECT 3497.580 4411.160 3497.860 4411.440 ;
        RECT 3498.200 4411.160 3498.480 4411.440 ;
        RECT 3498.820 4411.160 3499.100 4411.440 ;
        RECT 3499.440 4411.160 3499.720 4411.440 ;
        RECT 3500.060 4411.160 3500.340 4411.440 ;
        RECT 3500.680 4411.160 3500.960 4411.440 ;
        RECT 3496.960 4410.540 3497.240 4410.820 ;
        RECT 3497.580 4410.540 3497.860 4410.820 ;
        RECT 3498.200 4410.540 3498.480 4410.820 ;
        RECT 3498.820 4410.540 3499.100 4410.820 ;
        RECT 3499.440 4410.540 3499.720 4410.820 ;
        RECT 3500.060 4410.540 3500.340 4410.820 ;
        RECT 3500.680 4410.540 3500.960 4410.820 ;
        RECT 3496.960 4409.920 3497.240 4410.200 ;
        RECT 3497.580 4409.920 3497.860 4410.200 ;
        RECT 3498.200 4409.920 3498.480 4410.200 ;
        RECT 3498.820 4409.920 3499.100 4410.200 ;
        RECT 3499.440 4409.920 3499.720 4410.200 ;
        RECT 3500.060 4409.920 3500.340 4410.200 ;
        RECT 3500.680 4409.920 3500.960 4410.200 ;
        RECT 3496.960 4409.300 3497.240 4409.580 ;
        RECT 3497.580 4409.300 3497.860 4409.580 ;
        RECT 3498.200 4409.300 3498.480 4409.580 ;
        RECT 3498.820 4409.300 3499.100 4409.580 ;
        RECT 3499.440 4409.300 3499.720 4409.580 ;
        RECT 3500.060 4409.300 3500.340 4409.580 ;
        RECT 3500.680 4409.300 3500.960 4409.580 ;
        RECT 3539.350 4418.010 3539.630 4418.290 ;
        RECT 3539.350 4417.390 3539.630 4417.670 ;
        RECT 3539.350 4416.770 3539.630 4417.050 ;
        RECT 3539.350 4416.150 3539.630 4416.430 ;
        RECT 3539.350 4415.530 3539.630 4415.810 ;
        RECT 3539.350 4414.910 3539.630 4415.190 ;
        RECT 3539.350 4414.290 3539.630 4414.570 ;
        RECT 3539.350 4413.670 3539.630 4413.950 ;
        RECT 3539.350 4413.050 3539.630 4413.330 ;
        RECT 3539.350 4412.430 3539.630 4412.710 ;
        RECT 3539.350 4411.810 3539.630 4412.090 ;
        RECT 3539.350 4411.190 3539.630 4411.470 ;
        RECT 3539.350 4410.570 3539.630 4410.850 ;
        RECT 3539.350 4409.950 3539.630 4410.230 ;
        RECT 3539.350 4409.330 3539.630 4409.610 ;
        RECT 3496.960 4405.580 3497.240 4405.860 ;
        RECT 3497.580 4405.580 3497.860 4405.860 ;
        RECT 3498.200 4405.580 3498.480 4405.860 ;
        RECT 3498.820 4405.580 3499.100 4405.860 ;
        RECT 3499.440 4405.580 3499.720 4405.860 ;
        RECT 3500.060 4405.580 3500.340 4405.860 ;
        RECT 3500.680 4405.580 3500.960 4405.860 ;
        RECT 3496.960 4404.960 3497.240 4405.240 ;
        RECT 3497.580 4404.960 3497.860 4405.240 ;
        RECT 3498.200 4404.960 3498.480 4405.240 ;
        RECT 3498.820 4404.960 3499.100 4405.240 ;
        RECT 3499.440 4404.960 3499.720 4405.240 ;
        RECT 3500.060 4404.960 3500.340 4405.240 ;
        RECT 3500.680 4404.960 3500.960 4405.240 ;
        RECT 3496.960 4404.340 3497.240 4404.620 ;
        RECT 3497.580 4404.340 3497.860 4404.620 ;
        RECT 3498.200 4404.340 3498.480 4404.620 ;
        RECT 3498.820 4404.340 3499.100 4404.620 ;
        RECT 3499.440 4404.340 3499.720 4404.620 ;
        RECT 3500.060 4404.340 3500.340 4404.620 ;
        RECT 3500.680 4404.340 3500.960 4404.620 ;
        RECT 3496.960 4403.720 3497.240 4404.000 ;
        RECT 3497.580 4403.720 3497.860 4404.000 ;
        RECT 3498.200 4403.720 3498.480 4404.000 ;
        RECT 3498.820 4403.720 3499.100 4404.000 ;
        RECT 3499.440 4403.720 3499.720 4404.000 ;
        RECT 3500.060 4403.720 3500.340 4404.000 ;
        RECT 3500.680 4403.720 3500.960 4404.000 ;
        RECT 3496.960 4403.100 3497.240 4403.380 ;
        RECT 3497.580 4403.100 3497.860 4403.380 ;
        RECT 3498.200 4403.100 3498.480 4403.380 ;
        RECT 3498.820 4403.100 3499.100 4403.380 ;
        RECT 3499.440 4403.100 3499.720 4403.380 ;
        RECT 3500.060 4403.100 3500.340 4403.380 ;
        RECT 3500.680 4403.100 3500.960 4403.380 ;
        RECT 3496.960 4402.480 3497.240 4402.760 ;
        RECT 3497.580 4402.480 3497.860 4402.760 ;
        RECT 3498.200 4402.480 3498.480 4402.760 ;
        RECT 3498.820 4402.480 3499.100 4402.760 ;
        RECT 3499.440 4402.480 3499.720 4402.760 ;
        RECT 3500.060 4402.480 3500.340 4402.760 ;
        RECT 3500.680 4402.480 3500.960 4402.760 ;
        RECT 3496.960 4401.860 3497.240 4402.140 ;
        RECT 3497.580 4401.860 3497.860 4402.140 ;
        RECT 3498.200 4401.860 3498.480 4402.140 ;
        RECT 3498.820 4401.860 3499.100 4402.140 ;
        RECT 3499.440 4401.860 3499.720 4402.140 ;
        RECT 3500.060 4401.860 3500.340 4402.140 ;
        RECT 3500.680 4401.860 3500.960 4402.140 ;
        RECT 3496.960 4401.240 3497.240 4401.520 ;
        RECT 3497.580 4401.240 3497.860 4401.520 ;
        RECT 3498.200 4401.240 3498.480 4401.520 ;
        RECT 3498.820 4401.240 3499.100 4401.520 ;
        RECT 3499.440 4401.240 3499.720 4401.520 ;
        RECT 3500.060 4401.240 3500.340 4401.520 ;
        RECT 3500.680 4401.240 3500.960 4401.520 ;
        RECT 3496.960 4400.620 3497.240 4400.900 ;
        RECT 3497.580 4400.620 3497.860 4400.900 ;
        RECT 3498.200 4400.620 3498.480 4400.900 ;
        RECT 3498.820 4400.620 3499.100 4400.900 ;
        RECT 3499.440 4400.620 3499.720 4400.900 ;
        RECT 3500.060 4400.620 3500.340 4400.900 ;
        RECT 3500.680 4400.620 3500.960 4400.900 ;
        RECT 3496.960 4400.000 3497.240 4400.280 ;
        RECT 3497.580 4400.000 3497.860 4400.280 ;
        RECT 3498.200 4400.000 3498.480 4400.280 ;
        RECT 3498.820 4400.000 3499.100 4400.280 ;
        RECT 3499.440 4400.000 3499.720 4400.280 ;
        RECT 3500.060 4400.000 3500.340 4400.280 ;
        RECT 3500.680 4400.000 3500.960 4400.280 ;
        RECT 3496.960 4399.380 3497.240 4399.660 ;
        RECT 3497.580 4399.380 3497.860 4399.660 ;
        RECT 3498.200 4399.380 3498.480 4399.660 ;
        RECT 3498.820 4399.380 3499.100 4399.660 ;
        RECT 3499.440 4399.380 3499.720 4399.660 ;
        RECT 3500.060 4399.380 3500.340 4399.660 ;
        RECT 3500.680 4399.380 3500.960 4399.660 ;
        RECT 3496.960 4398.760 3497.240 4399.040 ;
        RECT 3497.580 4398.760 3497.860 4399.040 ;
        RECT 3498.200 4398.760 3498.480 4399.040 ;
        RECT 3498.820 4398.760 3499.100 4399.040 ;
        RECT 3499.440 4398.760 3499.720 4399.040 ;
        RECT 3500.060 4398.760 3500.340 4399.040 ;
        RECT 3500.680 4398.760 3500.960 4399.040 ;
        RECT 3496.960 4398.140 3497.240 4398.420 ;
        RECT 3497.580 4398.140 3497.860 4398.420 ;
        RECT 3498.200 4398.140 3498.480 4398.420 ;
        RECT 3498.820 4398.140 3499.100 4398.420 ;
        RECT 3499.440 4398.140 3499.720 4398.420 ;
        RECT 3500.060 4398.140 3500.340 4398.420 ;
        RECT 3500.680 4398.140 3500.960 4398.420 ;
        RECT 3496.960 4397.520 3497.240 4397.800 ;
        RECT 3497.580 4397.520 3497.860 4397.800 ;
        RECT 3498.200 4397.520 3498.480 4397.800 ;
        RECT 3498.820 4397.520 3499.100 4397.800 ;
        RECT 3499.440 4397.520 3499.720 4397.800 ;
        RECT 3500.060 4397.520 3500.340 4397.800 ;
        RECT 3500.680 4397.520 3500.960 4397.800 ;
        RECT 3496.960 4396.900 3497.240 4397.180 ;
        RECT 3497.580 4396.900 3497.860 4397.180 ;
        RECT 3498.200 4396.900 3498.480 4397.180 ;
        RECT 3498.820 4396.900 3499.100 4397.180 ;
        RECT 3499.440 4396.900 3499.720 4397.180 ;
        RECT 3500.060 4396.900 3500.340 4397.180 ;
        RECT 3500.680 4396.900 3500.960 4397.180 ;
        RECT 3496.960 4396.280 3497.240 4396.560 ;
        RECT 3497.580 4396.280 3497.860 4396.560 ;
        RECT 3498.200 4396.280 3498.480 4396.560 ;
        RECT 3498.820 4396.280 3499.100 4396.560 ;
        RECT 3499.440 4396.280 3499.720 4396.560 ;
        RECT 3500.060 4396.280 3500.340 4396.560 ;
        RECT 3500.680 4396.280 3500.960 4396.560 ;
        RECT 3539.350 4405.610 3539.630 4405.890 ;
        RECT 3539.350 4404.990 3539.630 4405.270 ;
        RECT 3539.350 4404.370 3539.630 4404.650 ;
        RECT 3539.350 4403.750 3539.630 4404.030 ;
        RECT 3539.350 4403.130 3539.630 4403.410 ;
        RECT 3539.350 4402.510 3539.630 4402.790 ;
        RECT 3539.350 4401.890 3539.630 4402.170 ;
        RECT 3539.350 4401.270 3539.630 4401.550 ;
        RECT 3539.350 4400.650 3539.630 4400.930 ;
        RECT 3539.350 4400.030 3539.630 4400.310 ;
        RECT 3539.350 4399.410 3539.630 4399.690 ;
        RECT 3539.350 4398.790 3539.630 4399.070 ;
        RECT 3539.350 4398.170 3539.630 4398.450 ;
        RECT 3539.350 4397.550 3539.630 4397.830 ;
        RECT 3539.350 4396.930 3539.630 4397.210 ;
        RECT 3539.350 4396.310 3539.630 4396.590 ;
        RECT 3496.960 4393.730 3497.240 4394.010 ;
        RECT 3497.580 4393.730 3497.860 4394.010 ;
        RECT 3498.200 4393.730 3498.480 4394.010 ;
        RECT 3498.820 4393.730 3499.100 4394.010 ;
        RECT 3499.440 4393.730 3499.720 4394.010 ;
        RECT 3500.060 4393.730 3500.340 4394.010 ;
        RECT 3500.680 4393.730 3500.960 4394.010 ;
        RECT 3496.960 4393.110 3497.240 4393.390 ;
        RECT 3497.580 4393.110 3497.860 4393.390 ;
        RECT 3498.200 4393.110 3498.480 4393.390 ;
        RECT 3498.820 4393.110 3499.100 4393.390 ;
        RECT 3499.440 4393.110 3499.720 4393.390 ;
        RECT 3500.060 4393.110 3500.340 4393.390 ;
        RECT 3500.680 4393.110 3500.960 4393.390 ;
        RECT 3496.960 4392.490 3497.240 4392.770 ;
        RECT 3497.580 4392.490 3497.860 4392.770 ;
        RECT 3498.200 4392.490 3498.480 4392.770 ;
        RECT 3498.820 4392.490 3499.100 4392.770 ;
        RECT 3499.440 4392.490 3499.720 4392.770 ;
        RECT 3500.060 4392.490 3500.340 4392.770 ;
        RECT 3500.680 4392.490 3500.960 4392.770 ;
        RECT 3496.960 4391.870 3497.240 4392.150 ;
        RECT 3497.580 4391.870 3497.860 4392.150 ;
        RECT 3498.200 4391.870 3498.480 4392.150 ;
        RECT 3498.820 4391.870 3499.100 4392.150 ;
        RECT 3499.440 4391.870 3499.720 4392.150 ;
        RECT 3500.060 4391.870 3500.340 4392.150 ;
        RECT 3500.680 4391.870 3500.960 4392.150 ;
        RECT 3496.960 4391.250 3497.240 4391.530 ;
        RECT 3497.580 4391.250 3497.860 4391.530 ;
        RECT 3498.200 4391.250 3498.480 4391.530 ;
        RECT 3498.820 4391.250 3499.100 4391.530 ;
        RECT 3499.440 4391.250 3499.720 4391.530 ;
        RECT 3500.060 4391.250 3500.340 4391.530 ;
        RECT 3500.680 4391.250 3500.960 4391.530 ;
        RECT 3496.960 4390.630 3497.240 4390.910 ;
        RECT 3497.580 4390.630 3497.860 4390.910 ;
        RECT 3498.200 4390.630 3498.480 4390.910 ;
        RECT 3498.820 4390.630 3499.100 4390.910 ;
        RECT 3499.440 4390.630 3499.720 4390.910 ;
        RECT 3500.060 4390.630 3500.340 4390.910 ;
        RECT 3500.680 4390.630 3500.960 4390.910 ;
        RECT 3496.960 4390.010 3497.240 4390.290 ;
        RECT 3497.580 4390.010 3497.860 4390.290 ;
        RECT 3498.200 4390.010 3498.480 4390.290 ;
        RECT 3498.820 4390.010 3499.100 4390.290 ;
        RECT 3499.440 4390.010 3499.720 4390.290 ;
        RECT 3500.060 4390.010 3500.340 4390.290 ;
        RECT 3500.680 4390.010 3500.960 4390.290 ;
        RECT 3496.960 4389.390 3497.240 4389.670 ;
        RECT 3497.580 4389.390 3497.860 4389.670 ;
        RECT 3498.200 4389.390 3498.480 4389.670 ;
        RECT 3498.820 4389.390 3499.100 4389.670 ;
        RECT 3499.440 4389.390 3499.720 4389.670 ;
        RECT 3500.060 4389.390 3500.340 4389.670 ;
        RECT 3500.680 4389.390 3500.960 4389.670 ;
        RECT 3496.960 4388.770 3497.240 4389.050 ;
        RECT 3497.580 4388.770 3497.860 4389.050 ;
        RECT 3498.200 4388.770 3498.480 4389.050 ;
        RECT 3498.820 4388.770 3499.100 4389.050 ;
        RECT 3499.440 4388.770 3499.720 4389.050 ;
        RECT 3500.060 4388.770 3500.340 4389.050 ;
        RECT 3500.680 4388.770 3500.960 4389.050 ;
        RECT 3496.960 4388.150 3497.240 4388.430 ;
        RECT 3497.580 4388.150 3497.860 4388.430 ;
        RECT 3498.200 4388.150 3498.480 4388.430 ;
        RECT 3498.820 4388.150 3499.100 4388.430 ;
        RECT 3499.440 4388.150 3499.720 4388.430 ;
        RECT 3500.060 4388.150 3500.340 4388.430 ;
        RECT 3500.680 4388.150 3500.960 4388.430 ;
        RECT 3496.960 4387.530 3497.240 4387.810 ;
        RECT 3497.580 4387.530 3497.860 4387.810 ;
        RECT 3498.200 4387.530 3498.480 4387.810 ;
        RECT 3498.820 4387.530 3499.100 4387.810 ;
        RECT 3499.440 4387.530 3499.720 4387.810 ;
        RECT 3500.060 4387.530 3500.340 4387.810 ;
        RECT 3500.680 4387.530 3500.960 4387.810 ;
        RECT 3496.960 4386.910 3497.240 4387.190 ;
        RECT 3497.580 4386.910 3497.860 4387.190 ;
        RECT 3498.200 4386.910 3498.480 4387.190 ;
        RECT 3498.820 4386.910 3499.100 4387.190 ;
        RECT 3499.440 4386.910 3499.720 4387.190 ;
        RECT 3500.060 4386.910 3500.340 4387.190 ;
        RECT 3500.680 4386.910 3500.960 4387.190 ;
        RECT 3496.960 4386.290 3497.240 4386.570 ;
        RECT 3497.580 4386.290 3497.860 4386.570 ;
        RECT 3498.200 4386.290 3498.480 4386.570 ;
        RECT 3498.820 4386.290 3499.100 4386.570 ;
        RECT 3499.440 4386.290 3499.720 4386.570 ;
        RECT 3500.060 4386.290 3500.340 4386.570 ;
        RECT 3500.680 4386.290 3500.960 4386.570 ;
        RECT 3496.960 4385.670 3497.240 4385.950 ;
        RECT 3497.580 4385.670 3497.860 4385.950 ;
        RECT 3498.200 4385.670 3498.480 4385.950 ;
        RECT 3498.820 4385.670 3499.100 4385.950 ;
        RECT 3499.440 4385.670 3499.720 4385.950 ;
        RECT 3500.060 4385.670 3500.340 4385.950 ;
        RECT 3500.680 4385.670 3500.960 4385.950 ;
        RECT 3496.960 4385.050 3497.240 4385.330 ;
        RECT 3497.580 4385.050 3497.860 4385.330 ;
        RECT 3498.200 4385.050 3498.480 4385.330 ;
        RECT 3498.820 4385.050 3499.100 4385.330 ;
        RECT 3499.440 4385.050 3499.720 4385.330 ;
        RECT 3500.060 4385.050 3500.340 4385.330 ;
        RECT 3500.680 4385.050 3500.960 4385.330 ;
        RECT 3496.960 4384.430 3497.240 4384.710 ;
        RECT 3497.580 4384.430 3497.860 4384.710 ;
        RECT 3498.200 4384.430 3498.480 4384.710 ;
        RECT 3498.820 4384.430 3499.100 4384.710 ;
        RECT 3499.440 4384.430 3499.720 4384.710 ;
        RECT 3500.060 4384.430 3500.340 4384.710 ;
        RECT 3500.680 4384.430 3500.960 4384.710 ;
        RECT 3539.350 4393.760 3539.630 4394.040 ;
        RECT 3539.350 4393.140 3539.630 4393.420 ;
        RECT 3539.350 4392.520 3539.630 4392.800 ;
        RECT 3539.350 4391.900 3539.630 4392.180 ;
        RECT 3539.350 4391.280 3539.630 4391.560 ;
        RECT 3539.350 4390.660 3539.630 4390.940 ;
        RECT 3539.350 4390.040 3539.630 4390.320 ;
        RECT 3539.350 4389.420 3539.630 4389.700 ;
        RECT 3539.350 4388.800 3539.630 4389.080 ;
        RECT 3539.350 4388.180 3539.630 4388.460 ;
        RECT 3539.350 4387.560 3539.630 4387.840 ;
        RECT 3539.350 4386.940 3539.630 4387.220 ;
        RECT 3539.350 4386.320 3539.630 4386.600 ;
        RECT 3539.350 4385.700 3539.630 4385.980 ;
        RECT 3539.350 4385.080 3539.630 4385.360 ;
        RECT 3539.350 4384.460 3539.630 4384.740 ;
        RECT 3496.960 4380.200 3497.240 4380.480 ;
        RECT 3497.580 4380.200 3497.860 4380.480 ;
        RECT 3498.200 4380.200 3498.480 4380.480 ;
        RECT 3498.820 4380.200 3499.100 4380.480 ;
        RECT 3499.440 4380.200 3499.720 4380.480 ;
        RECT 3500.060 4380.200 3500.340 4380.480 ;
        RECT 3500.680 4380.200 3500.960 4380.480 ;
        RECT 3496.960 4379.580 3497.240 4379.860 ;
        RECT 3497.580 4379.580 3497.860 4379.860 ;
        RECT 3498.200 4379.580 3498.480 4379.860 ;
        RECT 3498.820 4379.580 3499.100 4379.860 ;
        RECT 3499.440 4379.580 3499.720 4379.860 ;
        RECT 3500.060 4379.580 3500.340 4379.860 ;
        RECT 3500.680 4379.580 3500.960 4379.860 ;
        RECT 3496.960 4378.960 3497.240 4379.240 ;
        RECT 3497.580 4378.960 3497.860 4379.240 ;
        RECT 3498.200 4378.960 3498.480 4379.240 ;
        RECT 3498.820 4378.960 3499.100 4379.240 ;
        RECT 3499.440 4378.960 3499.720 4379.240 ;
        RECT 3500.060 4378.960 3500.340 4379.240 ;
        RECT 3500.680 4378.960 3500.960 4379.240 ;
        RECT 3496.960 4378.340 3497.240 4378.620 ;
        RECT 3497.580 4378.340 3497.860 4378.620 ;
        RECT 3498.200 4378.340 3498.480 4378.620 ;
        RECT 3498.820 4378.340 3499.100 4378.620 ;
        RECT 3499.440 4378.340 3499.720 4378.620 ;
        RECT 3500.060 4378.340 3500.340 4378.620 ;
        RECT 3500.680 4378.340 3500.960 4378.620 ;
        RECT 3496.960 4377.720 3497.240 4378.000 ;
        RECT 3497.580 4377.720 3497.860 4378.000 ;
        RECT 3498.200 4377.720 3498.480 4378.000 ;
        RECT 3498.820 4377.720 3499.100 4378.000 ;
        RECT 3499.440 4377.720 3499.720 4378.000 ;
        RECT 3500.060 4377.720 3500.340 4378.000 ;
        RECT 3500.680 4377.720 3500.960 4378.000 ;
        RECT 3496.960 4377.100 3497.240 4377.380 ;
        RECT 3497.580 4377.100 3497.860 4377.380 ;
        RECT 3498.200 4377.100 3498.480 4377.380 ;
        RECT 3498.820 4377.100 3499.100 4377.380 ;
        RECT 3499.440 4377.100 3499.720 4377.380 ;
        RECT 3500.060 4377.100 3500.340 4377.380 ;
        RECT 3500.680 4377.100 3500.960 4377.380 ;
        RECT 3496.960 4376.480 3497.240 4376.760 ;
        RECT 3497.580 4376.480 3497.860 4376.760 ;
        RECT 3498.200 4376.480 3498.480 4376.760 ;
        RECT 3498.820 4376.480 3499.100 4376.760 ;
        RECT 3499.440 4376.480 3499.720 4376.760 ;
        RECT 3500.060 4376.480 3500.340 4376.760 ;
        RECT 3500.680 4376.480 3500.960 4376.760 ;
        RECT 3496.960 4375.860 3497.240 4376.140 ;
        RECT 3497.580 4375.860 3497.860 4376.140 ;
        RECT 3498.200 4375.860 3498.480 4376.140 ;
        RECT 3498.820 4375.860 3499.100 4376.140 ;
        RECT 3499.440 4375.860 3499.720 4376.140 ;
        RECT 3500.060 4375.860 3500.340 4376.140 ;
        RECT 3500.680 4375.860 3500.960 4376.140 ;
        RECT 3496.960 4375.240 3497.240 4375.520 ;
        RECT 3497.580 4375.240 3497.860 4375.520 ;
        RECT 3498.200 4375.240 3498.480 4375.520 ;
        RECT 3498.820 4375.240 3499.100 4375.520 ;
        RECT 3499.440 4375.240 3499.720 4375.520 ;
        RECT 3500.060 4375.240 3500.340 4375.520 ;
        RECT 3500.680 4375.240 3500.960 4375.520 ;
        RECT 3496.960 4374.620 3497.240 4374.900 ;
        RECT 3497.580 4374.620 3497.860 4374.900 ;
        RECT 3498.200 4374.620 3498.480 4374.900 ;
        RECT 3498.820 4374.620 3499.100 4374.900 ;
        RECT 3499.440 4374.620 3499.720 4374.900 ;
        RECT 3500.060 4374.620 3500.340 4374.900 ;
        RECT 3500.680 4374.620 3500.960 4374.900 ;
        RECT 3496.960 4374.000 3497.240 4374.280 ;
        RECT 3497.580 4374.000 3497.860 4374.280 ;
        RECT 3498.200 4374.000 3498.480 4374.280 ;
        RECT 3498.820 4374.000 3499.100 4374.280 ;
        RECT 3499.440 4374.000 3499.720 4374.280 ;
        RECT 3500.060 4374.000 3500.340 4374.280 ;
        RECT 3500.680 4374.000 3500.960 4374.280 ;
        RECT 3496.960 4373.380 3497.240 4373.660 ;
        RECT 3497.580 4373.380 3497.860 4373.660 ;
        RECT 3498.200 4373.380 3498.480 4373.660 ;
        RECT 3498.820 4373.380 3499.100 4373.660 ;
        RECT 3499.440 4373.380 3499.720 4373.660 ;
        RECT 3500.060 4373.380 3500.340 4373.660 ;
        RECT 3500.680 4373.380 3500.960 4373.660 ;
        RECT 3496.960 4372.760 3497.240 4373.040 ;
        RECT 3497.580 4372.760 3497.860 4373.040 ;
        RECT 3498.200 4372.760 3498.480 4373.040 ;
        RECT 3498.820 4372.760 3499.100 4373.040 ;
        RECT 3499.440 4372.760 3499.720 4373.040 ;
        RECT 3500.060 4372.760 3500.340 4373.040 ;
        RECT 3500.680 4372.760 3500.960 4373.040 ;
        RECT 3496.960 4372.140 3497.240 4372.420 ;
        RECT 3497.580 4372.140 3497.860 4372.420 ;
        RECT 3498.200 4372.140 3498.480 4372.420 ;
        RECT 3498.820 4372.140 3499.100 4372.420 ;
        RECT 3499.440 4372.140 3499.720 4372.420 ;
        RECT 3500.060 4372.140 3500.340 4372.420 ;
        RECT 3500.680 4372.140 3500.960 4372.420 ;
        RECT 3496.960 4371.520 3497.240 4371.800 ;
        RECT 3497.580 4371.520 3497.860 4371.800 ;
        RECT 3498.200 4371.520 3498.480 4371.800 ;
        RECT 3498.820 4371.520 3499.100 4371.800 ;
        RECT 3499.440 4371.520 3499.720 4371.800 ;
        RECT 3500.060 4371.520 3500.340 4371.800 ;
        RECT 3500.680 4371.520 3500.960 4371.800 ;
        RECT 3496.960 4370.900 3497.240 4371.180 ;
        RECT 3497.580 4370.900 3497.860 4371.180 ;
        RECT 3498.200 4370.900 3498.480 4371.180 ;
        RECT 3498.820 4370.900 3499.100 4371.180 ;
        RECT 3499.440 4370.900 3499.720 4371.180 ;
        RECT 3500.060 4370.900 3500.340 4371.180 ;
        RECT 3500.680 4370.900 3500.960 4371.180 ;
        RECT 3539.350 4380.230 3539.630 4380.510 ;
        RECT 3539.350 4379.610 3539.630 4379.890 ;
        RECT 3539.350 4378.990 3539.630 4379.270 ;
        RECT 3539.350 4378.370 3539.630 4378.650 ;
        RECT 3539.350 4377.750 3539.630 4378.030 ;
        RECT 3539.350 4377.130 3539.630 4377.410 ;
        RECT 3539.350 4376.510 3539.630 4376.790 ;
        RECT 3539.350 4375.890 3539.630 4376.170 ;
        RECT 3539.350 4375.270 3539.630 4375.550 ;
        RECT 3539.350 4374.650 3539.630 4374.930 ;
        RECT 3539.350 4374.030 3539.630 4374.310 ;
        RECT 3539.350 4373.410 3539.630 4373.690 ;
        RECT 3539.350 4372.790 3539.630 4373.070 ;
        RECT 3539.350 4372.170 3539.630 4372.450 ;
        RECT 3539.350 4371.550 3539.630 4371.830 ;
        RECT 3539.350 4370.930 3539.630 4371.210 ;
        RECT 3496.960 4368.350 3497.240 4368.630 ;
        RECT 3497.580 4368.350 3497.860 4368.630 ;
        RECT 3498.200 4368.350 3498.480 4368.630 ;
        RECT 3498.820 4368.350 3499.100 4368.630 ;
        RECT 3499.440 4368.350 3499.720 4368.630 ;
        RECT 3500.060 4368.350 3500.340 4368.630 ;
        RECT 3500.680 4368.350 3500.960 4368.630 ;
        RECT 3496.960 4367.730 3497.240 4368.010 ;
        RECT 3497.580 4367.730 3497.860 4368.010 ;
        RECT 3498.200 4367.730 3498.480 4368.010 ;
        RECT 3498.820 4367.730 3499.100 4368.010 ;
        RECT 3499.440 4367.730 3499.720 4368.010 ;
        RECT 3500.060 4367.730 3500.340 4368.010 ;
        RECT 3500.680 4367.730 3500.960 4368.010 ;
        RECT 3496.960 4367.110 3497.240 4367.390 ;
        RECT 3497.580 4367.110 3497.860 4367.390 ;
        RECT 3498.200 4367.110 3498.480 4367.390 ;
        RECT 3498.820 4367.110 3499.100 4367.390 ;
        RECT 3499.440 4367.110 3499.720 4367.390 ;
        RECT 3500.060 4367.110 3500.340 4367.390 ;
        RECT 3500.680 4367.110 3500.960 4367.390 ;
        RECT 3496.960 4366.490 3497.240 4366.770 ;
        RECT 3497.580 4366.490 3497.860 4366.770 ;
        RECT 3498.200 4366.490 3498.480 4366.770 ;
        RECT 3498.820 4366.490 3499.100 4366.770 ;
        RECT 3499.440 4366.490 3499.720 4366.770 ;
        RECT 3500.060 4366.490 3500.340 4366.770 ;
        RECT 3500.680 4366.490 3500.960 4366.770 ;
        RECT 3496.960 4365.870 3497.240 4366.150 ;
        RECT 3497.580 4365.870 3497.860 4366.150 ;
        RECT 3498.200 4365.870 3498.480 4366.150 ;
        RECT 3498.820 4365.870 3499.100 4366.150 ;
        RECT 3499.440 4365.870 3499.720 4366.150 ;
        RECT 3500.060 4365.870 3500.340 4366.150 ;
        RECT 3500.680 4365.870 3500.960 4366.150 ;
        RECT 3496.960 4365.250 3497.240 4365.530 ;
        RECT 3497.580 4365.250 3497.860 4365.530 ;
        RECT 3498.200 4365.250 3498.480 4365.530 ;
        RECT 3498.820 4365.250 3499.100 4365.530 ;
        RECT 3499.440 4365.250 3499.720 4365.530 ;
        RECT 3500.060 4365.250 3500.340 4365.530 ;
        RECT 3500.680 4365.250 3500.960 4365.530 ;
        RECT 3496.960 4364.630 3497.240 4364.910 ;
        RECT 3497.580 4364.630 3497.860 4364.910 ;
        RECT 3498.200 4364.630 3498.480 4364.910 ;
        RECT 3498.820 4364.630 3499.100 4364.910 ;
        RECT 3499.440 4364.630 3499.720 4364.910 ;
        RECT 3500.060 4364.630 3500.340 4364.910 ;
        RECT 3500.680 4364.630 3500.960 4364.910 ;
        RECT 3496.960 4364.010 3497.240 4364.290 ;
        RECT 3497.580 4364.010 3497.860 4364.290 ;
        RECT 3498.200 4364.010 3498.480 4364.290 ;
        RECT 3498.820 4364.010 3499.100 4364.290 ;
        RECT 3499.440 4364.010 3499.720 4364.290 ;
        RECT 3500.060 4364.010 3500.340 4364.290 ;
        RECT 3500.680 4364.010 3500.960 4364.290 ;
        RECT 3496.960 4363.390 3497.240 4363.670 ;
        RECT 3497.580 4363.390 3497.860 4363.670 ;
        RECT 3498.200 4363.390 3498.480 4363.670 ;
        RECT 3498.820 4363.390 3499.100 4363.670 ;
        RECT 3499.440 4363.390 3499.720 4363.670 ;
        RECT 3500.060 4363.390 3500.340 4363.670 ;
        RECT 3500.680 4363.390 3500.960 4363.670 ;
        RECT 3496.960 4362.770 3497.240 4363.050 ;
        RECT 3497.580 4362.770 3497.860 4363.050 ;
        RECT 3498.200 4362.770 3498.480 4363.050 ;
        RECT 3498.820 4362.770 3499.100 4363.050 ;
        RECT 3499.440 4362.770 3499.720 4363.050 ;
        RECT 3500.060 4362.770 3500.340 4363.050 ;
        RECT 3500.680 4362.770 3500.960 4363.050 ;
        RECT 3496.960 4362.150 3497.240 4362.430 ;
        RECT 3497.580 4362.150 3497.860 4362.430 ;
        RECT 3498.200 4362.150 3498.480 4362.430 ;
        RECT 3498.820 4362.150 3499.100 4362.430 ;
        RECT 3499.440 4362.150 3499.720 4362.430 ;
        RECT 3500.060 4362.150 3500.340 4362.430 ;
        RECT 3500.680 4362.150 3500.960 4362.430 ;
        RECT 3496.960 4361.530 3497.240 4361.810 ;
        RECT 3497.580 4361.530 3497.860 4361.810 ;
        RECT 3498.200 4361.530 3498.480 4361.810 ;
        RECT 3498.820 4361.530 3499.100 4361.810 ;
        RECT 3499.440 4361.530 3499.720 4361.810 ;
        RECT 3500.060 4361.530 3500.340 4361.810 ;
        RECT 3500.680 4361.530 3500.960 4361.810 ;
        RECT 3496.960 4360.910 3497.240 4361.190 ;
        RECT 3497.580 4360.910 3497.860 4361.190 ;
        RECT 3498.200 4360.910 3498.480 4361.190 ;
        RECT 3498.820 4360.910 3499.100 4361.190 ;
        RECT 3499.440 4360.910 3499.720 4361.190 ;
        RECT 3500.060 4360.910 3500.340 4361.190 ;
        RECT 3500.680 4360.910 3500.960 4361.190 ;
        RECT 3496.960 4360.290 3497.240 4360.570 ;
        RECT 3497.580 4360.290 3497.860 4360.570 ;
        RECT 3498.200 4360.290 3498.480 4360.570 ;
        RECT 3498.820 4360.290 3499.100 4360.570 ;
        RECT 3499.440 4360.290 3499.720 4360.570 ;
        RECT 3500.060 4360.290 3500.340 4360.570 ;
        RECT 3500.680 4360.290 3500.960 4360.570 ;
        RECT 3496.960 4359.670 3497.240 4359.950 ;
        RECT 3497.580 4359.670 3497.860 4359.950 ;
        RECT 3498.200 4359.670 3498.480 4359.950 ;
        RECT 3498.820 4359.670 3499.100 4359.950 ;
        RECT 3499.440 4359.670 3499.720 4359.950 ;
        RECT 3500.060 4359.670 3500.340 4359.950 ;
        RECT 3500.680 4359.670 3500.960 4359.950 ;
        RECT 3496.960 4359.050 3497.240 4359.330 ;
        RECT 3497.580 4359.050 3497.860 4359.330 ;
        RECT 3498.200 4359.050 3498.480 4359.330 ;
        RECT 3498.820 4359.050 3499.100 4359.330 ;
        RECT 3499.440 4359.050 3499.720 4359.330 ;
        RECT 3500.060 4359.050 3500.340 4359.330 ;
        RECT 3500.680 4359.050 3500.960 4359.330 ;
        RECT 3539.350 4368.380 3539.630 4368.660 ;
        RECT 3539.350 4367.760 3539.630 4368.040 ;
        RECT 3539.350 4367.140 3539.630 4367.420 ;
        RECT 3539.350 4366.520 3539.630 4366.800 ;
        RECT 3539.350 4365.900 3539.630 4366.180 ;
        RECT 3539.350 4365.280 3539.630 4365.560 ;
        RECT 3539.350 4364.660 3539.630 4364.940 ;
        RECT 3539.350 4364.040 3539.630 4364.320 ;
        RECT 3539.350 4363.420 3539.630 4363.700 ;
        RECT 3539.350 4362.800 3539.630 4363.080 ;
        RECT 3539.350 4362.180 3539.630 4362.460 ;
        RECT 3539.350 4361.560 3539.630 4361.840 ;
        RECT 3539.350 4360.940 3539.630 4361.220 ;
        RECT 3539.350 4360.320 3539.630 4360.600 ;
        RECT 3539.350 4359.700 3539.630 4359.980 ;
        RECT 3539.350 4359.080 3539.630 4359.360 ;
        RECT 3496.960 4355.330 3497.240 4355.610 ;
        RECT 3497.580 4355.330 3497.860 4355.610 ;
        RECT 3498.200 4355.330 3498.480 4355.610 ;
        RECT 3498.820 4355.330 3499.100 4355.610 ;
        RECT 3499.440 4355.330 3499.720 4355.610 ;
        RECT 3500.060 4355.330 3500.340 4355.610 ;
        RECT 3500.680 4355.330 3500.960 4355.610 ;
        RECT 3496.960 4354.710 3497.240 4354.990 ;
        RECT 3497.580 4354.710 3497.860 4354.990 ;
        RECT 3498.200 4354.710 3498.480 4354.990 ;
        RECT 3498.820 4354.710 3499.100 4354.990 ;
        RECT 3499.440 4354.710 3499.720 4354.990 ;
        RECT 3500.060 4354.710 3500.340 4354.990 ;
        RECT 3500.680 4354.710 3500.960 4354.990 ;
        RECT 3496.960 4354.090 3497.240 4354.370 ;
        RECT 3497.580 4354.090 3497.860 4354.370 ;
        RECT 3498.200 4354.090 3498.480 4354.370 ;
        RECT 3498.820 4354.090 3499.100 4354.370 ;
        RECT 3499.440 4354.090 3499.720 4354.370 ;
        RECT 3500.060 4354.090 3500.340 4354.370 ;
        RECT 3500.680 4354.090 3500.960 4354.370 ;
        RECT 3496.960 4353.470 3497.240 4353.750 ;
        RECT 3497.580 4353.470 3497.860 4353.750 ;
        RECT 3498.200 4353.470 3498.480 4353.750 ;
        RECT 3498.820 4353.470 3499.100 4353.750 ;
        RECT 3499.440 4353.470 3499.720 4353.750 ;
        RECT 3500.060 4353.470 3500.340 4353.750 ;
        RECT 3500.680 4353.470 3500.960 4353.750 ;
        RECT 3496.960 4352.850 3497.240 4353.130 ;
        RECT 3497.580 4352.850 3497.860 4353.130 ;
        RECT 3498.200 4352.850 3498.480 4353.130 ;
        RECT 3498.820 4352.850 3499.100 4353.130 ;
        RECT 3499.440 4352.850 3499.720 4353.130 ;
        RECT 3500.060 4352.850 3500.340 4353.130 ;
        RECT 3500.680 4352.850 3500.960 4353.130 ;
        RECT 3496.960 4352.230 3497.240 4352.510 ;
        RECT 3497.580 4352.230 3497.860 4352.510 ;
        RECT 3498.200 4352.230 3498.480 4352.510 ;
        RECT 3498.820 4352.230 3499.100 4352.510 ;
        RECT 3499.440 4352.230 3499.720 4352.510 ;
        RECT 3500.060 4352.230 3500.340 4352.510 ;
        RECT 3500.680 4352.230 3500.960 4352.510 ;
        RECT 3496.960 4351.610 3497.240 4351.890 ;
        RECT 3497.580 4351.610 3497.860 4351.890 ;
        RECT 3498.200 4351.610 3498.480 4351.890 ;
        RECT 3498.820 4351.610 3499.100 4351.890 ;
        RECT 3499.440 4351.610 3499.720 4351.890 ;
        RECT 3500.060 4351.610 3500.340 4351.890 ;
        RECT 3500.680 4351.610 3500.960 4351.890 ;
        RECT 3496.960 4350.990 3497.240 4351.270 ;
        RECT 3497.580 4350.990 3497.860 4351.270 ;
        RECT 3498.200 4350.990 3498.480 4351.270 ;
        RECT 3498.820 4350.990 3499.100 4351.270 ;
        RECT 3499.440 4350.990 3499.720 4351.270 ;
        RECT 3500.060 4350.990 3500.340 4351.270 ;
        RECT 3500.680 4350.990 3500.960 4351.270 ;
        RECT 3496.960 4350.370 3497.240 4350.650 ;
        RECT 3497.580 4350.370 3497.860 4350.650 ;
        RECT 3498.200 4350.370 3498.480 4350.650 ;
        RECT 3498.820 4350.370 3499.100 4350.650 ;
        RECT 3499.440 4350.370 3499.720 4350.650 ;
        RECT 3500.060 4350.370 3500.340 4350.650 ;
        RECT 3500.680 4350.370 3500.960 4350.650 ;
        RECT 3496.960 4349.750 3497.240 4350.030 ;
        RECT 3497.580 4349.750 3497.860 4350.030 ;
        RECT 3498.200 4349.750 3498.480 4350.030 ;
        RECT 3498.820 4349.750 3499.100 4350.030 ;
        RECT 3499.440 4349.750 3499.720 4350.030 ;
        RECT 3500.060 4349.750 3500.340 4350.030 ;
        RECT 3500.680 4349.750 3500.960 4350.030 ;
        RECT 3496.960 4349.130 3497.240 4349.410 ;
        RECT 3497.580 4349.130 3497.860 4349.410 ;
        RECT 3498.200 4349.130 3498.480 4349.410 ;
        RECT 3498.820 4349.130 3499.100 4349.410 ;
        RECT 3499.440 4349.130 3499.720 4349.410 ;
        RECT 3500.060 4349.130 3500.340 4349.410 ;
        RECT 3500.680 4349.130 3500.960 4349.410 ;
        RECT 3496.960 4348.510 3497.240 4348.790 ;
        RECT 3497.580 4348.510 3497.860 4348.790 ;
        RECT 3498.200 4348.510 3498.480 4348.790 ;
        RECT 3498.820 4348.510 3499.100 4348.790 ;
        RECT 3499.440 4348.510 3499.720 4348.790 ;
        RECT 3500.060 4348.510 3500.340 4348.790 ;
        RECT 3500.680 4348.510 3500.960 4348.790 ;
        RECT 3496.960 4347.890 3497.240 4348.170 ;
        RECT 3497.580 4347.890 3497.860 4348.170 ;
        RECT 3498.200 4347.890 3498.480 4348.170 ;
        RECT 3498.820 4347.890 3499.100 4348.170 ;
        RECT 3499.440 4347.890 3499.720 4348.170 ;
        RECT 3500.060 4347.890 3500.340 4348.170 ;
        RECT 3500.680 4347.890 3500.960 4348.170 ;
        RECT 3496.960 4347.270 3497.240 4347.550 ;
        RECT 3497.580 4347.270 3497.860 4347.550 ;
        RECT 3498.200 4347.270 3498.480 4347.550 ;
        RECT 3498.820 4347.270 3499.100 4347.550 ;
        RECT 3499.440 4347.270 3499.720 4347.550 ;
        RECT 3500.060 4347.270 3500.340 4347.550 ;
        RECT 3500.680 4347.270 3500.960 4347.550 ;
        RECT 3496.960 4346.650 3497.240 4346.930 ;
        RECT 3497.580 4346.650 3497.860 4346.930 ;
        RECT 3498.200 4346.650 3498.480 4346.930 ;
        RECT 3498.820 4346.650 3499.100 4346.930 ;
        RECT 3499.440 4346.650 3499.720 4346.930 ;
        RECT 3500.060 4346.650 3500.340 4346.930 ;
        RECT 3500.680 4346.650 3500.960 4346.930 ;
        RECT 3539.350 4355.390 3539.630 4355.670 ;
        RECT 3539.350 4354.770 3539.630 4355.050 ;
        RECT 3539.350 4354.150 3539.630 4354.430 ;
        RECT 3539.350 4353.530 3539.630 4353.810 ;
        RECT 3539.350 4352.910 3539.630 4353.190 ;
        RECT 3539.350 4352.290 3539.630 4352.570 ;
        RECT 3539.350 4351.670 3539.630 4351.950 ;
        RECT 3539.350 4351.050 3539.630 4351.330 ;
        RECT 3539.350 4350.430 3539.630 4350.710 ;
        RECT 3539.350 4349.810 3539.630 4350.090 ;
        RECT 3539.350 4349.190 3539.630 4349.470 ;
        RECT 3539.350 4348.570 3539.630 4348.850 ;
        RECT 3539.350 4347.950 3539.630 4348.230 ;
        RECT 3539.350 4347.330 3539.630 4347.610 ;
        RECT 3539.350 4346.710 3539.630 4346.990 ;
        RECT 3497.720 4211.865 3498.000 4212.145 ;
        RECT 3499.220 4211.865 3499.500 4212.145 ;
        RECT 3500.720 4211.865 3501.000 4212.145 ;
        RECT 3497.720 4210.865 3498.000 4211.145 ;
        RECT 3499.220 4210.865 3499.500 4211.145 ;
        RECT 3500.720 4210.865 3501.000 4211.145 ;
        RECT 3497.220 4199.490 3497.500 4199.770 ;
        RECT 3498.720 4199.490 3499.000 4199.770 ;
        RECT 3500.220 4199.490 3500.500 4199.770 ;
        RECT 3497.220 4164.490 3497.500 4164.770 ;
        RECT 3498.720 4164.490 3499.000 4164.770 ;
        RECT 3500.220 4164.490 3500.500 4164.770 ;
        RECT 3497.220 4129.490 3497.500 4129.770 ;
        RECT 3498.720 4129.490 3499.000 4129.770 ;
        RECT 3500.220 4129.490 3500.500 4129.770 ;
        RECT 3497.485 4031.835 3497.765 4032.115 ;
        RECT 3498.985 4031.835 3499.265 4032.115 ;
        RECT 3500.485 4031.835 3500.765 4032.115 ;
        RECT 3496.960 3987.980 3497.240 3988.260 ;
        RECT 3497.580 3987.980 3497.860 3988.260 ;
        RECT 3498.200 3987.980 3498.480 3988.260 ;
        RECT 3498.820 3987.980 3499.100 3988.260 ;
        RECT 3499.440 3987.980 3499.720 3988.260 ;
        RECT 3500.060 3987.980 3500.340 3988.260 ;
        RECT 3500.680 3987.980 3500.960 3988.260 ;
        RECT 3496.960 3987.360 3497.240 3987.640 ;
        RECT 3497.580 3987.360 3497.860 3987.640 ;
        RECT 3498.200 3987.360 3498.480 3987.640 ;
        RECT 3498.820 3987.360 3499.100 3987.640 ;
        RECT 3499.440 3987.360 3499.720 3987.640 ;
        RECT 3500.060 3987.360 3500.340 3987.640 ;
        RECT 3500.680 3987.360 3500.960 3987.640 ;
        RECT 3496.960 3986.740 3497.240 3987.020 ;
        RECT 3497.580 3986.740 3497.860 3987.020 ;
        RECT 3498.200 3986.740 3498.480 3987.020 ;
        RECT 3498.820 3986.740 3499.100 3987.020 ;
        RECT 3499.440 3986.740 3499.720 3987.020 ;
        RECT 3500.060 3986.740 3500.340 3987.020 ;
        RECT 3500.680 3986.740 3500.960 3987.020 ;
        RECT 3496.960 3986.120 3497.240 3986.400 ;
        RECT 3497.580 3986.120 3497.860 3986.400 ;
        RECT 3498.200 3986.120 3498.480 3986.400 ;
        RECT 3498.820 3986.120 3499.100 3986.400 ;
        RECT 3499.440 3986.120 3499.720 3986.400 ;
        RECT 3500.060 3986.120 3500.340 3986.400 ;
        RECT 3500.680 3986.120 3500.960 3986.400 ;
        RECT 3496.960 3985.500 3497.240 3985.780 ;
        RECT 3497.580 3985.500 3497.860 3985.780 ;
        RECT 3498.200 3985.500 3498.480 3985.780 ;
        RECT 3498.820 3985.500 3499.100 3985.780 ;
        RECT 3499.440 3985.500 3499.720 3985.780 ;
        RECT 3500.060 3985.500 3500.340 3985.780 ;
        RECT 3500.680 3985.500 3500.960 3985.780 ;
        RECT 3496.960 3984.880 3497.240 3985.160 ;
        RECT 3497.580 3984.880 3497.860 3985.160 ;
        RECT 3498.200 3984.880 3498.480 3985.160 ;
        RECT 3498.820 3984.880 3499.100 3985.160 ;
        RECT 3499.440 3984.880 3499.720 3985.160 ;
        RECT 3500.060 3984.880 3500.340 3985.160 ;
        RECT 3500.680 3984.880 3500.960 3985.160 ;
        RECT 3496.960 3984.260 3497.240 3984.540 ;
        RECT 3497.580 3984.260 3497.860 3984.540 ;
        RECT 3498.200 3984.260 3498.480 3984.540 ;
        RECT 3498.820 3984.260 3499.100 3984.540 ;
        RECT 3499.440 3984.260 3499.720 3984.540 ;
        RECT 3500.060 3984.260 3500.340 3984.540 ;
        RECT 3500.680 3984.260 3500.960 3984.540 ;
        RECT 3496.960 3983.640 3497.240 3983.920 ;
        RECT 3497.580 3983.640 3497.860 3983.920 ;
        RECT 3498.200 3983.640 3498.480 3983.920 ;
        RECT 3498.820 3983.640 3499.100 3983.920 ;
        RECT 3499.440 3983.640 3499.720 3983.920 ;
        RECT 3500.060 3983.640 3500.340 3983.920 ;
        RECT 3500.680 3983.640 3500.960 3983.920 ;
        RECT 3496.960 3983.020 3497.240 3983.300 ;
        RECT 3497.580 3983.020 3497.860 3983.300 ;
        RECT 3498.200 3983.020 3498.480 3983.300 ;
        RECT 3498.820 3983.020 3499.100 3983.300 ;
        RECT 3499.440 3983.020 3499.720 3983.300 ;
        RECT 3500.060 3983.020 3500.340 3983.300 ;
        RECT 3500.680 3983.020 3500.960 3983.300 ;
        RECT 3496.960 3982.400 3497.240 3982.680 ;
        RECT 3497.580 3982.400 3497.860 3982.680 ;
        RECT 3498.200 3982.400 3498.480 3982.680 ;
        RECT 3498.820 3982.400 3499.100 3982.680 ;
        RECT 3499.440 3982.400 3499.720 3982.680 ;
        RECT 3500.060 3982.400 3500.340 3982.680 ;
        RECT 3500.680 3982.400 3500.960 3982.680 ;
        RECT 3496.960 3981.780 3497.240 3982.060 ;
        RECT 3497.580 3981.780 3497.860 3982.060 ;
        RECT 3498.200 3981.780 3498.480 3982.060 ;
        RECT 3498.820 3981.780 3499.100 3982.060 ;
        RECT 3499.440 3981.780 3499.720 3982.060 ;
        RECT 3500.060 3981.780 3500.340 3982.060 ;
        RECT 3500.680 3981.780 3500.960 3982.060 ;
        RECT 3496.960 3981.160 3497.240 3981.440 ;
        RECT 3497.580 3981.160 3497.860 3981.440 ;
        RECT 3498.200 3981.160 3498.480 3981.440 ;
        RECT 3498.820 3981.160 3499.100 3981.440 ;
        RECT 3499.440 3981.160 3499.720 3981.440 ;
        RECT 3500.060 3981.160 3500.340 3981.440 ;
        RECT 3500.680 3981.160 3500.960 3981.440 ;
        RECT 3496.960 3980.540 3497.240 3980.820 ;
        RECT 3497.580 3980.540 3497.860 3980.820 ;
        RECT 3498.200 3980.540 3498.480 3980.820 ;
        RECT 3498.820 3980.540 3499.100 3980.820 ;
        RECT 3499.440 3980.540 3499.720 3980.820 ;
        RECT 3500.060 3980.540 3500.340 3980.820 ;
        RECT 3500.680 3980.540 3500.960 3980.820 ;
        RECT 3496.960 3979.920 3497.240 3980.200 ;
        RECT 3497.580 3979.920 3497.860 3980.200 ;
        RECT 3498.200 3979.920 3498.480 3980.200 ;
        RECT 3498.820 3979.920 3499.100 3980.200 ;
        RECT 3499.440 3979.920 3499.720 3980.200 ;
        RECT 3500.060 3979.920 3500.340 3980.200 ;
        RECT 3500.680 3979.920 3500.960 3980.200 ;
        RECT 3496.960 3979.300 3497.240 3979.580 ;
        RECT 3497.580 3979.300 3497.860 3979.580 ;
        RECT 3498.200 3979.300 3498.480 3979.580 ;
        RECT 3498.820 3979.300 3499.100 3979.580 ;
        RECT 3499.440 3979.300 3499.720 3979.580 ;
        RECT 3500.060 3979.300 3500.340 3979.580 ;
        RECT 3500.680 3979.300 3500.960 3979.580 ;
        RECT 3539.350 3988.010 3539.630 3988.290 ;
        RECT 3539.350 3987.390 3539.630 3987.670 ;
        RECT 3539.350 3986.770 3539.630 3987.050 ;
        RECT 3539.350 3986.150 3539.630 3986.430 ;
        RECT 3539.350 3985.530 3539.630 3985.810 ;
        RECT 3539.350 3984.910 3539.630 3985.190 ;
        RECT 3539.350 3984.290 3539.630 3984.570 ;
        RECT 3539.350 3983.670 3539.630 3983.950 ;
        RECT 3539.350 3983.050 3539.630 3983.330 ;
        RECT 3539.350 3982.430 3539.630 3982.710 ;
        RECT 3539.350 3981.810 3539.630 3982.090 ;
        RECT 3539.350 3981.190 3539.630 3981.470 ;
        RECT 3539.350 3980.570 3539.630 3980.850 ;
        RECT 3539.350 3979.950 3539.630 3980.230 ;
        RECT 3539.350 3979.330 3539.630 3979.610 ;
        RECT 3496.960 3975.580 3497.240 3975.860 ;
        RECT 3497.580 3975.580 3497.860 3975.860 ;
        RECT 3498.200 3975.580 3498.480 3975.860 ;
        RECT 3498.820 3975.580 3499.100 3975.860 ;
        RECT 3499.440 3975.580 3499.720 3975.860 ;
        RECT 3500.060 3975.580 3500.340 3975.860 ;
        RECT 3500.680 3975.580 3500.960 3975.860 ;
        RECT 3496.960 3974.960 3497.240 3975.240 ;
        RECT 3497.580 3974.960 3497.860 3975.240 ;
        RECT 3498.200 3974.960 3498.480 3975.240 ;
        RECT 3498.820 3974.960 3499.100 3975.240 ;
        RECT 3499.440 3974.960 3499.720 3975.240 ;
        RECT 3500.060 3974.960 3500.340 3975.240 ;
        RECT 3500.680 3974.960 3500.960 3975.240 ;
        RECT 3496.960 3974.340 3497.240 3974.620 ;
        RECT 3497.580 3974.340 3497.860 3974.620 ;
        RECT 3498.200 3974.340 3498.480 3974.620 ;
        RECT 3498.820 3974.340 3499.100 3974.620 ;
        RECT 3499.440 3974.340 3499.720 3974.620 ;
        RECT 3500.060 3974.340 3500.340 3974.620 ;
        RECT 3500.680 3974.340 3500.960 3974.620 ;
        RECT 3496.960 3973.720 3497.240 3974.000 ;
        RECT 3497.580 3973.720 3497.860 3974.000 ;
        RECT 3498.200 3973.720 3498.480 3974.000 ;
        RECT 3498.820 3973.720 3499.100 3974.000 ;
        RECT 3499.440 3973.720 3499.720 3974.000 ;
        RECT 3500.060 3973.720 3500.340 3974.000 ;
        RECT 3500.680 3973.720 3500.960 3974.000 ;
        RECT 3496.960 3973.100 3497.240 3973.380 ;
        RECT 3497.580 3973.100 3497.860 3973.380 ;
        RECT 3498.200 3973.100 3498.480 3973.380 ;
        RECT 3498.820 3973.100 3499.100 3973.380 ;
        RECT 3499.440 3973.100 3499.720 3973.380 ;
        RECT 3500.060 3973.100 3500.340 3973.380 ;
        RECT 3500.680 3973.100 3500.960 3973.380 ;
        RECT 3496.960 3972.480 3497.240 3972.760 ;
        RECT 3497.580 3972.480 3497.860 3972.760 ;
        RECT 3498.200 3972.480 3498.480 3972.760 ;
        RECT 3498.820 3972.480 3499.100 3972.760 ;
        RECT 3499.440 3972.480 3499.720 3972.760 ;
        RECT 3500.060 3972.480 3500.340 3972.760 ;
        RECT 3500.680 3972.480 3500.960 3972.760 ;
        RECT 3496.960 3971.860 3497.240 3972.140 ;
        RECT 3497.580 3971.860 3497.860 3972.140 ;
        RECT 3498.200 3971.860 3498.480 3972.140 ;
        RECT 3498.820 3971.860 3499.100 3972.140 ;
        RECT 3499.440 3971.860 3499.720 3972.140 ;
        RECT 3500.060 3971.860 3500.340 3972.140 ;
        RECT 3500.680 3971.860 3500.960 3972.140 ;
        RECT 3496.960 3971.240 3497.240 3971.520 ;
        RECT 3497.580 3971.240 3497.860 3971.520 ;
        RECT 3498.200 3971.240 3498.480 3971.520 ;
        RECT 3498.820 3971.240 3499.100 3971.520 ;
        RECT 3499.440 3971.240 3499.720 3971.520 ;
        RECT 3500.060 3971.240 3500.340 3971.520 ;
        RECT 3500.680 3971.240 3500.960 3971.520 ;
        RECT 3496.960 3970.620 3497.240 3970.900 ;
        RECT 3497.580 3970.620 3497.860 3970.900 ;
        RECT 3498.200 3970.620 3498.480 3970.900 ;
        RECT 3498.820 3970.620 3499.100 3970.900 ;
        RECT 3499.440 3970.620 3499.720 3970.900 ;
        RECT 3500.060 3970.620 3500.340 3970.900 ;
        RECT 3500.680 3970.620 3500.960 3970.900 ;
        RECT 3496.960 3970.000 3497.240 3970.280 ;
        RECT 3497.580 3970.000 3497.860 3970.280 ;
        RECT 3498.200 3970.000 3498.480 3970.280 ;
        RECT 3498.820 3970.000 3499.100 3970.280 ;
        RECT 3499.440 3970.000 3499.720 3970.280 ;
        RECT 3500.060 3970.000 3500.340 3970.280 ;
        RECT 3500.680 3970.000 3500.960 3970.280 ;
        RECT 3496.960 3969.380 3497.240 3969.660 ;
        RECT 3497.580 3969.380 3497.860 3969.660 ;
        RECT 3498.200 3969.380 3498.480 3969.660 ;
        RECT 3498.820 3969.380 3499.100 3969.660 ;
        RECT 3499.440 3969.380 3499.720 3969.660 ;
        RECT 3500.060 3969.380 3500.340 3969.660 ;
        RECT 3500.680 3969.380 3500.960 3969.660 ;
        RECT 3496.960 3968.760 3497.240 3969.040 ;
        RECT 3497.580 3968.760 3497.860 3969.040 ;
        RECT 3498.200 3968.760 3498.480 3969.040 ;
        RECT 3498.820 3968.760 3499.100 3969.040 ;
        RECT 3499.440 3968.760 3499.720 3969.040 ;
        RECT 3500.060 3968.760 3500.340 3969.040 ;
        RECT 3500.680 3968.760 3500.960 3969.040 ;
        RECT 3496.960 3968.140 3497.240 3968.420 ;
        RECT 3497.580 3968.140 3497.860 3968.420 ;
        RECT 3498.200 3968.140 3498.480 3968.420 ;
        RECT 3498.820 3968.140 3499.100 3968.420 ;
        RECT 3499.440 3968.140 3499.720 3968.420 ;
        RECT 3500.060 3968.140 3500.340 3968.420 ;
        RECT 3500.680 3968.140 3500.960 3968.420 ;
        RECT 3496.960 3967.520 3497.240 3967.800 ;
        RECT 3497.580 3967.520 3497.860 3967.800 ;
        RECT 3498.200 3967.520 3498.480 3967.800 ;
        RECT 3498.820 3967.520 3499.100 3967.800 ;
        RECT 3499.440 3967.520 3499.720 3967.800 ;
        RECT 3500.060 3967.520 3500.340 3967.800 ;
        RECT 3500.680 3967.520 3500.960 3967.800 ;
        RECT 3496.960 3966.900 3497.240 3967.180 ;
        RECT 3497.580 3966.900 3497.860 3967.180 ;
        RECT 3498.200 3966.900 3498.480 3967.180 ;
        RECT 3498.820 3966.900 3499.100 3967.180 ;
        RECT 3499.440 3966.900 3499.720 3967.180 ;
        RECT 3500.060 3966.900 3500.340 3967.180 ;
        RECT 3500.680 3966.900 3500.960 3967.180 ;
        RECT 3496.960 3966.280 3497.240 3966.560 ;
        RECT 3497.580 3966.280 3497.860 3966.560 ;
        RECT 3498.200 3966.280 3498.480 3966.560 ;
        RECT 3498.820 3966.280 3499.100 3966.560 ;
        RECT 3499.440 3966.280 3499.720 3966.560 ;
        RECT 3500.060 3966.280 3500.340 3966.560 ;
        RECT 3500.680 3966.280 3500.960 3966.560 ;
        RECT 3539.350 3975.610 3539.630 3975.890 ;
        RECT 3539.350 3974.990 3539.630 3975.270 ;
        RECT 3539.350 3974.370 3539.630 3974.650 ;
        RECT 3539.350 3973.750 3539.630 3974.030 ;
        RECT 3539.350 3973.130 3539.630 3973.410 ;
        RECT 3539.350 3972.510 3539.630 3972.790 ;
        RECT 3539.350 3971.890 3539.630 3972.170 ;
        RECT 3539.350 3971.270 3539.630 3971.550 ;
        RECT 3539.350 3970.650 3539.630 3970.930 ;
        RECT 3539.350 3970.030 3539.630 3970.310 ;
        RECT 3539.350 3969.410 3539.630 3969.690 ;
        RECT 3539.350 3968.790 3539.630 3969.070 ;
        RECT 3539.350 3968.170 3539.630 3968.450 ;
        RECT 3539.350 3967.550 3539.630 3967.830 ;
        RECT 3539.350 3966.930 3539.630 3967.210 ;
        RECT 3539.350 3966.310 3539.630 3966.590 ;
        RECT 3496.960 3963.730 3497.240 3964.010 ;
        RECT 3497.580 3963.730 3497.860 3964.010 ;
        RECT 3498.200 3963.730 3498.480 3964.010 ;
        RECT 3498.820 3963.730 3499.100 3964.010 ;
        RECT 3499.440 3963.730 3499.720 3964.010 ;
        RECT 3500.060 3963.730 3500.340 3964.010 ;
        RECT 3500.680 3963.730 3500.960 3964.010 ;
        RECT 3496.960 3963.110 3497.240 3963.390 ;
        RECT 3497.580 3963.110 3497.860 3963.390 ;
        RECT 3498.200 3963.110 3498.480 3963.390 ;
        RECT 3498.820 3963.110 3499.100 3963.390 ;
        RECT 3499.440 3963.110 3499.720 3963.390 ;
        RECT 3500.060 3963.110 3500.340 3963.390 ;
        RECT 3500.680 3963.110 3500.960 3963.390 ;
        RECT 3496.960 3962.490 3497.240 3962.770 ;
        RECT 3497.580 3962.490 3497.860 3962.770 ;
        RECT 3498.200 3962.490 3498.480 3962.770 ;
        RECT 3498.820 3962.490 3499.100 3962.770 ;
        RECT 3499.440 3962.490 3499.720 3962.770 ;
        RECT 3500.060 3962.490 3500.340 3962.770 ;
        RECT 3500.680 3962.490 3500.960 3962.770 ;
        RECT 3496.960 3961.870 3497.240 3962.150 ;
        RECT 3497.580 3961.870 3497.860 3962.150 ;
        RECT 3498.200 3961.870 3498.480 3962.150 ;
        RECT 3498.820 3961.870 3499.100 3962.150 ;
        RECT 3499.440 3961.870 3499.720 3962.150 ;
        RECT 3500.060 3961.870 3500.340 3962.150 ;
        RECT 3500.680 3961.870 3500.960 3962.150 ;
        RECT 3496.960 3961.250 3497.240 3961.530 ;
        RECT 3497.580 3961.250 3497.860 3961.530 ;
        RECT 3498.200 3961.250 3498.480 3961.530 ;
        RECT 3498.820 3961.250 3499.100 3961.530 ;
        RECT 3499.440 3961.250 3499.720 3961.530 ;
        RECT 3500.060 3961.250 3500.340 3961.530 ;
        RECT 3500.680 3961.250 3500.960 3961.530 ;
        RECT 3496.960 3960.630 3497.240 3960.910 ;
        RECT 3497.580 3960.630 3497.860 3960.910 ;
        RECT 3498.200 3960.630 3498.480 3960.910 ;
        RECT 3498.820 3960.630 3499.100 3960.910 ;
        RECT 3499.440 3960.630 3499.720 3960.910 ;
        RECT 3500.060 3960.630 3500.340 3960.910 ;
        RECT 3500.680 3960.630 3500.960 3960.910 ;
        RECT 3496.960 3960.010 3497.240 3960.290 ;
        RECT 3497.580 3960.010 3497.860 3960.290 ;
        RECT 3498.200 3960.010 3498.480 3960.290 ;
        RECT 3498.820 3960.010 3499.100 3960.290 ;
        RECT 3499.440 3960.010 3499.720 3960.290 ;
        RECT 3500.060 3960.010 3500.340 3960.290 ;
        RECT 3500.680 3960.010 3500.960 3960.290 ;
        RECT 3496.960 3959.390 3497.240 3959.670 ;
        RECT 3497.580 3959.390 3497.860 3959.670 ;
        RECT 3498.200 3959.390 3498.480 3959.670 ;
        RECT 3498.820 3959.390 3499.100 3959.670 ;
        RECT 3499.440 3959.390 3499.720 3959.670 ;
        RECT 3500.060 3959.390 3500.340 3959.670 ;
        RECT 3500.680 3959.390 3500.960 3959.670 ;
        RECT 3496.960 3958.770 3497.240 3959.050 ;
        RECT 3497.580 3958.770 3497.860 3959.050 ;
        RECT 3498.200 3958.770 3498.480 3959.050 ;
        RECT 3498.820 3958.770 3499.100 3959.050 ;
        RECT 3499.440 3958.770 3499.720 3959.050 ;
        RECT 3500.060 3958.770 3500.340 3959.050 ;
        RECT 3500.680 3958.770 3500.960 3959.050 ;
        RECT 3496.960 3958.150 3497.240 3958.430 ;
        RECT 3497.580 3958.150 3497.860 3958.430 ;
        RECT 3498.200 3958.150 3498.480 3958.430 ;
        RECT 3498.820 3958.150 3499.100 3958.430 ;
        RECT 3499.440 3958.150 3499.720 3958.430 ;
        RECT 3500.060 3958.150 3500.340 3958.430 ;
        RECT 3500.680 3958.150 3500.960 3958.430 ;
        RECT 3496.960 3957.530 3497.240 3957.810 ;
        RECT 3497.580 3957.530 3497.860 3957.810 ;
        RECT 3498.200 3957.530 3498.480 3957.810 ;
        RECT 3498.820 3957.530 3499.100 3957.810 ;
        RECT 3499.440 3957.530 3499.720 3957.810 ;
        RECT 3500.060 3957.530 3500.340 3957.810 ;
        RECT 3500.680 3957.530 3500.960 3957.810 ;
        RECT 3496.960 3956.910 3497.240 3957.190 ;
        RECT 3497.580 3956.910 3497.860 3957.190 ;
        RECT 3498.200 3956.910 3498.480 3957.190 ;
        RECT 3498.820 3956.910 3499.100 3957.190 ;
        RECT 3499.440 3956.910 3499.720 3957.190 ;
        RECT 3500.060 3956.910 3500.340 3957.190 ;
        RECT 3500.680 3956.910 3500.960 3957.190 ;
        RECT 3496.960 3956.290 3497.240 3956.570 ;
        RECT 3497.580 3956.290 3497.860 3956.570 ;
        RECT 3498.200 3956.290 3498.480 3956.570 ;
        RECT 3498.820 3956.290 3499.100 3956.570 ;
        RECT 3499.440 3956.290 3499.720 3956.570 ;
        RECT 3500.060 3956.290 3500.340 3956.570 ;
        RECT 3500.680 3956.290 3500.960 3956.570 ;
        RECT 3496.960 3955.670 3497.240 3955.950 ;
        RECT 3497.580 3955.670 3497.860 3955.950 ;
        RECT 3498.200 3955.670 3498.480 3955.950 ;
        RECT 3498.820 3955.670 3499.100 3955.950 ;
        RECT 3499.440 3955.670 3499.720 3955.950 ;
        RECT 3500.060 3955.670 3500.340 3955.950 ;
        RECT 3500.680 3955.670 3500.960 3955.950 ;
        RECT 3496.960 3955.050 3497.240 3955.330 ;
        RECT 3497.580 3955.050 3497.860 3955.330 ;
        RECT 3498.200 3955.050 3498.480 3955.330 ;
        RECT 3498.820 3955.050 3499.100 3955.330 ;
        RECT 3499.440 3955.050 3499.720 3955.330 ;
        RECT 3500.060 3955.050 3500.340 3955.330 ;
        RECT 3500.680 3955.050 3500.960 3955.330 ;
        RECT 3496.960 3954.430 3497.240 3954.710 ;
        RECT 3497.580 3954.430 3497.860 3954.710 ;
        RECT 3498.200 3954.430 3498.480 3954.710 ;
        RECT 3498.820 3954.430 3499.100 3954.710 ;
        RECT 3499.440 3954.430 3499.720 3954.710 ;
        RECT 3500.060 3954.430 3500.340 3954.710 ;
        RECT 3500.680 3954.430 3500.960 3954.710 ;
        RECT 3539.350 3963.760 3539.630 3964.040 ;
        RECT 3539.350 3963.140 3539.630 3963.420 ;
        RECT 3539.350 3962.520 3539.630 3962.800 ;
        RECT 3539.350 3961.900 3539.630 3962.180 ;
        RECT 3539.350 3961.280 3539.630 3961.560 ;
        RECT 3539.350 3960.660 3539.630 3960.940 ;
        RECT 3539.350 3960.040 3539.630 3960.320 ;
        RECT 3539.350 3959.420 3539.630 3959.700 ;
        RECT 3539.350 3958.800 3539.630 3959.080 ;
        RECT 3539.350 3958.180 3539.630 3958.460 ;
        RECT 3539.350 3957.560 3539.630 3957.840 ;
        RECT 3539.350 3956.940 3539.630 3957.220 ;
        RECT 3539.350 3956.320 3539.630 3956.600 ;
        RECT 3539.350 3955.700 3539.630 3955.980 ;
        RECT 3539.350 3955.080 3539.630 3955.360 ;
        RECT 3539.350 3954.460 3539.630 3954.740 ;
        RECT 3496.960 3950.200 3497.240 3950.480 ;
        RECT 3497.580 3950.200 3497.860 3950.480 ;
        RECT 3498.200 3950.200 3498.480 3950.480 ;
        RECT 3498.820 3950.200 3499.100 3950.480 ;
        RECT 3499.440 3950.200 3499.720 3950.480 ;
        RECT 3500.060 3950.200 3500.340 3950.480 ;
        RECT 3500.680 3950.200 3500.960 3950.480 ;
        RECT 3496.960 3949.580 3497.240 3949.860 ;
        RECT 3497.580 3949.580 3497.860 3949.860 ;
        RECT 3498.200 3949.580 3498.480 3949.860 ;
        RECT 3498.820 3949.580 3499.100 3949.860 ;
        RECT 3499.440 3949.580 3499.720 3949.860 ;
        RECT 3500.060 3949.580 3500.340 3949.860 ;
        RECT 3500.680 3949.580 3500.960 3949.860 ;
        RECT 3496.960 3948.960 3497.240 3949.240 ;
        RECT 3497.580 3948.960 3497.860 3949.240 ;
        RECT 3498.200 3948.960 3498.480 3949.240 ;
        RECT 3498.820 3948.960 3499.100 3949.240 ;
        RECT 3499.440 3948.960 3499.720 3949.240 ;
        RECT 3500.060 3948.960 3500.340 3949.240 ;
        RECT 3500.680 3948.960 3500.960 3949.240 ;
        RECT 3496.960 3948.340 3497.240 3948.620 ;
        RECT 3497.580 3948.340 3497.860 3948.620 ;
        RECT 3498.200 3948.340 3498.480 3948.620 ;
        RECT 3498.820 3948.340 3499.100 3948.620 ;
        RECT 3499.440 3948.340 3499.720 3948.620 ;
        RECT 3500.060 3948.340 3500.340 3948.620 ;
        RECT 3500.680 3948.340 3500.960 3948.620 ;
        RECT 3496.960 3947.720 3497.240 3948.000 ;
        RECT 3497.580 3947.720 3497.860 3948.000 ;
        RECT 3498.200 3947.720 3498.480 3948.000 ;
        RECT 3498.820 3947.720 3499.100 3948.000 ;
        RECT 3499.440 3947.720 3499.720 3948.000 ;
        RECT 3500.060 3947.720 3500.340 3948.000 ;
        RECT 3500.680 3947.720 3500.960 3948.000 ;
        RECT 3496.960 3947.100 3497.240 3947.380 ;
        RECT 3497.580 3947.100 3497.860 3947.380 ;
        RECT 3498.200 3947.100 3498.480 3947.380 ;
        RECT 3498.820 3947.100 3499.100 3947.380 ;
        RECT 3499.440 3947.100 3499.720 3947.380 ;
        RECT 3500.060 3947.100 3500.340 3947.380 ;
        RECT 3500.680 3947.100 3500.960 3947.380 ;
        RECT 3496.960 3946.480 3497.240 3946.760 ;
        RECT 3497.580 3946.480 3497.860 3946.760 ;
        RECT 3498.200 3946.480 3498.480 3946.760 ;
        RECT 3498.820 3946.480 3499.100 3946.760 ;
        RECT 3499.440 3946.480 3499.720 3946.760 ;
        RECT 3500.060 3946.480 3500.340 3946.760 ;
        RECT 3500.680 3946.480 3500.960 3946.760 ;
        RECT 3496.960 3945.860 3497.240 3946.140 ;
        RECT 3497.580 3945.860 3497.860 3946.140 ;
        RECT 3498.200 3945.860 3498.480 3946.140 ;
        RECT 3498.820 3945.860 3499.100 3946.140 ;
        RECT 3499.440 3945.860 3499.720 3946.140 ;
        RECT 3500.060 3945.860 3500.340 3946.140 ;
        RECT 3500.680 3945.860 3500.960 3946.140 ;
        RECT 3496.960 3945.240 3497.240 3945.520 ;
        RECT 3497.580 3945.240 3497.860 3945.520 ;
        RECT 3498.200 3945.240 3498.480 3945.520 ;
        RECT 3498.820 3945.240 3499.100 3945.520 ;
        RECT 3499.440 3945.240 3499.720 3945.520 ;
        RECT 3500.060 3945.240 3500.340 3945.520 ;
        RECT 3500.680 3945.240 3500.960 3945.520 ;
        RECT 3496.960 3944.620 3497.240 3944.900 ;
        RECT 3497.580 3944.620 3497.860 3944.900 ;
        RECT 3498.200 3944.620 3498.480 3944.900 ;
        RECT 3498.820 3944.620 3499.100 3944.900 ;
        RECT 3499.440 3944.620 3499.720 3944.900 ;
        RECT 3500.060 3944.620 3500.340 3944.900 ;
        RECT 3500.680 3944.620 3500.960 3944.900 ;
        RECT 3496.960 3944.000 3497.240 3944.280 ;
        RECT 3497.580 3944.000 3497.860 3944.280 ;
        RECT 3498.200 3944.000 3498.480 3944.280 ;
        RECT 3498.820 3944.000 3499.100 3944.280 ;
        RECT 3499.440 3944.000 3499.720 3944.280 ;
        RECT 3500.060 3944.000 3500.340 3944.280 ;
        RECT 3500.680 3944.000 3500.960 3944.280 ;
        RECT 3496.960 3943.380 3497.240 3943.660 ;
        RECT 3497.580 3943.380 3497.860 3943.660 ;
        RECT 3498.200 3943.380 3498.480 3943.660 ;
        RECT 3498.820 3943.380 3499.100 3943.660 ;
        RECT 3499.440 3943.380 3499.720 3943.660 ;
        RECT 3500.060 3943.380 3500.340 3943.660 ;
        RECT 3500.680 3943.380 3500.960 3943.660 ;
        RECT 3496.960 3942.760 3497.240 3943.040 ;
        RECT 3497.580 3942.760 3497.860 3943.040 ;
        RECT 3498.200 3942.760 3498.480 3943.040 ;
        RECT 3498.820 3942.760 3499.100 3943.040 ;
        RECT 3499.440 3942.760 3499.720 3943.040 ;
        RECT 3500.060 3942.760 3500.340 3943.040 ;
        RECT 3500.680 3942.760 3500.960 3943.040 ;
        RECT 3496.960 3942.140 3497.240 3942.420 ;
        RECT 3497.580 3942.140 3497.860 3942.420 ;
        RECT 3498.200 3942.140 3498.480 3942.420 ;
        RECT 3498.820 3942.140 3499.100 3942.420 ;
        RECT 3499.440 3942.140 3499.720 3942.420 ;
        RECT 3500.060 3942.140 3500.340 3942.420 ;
        RECT 3500.680 3942.140 3500.960 3942.420 ;
        RECT 3496.960 3941.520 3497.240 3941.800 ;
        RECT 3497.580 3941.520 3497.860 3941.800 ;
        RECT 3498.200 3941.520 3498.480 3941.800 ;
        RECT 3498.820 3941.520 3499.100 3941.800 ;
        RECT 3499.440 3941.520 3499.720 3941.800 ;
        RECT 3500.060 3941.520 3500.340 3941.800 ;
        RECT 3500.680 3941.520 3500.960 3941.800 ;
        RECT 3496.960 3940.900 3497.240 3941.180 ;
        RECT 3497.580 3940.900 3497.860 3941.180 ;
        RECT 3498.200 3940.900 3498.480 3941.180 ;
        RECT 3498.820 3940.900 3499.100 3941.180 ;
        RECT 3499.440 3940.900 3499.720 3941.180 ;
        RECT 3500.060 3940.900 3500.340 3941.180 ;
        RECT 3500.680 3940.900 3500.960 3941.180 ;
        RECT 3539.350 3950.230 3539.630 3950.510 ;
        RECT 3539.350 3949.610 3539.630 3949.890 ;
        RECT 3539.350 3948.990 3539.630 3949.270 ;
        RECT 3539.350 3948.370 3539.630 3948.650 ;
        RECT 3539.350 3947.750 3539.630 3948.030 ;
        RECT 3539.350 3947.130 3539.630 3947.410 ;
        RECT 3539.350 3946.510 3539.630 3946.790 ;
        RECT 3539.350 3945.890 3539.630 3946.170 ;
        RECT 3539.350 3945.270 3539.630 3945.550 ;
        RECT 3539.350 3944.650 3539.630 3944.930 ;
        RECT 3539.350 3944.030 3539.630 3944.310 ;
        RECT 3539.350 3943.410 3539.630 3943.690 ;
        RECT 3539.350 3942.790 3539.630 3943.070 ;
        RECT 3539.350 3942.170 3539.630 3942.450 ;
        RECT 3539.350 3941.550 3539.630 3941.830 ;
        RECT 3539.350 3940.930 3539.630 3941.210 ;
        RECT 3496.960 3938.350 3497.240 3938.630 ;
        RECT 3497.580 3938.350 3497.860 3938.630 ;
        RECT 3498.200 3938.350 3498.480 3938.630 ;
        RECT 3498.820 3938.350 3499.100 3938.630 ;
        RECT 3499.440 3938.350 3499.720 3938.630 ;
        RECT 3500.060 3938.350 3500.340 3938.630 ;
        RECT 3500.680 3938.350 3500.960 3938.630 ;
        RECT 3496.960 3937.730 3497.240 3938.010 ;
        RECT 3497.580 3937.730 3497.860 3938.010 ;
        RECT 3498.200 3937.730 3498.480 3938.010 ;
        RECT 3498.820 3937.730 3499.100 3938.010 ;
        RECT 3499.440 3937.730 3499.720 3938.010 ;
        RECT 3500.060 3937.730 3500.340 3938.010 ;
        RECT 3500.680 3937.730 3500.960 3938.010 ;
        RECT 3496.960 3937.110 3497.240 3937.390 ;
        RECT 3497.580 3937.110 3497.860 3937.390 ;
        RECT 3498.200 3937.110 3498.480 3937.390 ;
        RECT 3498.820 3937.110 3499.100 3937.390 ;
        RECT 3499.440 3937.110 3499.720 3937.390 ;
        RECT 3500.060 3937.110 3500.340 3937.390 ;
        RECT 3500.680 3937.110 3500.960 3937.390 ;
        RECT 3496.960 3936.490 3497.240 3936.770 ;
        RECT 3497.580 3936.490 3497.860 3936.770 ;
        RECT 3498.200 3936.490 3498.480 3936.770 ;
        RECT 3498.820 3936.490 3499.100 3936.770 ;
        RECT 3499.440 3936.490 3499.720 3936.770 ;
        RECT 3500.060 3936.490 3500.340 3936.770 ;
        RECT 3500.680 3936.490 3500.960 3936.770 ;
        RECT 3496.960 3935.870 3497.240 3936.150 ;
        RECT 3497.580 3935.870 3497.860 3936.150 ;
        RECT 3498.200 3935.870 3498.480 3936.150 ;
        RECT 3498.820 3935.870 3499.100 3936.150 ;
        RECT 3499.440 3935.870 3499.720 3936.150 ;
        RECT 3500.060 3935.870 3500.340 3936.150 ;
        RECT 3500.680 3935.870 3500.960 3936.150 ;
        RECT 3496.960 3935.250 3497.240 3935.530 ;
        RECT 3497.580 3935.250 3497.860 3935.530 ;
        RECT 3498.200 3935.250 3498.480 3935.530 ;
        RECT 3498.820 3935.250 3499.100 3935.530 ;
        RECT 3499.440 3935.250 3499.720 3935.530 ;
        RECT 3500.060 3935.250 3500.340 3935.530 ;
        RECT 3500.680 3935.250 3500.960 3935.530 ;
        RECT 3496.960 3934.630 3497.240 3934.910 ;
        RECT 3497.580 3934.630 3497.860 3934.910 ;
        RECT 3498.200 3934.630 3498.480 3934.910 ;
        RECT 3498.820 3934.630 3499.100 3934.910 ;
        RECT 3499.440 3934.630 3499.720 3934.910 ;
        RECT 3500.060 3934.630 3500.340 3934.910 ;
        RECT 3500.680 3934.630 3500.960 3934.910 ;
        RECT 3496.960 3934.010 3497.240 3934.290 ;
        RECT 3497.580 3934.010 3497.860 3934.290 ;
        RECT 3498.200 3934.010 3498.480 3934.290 ;
        RECT 3498.820 3934.010 3499.100 3934.290 ;
        RECT 3499.440 3934.010 3499.720 3934.290 ;
        RECT 3500.060 3934.010 3500.340 3934.290 ;
        RECT 3500.680 3934.010 3500.960 3934.290 ;
        RECT 3496.960 3933.390 3497.240 3933.670 ;
        RECT 3497.580 3933.390 3497.860 3933.670 ;
        RECT 3498.200 3933.390 3498.480 3933.670 ;
        RECT 3498.820 3933.390 3499.100 3933.670 ;
        RECT 3499.440 3933.390 3499.720 3933.670 ;
        RECT 3500.060 3933.390 3500.340 3933.670 ;
        RECT 3500.680 3933.390 3500.960 3933.670 ;
        RECT 3496.960 3932.770 3497.240 3933.050 ;
        RECT 3497.580 3932.770 3497.860 3933.050 ;
        RECT 3498.200 3932.770 3498.480 3933.050 ;
        RECT 3498.820 3932.770 3499.100 3933.050 ;
        RECT 3499.440 3932.770 3499.720 3933.050 ;
        RECT 3500.060 3932.770 3500.340 3933.050 ;
        RECT 3500.680 3932.770 3500.960 3933.050 ;
        RECT 3496.960 3932.150 3497.240 3932.430 ;
        RECT 3497.580 3932.150 3497.860 3932.430 ;
        RECT 3498.200 3932.150 3498.480 3932.430 ;
        RECT 3498.820 3932.150 3499.100 3932.430 ;
        RECT 3499.440 3932.150 3499.720 3932.430 ;
        RECT 3500.060 3932.150 3500.340 3932.430 ;
        RECT 3500.680 3932.150 3500.960 3932.430 ;
        RECT 3496.960 3931.530 3497.240 3931.810 ;
        RECT 3497.580 3931.530 3497.860 3931.810 ;
        RECT 3498.200 3931.530 3498.480 3931.810 ;
        RECT 3498.820 3931.530 3499.100 3931.810 ;
        RECT 3499.440 3931.530 3499.720 3931.810 ;
        RECT 3500.060 3931.530 3500.340 3931.810 ;
        RECT 3500.680 3931.530 3500.960 3931.810 ;
        RECT 3496.960 3930.910 3497.240 3931.190 ;
        RECT 3497.580 3930.910 3497.860 3931.190 ;
        RECT 3498.200 3930.910 3498.480 3931.190 ;
        RECT 3498.820 3930.910 3499.100 3931.190 ;
        RECT 3499.440 3930.910 3499.720 3931.190 ;
        RECT 3500.060 3930.910 3500.340 3931.190 ;
        RECT 3500.680 3930.910 3500.960 3931.190 ;
        RECT 3496.960 3930.290 3497.240 3930.570 ;
        RECT 3497.580 3930.290 3497.860 3930.570 ;
        RECT 3498.200 3930.290 3498.480 3930.570 ;
        RECT 3498.820 3930.290 3499.100 3930.570 ;
        RECT 3499.440 3930.290 3499.720 3930.570 ;
        RECT 3500.060 3930.290 3500.340 3930.570 ;
        RECT 3500.680 3930.290 3500.960 3930.570 ;
        RECT 3496.960 3929.670 3497.240 3929.950 ;
        RECT 3497.580 3929.670 3497.860 3929.950 ;
        RECT 3498.200 3929.670 3498.480 3929.950 ;
        RECT 3498.820 3929.670 3499.100 3929.950 ;
        RECT 3499.440 3929.670 3499.720 3929.950 ;
        RECT 3500.060 3929.670 3500.340 3929.950 ;
        RECT 3500.680 3929.670 3500.960 3929.950 ;
        RECT 3496.960 3929.050 3497.240 3929.330 ;
        RECT 3497.580 3929.050 3497.860 3929.330 ;
        RECT 3498.200 3929.050 3498.480 3929.330 ;
        RECT 3498.820 3929.050 3499.100 3929.330 ;
        RECT 3499.440 3929.050 3499.720 3929.330 ;
        RECT 3500.060 3929.050 3500.340 3929.330 ;
        RECT 3500.680 3929.050 3500.960 3929.330 ;
        RECT 3539.350 3938.380 3539.630 3938.660 ;
        RECT 3539.350 3937.760 3539.630 3938.040 ;
        RECT 3539.350 3937.140 3539.630 3937.420 ;
        RECT 3539.350 3936.520 3539.630 3936.800 ;
        RECT 3539.350 3935.900 3539.630 3936.180 ;
        RECT 3539.350 3935.280 3539.630 3935.560 ;
        RECT 3539.350 3934.660 3539.630 3934.940 ;
        RECT 3539.350 3934.040 3539.630 3934.320 ;
        RECT 3539.350 3933.420 3539.630 3933.700 ;
        RECT 3539.350 3932.800 3539.630 3933.080 ;
        RECT 3539.350 3932.180 3539.630 3932.460 ;
        RECT 3539.350 3931.560 3539.630 3931.840 ;
        RECT 3539.350 3930.940 3539.630 3931.220 ;
        RECT 3539.350 3930.320 3539.630 3930.600 ;
        RECT 3539.350 3929.700 3539.630 3929.980 ;
        RECT 3539.350 3929.080 3539.630 3929.360 ;
        RECT 3496.960 3925.330 3497.240 3925.610 ;
        RECT 3497.580 3925.330 3497.860 3925.610 ;
        RECT 3498.200 3925.330 3498.480 3925.610 ;
        RECT 3498.820 3925.330 3499.100 3925.610 ;
        RECT 3499.440 3925.330 3499.720 3925.610 ;
        RECT 3500.060 3925.330 3500.340 3925.610 ;
        RECT 3500.680 3925.330 3500.960 3925.610 ;
        RECT 3496.960 3924.710 3497.240 3924.990 ;
        RECT 3497.580 3924.710 3497.860 3924.990 ;
        RECT 3498.200 3924.710 3498.480 3924.990 ;
        RECT 3498.820 3924.710 3499.100 3924.990 ;
        RECT 3499.440 3924.710 3499.720 3924.990 ;
        RECT 3500.060 3924.710 3500.340 3924.990 ;
        RECT 3500.680 3924.710 3500.960 3924.990 ;
        RECT 3496.960 3924.090 3497.240 3924.370 ;
        RECT 3497.580 3924.090 3497.860 3924.370 ;
        RECT 3498.200 3924.090 3498.480 3924.370 ;
        RECT 3498.820 3924.090 3499.100 3924.370 ;
        RECT 3499.440 3924.090 3499.720 3924.370 ;
        RECT 3500.060 3924.090 3500.340 3924.370 ;
        RECT 3500.680 3924.090 3500.960 3924.370 ;
        RECT 3496.960 3923.470 3497.240 3923.750 ;
        RECT 3497.580 3923.470 3497.860 3923.750 ;
        RECT 3498.200 3923.470 3498.480 3923.750 ;
        RECT 3498.820 3923.470 3499.100 3923.750 ;
        RECT 3499.440 3923.470 3499.720 3923.750 ;
        RECT 3500.060 3923.470 3500.340 3923.750 ;
        RECT 3500.680 3923.470 3500.960 3923.750 ;
        RECT 3496.960 3922.850 3497.240 3923.130 ;
        RECT 3497.580 3922.850 3497.860 3923.130 ;
        RECT 3498.200 3922.850 3498.480 3923.130 ;
        RECT 3498.820 3922.850 3499.100 3923.130 ;
        RECT 3499.440 3922.850 3499.720 3923.130 ;
        RECT 3500.060 3922.850 3500.340 3923.130 ;
        RECT 3500.680 3922.850 3500.960 3923.130 ;
        RECT 3496.960 3922.230 3497.240 3922.510 ;
        RECT 3497.580 3922.230 3497.860 3922.510 ;
        RECT 3498.200 3922.230 3498.480 3922.510 ;
        RECT 3498.820 3922.230 3499.100 3922.510 ;
        RECT 3499.440 3922.230 3499.720 3922.510 ;
        RECT 3500.060 3922.230 3500.340 3922.510 ;
        RECT 3500.680 3922.230 3500.960 3922.510 ;
        RECT 3496.960 3921.610 3497.240 3921.890 ;
        RECT 3497.580 3921.610 3497.860 3921.890 ;
        RECT 3498.200 3921.610 3498.480 3921.890 ;
        RECT 3498.820 3921.610 3499.100 3921.890 ;
        RECT 3499.440 3921.610 3499.720 3921.890 ;
        RECT 3500.060 3921.610 3500.340 3921.890 ;
        RECT 3500.680 3921.610 3500.960 3921.890 ;
        RECT 3496.960 3920.990 3497.240 3921.270 ;
        RECT 3497.580 3920.990 3497.860 3921.270 ;
        RECT 3498.200 3920.990 3498.480 3921.270 ;
        RECT 3498.820 3920.990 3499.100 3921.270 ;
        RECT 3499.440 3920.990 3499.720 3921.270 ;
        RECT 3500.060 3920.990 3500.340 3921.270 ;
        RECT 3500.680 3920.990 3500.960 3921.270 ;
        RECT 3496.960 3920.370 3497.240 3920.650 ;
        RECT 3497.580 3920.370 3497.860 3920.650 ;
        RECT 3498.200 3920.370 3498.480 3920.650 ;
        RECT 3498.820 3920.370 3499.100 3920.650 ;
        RECT 3499.440 3920.370 3499.720 3920.650 ;
        RECT 3500.060 3920.370 3500.340 3920.650 ;
        RECT 3500.680 3920.370 3500.960 3920.650 ;
        RECT 3496.960 3919.750 3497.240 3920.030 ;
        RECT 3497.580 3919.750 3497.860 3920.030 ;
        RECT 3498.200 3919.750 3498.480 3920.030 ;
        RECT 3498.820 3919.750 3499.100 3920.030 ;
        RECT 3499.440 3919.750 3499.720 3920.030 ;
        RECT 3500.060 3919.750 3500.340 3920.030 ;
        RECT 3500.680 3919.750 3500.960 3920.030 ;
        RECT 3496.960 3919.130 3497.240 3919.410 ;
        RECT 3497.580 3919.130 3497.860 3919.410 ;
        RECT 3498.200 3919.130 3498.480 3919.410 ;
        RECT 3498.820 3919.130 3499.100 3919.410 ;
        RECT 3499.440 3919.130 3499.720 3919.410 ;
        RECT 3500.060 3919.130 3500.340 3919.410 ;
        RECT 3500.680 3919.130 3500.960 3919.410 ;
        RECT 3496.960 3918.510 3497.240 3918.790 ;
        RECT 3497.580 3918.510 3497.860 3918.790 ;
        RECT 3498.200 3918.510 3498.480 3918.790 ;
        RECT 3498.820 3918.510 3499.100 3918.790 ;
        RECT 3499.440 3918.510 3499.720 3918.790 ;
        RECT 3500.060 3918.510 3500.340 3918.790 ;
        RECT 3500.680 3918.510 3500.960 3918.790 ;
        RECT 3496.960 3917.890 3497.240 3918.170 ;
        RECT 3497.580 3917.890 3497.860 3918.170 ;
        RECT 3498.200 3917.890 3498.480 3918.170 ;
        RECT 3498.820 3917.890 3499.100 3918.170 ;
        RECT 3499.440 3917.890 3499.720 3918.170 ;
        RECT 3500.060 3917.890 3500.340 3918.170 ;
        RECT 3500.680 3917.890 3500.960 3918.170 ;
        RECT 3496.960 3917.270 3497.240 3917.550 ;
        RECT 3497.580 3917.270 3497.860 3917.550 ;
        RECT 3498.200 3917.270 3498.480 3917.550 ;
        RECT 3498.820 3917.270 3499.100 3917.550 ;
        RECT 3499.440 3917.270 3499.720 3917.550 ;
        RECT 3500.060 3917.270 3500.340 3917.550 ;
        RECT 3500.680 3917.270 3500.960 3917.550 ;
        RECT 3496.960 3916.650 3497.240 3916.930 ;
        RECT 3497.580 3916.650 3497.860 3916.930 ;
        RECT 3498.200 3916.650 3498.480 3916.930 ;
        RECT 3498.820 3916.650 3499.100 3916.930 ;
        RECT 3499.440 3916.650 3499.720 3916.930 ;
        RECT 3500.060 3916.650 3500.340 3916.930 ;
        RECT 3500.680 3916.650 3500.960 3916.930 ;
        RECT 3539.350 3925.390 3539.630 3925.670 ;
        RECT 3539.350 3924.770 3539.630 3925.050 ;
        RECT 3539.350 3924.150 3539.630 3924.430 ;
        RECT 3539.350 3923.530 3539.630 3923.810 ;
        RECT 3539.350 3922.910 3539.630 3923.190 ;
        RECT 3539.350 3922.290 3539.630 3922.570 ;
        RECT 3539.350 3921.670 3539.630 3921.950 ;
        RECT 3539.350 3921.050 3539.630 3921.330 ;
        RECT 3539.350 3920.430 3539.630 3920.710 ;
        RECT 3539.350 3919.810 3539.630 3920.090 ;
        RECT 3539.350 3919.190 3539.630 3919.470 ;
        RECT 3539.350 3918.570 3539.630 3918.850 ;
        RECT 3539.350 3917.950 3539.630 3918.230 ;
        RECT 3539.350 3917.330 3539.630 3917.610 ;
        RECT 3539.350 3916.710 3539.630 3916.990 ;
        RECT 3497.720 3851.865 3498.000 3852.145 ;
        RECT 3499.220 3851.865 3499.500 3852.145 ;
        RECT 3500.720 3851.865 3501.000 3852.145 ;
        RECT 3497.720 3850.865 3498.000 3851.145 ;
        RECT 3499.220 3850.865 3499.500 3851.145 ;
        RECT 3500.720 3850.865 3501.000 3851.145 ;
        RECT 3497.220 3769.490 3497.500 3769.770 ;
        RECT 3498.720 3769.490 3499.000 3769.770 ;
        RECT 3500.220 3769.490 3500.500 3769.770 ;
        RECT 3497.220 3734.490 3497.500 3734.770 ;
        RECT 3498.720 3734.490 3499.000 3734.770 ;
        RECT 3500.220 3734.490 3500.500 3734.770 ;
        RECT 3497.220 3699.490 3497.500 3699.770 ;
        RECT 3498.720 3699.490 3499.000 3699.770 ;
        RECT 3500.220 3699.490 3500.500 3699.770 ;
        RECT 3497.720 3671.865 3498.000 3672.145 ;
        RECT 3499.220 3671.865 3499.500 3672.145 ;
        RECT 3500.720 3671.865 3501.000 3672.145 ;
        RECT 3497.720 3670.865 3498.000 3671.145 ;
        RECT 3499.220 3670.865 3499.500 3671.145 ;
        RECT 3500.720 3670.865 3501.000 3671.145 ;
        RECT 3497.485 3601.835 3497.765 3602.115 ;
        RECT 3498.985 3601.835 3499.265 3602.115 ;
        RECT 3500.485 3601.835 3500.765 3602.115 ;
        RECT 3497.220 3554.490 3497.500 3554.770 ;
        RECT 3498.720 3554.490 3499.000 3554.770 ;
        RECT 3500.220 3554.490 3500.500 3554.770 ;
        RECT 3497.220 3519.490 3497.500 3519.770 ;
        RECT 3498.720 3519.490 3499.000 3519.770 ;
        RECT 3500.220 3519.490 3500.500 3519.770 ;
        RECT 3497.720 3491.865 3498.000 3492.145 ;
        RECT 3499.220 3491.865 3499.500 3492.145 ;
        RECT 3500.720 3491.865 3501.000 3492.145 ;
        RECT 3497.720 3490.865 3498.000 3491.145 ;
        RECT 3499.220 3490.865 3499.500 3491.145 ;
        RECT 3500.720 3490.865 3501.000 3491.145 ;
        RECT 3497.220 3484.490 3497.500 3484.770 ;
        RECT 3498.720 3484.490 3499.000 3484.770 ;
        RECT 3500.220 3484.490 3500.500 3484.770 ;
        RECT 3497.485 3386.835 3497.765 3387.115 ;
        RECT 3498.985 3386.835 3499.265 3387.115 ;
        RECT 3500.485 3386.835 3500.765 3387.115 ;
        RECT 3497.220 3339.490 3497.500 3339.770 ;
        RECT 3498.720 3339.490 3499.000 3339.770 ;
        RECT 3500.220 3339.490 3500.500 3339.770 ;
        RECT 3497.720 3311.865 3498.000 3312.145 ;
        RECT 3499.220 3311.865 3499.500 3312.145 ;
        RECT 3500.720 3311.865 3501.000 3312.145 ;
        RECT 3497.720 3310.865 3498.000 3311.145 ;
        RECT 3499.220 3310.865 3499.500 3311.145 ;
        RECT 3500.720 3310.865 3501.000 3311.145 ;
        RECT 3497.220 3304.490 3497.500 3304.770 ;
        RECT 3498.720 3304.490 3499.000 3304.770 ;
        RECT 3500.220 3304.490 3500.500 3304.770 ;
        RECT 3497.220 3269.490 3497.500 3269.770 ;
        RECT 3498.720 3269.490 3499.000 3269.770 ;
        RECT 3500.220 3269.490 3500.500 3269.770 ;
        RECT 3497.485 3171.835 3497.765 3172.115 ;
        RECT 3498.985 3171.835 3499.265 3172.115 ;
        RECT 3500.485 3171.835 3500.765 3172.115 ;
        RECT 3497.720 3131.865 3498.000 3132.145 ;
        RECT 3499.220 3131.865 3499.500 3132.145 ;
        RECT 3500.720 3131.865 3501.000 3132.145 ;
        RECT 3497.720 3130.865 3498.000 3131.145 ;
        RECT 3499.220 3130.865 3499.500 3131.145 ;
        RECT 3500.720 3130.865 3501.000 3131.145 ;
        RECT 3497.220 3124.490 3497.500 3124.770 ;
        RECT 3498.720 3124.490 3499.000 3124.770 ;
        RECT 3500.220 3124.490 3500.500 3124.770 ;
        RECT 3497.220 3089.490 3497.500 3089.770 ;
        RECT 3498.720 3089.490 3499.000 3089.770 ;
        RECT 3500.220 3089.490 3500.500 3089.770 ;
        RECT 3497.220 3054.490 3497.500 3054.770 ;
        RECT 3498.720 3054.490 3499.000 3054.770 ;
        RECT 3500.220 3054.490 3500.500 3054.770 ;
        RECT 3497.485 2956.835 3497.765 2957.115 ;
        RECT 3498.985 2956.835 3499.265 2957.115 ;
        RECT 3500.485 2956.835 3500.765 2957.115 ;
        RECT 3497.720 2951.865 3498.000 2952.145 ;
        RECT 3499.220 2951.865 3499.500 2952.145 ;
        RECT 3500.720 2951.865 3501.000 2952.145 ;
        RECT 3497.720 2950.865 3498.000 2951.145 ;
        RECT 3499.220 2950.865 3499.500 2951.145 ;
        RECT 3500.720 2950.865 3501.000 2951.145 ;
        RECT 3497.220 2909.490 3497.500 2909.770 ;
        RECT 3498.720 2909.490 3499.000 2909.770 ;
        RECT 3500.220 2909.490 3500.500 2909.770 ;
        RECT 3497.220 2874.490 3497.500 2874.770 ;
        RECT 3498.720 2874.490 3499.000 2874.770 ;
        RECT 3500.220 2874.490 3500.500 2874.770 ;
        RECT 3497.220 2839.490 3497.500 2839.770 ;
        RECT 3498.720 2839.490 3499.000 2839.770 ;
        RECT 3500.220 2839.490 3500.500 2839.770 ;
        RECT 3497.720 2771.865 3498.000 2772.145 ;
        RECT 3499.220 2771.865 3499.500 2772.145 ;
        RECT 3500.720 2771.865 3501.000 2772.145 ;
        RECT 3497.720 2770.865 3498.000 2771.145 ;
        RECT 3499.220 2770.865 3499.500 2771.145 ;
        RECT 3500.720 2770.865 3501.000 2771.145 ;
        RECT 3497.485 2741.835 3497.765 2742.115 ;
        RECT 3498.985 2741.835 3499.265 2742.115 ;
        RECT 3500.485 2741.835 3500.765 2742.115 ;
        RECT 3497.220 2694.490 3497.500 2694.770 ;
        RECT 3498.720 2694.490 3499.000 2694.770 ;
        RECT 3500.220 2694.490 3500.500 2694.770 ;
        RECT 3497.220 2659.490 3497.500 2659.770 ;
        RECT 3498.720 2659.490 3499.000 2659.770 ;
        RECT 3500.220 2659.490 3500.500 2659.770 ;
        RECT 3497.220 2624.490 3497.500 2624.770 ;
        RECT 3498.720 2624.490 3499.000 2624.770 ;
        RECT 3500.220 2624.490 3500.500 2624.770 ;
        RECT 3497.720 2591.865 3498.000 2592.145 ;
        RECT 3499.220 2591.865 3499.500 2592.145 ;
        RECT 3500.720 2591.865 3501.000 2592.145 ;
        RECT 3497.720 2590.865 3498.000 2591.145 ;
        RECT 3499.220 2590.865 3499.500 2591.145 ;
        RECT 3500.720 2590.865 3501.000 2591.145 ;
        RECT 3497.485 2526.835 3497.765 2527.115 ;
        RECT 3498.985 2526.835 3499.265 2527.115 ;
        RECT 3500.485 2526.835 3500.765 2527.115 ;
        RECT 3496.960 2482.980 3497.240 2483.260 ;
        RECT 3497.580 2482.980 3497.860 2483.260 ;
        RECT 3498.200 2482.980 3498.480 2483.260 ;
        RECT 3498.820 2482.980 3499.100 2483.260 ;
        RECT 3499.440 2482.980 3499.720 2483.260 ;
        RECT 3500.060 2482.980 3500.340 2483.260 ;
        RECT 3500.680 2482.980 3500.960 2483.260 ;
        RECT 3496.960 2482.360 3497.240 2482.640 ;
        RECT 3497.580 2482.360 3497.860 2482.640 ;
        RECT 3498.200 2482.360 3498.480 2482.640 ;
        RECT 3498.820 2482.360 3499.100 2482.640 ;
        RECT 3499.440 2482.360 3499.720 2482.640 ;
        RECT 3500.060 2482.360 3500.340 2482.640 ;
        RECT 3500.680 2482.360 3500.960 2482.640 ;
        RECT 3496.960 2481.740 3497.240 2482.020 ;
        RECT 3497.580 2481.740 3497.860 2482.020 ;
        RECT 3498.200 2481.740 3498.480 2482.020 ;
        RECT 3498.820 2481.740 3499.100 2482.020 ;
        RECT 3499.440 2481.740 3499.720 2482.020 ;
        RECT 3500.060 2481.740 3500.340 2482.020 ;
        RECT 3500.680 2481.740 3500.960 2482.020 ;
        RECT 3496.960 2481.120 3497.240 2481.400 ;
        RECT 3497.580 2481.120 3497.860 2481.400 ;
        RECT 3498.200 2481.120 3498.480 2481.400 ;
        RECT 3498.820 2481.120 3499.100 2481.400 ;
        RECT 3499.440 2481.120 3499.720 2481.400 ;
        RECT 3500.060 2481.120 3500.340 2481.400 ;
        RECT 3500.680 2481.120 3500.960 2481.400 ;
        RECT 3496.960 2480.500 3497.240 2480.780 ;
        RECT 3497.580 2480.500 3497.860 2480.780 ;
        RECT 3498.200 2480.500 3498.480 2480.780 ;
        RECT 3498.820 2480.500 3499.100 2480.780 ;
        RECT 3499.440 2480.500 3499.720 2480.780 ;
        RECT 3500.060 2480.500 3500.340 2480.780 ;
        RECT 3500.680 2480.500 3500.960 2480.780 ;
        RECT 3496.960 2479.880 3497.240 2480.160 ;
        RECT 3497.580 2479.880 3497.860 2480.160 ;
        RECT 3498.200 2479.880 3498.480 2480.160 ;
        RECT 3498.820 2479.880 3499.100 2480.160 ;
        RECT 3499.440 2479.880 3499.720 2480.160 ;
        RECT 3500.060 2479.880 3500.340 2480.160 ;
        RECT 3500.680 2479.880 3500.960 2480.160 ;
        RECT 3496.960 2479.260 3497.240 2479.540 ;
        RECT 3497.580 2479.260 3497.860 2479.540 ;
        RECT 3498.200 2479.260 3498.480 2479.540 ;
        RECT 3498.820 2479.260 3499.100 2479.540 ;
        RECT 3499.440 2479.260 3499.720 2479.540 ;
        RECT 3500.060 2479.260 3500.340 2479.540 ;
        RECT 3500.680 2479.260 3500.960 2479.540 ;
        RECT 3496.960 2478.640 3497.240 2478.920 ;
        RECT 3497.580 2478.640 3497.860 2478.920 ;
        RECT 3498.200 2478.640 3498.480 2478.920 ;
        RECT 3498.820 2478.640 3499.100 2478.920 ;
        RECT 3499.440 2478.640 3499.720 2478.920 ;
        RECT 3500.060 2478.640 3500.340 2478.920 ;
        RECT 3500.680 2478.640 3500.960 2478.920 ;
        RECT 3496.960 2478.020 3497.240 2478.300 ;
        RECT 3497.580 2478.020 3497.860 2478.300 ;
        RECT 3498.200 2478.020 3498.480 2478.300 ;
        RECT 3498.820 2478.020 3499.100 2478.300 ;
        RECT 3499.440 2478.020 3499.720 2478.300 ;
        RECT 3500.060 2478.020 3500.340 2478.300 ;
        RECT 3500.680 2478.020 3500.960 2478.300 ;
        RECT 3496.960 2477.400 3497.240 2477.680 ;
        RECT 3497.580 2477.400 3497.860 2477.680 ;
        RECT 3498.200 2477.400 3498.480 2477.680 ;
        RECT 3498.820 2477.400 3499.100 2477.680 ;
        RECT 3499.440 2477.400 3499.720 2477.680 ;
        RECT 3500.060 2477.400 3500.340 2477.680 ;
        RECT 3500.680 2477.400 3500.960 2477.680 ;
        RECT 3496.960 2476.780 3497.240 2477.060 ;
        RECT 3497.580 2476.780 3497.860 2477.060 ;
        RECT 3498.200 2476.780 3498.480 2477.060 ;
        RECT 3498.820 2476.780 3499.100 2477.060 ;
        RECT 3499.440 2476.780 3499.720 2477.060 ;
        RECT 3500.060 2476.780 3500.340 2477.060 ;
        RECT 3500.680 2476.780 3500.960 2477.060 ;
        RECT 3496.960 2476.160 3497.240 2476.440 ;
        RECT 3497.580 2476.160 3497.860 2476.440 ;
        RECT 3498.200 2476.160 3498.480 2476.440 ;
        RECT 3498.820 2476.160 3499.100 2476.440 ;
        RECT 3499.440 2476.160 3499.720 2476.440 ;
        RECT 3500.060 2476.160 3500.340 2476.440 ;
        RECT 3500.680 2476.160 3500.960 2476.440 ;
        RECT 3496.960 2475.540 3497.240 2475.820 ;
        RECT 3497.580 2475.540 3497.860 2475.820 ;
        RECT 3498.200 2475.540 3498.480 2475.820 ;
        RECT 3498.820 2475.540 3499.100 2475.820 ;
        RECT 3499.440 2475.540 3499.720 2475.820 ;
        RECT 3500.060 2475.540 3500.340 2475.820 ;
        RECT 3500.680 2475.540 3500.960 2475.820 ;
        RECT 3496.960 2474.920 3497.240 2475.200 ;
        RECT 3497.580 2474.920 3497.860 2475.200 ;
        RECT 3498.200 2474.920 3498.480 2475.200 ;
        RECT 3498.820 2474.920 3499.100 2475.200 ;
        RECT 3499.440 2474.920 3499.720 2475.200 ;
        RECT 3500.060 2474.920 3500.340 2475.200 ;
        RECT 3500.680 2474.920 3500.960 2475.200 ;
        RECT 3496.960 2474.300 3497.240 2474.580 ;
        RECT 3497.580 2474.300 3497.860 2474.580 ;
        RECT 3498.200 2474.300 3498.480 2474.580 ;
        RECT 3498.820 2474.300 3499.100 2474.580 ;
        RECT 3499.440 2474.300 3499.720 2474.580 ;
        RECT 3500.060 2474.300 3500.340 2474.580 ;
        RECT 3500.680 2474.300 3500.960 2474.580 ;
        RECT 3539.350 2483.010 3539.630 2483.290 ;
        RECT 3539.350 2482.390 3539.630 2482.670 ;
        RECT 3539.350 2481.770 3539.630 2482.050 ;
        RECT 3539.350 2481.150 3539.630 2481.430 ;
        RECT 3539.350 2480.530 3539.630 2480.810 ;
        RECT 3539.350 2479.910 3539.630 2480.190 ;
        RECT 3539.350 2479.290 3539.630 2479.570 ;
        RECT 3539.350 2478.670 3539.630 2478.950 ;
        RECT 3539.350 2478.050 3539.630 2478.330 ;
        RECT 3539.350 2477.430 3539.630 2477.710 ;
        RECT 3539.350 2476.810 3539.630 2477.090 ;
        RECT 3539.350 2476.190 3539.630 2476.470 ;
        RECT 3539.350 2475.570 3539.630 2475.850 ;
        RECT 3539.350 2474.950 3539.630 2475.230 ;
        RECT 3539.350 2474.330 3539.630 2474.610 ;
        RECT 3496.960 2470.580 3497.240 2470.860 ;
        RECT 3497.580 2470.580 3497.860 2470.860 ;
        RECT 3498.200 2470.580 3498.480 2470.860 ;
        RECT 3498.820 2470.580 3499.100 2470.860 ;
        RECT 3499.440 2470.580 3499.720 2470.860 ;
        RECT 3500.060 2470.580 3500.340 2470.860 ;
        RECT 3500.680 2470.580 3500.960 2470.860 ;
        RECT 3496.960 2469.960 3497.240 2470.240 ;
        RECT 3497.580 2469.960 3497.860 2470.240 ;
        RECT 3498.200 2469.960 3498.480 2470.240 ;
        RECT 3498.820 2469.960 3499.100 2470.240 ;
        RECT 3499.440 2469.960 3499.720 2470.240 ;
        RECT 3500.060 2469.960 3500.340 2470.240 ;
        RECT 3500.680 2469.960 3500.960 2470.240 ;
        RECT 3496.960 2469.340 3497.240 2469.620 ;
        RECT 3497.580 2469.340 3497.860 2469.620 ;
        RECT 3498.200 2469.340 3498.480 2469.620 ;
        RECT 3498.820 2469.340 3499.100 2469.620 ;
        RECT 3499.440 2469.340 3499.720 2469.620 ;
        RECT 3500.060 2469.340 3500.340 2469.620 ;
        RECT 3500.680 2469.340 3500.960 2469.620 ;
        RECT 3496.960 2468.720 3497.240 2469.000 ;
        RECT 3497.580 2468.720 3497.860 2469.000 ;
        RECT 3498.200 2468.720 3498.480 2469.000 ;
        RECT 3498.820 2468.720 3499.100 2469.000 ;
        RECT 3499.440 2468.720 3499.720 2469.000 ;
        RECT 3500.060 2468.720 3500.340 2469.000 ;
        RECT 3500.680 2468.720 3500.960 2469.000 ;
        RECT 3496.960 2468.100 3497.240 2468.380 ;
        RECT 3497.580 2468.100 3497.860 2468.380 ;
        RECT 3498.200 2468.100 3498.480 2468.380 ;
        RECT 3498.820 2468.100 3499.100 2468.380 ;
        RECT 3499.440 2468.100 3499.720 2468.380 ;
        RECT 3500.060 2468.100 3500.340 2468.380 ;
        RECT 3500.680 2468.100 3500.960 2468.380 ;
        RECT 3496.960 2467.480 3497.240 2467.760 ;
        RECT 3497.580 2467.480 3497.860 2467.760 ;
        RECT 3498.200 2467.480 3498.480 2467.760 ;
        RECT 3498.820 2467.480 3499.100 2467.760 ;
        RECT 3499.440 2467.480 3499.720 2467.760 ;
        RECT 3500.060 2467.480 3500.340 2467.760 ;
        RECT 3500.680 2467.480 3500.960 2467.760 ;
        RECT 3496.960 2466.860 3497.240 2467.140 ;
        RECT 3497.580 2466.860 3497.860 2467.140 ;
        RECT 3498.200 2466.860 3498.480 2467.140 ;
        RECT 3498.820 2466.860 3499.100 2467.140 ;
        RECT 3499.440 2466.860 3499.720 2467.140 ;
        RECT 3500.060 2466.860 3500.340 2467.140 ;
        RECT 3500.680 2466.860 3500.960 2467.140 ;
        RECT 3496.960 2466.240 3497.240 2466.520 ;
        RECT 3497.580 2466.240 3497.860 2466.520 ;
        RECT 3498.200 2466.240 3498.480 2466.520 ;
        RECT 3498.820 2466.240 3499.100 2466.520 ;
        RECT 3499.440 2466.240 3499.720 2466.520 ;
        RECT 3500.060 2466.240 3500.340 2466.520 ;
        RECT 3500.680 2466.240 3500.960 2466.520 ;
        RECT 3496.960 2465.620 3497.240 2465.900 ;
        RECT 3497.580 2465.620 3497.860 2465.900 ;
        RECT 3498.200 2465.620 3498.480 2465.900 ;
        RECT 3498.820 2465.620 3499.100 2465.900 ;
        RECT 3499.440 2465.620 3499.720 2465.900 ;
        RECT 3500.060 2465.620 3500.340 2465.900 ;
        RECT 3500.680 2465.620 3500.960 2465.900 ;
        RECT 3496.960 2465.000 3497.240 2465.280 ;
        RECT 3497.580 2465.000 3497.860 2465.280 ;
        RECT 3498.200 2465.000 3498.480 2465.280 ;
        RECT 3498.820 2465.000 3499.100 2465.280 ;
        RECT 3499.440 2465.000 3499.720 2465.280 ;
        RECT 3500.060 2465.000 3500.340 2465.280 ;
        RECT 3500.680 2465.000 3500.960 2465.280 ;
        RECT 3496.960 2464.380 3497.240 2464.660 ;
        RECT 3497.580 2464.380 3497.860 2464.660 ;
        RECT 3498.200 2464.380 3498.480 2464.660 ;
        RECT 3498.820 2464.380 3499.100 2464.660 ;
        RECT 3499.440 2464.380 3499.720 2464.660 ;
        RECT 3500.060 2464.380 3500.340 2464.660 ;
        RECT 3500.680 2464.380 3500.960 2464.660 ;
        RECT 3496.960 2463.760 3497.240 2464.040 ;
        RECT 3497.580 2463.760 3497.860 2464.040 ;
        RECT 3498.200 2463.760 3498.480 2464.040 ;
        RECT 3498.820 2463.760 3499.100 2464.040 ;
        RECT 3499.440 2463.760 3499.720 2464.040 ;
        RECT 3500.060 2463.760 3500.340 2464.040 ;
        RECT 3500.680 2463.760 3500.960 2464.040 ;
        RECT 3496.960 2463.140 3497.240 2463.420 ;
        RECT 3497.580 2463.140 3497.860 2463.420 ;
        RECT 3498.200 2463.140 3498.480 2463.420 ;
        RECT 3498.820 2463.140 3499.100 2463.420 ;
        RECT 3499.440 2463.140 3499.720 2463.420 ;
        RECT 3500.060 2463.140 3500.340 2463.420 ;
        RECT 3500.680 2463.140 3500.960 2463.420 ;
        RECT 3496.960 2462.520 3497.240 2462.800 ;
        RECT 3497.580 2462.520 3497.860 2462.800 ;
        RECT 3498.200 2462.520 3498.480 2462.800 ;
        RECT 3498.820 2462.520 3499.100 2462.800 ;
        RECT 3499.440 2462.520 3499.720 2462.800 ;
        RECT 3500.060 2462.520 3500.340 2462.800 ;
        RECT 3500.680 2462.520 3500.960 2462.800 ;
        RECT 3496.960 2461.900 3497.240 2462.180 ;
        RECT 3497.580 2461.900 3497.860 2462.180 ;
        RECT 3498.200 2461.900 3498.480 2462.180 ;
        RECT 3498.820 2461.900 3499.100 2462.180 ;
        RECT 3499.440 2461.900 3499.720 2462.180 ;
        RECT 3500.060 2461.900 3500.340 2462.180 ;
        RECT 3500.680 2461.900 3500.960 2462.180 ;
        RECT 3496.960 2461.280 3497.240 2461.560 ;
        RECT 3497.580 2461.280 3497.860 2461.560 ;
        RECT 3498.200 2461.280 3498.480 2461.560 ;
        RECT 3498.820 2461.280 3499.100 2461.560 ;
        RECT 3499.440 2461.280 3499.720 2461.560 ;
        RECT 3500.060 2461.280 3500.340 2461.560 ;
        RECT 3500.680 2461.280 3500.960 2461.560 ;
        RECT 3539.350 2470.610 3539.630 2470.890 ;
        RECT 3539.350 2469.990 3539.630 2470.270 ;
        RECT 3539.350 2469.370 3539.630 2469.650 ;
        RECT 3539.350 2468.750 3539.630 2469.030 ;
        RECT 3539.350 2468.130 3539.630 2468.410 ;
        RECT 3539.350 2467.510 3539.630 2467.790 ;
        RECT 3539.350 2466.890 3539.630 2467.170 ;
        RECT 3539.350 2466.270 3539.630 2466.550 ;
        RECT 3539.350 2465.650 3539.630 2465.930 ;
        RECT 3539.350 2465.030 3539.630 2465.310 ;
        RECT 3539.350 2464.410 3539.630 2464.690 ;
        RECT 3539.350 2463.790 3539.630 2464.070 ;
        RECT 3539.350 2463.170 3539.630 2463.450 ;
        RECT 3539.350 2462.550 3539.630 2462.830 ;
        RECT 3539.350 2461.930 3539.630 2462.210 ;
        RECT 3539.350 2461.310 3539.630 2461.590 ;
        RECT 3496.960 2458.730 3497.240 2459.010 ;
        RECT 3497.580 2458.730 3497.860 2459.010 ;
        RECT 3498.200 2458.730 3498.480 2459.010 ;
        RECT 3498.820 2458.730 3499.100 2459.010 ;
        RECT 3499.440 2458.730 3499.720 2459.010 ;
        RECT 3500.060 2458.730 3500.340 2459.010 ;
        RECT 3500.680 2458.730 3500.960 2459.010 ;
        RECT 3496.960 2458.110 3497.240 2458.390 ;
        RECT 3497.580 2458.110 3497.860 2458.390 ;
        RECT 3498.200 2458.110 3498.480 2458.390 ;
        RECT 3498.820 2458.110 3499.100 2458.390 ;
        RECT 3499.440 2458.110 3499.720 2458.390 ;
        RECT 3500.060 2458.110 3500.340 2458.390 ;
        RECT 3500.680 2458.110 3500.960 2458.390 ;
        RECT 3496.960 2457.490 3497.240 2457.770 ;
        RECT 3497.580 2457.490 3497.860 2457.770 ;
        RECT 3498.200 2457.490 3498.480 2457.770 ;
        RECT 3498.820 2457.490 3499.100 2457.770 ;
        RECT 3499.440 2457.490 3499.720 2457.770 ;
        RECT 3500.060 2457.490 3500.340 2457.770 ;
        RECT 3500.680 2457.490 3500.960 2457.770 ;
        RECT 3496.960 2456.870 3497.240 2457.150 ;
        RECT 3497.580 2456.870 3497.860 2457.150 ;
        RECT 3498.200 2456.870 3498.480 2457.150 ;
        RECT 3498.820 2456.870 3499.100 2457.150 ;
        RECT 3499.440 2456.870 3499.720 2457.150 ;
        RECT 3500.060 2456.870 3500.340 2457.150 ;
        RECT 3500.680 2456.870 3500.960 2457.150 ;
        RECT 3496.960 2456.250 3497.240 2456.530 ;
        RECT 3497.580 2456.250 3497.860 2456.530 ;
        RECT 3498.200 2456.250 3498.480 2456.530 ;
        RECT 3498.820 2456.250 3499.100 2456.530 ;
        RECT 3499.440 2456.250 3499.720 2456.530 ;
        RECT 3500.060 2456.250 3500.340 2456.530 ;
        RECT 3500.680 2456.250 3500.960 2456.530 ;
        RECT 3496.960 2455.630 3497.240 2455.910 ;
        RECT 3497.580 2455.630 3497.860 2455.910 ;
        RECT 3498.200 2455.630 3498.480 2455.910 ;
        RECT 3498.820 2455.630 3499.100 2455.910 ;
        RECT 3499.440 2455.630 3499.720 2455.910 ;
        RECT 3500.060 2455.630 3500.340 2455.910 ;
        RECT 3500.680 2455.630 3500.960 2455.910 ;
        RECT 3496.960 2455.010 3497.240 2455.290 ;
        RECT 3497.580 2455.010 3497.860 2455.290 ;
        RECT 3498.200 2455.010 3498.480 2455.290 ;
        RECT 3498.820 2455.010 3499.100 2455.290 ;
        RECT 3499.440 2455.010 3499.720 2455.290 ;
        RECT 3500.060 2455.010 3500.340 2455.290 ;
        RECT 3500.680 2455.010 3500.960 2455.290 ;
        RECT 3496.960 2454.390 3497.240 2454.670 ;
        RECT 3497.580 2454.390 3497.860 2454.670 ;
        RECT 3498.200 2454.390 3498.480 2454.670 ;
        RECT 3498.820 2454.390 3499.100 2454.670 ;
        RECT 3499.440 2454.390 3499.720 2454.670 ;
        RECT 3500.060 2454.390 3500.340 2454.670 ;
        RECT 3500.680 2454.390 3500.960 2454.670 ;
        RECT 3496.960 2453.770 3497.240 2454.050 ;
        RECT 3497.580 2453.770 3497.860 2454.050 ;
        RECT 3498.200 2453.770 3498.480 2454.050 ;
        RECT 3498.820 2453.770 3499.100 2454.050 ;
        RECT 3499.440 2453.770 3499.720 2454.050 ;
        RECT 3500.060 2453.770 3500.340 2454.050 ;
        RECT 3500.680 2453.770 3500.960 2454.050 ;
        RECT 3496.960 2453.150 3497.240 2453.430 ;
        RECT 3497.580 2453.150 3497.860 2453.430 ;
        RECT 3498.200 2453.150 3498.480 2453.430 ;
        RECT 3498.820 2453.150 3499.100 2453.430 ;
        RECT 3499.440 2453.150 3499.720 2453.430 ;
        RECT 3500.060 2453.150 3500.340 2453.430 ;
        RECT 3500.680 2453.150 3500.960 2453.430 ;
        RECT 3496.960 2452.530 3497.240 2452.810 ;
        RECT 3497.580 2452.530 3497.860 2452.810 ;
        RECT 3498.200 2452.530 3498.480 2452.810 ;
        RECT 3498.820 2452.530 3499.100 2452.810 ;
        RECT 3499.440 2452.530 3499.720 2452.810 ;
        RECT 3500.060 2452.530 3500.340 2452.810 ;
        RECT 3500.680 2452.530 3500.960 2452.810 ;
        RECT 3496.960 2451.910 3497.240 2452.190 ;
        RECT 3497.580 2451.910 3497.860 2452.190 ;
        RECT 3498.200 2451.910 3498.480 2452.190 ;
        RECT 3498.820 2451.910 3499.100 2452.190 ;
        RECT 3499.440 2451.910 3499.720 2452.190 ;
        RECT 3500.060 2451.910 3500.340 2452.190 ;
        RECT 3500.680 2451.910 3500.960 2452.190 ;
        RECT 3496.960 2451.290 3497.240 2451.570 ;
        RECT 3497.580 2451.290 3497.860 2451.570 ;
        RECT 3498.200 2451.290 3498.480 2451.570 ;
        RECT 3498.820 2451.290 3499.100 2451.570 ;
        RECT 3499.440 2451.290 3499.720 2451.570 ;
        RECT 3500.060 2451.290 3500.340 2451.570 ;
        RECT 3500.680 2451.290 3500.960 2451.570 ;
        RECT 3496.960 2450.670 3497.240 2450.950 ;
        RECT 3497.580 2450.670 3497.860 2450.950 ;
        RECT 3498.200 2450.670 3498.480 2450.950 ;
        RECT 3498.820 2450.670 3499.100 2450.950 ;
        RECT 3499.440 2450.670 3499.720 2450.950 ;
        RECT 3500.060 2450.670 3500.340 2450.950 ;
        RECT 3500.680 2450.670 3500.960 2450.950 ;
        RECT 3496.960 2450.050 3497.240 2450.330 ;
        RECT 3497.580 2450.050 3497.860 2450.330 ;
        RECT 3498.200 2450.050 3498.480 2450.330 ;
        RECT 3498.820 2450.050 3499.100 2450.330 ;
        RECT 3499.440 2450.050 3499.720 2450.330 ;
        RECT 3500.060 2450.050 3500.340 2450.330 ;
        RECT 3500.680 2450.050 3500.960 2450.330 ;
        RECT 3496.960 2449.430 3497.240 2449.710 ;
        RECT 3497.580 2449.430 3497.860 2449.710 ;
        RECT 3498.200 2449.430 3498.480 2449.710 ;
        RECT 3498.820 2449.430 3499.100 2449.710 ;
        RECT 3499.440 2449.430 3499.720 2449.710 ;
        RECT 3500.060 2449.430 3500.340 2449.710 ;
        RECT 3500.680 2449.430 3500.960 2449.710 ;
        RECT 3539.350 2458.760 3539.630 2459.040 ;
        RECT 3539.350 2458.140 3539.630 2458.420 ;
        RECT 3539.350 2457.520 3539.630 2457.800 ;
        RECT 3539.350 2456.900 3539.630 2457.180 ;
        RECT 3539.350 2456.280 3539.630 2456.560 ;
        RECT 3539.350 2455.660 3539.630 2455.940 ;
        RECT 3539.350 2455.040 3539.630 2455.320 ;
        RECT 3539.350 2454.420 3539.630 2454.700 ;
        RECT 3539.350 2453.800 3539.630 2454.080 ;
        RECT 3539.350 2453.180 3539.630 2453.460 ;
        RECT 3539.350 2452.560 3539.630 2452.840 ;
        RECT 3539.350 2451.940 3539.630 2452.220 ;
        RECT 3539.350 2451.320 3539.630 2451.600 ;
        RECT 3539.350 2450.700 3539.630 2450.980 ;
        RECT 3539.350 2450.080 3539.630 2450.360 ;
        RECT 3539.350 2449.460 3539.630 2449.740 ;
        RECT 3496.960 2445.200 3497.240 2445.480 ;
        RECT 3497.580 2445.200 3497.860 2445.480 ;
        RECT 3498.200 2445.200 3498.480 2445.480 ;
        RECT 3498.820 2445.200 3499.100 2445.480 ;
        RECT 3499.440 2445.200 3499.720 2445.480 ;
        RECT 3500.060 2445.200 3500.340 2445.480 ;
        RECT 3500.680 2445.200 3500.960 2445.480 ;
        RECT 3496.960 2444.580 3497.240 2444.860 ;
        RECT 3497.580 2444.580 3497.860 2444.860 ;
        RECT 3498.200 2444.580 3498.480 2444.860 ;
        RECT 3498.820 2444.580 3499.100 2444.860 ;
        RECT 3499.440 2444.580 3499.720 2444.860 ;
        RECT 3500.060 2444.580 3500.340 2444.860 ;
        RECT 3500.680 2444.580 3500.960 2444.860 ;
        RECT 3496.960 2443.960 3497.240 2444.240 ;
        RECT 3497.580 2443.960 3497.860 2444.240 ;
        RECT 3498.200 2443.960 3498.480 2444.240 ;
        RECT 3498.820 2443.960 3499.100 2444.240 ;
        RECT 3499.440 2443.960 3499.720 2444.240 ;
        RECT 3500.060 2443.960 3500.340 2444.240 ;
        RECT 3500.680 2443.960 3500.960 2444.240 ;
        RECT 3496.960 2443.340 3497.240 2443.620 ;
        RECT 3497.580 2443.340 3497.860 2443.620 ;
        RECT 3498.200 2443.340 3498.480 2443.620 ;
        RECT 3498.820 2443.340 3499.100 2443.620 ;
        RECT 3499.440 2443.340 3499.720 2443.620 ;
        RECT 3500.060 2443.340 3500.340 2443.620 ;
        RECT 3500.680 2443.340 3500.960 2443.620 ;
        RECT 3496.960 2442.720 3497.240 2443.000 ;
        RECT 3497.580 2442.720 3497.860 2443.000 ;
        RECT 3498.200 2442.720 3498.480 2443.000 ;
        RECT 3498.820 2442.720 3499.100 2443.000 ;
        RECT 3499.440 2442.720 3499.720 2443.000 ;
        RECT 3500.060 2442.720 3500.340 2443.000 ;
        RECT 3500.680 2442.720 3500.960 2443.000 ;
        RECT 3496.960 2442.100 3497.240 2442.380 ;
        RECT 3497.580 2442.100 3497.860 2442.380 ;
        RECT 3498.200 2442.100 3498.480 2442.380 ;
        RECT 3498.820 2442.100 3499.100 2442.380 ;
        RECT 3499.440 2442.100 3499.720 2442.380 ;
        RECT 3500.060 2442.100 3500.340 2442.380 ;
        RECT 3500.680 2442.100 3500.960 2442.380 ;
        RECT 3496.960 2441.480 3497.240 2441.760 ;
        RECT 3497.580 2441.480 3497.860 2441.760 ;
        RECT 3498.200 2441.480 3498.480 2441.760 ;
        RECT 3498.820 2441.480 3499.100 2441.760 ;
        RECT 3499.440 2441.480 3499.720 2441.760 ;
        RECT 3500.060 2441.480 3500.340 2441.760 ;
        RECT 3500.680 2441.480 3500.960 2441.760 ;
        RECT 3496.960 2440.860 3497.240 2441.140 ;
        RECT 3497.580 2440.860 3497.860 2441.140 ;
        RECT 3498.200 2440.860 3498.480 2441.140 ;
        RECT 3498.820 2440.860 3499.100 2441.140 ;
        RECT 3499.440 2440.860 3499.720 2441.140 ;
        RECT 3500.060 2440.860 3500.340 2441.140 ;
        RECT 3500.680 2440.860 3500.960 2441.140 ;
        RECT 3496.960 2440.240 3497.240 2440.520 ;
        RECT 3497.580 2440.240 3497.860 2440.520 ;
        RECT 3498.200 2440.240 3498.480 2440.520 ;
        RECT 3498.820 2440.240 3499.100 2440.520 ;
        RECT 3499.440 2440.240 3499.720 2440.520 ;
        RECT 3500.060 2440.240 3500.340 2440.520 ;
        RECT 3500.680 2440.240 3500.960 2440.520 ;
        RECT 3496.960 2439.620 3497.240 2439.900 ;
        RECT 3497.580 2439.620 3497.860 2439.900 ;
        RECT 3498.200 2439.620 3498.480 2439.900 ;
        RECT 3498.820 2439.620 3499.100 2439.900 ;
        RECT 3499.440 2439.620 3499.720 2439.900 ;
        RECT 3500.060 2439.620 3500.340 2439.900 ;
        RECT 3500.680 2439.620 3500.960 2439.900 ;
        RECT 3496.960 2439.000 3497.240 2439.280 ;
        RECT 3497.580 2439.000 3497.860 2439.280 ;
        RECT 3498.200 2439.000 3498.480 2439.280 ;
        RECT 3498.820 2439.000 3499.100 2439.280 ;
        RECT 3499.440 2439.000 3499.720 2439.280 ;
        RECT 3500.060 2439.000 3500.340 2439.280 ;
        RECT 3500.680 2439.000 3500.960 2439.280 ;
        RECT 3496.960 2438.380 3497.240 2438.660 ;
        RECT 3497.580 2438.380 3497.860 2438.660 ;
        RECT 3498.200 2438.380 3498.480 2438.660 ;
        RECT 3498.820 2438.380 3499.100 2438.660 ;
        RECT 3499.440 2438.380 3499.720 2438.660 ;
        RECT 3500.060 2438.380 3500.340 2438.660 ;
        RECT 3500.680 2438.380 3500.960 2438.660 ;
        RECT 3496.960 2437.760 3497.240 2438.040 ;
        RECT 3497.580 2437.760 3497.860 2438.040 ;
        RECT 3498.200 2437.760 3498.480 2438.040 ;
        RECT 3498.820 2437.760 3499.100 2438.040 ;
        RECT 3499.440 2437.760 3499.720 2438.040 ;
        RECT 3500.060 2437.760 3500.340 2438.040 ;
        RECT 3500.680 2437.760 3500.960 2438.040 ;
        RECT 3496.960 2437.140 3497.240 2437.420 ;
        RECT 3497.580 2437.140 3497.860 2437.420 ;
        RECT 3498.200 2437.140 3498.480 2437.420 ;
        RECT 3498.820 2437.140 3499.100 2437.420 ;
        RECT 3499.440 2437.140 3499.720 2437.420 ;
        RECT 3500.060 2437.140 3500.340 2437.420 ;
        RECT 3500.680 2437.140 3500.960 2437.420 ;
        RECT 3496.960 2436.520 3497.240 2436.800 ;
        RECT 3497.580 2436.520 3497.860 2436.800 ;
        RECT 3498.200 2436.520 3498.480 2436.800 ;
        RECT 3498.820 2436.520 3499.100 2436.800 ;
        RECT 3499.440 2436.520 3499.720 2436.800 ;
        RECT 3500.060 2436.520 3500.340 2436.800 ;
        RECT 3500.680 2436.520 3500.960 2436.800 ;
        RECT 3496.960 2435.900 3497.240 2436.180 ;
        RECT 3497.580 2435.900 3497.860 2436.180 ;
        RECT 3498.200 2435.900 3498.480 2436.180 ;
        RECT 3498.820 2435.900 3499.100 2436.180 ;
        RECT 3499.440 2435.900 3499.720 2436.180 ;
        RECT 3500.060 2435.900 3500.340 2436.180 ;
        RECT 3500.680 2435.900 3500.960 2436.180 ;
        RECT 3539.350 2445.230 3539.630 2445.510 ;
        RECT 3539.350 2444.610 3539.630 2444.890 ;
        RECT 3539.350 2443.990 3539.630 2444.270 ;
        RECT 3539.350 2443.370 3539.630 2443.650 ;
        RECT 3539.350 2442.750 3539.630 2443.030 ;
        RECT 3539.350 2442.130 3539.630 2442.410 ;
        RECT 3539.350 2441.510 3539.630 2441.790 ;
        RECT 3539.350 2440.890 3539.630 2441.170 ;
        RECT 3539.350 2440.270 3539.630 2440.550 ;
        RECT 3539.350 2439.650 3539.630 2439.930 ;
        RECT 3539.350 2439.030 3539.630 2439.310 ;
        RECT 3539.350 2438.410 3539.630 2438.690 ;
        RECT 3539.350 2437.790 3539.630 2438.070 ;
        RECT 3539.350 2437.170 3539.630 2437.450 ;
        RECT 3539.350 2436.550 3539.630 2436.830 ;
        RECT 3539.350 2435.930 3539.630 2436.210 ;
        RECT 3496.960 2433.350 3497.240 2433.630 ;
        RECT 3497.580 2433.350 3497.860 2433.630 ;
        RECT 3498.200 2433.350 3498.480 2433.630 ;
        RECT 3498.820 2433.350 3499.100 2433.630 ;
        RECT 3499.440 2433.350 3499.720 2433.630 ;
        RECT 3500.060 2433.350 3500.340 2433.630 ;
        RECT 3500.680 2433.350 3500.960 2433.630 ;
        RECT 3496.960 2432.730 3497.240 2433.010 ;
        RECT 3497.580 2432.730 3497.860 2433.010 ;
        RECT 3498.200 2432.730 3498.480 2433.010 ;
        RECT 3498.820 2432.730 3499.100 2433.010 ;
        RECT 3499.440 2432.730 3499.720 2433.010 ;
        RECT 3500.060 2432.730 3500.340 2433.010 ;
        RECT 3500.680 2432.730 3500.960 2433.010 ;
        RECT 3496.960 2432.110 3497.240 2432.390 ;
        RECT 3497.580 2432.110 3497.860 2432.390 ;
        RECT 3498.200 2432.110 3498.480 2432.390 ;
        RECT 3498.820 2432.110 3499.100 2432.390 ;
        RECT 3499.440 2432.110 3499.720 2432.390 ;
        RECT 3500.060 2432.110 3500.340 2432.390 ;
        RECT 3500.680 2432.110 3500.960 2432.390 ;
        RECT 3496.960 2431.490 3497.240 2431.770 ;
        RECT 3497.580 2431.490 3497.860 2431.770 ;
        RECT 3498.200 2431.490 3498.480 2431.770 ;
        RECT 3498.820 2431.490 3499.100 2431.770 ;
        RECT 3499.440 2431.490 3499.720 2431.770 ;
        RECT 3500.060 2431.490 3500.340 2431.770 ;
        RECT 3500.680 2431.490 3500.960 2431.770 ;
        RECT 3496.960 2430.870 3497.240 2431.150 ;
        RECT 3497.580 2430.870 3497.860 2431.150 ;
        RECT 3498.200 2430.870 3498.480 2431.150 ;
        RECT 3498.820 2430.870 3499.100 2431.150 ;
        RECT 3499.440 2430.870 3499.720 2431.150 ;
        RECT 3500.060 2430.870 3500.340 2431.150 ;
        RECT 3500.680 2430.870 3500.960 2431.150 ;
        RECT 3496.960 2430.250 3497.240 2430.530 ;
        RECT 3497.580 2430.250 3497.860 2430.530 ;
        RECT 3498.200 2430.250 3498.480 2430.530 ;
        RECT 3498.820 2430.250 3499.100 2430.530 ;
        RECT 3499.440 2430.250 3499.720 2430.530 ;
        RECT 3500.060 2430.250 3500.340 2430.530 ;
        RECT 3500.680 2430.250 3500.960 2430.530 ;
        RECT 3496.960 2429.630 3497.240 2429.910 ;
        RECT 3497.580 2429.630 3497.860 2429.910 ;
        RECT 3498.200 2429.630 3498.480 2429.910 ;
        RECT 3498.820 2429.630 3499.100 2429.910 ;
        RECT 3499.440 2429.630 3499.720 2429.910 ;
        RECT 3500.060 2429.630 3500.340 2429.910 ;
        RECT 3500.680 2429.630 3500.960 2429.910 ;
        RECT 3496.960 2429.010 3497.240 2429.290 ;
        RECT 3497.580 2429.010 3497.860 2429.290 ;
        RECT 3498.200 2429.010 3498.480 2429.290 ;
        RECT 3498.820 2429.010 3499.100 2429.290 ;
        RECT 3499.440 2429.010 3499.720 2429.290 ;
        RECT 3500.060 2429.010 3500.340 2429.290 ;
        RECT 3500.680 2429.010 3500.960 2429.290 ;
        RECT 3496.960 2428.390 3497.240 2428.670 ;
        RECT 3497.580 2428.390 3497.860 2428.670 ;
        RECT 3498.200 2428.390 3498.480 2428.670 ;
        RECT 3498.820 2428.390 3499.100 2428.670 ;
        RECT 3499.440 2428.390 3499.720 2428.670 ;
        RECT 3500.060 2428.390 3500.340 2428.670 ;
        RECT 3500.680 2428.390 3500.960 2428.670 ;
        RECT 3496.960 2427.770 3497.240 2428.050 ;
        RECT 3497.580 2427.770 3497.860 2428.050 ;
        RECT 3498.200 2427.770 3498.480 2428.050 ;
        RECT 3498.820 2427.770 3499.100 2428.050 ;
        RECT 3499.440 2427.770 3499.720 2428.050 ;
        RECT 3500.060 2427.770 3500.340 2428.050 ;
        RECT 3500.680 2427.770 3500.960 2428.050 ;
        RECT 3496.960 2427.150 3497.240 2427.430 ;
        RECT 3497.580 2427.150 3497.860 2427.430 ;
        RECT 3498.200 2427.150 3498.480 2427.430 ;
        RECT 3498.820 2427.150 3499.100 2427.430 ;
        RECT 3499.440 2427.150 3499.720 2427.430 ;
        RECT 3500.060 2427.150 3500.340 2427.430 ;
        RECT 3500.680 2427.150 3500.960 2427.430 ;
        RECT 3496.960 2426.530 3497.240 2426.810 ;
        RECT 3497.580 2426.530 3497.860 2426.810 ;
        RECT 3498.200 2426.530 3498.480 2426.810 ;
        RECT 3498.820 2426.530 3499.100 2426.810 ;
        RECT 3499.440 2426.530 3499.720 2426.810 ;
        RECT 3500.060 2426.530 3500.340 2426.810 ;
        RECT 3500.680 2426.530 3500.960 2426.810 ;
        RECT 3496.960 2425.910 3497.240 2426.190 ;
        RECT 3497.580 2425.910 3497.860 2426.190 ;
        RECT 3498.200 2425.910 3498.480 2426.190 ;
        RECT 3498.820 2425.910 3499.100 2426.190 ;
        RECT 3499.440 2425.910 3499.720 2426.190 ;
        RECT 3500.060 2425.910 3500.340 2426.190 ;
        RECT 3500.680 2425.910 3500.960 2426.190 ;
        RECT 3496.960 2425.290 3497.240 2425.570 ;
        RECT 3497.580 2425.290 3497.860 2425.570 ;
        RECT 3498.200 2425.290 3498.480 2425.570 ;
        RECT 3498.820 2425.290 3499.100 2425.570 ;
        RECT 3499.440 2425.290 3499.720 2425.570 ;
        RECT 3500.060 2425.290 3500.340 2425.570 ;
        RECT 3500.680 2425.290 3500.960 2425.570 ;
        RECT 3496.960 2424.670 3497.240 2424.950 ;
        RECT 3497.580 2424.670 3497.860 2424.950 ;
        RECT 3498.200 2424.670 3498.480 2424.950 ;
        RECT 3498.820 2424.670 3499.100 2424.950 ;
        RECT 3499.440 2424.670 3499.720 2424.950 ;
        RECT 3500.060 2424.670 3500.340 2424.950 ;
        RECT 3500.680 2424.670 3500.960 2424.950 ;
        RECT 3496.960 2424.050 3497.240 2424.330 ;
        RECT 3497.580 2424.050 3497.860 2424.330 ;
        RECT 3498.200 2424.050 3498.480 2424.330 ;
        RECT 3498.820 2424.050 3499.100 2424.330 ;
        RECT 3499.440 2424.050 3499.720 2424.330 ;
        RECT 3500.060 2424.050 3500.340 2424.330 ;
        RECT 3500.680 2424.050 3500.960 2424.330 ;
        RECT 3539.350 2433.380 3539.630 2433.660 ;
        RECT 3539.350 2432.760 3539.630 2433.040 ;
        RECT 3539.350 2432.140 3539.630 2432.420 ;
        RECT 3539.350 2431.520 3539.630 2431.800 ;
        RECT 3539.350 2430.900 3539.630 2431.180 ;
        RECT 3539.350 2430.280 3539.630 2430.560 ;
        RECT 3539.350 2429.660 3539.630 2429.940 ;
        RECT 3539.350 2429.040 3539.630 2429.320 ;
        RECT 3539.350 2428.420 3539.630 2428.700 ;
        RECT 3539.350 2427.800 3539.630 2428.080 ;
        RECT 3539.350 2427.180 3539.630 2427.460 ;
        RECT 3539.350 2426.560 3539.630 2426.840 ;
        RECT 3539.350 2425.940 3539.630 2426.220 ;
        RECT 3539.350 2425.320 3539.630 2425.600 ;
        RECT 3539.350 2424.700 3539.630 2424.980 ;
        RECT 3539.350 2424.080 3539.630 2424.360 ;
        RECT 3496.960 2420.330 3497.240 2420.610 ;
        RECT 3497.580 2420.330 3497.860 2420.610 ;
        RECT 3498.200 2420.330 3498.480 2420.610 ;
        RECT 3498.820 2420.330 3499.100 2420.610 ;
        RECT 3499.440 2420.330 3499.720 2420.610 ;
        RECT 3500.060 2420.330 3500.340 2420.610 ;
        RECT 3500.680 2420.330 3500.960 2420.610 ;
        RECT 3496.960 2419.710 3497.240 2419.990 ;
        RECT 3497.580 2419.710 3497.860 2419.990 ;
        RECT 3498.200 2419.710 3498.480 2419.990 ;
        RECT 3498.820 2419.710 3499.100 2419.990 ;
        RECT 3499.440 2419.710 3499.720 2419.990 ;
        RECT 3500.060 2419.710 3500.340 2419.990 ;
        RECT 3500.680 2419.710 3500.960 2419.990 ;
        RECT 3496.960 2419.090 3497.240 2419.370 ;
        RECT 3497.580 2419.090 3497.860 2419.370 ;
        RECT 3498.200 2419.090 3498.480 2419.370 ;
        RECT 3498.820 2419.090 3499.100 2419.370 ;
        RECT 3499.440 2419.090 3499.720 2419.370 ;
        RECT 3500.060 2419.090 3500.340 2419.370 ;
        RECT 3500.680 2419.090 3500.960 2419.370 ;
        RECT 3496.960 2418.470 3497.240 2418.750 ;
        RECT 3497.580 2418.470 3497.860 2418.750 ;
        RECT 3498.200 2418.470 3498.480 2418.750 ;
        RECT 3498.820 2418.470 3499.100 2418.750 ;
        RECT 3499.440 2418.470 3499.720 2418.750 ;
        RECT 3500.060 2418.470 3500.340 2418.750 ;
        RECT 3500.680 2418.470 3500.960 2418.750 ;
        RECT 3496.960 2417.850 3497.240 2418.130 ;
        RECT 3497.580 2417.850 3497.860 2418.130 ;
        RECT 3498.200 2417.850 3498.480 2418.130 ;
        RECT 3498.820 2417.850 3499.100 2418.130 ;
        RECT 3499.440 2417.850 3499.720 2418.130 ;
        RECT 3500.060 2417.850 3500.340 2418.130 ;
        RECT 3500.680 2417.850 3500.960 2418.130 ;
        RECT 3496.960 2417.230 3497.240 2417.510 ;
        RECT 3497.580 2417.230 3497.860 2417.510 ;
        RECT 3498.200 2417.230 3498.480 2417.510 ;
        RECT 3498.820 2417.230 3499.100 2417.510 ;
        RECT 3499.440 2417.230 3499.720 2417.510 ;
        RECT 3500.060 2417.230 3500.340 2417.510 ;
        RECT 3500.680 2417.230 3500.960 2417.510 ;
        RECT 3496.960 2416.610 3497.240 2416.890 ;
        RECT 3497.580 2416.610 3497.860 2416.890 ;
        RECT 3498.200 2416.610 3498.480 2416.890 ;
        RECT 3498.820 2416.610 3499.100 2416.890 ;
        RECT 3499.440 2416.610 3499.720 2416.890 ;
        RECT 3500.060 2416.610 3500.340 2416.890 ;
        RECT 3500.680 2416.610 3500.960 2416.890 ;
        RECT 3496.960 2415.990 3497.240 2416.270 ;
        RECT 3497.580 2415.990 3497.860 2416.270 ;
        RECT 3498.200 2415.990 3498.480 2416.270 ;
        RECT 3498.820 2415.990 3499.100 2416.270 ;
        RECT 3499.440 2415.990 3499.720 2416.270 ;
        RECT 3500.060 2415.990 3500.340 2416.270 ;
        RECT 3500.680 2415.990 3500.960 2416.270 ;
        RECT 3496.960 2415.370 3497.240 2415.650 ;
        RECT 3497.580 2415.370 3497.860 2415.650 ;
        RECT 3498.200 2415.370 3498.480 2415.650 ;
        RECT 3498.820 2415.370 3499.100 2415.650 ;
        RECT 3499.440 2415.370 3499.720 2415.650 ;
        RECT 3500.060 2415.370 3500.340 2415.650 ;
        RECT 3500.680 2415.370 3500.960 2415.650 ;
        RECT 3496.960 2414.750 3497.240 2415.030 ;
        RECT 3497.580 2414.750 3497.860 2415.030 ;
        RECT 3498.200 2414.750 3498.480 2415.030 ;
        RECT 3498.820 2414.750 3499.100 2415.030 ;
        RECT 3499.440 2414.750 3499.720 2415.030 ;
        RECT 3500.060 2414.750 3500.340 2415.030 ;
        RECT 3500.680 2414.750 3500.960 2415.030 ;
        RECT 3496.960 2414.130 3497.240 2414.410 ;
        RECT 3497.580 2414.130 3497.860 2414.410 ;
        RECT 3498.200 2414.130 3498.480 2414.410 ;
        RECT 3498.820 2414.130 3499.100 2414.410 ;
        RECT 3499.440 2414.130 3499.720 2414.410 ;
        RECT 3500.060 2414.130 3500.340 2414.410 ;
        RECT 3500.680 2414.130 3500.960 2414.410 ;
        RECT 3496.960 2413.510 3497.240 2413.790 ;
        RECT 3497.580 2413.510 3497.860 2413.790 ;
        RECT 3498.200 2413.510 3498.480 2413.790 ;
        RECT 3498.820 2413.510 3499.100 2413.790 ;
        RECT 3499.440 2413.510 3499.720 2413.790 ;
        RECT 3500.060 2413.510 3500.340 2413.790 ;
        RECT 3500.680 2413.510 3500.960 2413.790 ;
        RECT 3496.960 2412.890 3497.240 2413.170 ;
        RECT 3497.580 2412.890 3497.860 2413.170 ;
        RECT 3498.200 2412.890 3498.480 2413.170 ;
        RECT 3498.820 2412.890 3499.100 2413.170 ;
        RECT 3499.440 2412.890 3499.720 2413.170 ;
        RECT 3500.060 2412.890 3500.340 2413.170 ;
        RECT 3500.680 2412.890 3500.960 2413.170 ;
        RECT 3496.960 2412.270 3497.240 2412.550 ;
        RECT 3497.580 2412.270 3497.860 2412.550 ;
        RECT 3498.200 2412.270 3498.480 2412.550 ;
        RECT 3498.820 2412.270 3499.100 2412.550 ;
        RECT 3499.440 2412.270 3499.720 2412.550 ;
        RECT 3500.060 2412.270 3500.340 2412.550 ;
        RECT 3500.680 2412.270 3500.960 2412.550 ;
        RECT 3496.960 2411.650 3497.240 2411.930 ;
        RECT 3497.580 2411.650 3497.860 2411.930 ;
        RECT 3498.200 2411.650 3498.480 2411.930 ;
        RECT 3498.820 2411.650 3499.100 2411.930 ;
        RECT 3499.440 2411.650 3499.720 2411.930 ;
        RECT 3500.060 2411.650 3500.340 2411.930 ;
        RECT 3500.680 2411.650 3500.960 2411.930 ;
        RECT 3539.350 2420.390 3539.630 2420.670 ;
        RECT 3539.350 2419.770 3539.630 2420.050 ;
        RECT 3539.350 2419.150 3539.630 2419.430 ;
        RECT 3539.350 2418.530 3539.630 2418.810 ;
        RECT 3539.350 2417.910 3539.630 2418.190 ;
        RECT 3539.350 2417.290 3539.630 2417.570 ;
        RECT 3539.350 2416.670 3539.630 2416.950 ;
        RECT 3539.350 2416.050 3539.630 2416.330 ;
        RECT 3539.350 2415.430 3539.630 2415.710 ;
        RECT 3539.350 2414.810 3539.630 2415.090 ;
        RECT 3539.350 2414.190 3539.630 2414.470 ;
        RECT 3539.350 2413.570 3539.630 2413.850 ;
        RECT 3539.350 2412.950 3539.630 2413.230 ;
        RECT 3539.350 2412.330 3539.630 2412.610 ;
        RECT 3539.350 2411.710 3539.630 2411.990 ;
        RECT 3539.350 2268.010 3539.630 2268.290 ;
        RECT 3539.350 2267.390 3539.630 2267.670 ;
        RECT 3539.350 2266.770 3539.630 2267.050 ;
        RECT 3539.350 2266.150 3539.630 2266.430 ;
        RECT 3539.350 2265.530 3539.630 2265.810 ;
        RECT 3539.350 2264.910 3539.630 2265.190 ;
        RECT 3539.350 2264.290 3539.630 2264.570 ;
        RECT 3539.350 2263.670 3539.630 2263.950 ;
        RECT 3539.350 2263.050 3539.630 2263.330 ;
        RECT 3539.350 2262.430 3539.630 2262.710 ;
        RECT 3539.350 2261.810 3539.630 2262.090 ;
        RECT 3539.350 2261.190 3539.630 2261.470 ;
        RECT 3539.350 2260.570 3539.630 2260.850 ;
        RECT 3539.350 2259.950 3539.630 2260.230 ;
        RECT 3539.350 2259.330 3539.630 2259.610 ;
        RECT 3539.350 2255.610 3539.630 2255.890 ;
        RECT 3539.350 2254.990 3539.630 2255.270 ;
        RECT 3539.350 2254.370 3539.630 2254.650 ;
        RECT 3539.350 2253.750 3539.630 2254.030 ;
        RECT 3539.350 2253.130 3539.630 2253.410 ;
        RECT 3539.350 2252.510 3539.630 2252.790 ;
        RECT 3539.350 2251.890 3539.630 2252.170 ;
        RECT 3539.350 2251.270 3539.630 2251.550 ;
        RECT 3539.350 2250.650 3539.630 2250.930 ;
        RECT 3539.350 2250.030 3539.630 2250.310 ;
        RECT 3539.350 2249.410 3539.630 2249.690 ;
        RECT 3539.350 2248.790 3539.630 2249.070 ;
        RECT 3539.350 2248.170 3539.630 2248.450 ;
        RECT 3539.350 2247.550 3539.630 2247.830 ;
        RECT 3539.350 2246.930 3539.630 2247.210 ;
        RECT 3539.350 2246.310 3539.630 2246.590 ;
        RECT 3539.350 2243.760 3539.630 2244.040 ;
        RECT 3539.350 2243.140 3539.630 2243.420 ;
        RECT 3539.350 2242.520 3539.630 2242.800 ;
        RECT 3539.350 2241.900 3539.630 2242.180 ;
        RECT 3539.350 2241.280 3539.630 2241.560 ;
        RECT 3539.350 2240.660 3539.630 2240.940 ;
        RECT 3539.350 2240.040 3539.630 2240.320 ;
        RECT 3539.350 2239.420 3539.630 2239.700 ;
        RECT 3539.350 2238.800 3539.630 2239.080 ;
        RECT 3539.350 2238.180 3539.630 2238.460 ;
        RECT 3539.350 2237.560 3539.630 2237.840 ;
        RECT 3539.350 2236.940 3539.630 2237.220 ;
        RECT 3539.350 2236.320 3539.630 2236.600 ;
        RECT 3539.350 2235.700 3539.630 2235.980 ;
        RECT 3539.350 2235.080 3539.630 2235.360 ;
        RECT 3539.350 2234.460 3539.630 2234.740 ;
        RECT 3539.350 2230.230 3539.630 2230.510 ;
        RECT 3539.350 2229.610 3539.630 2229.890 ;
        RECT 3539.350 2228.990 3539.630 2229.270 ;
        RECT 3539.350 2228.370 3539.630 2228.650 ;
        RECT 3539.350 2227.750 3539.630 2228.030 ;
        RECT 3539.350 2227.130 3539.630 2227.410 ;
        RECT 3539.350 2226.510 3539.630 2226.790 ;
        RECT 3539.350 2225.890 3539.630 2226.170 ;
        RECT 3539.350 2225.270 3539.630 2225.550 ;
        RECT 3539.350 2224.650 3539.630 2224.930 ;
        RECT 3539.350 2224.030 3539.630 2224.310 ;
        RECT 3539.350 2223.410 3539.630 2223.690 ;
        RECT 3539.350 2222.790 3539.630 2223.070 ;
        RECT 3539.350 2222.170 3539.630 2222.450 ;
        RECT 3539.350 2221.550 3539.630 2221.830 ;
        RECT 3539.350 2220.930 3539.630 2221.210 ;
        RECT 3539.350 2218.380 3539.630 2218.660 ;
        RECT 3539.350 2217.760 3539.630 2218.040 ;
        RECT 3539.350 2217.140 3539.630 2217.420 ;
        RECT 3539.350 2216.520 3539.630 2216.800 ;
        RECT 3539.350 2215.900 3539.630 2216.180 ;
        RECT 3539.350 2215.280 3539.630 2215.560 ;
        RECT 3539.350 2214.660 3539.630 2214.940 ;
        RECT 3539.350 2214.040 3539.630 2214.320 ;
        RECT 3539.350 2213.420 3539.630 2213.700 ;
        RECT 3539.350 2212.800 3539.630 2213.080 ;
        RECT 3539.350 2212.180 3539.630 2212.460 ;
        RECT 3539.350 2211.560 3539.630 2211.840 ;
        RECT 3539.350 2210.940 3539.630 2211.220 ;
        RECT 3539.350 2210.320 3539.630 2210.600 ;
        RECT 3539.350 2209.700 3539.630 2209.980 ;
        RECT 3539.350 2209.080 3539.630 2209.360 ;
        RECT 3539.350 2205.390 3539.630 2205.670 ;
        RECT 3539.350 2204.770 3539.630 2205.050 ;
        RECT 3539.350 2204.150 3539.630 2204.430 ;
        RECT 3539.350 2203.530 3539.630 2203.810 ;
        RECT 3539.350 2202.910 3539.630 2203.190 ;
        RECT 3539.350 2202.290 3539.630 2202.570 ;
        RECT 3539.350 2201.670 3539.630 2201.950 ;
        RECT 3539.350 2201.050 3539.630 2201.330 ;
        RECT 3539.350 2200.430 3539.630 2200.710 ;
        RECT 3539.350 2199.810 3539.630 2200.090 ;
        RECT 3539.350 2199.190 3539.630 2199.470 ;
        RECT 3539.350 2198.570 3539.630 2198.850 ;
        RECT 3539.350 2197.950 3539.630 2198.230 ;
        RECT 3539.350 2197.330 3539.630 2197.610 ;
        RECT 3539.350 2196.710 3539.630 2196.990 ;
        RECT 3539.350 2053.010 3539.630 2053.290 ;
        RECT 3539.350 2052.390 3539.630 2052.670 ;
        RECT 3539.350 2051.770 3539.630 2052.050 ;
        RECT 3539.350 2051.150 3539.630 2051.430 ;
        RECT 3539.350 2050.530 3539.630 2050.810 ;
        RECT 3539.350 2049.910 3539.630 2050.190 ;
        RECT 3539.350 2049.290 3539.630 2049.570 ;
        RECT 3539.350 2048.670 3539.630 2048.950 ;
        RECT 3539.350 2048.050 3539.630 2048.330 ;
        RECT 3539.350 2047.430 3539.630 2047.710 ;
        RECT 3539.350 2046.810 3539.630 2047.090 ;
        RECT 3539.350 2046.190 3539.630 2046.470 ;
        RECT 3539.350 2045.570 3539.630 2045.850 ;
        RECT 3539.350 2044.950 3539.630 2045.230 ;
        RECT 3539.350 2044.330 3539.630 2044.610 ;
        RECT 3539.350 2040.610 3539.630 2040.890 ;
        RECT 3539.350 2039.990 3539.630 2040.270 ;
        RECT 3539.350 2039.370 3539.630 2039.650 ;
        RECT 3539.350 2038.750 3539.630 2039.030 ;
        RECT 3539.350 2038.130 3539.630 2038.410 ;
        RECT 3539.350 2037.510 3539.630 2037.790 ;
        RECT 3539.350 2036.890 3539.630 2037.170 ;
        RECT 3539.350 2036.270 3539.630 2036.550 ;
        RECT 3539.350 2035.650 3539.630 2035.930 ;
        RECT 3539.350 2035.030 3539.630 2035.310 ;
        RECT 3539.350 2034.410 3539.630 2034.690 ;
        RECT 3539.350 2033.790 3539.630 2034.070 ;
        RECT 3539.350 2033.170 3539.630 2033.450 ;
        RECT 3539.350 2032.550 3539.630 2032.830 ;
        RECT 3539.350 2031.930 3539.630 2032.210 ;
        RECT 3539.350 2031.310 3539.630 2031.590 ;
        RECT 3539.350 2028.760 3539.630 2029.040 ;
        RECT 3539.350 2028.140 3539.630 2028.420 ;
        RECT 3539.350 2027.520 3539.630 2027.800 ;
        RECT 3539.350 2026.900 3539.630 2027.180 ;
        RECT 3539.350 2026.280 3539.630 2026.560 ;
        RECT 3539.350 2025.660 3539.630 2025.940 ;
        RECT 3539.350 2025.040 3539.630 2025.320 ;
        RECT 3539.350 2024.420 3539.630 2024.700 ;
        RECT 3539.350 2023.800 3539.630 2024.080 ;
        RECT 3539.350 2023.180 3539.630 2023.460 ;
        RECT 3539.350 2022.560 3539.630 2022.840 ;
        RECT 3539.350 2021.940 3539.630 2022.220 ;
        RECT 3539.350 2021.320 3539.630 2021.600 ;
        RECT 3539.350 2020.700 3539.630 2020.980 ;
        RECT 3539.350 2020.080 3539.630 2020.360 ;
        RECT 3539.350 2019.460 3539.630 2019.740 ;
        RECT 3539.350 2015.230 3539.630 2015.510 ;
        RECT 3539.350 2014.610 3539.630 2014.890 ;
        RECT 3539.350 2013.990 3539.630 2014.270 ;
        RECT 3539.350 2013.370 3539.630 2013.650 ;
        RECT 3539.350 2012.750 3539.630 2013.030 ;
        RECT 3539.350 2012.130 3539.630 2012.410 ;
        RECT 3539.350 2011.510 3539.630 2011.790 ;
        RECT 3539.350 2010.890 3539.630 2011.170 ;
        RECT 3539.350 2010.270 3539.630 2010.550 ;
        RECT 3539.350 2009.650 3539.630 2009.930 ;
        RECT 3539.350 2009.030 3539.630 2009.310 ;
        RECT 3539.350 2008.410 3539.630 2008.690 ;
        RECT 3539.350 2007.790 3539.630 2008.070 ;
        RECT 3539.350 2007.170 3539.630 2007.450 ;
        RECT 3539.350 2006.550 3539.630 2006.830 ;
        RECT 3539.350 2005.930 3539.630 2006.210 ;
        RECT 3539.350 2003.380 3539.630 2003.660 ;
        RECT 3539.350 2002.760 3539.630 2003.040 ;
        RECT 3539.350 2002.140 3539.630 2002.420 ;
        RECT 3539.350 2001.520 3539.630 2001.800 ;
        RECT 3539.350 2000.900 3539.630 2001.180 ;
        RECT 3539.350 2000.280 3539.630 2000.560 ;
        RECT 3539.350 1999.660 3539.630 1999.940 ;
        RECT 3539.350 1999.040 3539.630 1999.320 ;
        RECT 3539.350 1998.420 3539.630 1998.700 ;
        RECT 3539.350 1997.800 3539.630 1998.080 ;
        RECT 3539.350 1997.180 3539.630 1997.460 ;
        RECT 3539.350 1996.560 3539.630 1996.840 ;
        RECT 3539.350 1995.940 3539.630 1996.220 ;
        RECT 3539.350 1995.320 3539.630 1995.600 ;
        RECT 3539.350 1994.700 3539.630 1994.980 ;
        RECT 3539.350 1994.080 3539.630 1994.360 ;
        RECT 3539.350 1990.390 3539.630 1990.670 ;
        RECT 3539.350 1989.770 3539.630 1990.050 ;
        RECT 3539.350 1989.150 3539.630 1989.430 ;
        RECT 3539.350 1988.530 3539.630 1988.810 ;
        RECT 3539.350 1987.910 3539.630 1988.190 ;
        RECT 3539.350 1987.290 3539.630 1987.570 ;
        RECT 3539.350 1986.670 3539.630 1986.950 ;
        RECT 3539.350 1986.050 3539.630 1986.330 ;
        RECT 3539.350 1985.430 3539.630 1985.710 ;
        RECT 3539.350 1984.810 3539.630 1985.090 ;
        RECT 3539.350 1984.190 3539.630 1984.470 ;
        RECT 3539.350 1983.570 3539.630 1983.850 ;
        RECT 3539.350 1982.950 3539.630 1983.230 ;
        RECT 3539.350 1982.330 3539.630 1982.610 ;
        RECT 3539.350 1981.710 3539.630 1981.990 ;
        RECT 3497.720 1871.865 3498.000 1872.145 ;
        RECT 3499.220 1871.865 3499.500 1872.145 ;
        RECT 3500.720 1871.865 3501.000 1872.145 ;
        RECT 3497.720 1870.865 3498.000 1871.145 ;
        RECT 3499.220 1870.865 3499.500 1871.145 ;
        RECT 3500.720 1870.865 3501.000 1871.145 ;
        RECT 3497.220 1834.490 3497.500 1834.770 ;
        RECT 3498.720 1834.490 3499.000 1834.770 ;
        RECT 3500.220 1834.490 3500.500 1834.770 ;
        RECT 3497.220 1799.490 3497.500 1799.770 ;
        RECT 3498.720 1799.490 3499.000 1799.770 ;
        RECT 3500.220 1799.490 3500.500 1799.770 ;
        RECT 3497.220 1764.490 3497.500 1764.770 ;
        RECT 3498.720 1764.490 3499.000 1764.770 ;
        RECT 3500.220 1764.490 3500.500 1764.770 ;
        RECT 3497.720 1691.865 3498.000 1692.145 ;
        RECT 3499.220 1691.865 3499.500 1692.145 ;
        RECT 3500.720 1691.865 3501.000 1692.145 ;
        RECT 3497.720 1690.865 3498.000 1691.145 ;
        RECT 3499.220 1690.865 3499.500 1691.145 ;
        RECT 3500.720 1690.865 3501.000 1691.145 ;
        RECT 3497.485 1666.835 3497.765 1667.115 ;
        RECT 3498.985 1666.835 3499.265 1667.115 ;
        RECT 3500.485 1666.835 3500.765 1667.115 ;
        RECT 3497.260 1647.920 3497.540 1648.200 ;
        RECT 3497.880 1647.920 3498.160 1648.200 ;
        RECT 3498.500 1647.920 3498.780 1648.200 ;
        RECT 3499.120 1647.920 3499.400 1648.200 ;
        RECT 3499.740 1647.920 3500.020 1648.200 ;
        RECT 3500.360 1647.920 3500.640 1648.200 ;
        RECT 3500.980 1647.920 3501.260 1648.200 ;
        RECT 3497.260 1647.300 3497.540 1647.580 ;
        RECT 3497.880 1647.300 3498.160 1647.580 ;
        RECT 3498.500 1647.300 3498.780 1647.580 ;
        RECT 3499.120 1647.300 3499.400 1647.580 ;
        RECT 3499.740 1647.300 3500.020 1647.580 ;
        RECT 3500.360 1647.300 3500.640 1647.580 ;
        RECT 3500.980 1647.300 3501.260 1647.580 ;
        RECT 3497.260 1646.680 3497.540 1646.960 ;
        RECT 3497.880 1646.680 3498.160 1646.960 ;
        RECT 3498.500 1646.680 3498.780 1646.960 ;
        RECT 3499.120 1646.680 3499.400 1646.960 ;
        RECT 3499.740 1646.680 3500.020 1646.960 ;
        RECT 3500.360 1646.680 3500.640 1646.960 ;
        RECT 3500.980 1646.680 3501.260 1646.960 ;
        RECT 3497.260 1646.060 3497.540 1646.340 ;
        RECT 3497.880 1646.060 3498.160 1646.340 ;
        RECT 3498.500 1646.060 3498.780 1646.340 ;
        RECT 3499.120 1646.060 3499.400 1646.340 ;
        RECT 3499.740 1646.060 3500.020 1646.340 ;
        RECT 3500.360 1646.060 3500.640 1646.340 ;
        RECT 3500.980 1646.060 3501.260 1646.340 ;
        RECT 3497.260 1645.440 3497.540 1645.720 ;
        RECT 3497.880 1645.440 3498.160 1645.720 ;
        RECT 3498.500 1645.440 3498.780 1645.720 ;
        RECT 3499.120 1645.440 3499.400 1645.720 ;
        RECT 3499.740 1645.440 3500.020 1645.720 ;
        RECT 3500.360 1645.440 3500.640 1645.720 ;
        RECT 3500.980 1645.440 3501.260 1645.720 ;
        RECT 3497.260 1644.820 3497.540 1645.100 ;
        RECT 3497.880 1644.820 3498.160 1645.100 ;
        RECT 3498.500 1644.820 3498.780 1645.100 ;
        RECT 3499.120 1644.820 3499.400 1645.100 ;
        RECT 3499.740 1644.820 3500.020 1645.100 ;
        RECT 3500.360 1644.820 3500.640 1645.100 ;
        RECT 3500.980 1644.820 3501.260 1645.100 ;
        RECT 3497.260 1644.200 3497.540 1644.480 ;
        RECT 3497.880 1644.200 3498.160 1644.480 ;
        RECT 3498.500 1644.200 3498.780 1644.480 ;
        RECT 3499.120 1644.200 3499.400 1644.480 ;
        RECT 3499.740 1644.200 3500.020 1644.480 ;
        RECT 3500.360 1644.200 3500.640 1644.480 ;
        RECT 3500.980 1644.200 3501.260 1644.480 ;
        RECT 3497.220 1619.490 3497.500 1619.770 ;
        RECT 3498.720 1619.490 3499.000 1619.770 ;
        RECT 3500.220 1619.490 3500.500 1619.770 ;
        RECT 3497.220 1584.490 3497.500 1584.770 ;
        RECT 3498.720 1584.490 3499.000 1584.770 ;
        RECT 3500.220 1584.490 3500.500 1584.770 ;
        RECT 3497.220 1549.490 3497.500 1549.770 ;
        RECT 3498.720 1549.490 3499.000 1549.770 ;
        RECT 3500.220 1549.490 3500.500 1549.770 ;
        RECT 3497.260 1528.650 3497.540 1528.930 ;
        RECT 3497.880 1528.650 3498.160 1528.930 ;
        RECT 3498.500 1528.650 3498.780 1528.930 ;
        RECT 3499.120 1528.650 3499.400 1528.930 ;
        RECT 3499.740 1528.650 3500.020 1528.930 ;
        RECT 3500.360 1528.650 3500.640 1528.930 ;
        RECT 3500.980 1528.650 3501.260 1528.930 ;
        RECT 3497.260 1528.030 3497.540 1528.310 ;
        RECT 3497.880 1528.030 3498.160 1528.310 ;
        RECT 3498.500 1528.030 3498.780 1528.310 ;
        RECT 3499.120 1528.030 3499.400 1528.310 ;
        RECT 3499.740 1528.030 3500.020 1528.310 ;
        RECT 3500.360 1528.030 3500.640 1528.310 ;
        RECT 3500.980 1528.030 3501.260 1528.310 ;
        RECT 3497.260 1527.410 3497.540 1527.690 ;
        RECT 3497.880 1527.410 3498.160 1527.690 ;
        RECT 3498.500 1527.410 3498.780 1527.690 ;
        RECT 3499.120 1527.410 3499.400 1527.690 ;
        RECT 3499.740 1527.410 3500.020 1527.690 ;
        RECT 3500.360 1527.410 3500.640 1527.690 ;
        RECT 3500.980 1527.410 3501.260 1527.690 ;
        RECT 3497.260 1526.790 3497.540 1527.070 ;
        RECT 3497.880 1526.790 3498.160 1527.070 ;
        RECT 3498.500 1526.790 3498.780 1527.070 ;
        RECT 3499.120 1526.790 3499.400 1527.070 ;
        RECT 3499.740 1526.790 3500.020 1527.070 ;
        RECT 3500.360 1526.790 3500.640 1527.070 ;
        RECT 3500.980 1526.790 3501.260 1527.070 ;
        RECT 3497.260 1526.170 3497.540 1526.450 ;
        RECT 3497.880 1526.170 3498.160 1526.450 ;
        RECT 3498.500 1526.170 3498.780 1526.450 ;
        RECT 3499.120 1526.170 3499.400 1526.450 ;
        RECT 3499.740 1526.170 3500.020 1526.450 ;
        RECT 3500.360 1526.170 3500.640 1526.450 ;
        RECT 3500.980 1526.170 3501.260 1526.450 ;
        RECT 3497.260 1525.550 3497.540 1525.830 ;
        RECT 3497.880 1525.550 3498.160 1525.830 ;
        RECT 3498.500 1525.550 3498.780 1525.830 ;
        RECT 3499.120 1525.550 3499.400 1525.830 ;
        RECT 3499.740 1525.550 3500.020 1525.830 ;
        RECT 3500.360 1525.550 3500.640 1525.830 ;
        RECT 3500.980 1525.550 3501.260 1525.830 ;
        RECT 3497.260 1524.930 3497.540 1525.210 ;
        RECT 3497.880 1524.930 3498.160 1525.210 ;
        RECT 3498.500 1524.930 3498.780 1525.210 ;
        RECT 3499.120 1524.930 3499.400 1525.210 ;
        RECT 3499.740 1524.930 3500.020 1525.210 ;
        RECT 3500.360 1524.930 3500.640 1525.210 ;
        RECT 3500.980 1524.930 3501.260 1525.210 ;
        RECT 3497.485 1451.835 3497.765 1452.115 ;
        RECT 3498.985 1451.835 3499.265 1452.115 ;
        RECT 3500.485 1451.835 3500.765 1452.115 ;
        RECT 3497.220 1404.490 3497.500 1404.770 ;
        RECT 3498.720 1404.490 3499.000 1404.770 ;
        RECT 3500.220 1404.490 3500.500 1404.770 ;
        RECT 3497.220 1369.490 3497.500 1369.770 ;
        RECT 3498.720 1369.490 3499.000 1369.770 ;
        RECT 3500.220 1369.490 3500.500 1369.770 ;
        RECT 3497.220 1342.755 3497.500 1343.035 ;
        RECT 3498.720 1342.755 3499.000 1343.035 ;
        RECT 3500.220 1342.755 3500.500 1343.035 ;
        RECT 3497.220 1334.490 3497.500 1334.770 ;
        RECT 3498.720 1334.490 3499.000 1334.770 ;
        RECT 3500.220 1334.490 3500.500 1334.770 ;
        RECT 3497.485 1236.835 3497.765 1237.115 ;
        RECT 3498.985 1236.835 3499.265 1237.115 ;
        RECT 3500.485 1236.835 3500.765 1237.115 ;
        RECT 3497.220 1189.575 3497.500 1189.855 ;
        RECT 3498.720 1189.575 3499.000 1189.855 ;
        RECT 3500.220 1189.575 3500.500 1189.855 ;
        RECT 3497.220 1154.490 3497.500 1154.770 ;
        RECT 3498.720 1154.490 3499.000 1154.770 ;
        RECT 3500.220 1154.490 3500.500 1154.770 ;
        RECT 3497.220 1119.490 3497.500 1119.770 ;
        RECT 3498.720 1119.490 3499.000 1119.770 ;
        RECT 3500.220 1119.490 3500.500 1119.770 ;
        RECT 3497.220 1036.395 3497.500 1036.675 ;
        RECT 3498.720 1036.395 3499.000 1036.675 ;
        RECT 3500.220 1036.395 3500.500 1036.675 ;
        RECT 3497.485 1021.835 3497.765 1022.115 ;
        RECT 3498.985 1021.835 3499.265 1022.115 ;
        RECT 3500.485 1021.835 3500.765 1022.115 ;
        RECT 3497.220 974.490 3497.500 974.770 ;
        RECT 3498.720 974.490 3499.000 974.770 ;
        RECT 3500.220 974.490 3500.500 974.770 ;
        RECT 3497.220 939.490 3497.500 939.770 ;
        RECT 3498.720 939.490 3499.000 939.770 ;
        RECT 3500.220 939.490 3500.500 939.770 ;
        RECT 3497.220 904.490 3497.500 904.770 ;
        RECT 3498.720 904.490 3499.000 904.770 ;
        RECT 3500.220 904.490 3500.500 904.770 ;
        RECT 3497.220 883.215 3497.500 883.495 ;
        RECT 3498.720 883.215 3499.000 883.495 ;
        RECT 3500.220 883.215 3500.500 883.495 ;
        RECT 3497.485 806.835 3497.765 807.115 ;
        RECT 3498.985 806.835 3499.265 807.115 ;
        RECT 3500.485 806.835 3500.765 807.115 ;
        RECT 3497.220 759.490 3497.500 759.770 ;
        RECT 3498.720 759.490 3499.000 759.770 ;
        RECT 3500.220 759.490 3500.500 759.770 ;
        RECT 3497.220 730.035 3497.500 730.315 ;
        RECT 3498.720 730.035 3499.000 730.315 ;
        RECT 3500.220 730.035 3500.500 730.315 ;
        RECT 3497.220 724.490 3497.500 724.770 ;
        RECT 3498.720 724.490 3499.000 724.770 ;
        RECT 3500.220 724.490 3500.500 724.770 ;
        RECT 3497.220 689.490 3497.500 689.770 ;
        RECT 3498.720 689.490 3499.000 689.770 ;
        RECT 3500.220 689.490 3500.500 689.770 ;
        RECT 3497.220 668.735 3497.500 669.015 ;
        RECT 3498.720 668.735 3499.000 669.015 ;
        RECT 3500.220 668.735 3500.500 669.015 ;
        RECT 3497.485 591.835 3497.765 592.115 ;
        RECT 3498.985 591.835 3499.265 592.115 ;
        RECT 3500.485 591.835 3500.765 592.115 ;
        RECT 3497.220 544.490 3497.500 544.770 ;
        RECT 3498.720 544.490 3499.000 544.770 ;
        RECT 3500.220 544.490 3500.500 544.770 ;
        RECT 3497.220 509.490 3497.500 509.770 ;
        RECT 3498.720 509.490 3499.000 509.770 ;
        RECT 3500.220 509.490 3500.500 509.770 ;
        RECT 3497.220 474.490 3497.500 474.770 ;
        RECT 3498.720 474.490 3499.000 474.770 ;
        RECT 3500.220 474.490 3500.500 474.770 ;
        RECT 3497.260 392.760 3497.540 393.040 ;
        RECT 3497.880 392.760 3498.160 393.040 ;
        RECT 3498.500 392.760 3498.780 393.040 ;
        RECT 3499.120 392.760 3499.400 393.040 ;
        RECT 3499.740 392.760 3500.020 393.040 ;
        RECT 3500.360 392.760 3500.640 393.040 ;
        RECT 3500.980 392.760 3501.260 393.040 ;
        RECT 3497.260 392.140 3497.540 392.420 ;
        RECT 3497.880 392.140 3498.160 392.420 ;
        RECT 3498.500 392.140 3498.780 392.420 ;
        RECT 3499.120 392.140 3499.400 392.420 ;
        RECT 3499.740 392.140 3500.020 392.420 ;
        RECT 3500.360 392.140 3500.640 392.420 ;
        RECT 3500.980 392.140 3501.260 392.420 ;
        RECT 3497.260 391.520 3497.540 391.800 ;
        RECT 3497.880 391.520 3498.160 391.800 ;
        RECT 3498.500 391.520 3498.780 391.800 ;
        RECT 3499.120 391.520 3499.400 391.800 ;
        RECT 3499.740 391.520 3500.020 391.800 ;
        RECT 3500.360 391.520 3500.640 391.800 ;
        RECT 3500.980 391.520 3501.260 391.800 ;
        RECT 3497.260 390.900 3497.540 391.180 ;
        RECT 3497.880 390.900 3498.160 391.180 ;
        RECT 3498.500 390.900 3498.780 391.180 ;
        RECT 3499.120 390.900 3499.400 391.180 ;
        RECT 3499.740 390.900 3500.020 391.180 ;
        RECT 3500.360 390.900 3500.640 391.180 ;
        RECT 3500.980 390.900 3501.260 391.180 ;
        RECT 3497.260 390.280 3497.540 390.560 ;
        RECT 3497.880 390.280 3498.160 390.560 ;
        RECT 3498.500 390.280 3498.780 390.560 ;
        RECT 3499.120 390.280 3499.400 390.560 ;
        RECT 3499.740 390.280 3500.020 390.560 ;
        RECT 3500.360 390.280 3500.640 390.560 ;
        RECT 3500.980 390.280 3501.260 390.560 ;
        RECT 3497.260 389.660 3497.540 389.940 ;
        RECT 3497.880 389.660 3498.160 389.940 ;
        RECT 3498.500 389.660 3498.780 389.940 ;
        RECT 3499.120 389.660 3499.400 389.940 ;
        RECT 3499.740 389.660 3500.020 389.940 ;
        RECT 3500.360 389.660 3500.640 389.940 ;
        RECT 3500.980 389.660 3501.260 389.940 ;
        RECT 3497.260 389.040 3497.540 389.320 ;
        RECT 3497.880 389.040 3498.160 389.320 ;
        RECT 3498.500 389.040 3498.780 389.320 ;
        RECT 3499.120 389.040 3499.400 389.320 ;
        RECT 3499.740 389.040 3500.020 389.320 ;
        RECT 3500.360 389.040 3500.640 389.320 ;
        RECT 3500.980 389.040 3501.260 389.320 ;
        RECT 3497.485 376.835 3497.765 377.115 ;
        RECT 3498.985 376.835 3499.265 377.115 ;
        RECT 3500.485 376.835 3500.765 377.115 ;
        RECT 3490.300 374.760 3490.580 375.040 ;
        RECT 3491.800 374.760 3492.080 375.040 ;
        RECT 3493.300 374.760 3493.580 375.040 ;
      LAYER Metal5 ;
        RECT 380.575 4729.550 400.390 4730.550 ;
        RECT 380.575 4727.550 382.175 4729.550 ;
        RECT 384.575 4727.550 393.390 4728.550 ;
        RECT 534.620 4711.610 536.220 4723.440 ;
        RECT 552.120 4716.520 553.720 4723.120 ;
        RECT 569.620 4711.610 571.220 4723.440 ;
        RECT 587.120 4716.520 588.720 4723.120 ;
        RECT 604.620 4711.610 606.220 4723.440 ;
        RECT 622.120 4716.520 623.720 4723.120 ;
        RECT 809.620 4711.610 811.220 4723.440 ;
        RECT 827.120 4716.520 828.720 4723.120 ;
        RECT 844.620 4711.610 846.220 4723.440 ;
        RECT 862.120 4716.520 863.720 4723.120 ;
        RECT 879.620 4711.610 881.220 4723.440 ;
        RECT 897.120 4716.520 898.720 4723.120 ;
        RECT 1084.620 4711.610 1086.220 4723.440 ;
        RECT 1102.120 4716.520 1103.720 4723.120 ;
        RECT 1119.620 4711.610 1121.220 4723.440 ;
        RECT 1137.120 4716.520 1138.720 4723.120 ;
        RECT 1154.620 4711.610 1156.220 4723.440 ;
        RECT 1172.120 4716.520 1173.720 4723.120 ;
        RECT 1359.620 4711.610 1361.220 4723.440 ;
        RECT 1377.120 4716.520 1378.720 4723.120 ;
        RECT 1394.620 4711.610 1396.220 4723.440 ;
        RECT 1412.120 4716.520 1413.720 4723.120 ;
        RECT 1429.620 4711.610 1431.220 4723.440 ;
        RECT 1447.120 4716.520 1448.720 4723.120 ;
        RECT 1634.620 4711.610 1636.220 4723.440 ;
        RECT 1652.120 4716.520 1653.720 4723.120 ;
        RECT 1669.620 4711.610 1671.220 4723.440 ;
        RECT 1687.120 4716.520 1688.720 4723.120 ;
        RECT 1704.620 4711.610 1706.220 4723.440 ;
        RECT 1722.120 4716.520 1723.720 4723.120 ;
        RECT 2184.620 4711.610 2186.220 4723.440 ;
        RECT 2202.120 4716.520 2203.720 4723.120 ;
        RECT 2219.620 4711.610 2221.220 4723.440 ;
        RECT 2237.120 4716.520 2238.720 4723.120 ;
        RECT 2254.620 4711.610 2256.220 4723.440 ;
        RECT 2272.120 4716.520 2273.720 4723.120 ;
        RECT 2459.620 4711.610 2461.220 4723.440 ;
        RECT 2477.120 4716.520 2478.720 4723.120 ;
        RECT 2494.620 4711.610 2496.220 4723.440 ;
        RECT 2512.120 4716.520 2513.720 4723.120 ;
        RECT 2529.620 4711.610 2531.220 4723.440 ;
        RECT 2547.120 4716.520 2548.720 4723.120 ;
        RECT 2734.620 4711.610 2736.220 4723.440 ;
        RECT 2752.120 4716.520 2753.720 4723.120 ;
        RECT 2769.620 4711.610 2771.220 4723.440 ;
        RECT 2787.120 4716.520 2788.720 4723.120 ;
        RECT 2804.620 4711.610 2806.220 4723.440 ;
        RECT 2822.120 4716.520 2823.720 4723.120 ;
        RECT 3284.620 4711.610 3286.220 4723.440 ;
        RECT 3302.120 4716.520 3303.720 4723.120 ;
        RECT 3319.620 4711.610 3321.220 4723.440 ;
        RECT 3337.120 4716.520 3338.720 4723.120 ;
        RECT 3354.620 4711.610 3356.220 4723.440 ;
        RECT 3372.120 4716.520 3373.720 4723.120 ;
        RECT 388.390 4706.610 3501.610 4711.610 ;
        RECT 395.390 4699.610 3494.610 4704.610 ;
        RECT 376.880 4647.120 400.390 4648.720 ;
        RECT 376.560 4629.620 393.390 4631.220 ;
        RECT 3496.610 4628.780 3513.440 4630.380 ;
        RECT 376.880 4612.120 400.390 4613.720 ;
        RECT 3489.610 4611.280 3513.120 4612.880 ;
        RECT 376.560 4594.620 393.390 4596.220 ;
        RECT 3496.610 4593.780 3513.440 4595.380 ;
        RECT 376.880 4577.120 400.390 4578.720 ;
        RECT 3489.610 4576.280 3513.120 4577.880 ;
        RECT 388.390 4570.050 422.580 4573.150 ;
        RECT 3437.060 4570.050 3501.610 4573.150 ;
        RECT 376.560 4559.620 393.390 4561.220 ;
        RECT 3496.610 4558.780 3513.440 4560.380 ;
        RECT 3489.610 4541.280 3513.120 4542.880 ;
        RECT 395.390 4480.050 417.780 4483.150 ;
        RECT 3441.860 4480.050 3494.610 4483.150 ;
        RECT 3496.610 4461.450 3505.425 4462.450 ;
        RECT 3507.825 4460.450 3509.425 4462.450 ;
        RECT 3489.610 4459.450 3509.425 4460.450 ;
        RECT 350.000 4414.140 393.390 4423.640 ;
        RECT 350.000 4400.990 393.390 4411.240 ;
        RECT 3496.610 4409.140 3540.000 4418.640 ;
        RECT 350.000 4389.140 393.390 4399.390 ;
        RECT 3496.610 4395.990 3540.000 4406.240 ;
        RECT 350.000 4375.610 393.390 4385.860 ;
        RECT 3496.610 4384.140 3540.000 4394.390 ;
        RECT 350.000 4363.760 393.390 4374.010 ;
        RECT 3496.610 4370.610 3540.000 4380.860 ;
        RECT 350.000 4351.360 393.390 4360.860 ;
        RECT 3496.610 4358.760 3540.000 4369.010 ;
        RECT 3496.610 4346.360 3540.000 4355.860 ;
        RECT 395.390 4300.050 417.780 4303.150 ;
        RECT 3441.860 4300.050 3494.610 4303.150 ;
        RECT 350.000 4213.150 393.390 4218.640 ;
        RECT 350.000 4210.050 422.580 4213.150 ;
        RECT 3437.060 4210.050 3501.610 4213.150 ;
        RECT 350.000 4209.140 393.390 4210.050 ;
        RECT 350.000 4195.990 393.390 4206.240 ;
        RECT 3496.610 4198.780 3513.440 4200.380 ;
        RECT 350.000 4184.140 393.390 4194.390 ;
        RECT 3489.610 4181.280 3513.120 4182.880 ;
        RECT 350.000 4170.610 393.390 4180.860 ;
        RECT 350.000 4158.760 393.390 4169.010 ;
        RECT 3496.610 4163.780 3513.440 4165.380 ;
        RECT 350.000 4146.360 393.390 4155.860 ;
        RECT 3489.610 4146.280 3513.120 4147.880 ;
        RECT 3496.610 4128.780 3513.440 4130.380 ;
        RECT 395.390 4120.050 417.780 4123.150 ;
        RECT 3441.860 4120.050 3494.610 4123.150 ;
        RECT 3489.610 4111.280 3513.120 4112.880 ;
        RECT 388.390 4030.050 422.580 4033.150 ;
        RECT 3496.610 4031.450 3505.425 4032.450 ;
        RECT 3507.825 4030.450 3509.425 4032.450 ;
        RECT 3489.610 4029.450 3509.425 4030.450 ;
        RECT 350.000 4004.140 400.390 4013.640 ;
        RECT 350.000 3990.990 400.390 4001.240 ;
        RECT 350.000 3979.140 400.390 3989.390 ;
        RECT 3496.610 3979.140 3540.000 3988.640 ;
        RECT 350.000 3965.610 400.390 3975.860 ;
        RECT 3496.610 3965.990 3540.000 3976.240 ;
        RECT 350.000 3953.760 400.390 3964.010 ;
        RECT 3496.610 3954.140 3540.000 3964.390 ;
        RECT 350.000 3943.150 400.390 3950.860 ;
        RECT 350.000 3941.360 417.780 3943.150 ;
        RECT 395.390 3940.050 417.780 3941.360 ;
        RECT 3496.610 3940.610 3540.000 3950.860 ;
        RECT 3496.610 3928.760 3540.000 3939.010 ;
        RECT 3496.610 3916.360 3540.000 3925.860 ;
        RECT 380.575 3909.550 400.390 3910.550 ;
        RECT 380.575 3907.550 382.175 3909.550 ;
        RECT 384.575 3907.550 393.390 3908.550 ;
        RECT 388.390 3850.050 422.580 3853.150 ;
        RECT 3437.060 3850.050 3501.610 3853.150 ;
        RECT 376.880 3827.120 400.390 3828.720 ;
        RECT 376.560 3809.620 393.390 3811.220 ;
        RECT 376.880 3792.120 400.390 3793.720 ;
        RECT 376.560 3774.620 393.390 3776.220 ;
        RECT 3496.610 3768.780 3513.440 3770.380 ;
        RECT 395.390 3760.050 417.780 3763.150 ;
        RECT 3441.860 3760.050 3494.610 3763.150 ;
        RECT 376.880 3757.120 400.390 3758.720 ;
        RECT 3489.610 3751.280 3513.120 3752.880 ;
        RECT 376.560 3739.620 393.390 3741.220 ;
        RECT 3496.610 3733.780 3513.440 3735.380 ;
        RECT 3489.610 3716.280 3513.120 3717.880 ;
        RECT 380.575 3704.550 400.390 3705.550 ;
        RECT 380.575 3702.550 382.175 3704.550 ;
        RECT 384.575 3702.550 393.390 3703.550 ;
        RECT 3496.610 3698.780 3513.440 3700.380 ;
        RECT 3489.610 3681.280 3513.120 3682.880 ;
        RECT 388.390 3670.050 422.580 3673.150 ;
        RECT 3437.060 3670.050 3501.610 3673.150 ;
        RECT 376.880 3622.120 400.390 3623.720 ;
        RECT 376.560 3604.620 393.390 3606.220 ;
        RECT 3496.610 3601.450 3505.425 3602.450 ;
        RECT 3507.825 3600.450 3509.425 3602.450 ;
        RECT 3489.610 3599.450 3509.425 3600.450 ;
        RECT 376.880 3587.120 400.390 3588.720 ;
        RECT 395.390 3580.050 417.780 3583.150 ;
        RECT 3441.860 3580.050 3494.610 3583.150 ;
        RECT 376.560 3569.620 393.390 3571.220 ;
        RECT 3496.610 3553.780 3513.440 3555.380 ;
        RECT 376.880 3552.120 400.390 3553.720 ;
        RECT 3489.610 3536.280 3513.120 3537.880 ;
        RECT 376.560 3534.620 393.390 3536.220 ;
        RECT 3496.610 3518.780 3513.440 3520.380 ;
        RECT 3489.610 3501.280 3513.120 3502.880 ;
        RECT 380.575 3499.550 400.390 3500.550 ;
        RECT 380.575 3497.550 382.175 3499.550 ;
        RECT 384.575 3497.550 393.390 3498.550 ;
        RECT 388.390 3490.050 422.580 3493.150 ;
        RECT 3437.060 3490.050 3501.610 3493.150 ;
        RECT 3496.610 3483.780 3513.440 3485.380 ;
        RECT 3489.610 3466.280 3513.120 3467.880 ;
        RECT 376.880 3417.120 400.390 3418.720 ;
        RECT 376.560 3399.620 393.390 3401.220 ;
        RECT 395.390 3400.050 417.780 3403.150 ;
        RECT 3441.860 3400.050 3494.610 3403.150 ;
        RECT 3496.610 3386.450 3505.425 3387.450 ;
        RECT 3507.825 3385.450 3509.425 3387.450 ;
        RECT 3489.610 3384.450 3509.425 3385.450 ;
        RECT 376.880 3382.120 400.390 3383.720 ;
        RECT 376.560 3364.620 393.390 3366.220 ;
        RECT 376.880 3347.120 400.390 3348.720 ;
        RECT 3496.610 3338.780 3513.440 3340.380 ;
        RECT 376.560 3329.620 393.390 3331.220 ;
        RECT 3489.610 3321.280 3513.120 3322.880 ;
        RECT 388.390 3310.050 422.580 3313.150 ;
        RECT 3437.060 3310.050 3501.610 3313.150 ;
        RECT 3496.610 3303.780 3513.440 3305.380 ;
        RECT 380.575 3294.550 400.390 3295.550 ;
        RECT 380.575 3292.550 382.175 3294.550 ;
        RECT 384.575 3292.550 393.390 3293.550 ;
        RECT 3489.610 3286.280 3513.120 3287.880 ;
        RECT 3496.610 3268.780 3513.440 3270.380 ;
        RECT 3489.610 3251.280 3513.120 3252.880 ;
        RECT 395.390 3220.050 417.780 3223.150 ;
        RECT 3441.860 3220.050 3494.610 3223.150 ;
        RECT 376.880 3212.120 400.390 3213.720 ;
        RECT 376.560 3194.620 393.390 3196.220 ;
        RECT 376.880 3177.120 400.390 3178.720 ;
        RECT 3496.610 3171.450 3505.425 3172.450 ;
        RECT 3507.825 3170.450 3509.425 3172.450 ;
        RECT 3489.610 3169.450 3509.425 3170.450 ;
        RECT 376.560 3159.620 393.390 3161.220 ;
        RECT 376.880 3142.120 400.390 3143.720 ;
        RECT 388.390 3130.050 422.580 3133.150 ;
        RECT 3437.060 3130.050 3501.610 3133.150 ;
        RECT 376.560 3124.620 393.390 3126.220 ;
        RECT 3496.610 3123.780 3513.440 3125.380 ;
        RECT 3489.610 3106.280 3513.120 3107.880 ;
        RECT 380.575 3089.550 400.390 3090.550 ;
        RECT 380.575 3087.550 382.175 3089.550 ;
        RECT 3496.610 3088.780 3513.440 3090.380 ;
        RECT 384.575 3087.550 393.390 3088.550 ;
        RECT 3489.610 3071.280 3513.120 3072.880 ;
        RECT 3496.610 3053.780 3513.440 3055.380 ;
        RECT 395.390 3040.050 417.780 3043.150 ;
        RECT 3441.860 3040.050 3494.610 3043.150 ;
        RECT 3489.610 3036.280 3513.120 3037.880 ;
        RECT 376.880 3007.120 400.390 3008.720 ;
        RECT 376.560 2989.620 393.390 2991.220 ;
        RECT 376.880 2972.120 400.390 2973.720 ;
        RECT 3496.610 2956.450 3505.425 2957.450 ;
        RECT 376.560 2954.620 393.390 2956.220 ;
        RECT 3507.825 2955.450 3509.425 2957.450 ;
        RECT 3489.610 2954.450 3509.425 2955.450 ;
        RECT 388.390 2950.050 422.580 2953.150 ;
        RECT 3437.060 2950.050 3501.610 2953.150 ;
        RECT 376.880 2937.120 400.390 2938.720 ;
        RECT 376.560 2919.620 393.390 2921.220 ;
        RECT 3496.610 2908.780 3513.440 2910.380 ;
        RECT 3489.610 2891.280 3513.120 2892.880 ;
        RECT 380.575 2884.550 400.390 2885.550 ;
        RECT 380.575 2882.550 382.175 2884.550 ;
        RECT 384.575 2882.550 393.390 2883.550 ;
        RECT 3496.610 2873.780 3513.440 2875.380 ;
        RECT 395.390 2860.050 417.780 2863.150 ;
        RECT 3441.860 2860.050 3494.610 2863.150 ;
        RECT 3489.610 2856.280 3513.120 2857.880 ;
        RECT 3496.610 2838.780 3513.440 2840.380 ;
        RECT 3489.610 2821.280 3513.120 2822.880 ;
        RECT 376.880 2802.120 400.390 2803.720 ;
        RECT 376.560 2784.620 393.390 2786.220 ;
        RECT 388.390 2770.050 422.580 2773.150 ;
        RECT 3437.060 2770.050 3501.610 2773.150 ;
        RECT 376.880 2767.120 400.390 2768.720 ;
        RECT 376.560 2749.620 393.390 2751.220 ;
        RECT 3496.610 2741.450 3505.425 2742.450 ;
        RECT 3507.825 2740.450 3509.425 2742.450 ;
        RECT 3489.610 2739.450 3509.425 2740.450 ;
        RECT 376.880 2732.120 400.390 2733.720 ;
        RECT 376.560 2714.620 393.390 2716.220 ;
        RECT 3496.610 2693.780 3513.440 2695.380 ;
        RECT 395.390 2680.550 417.780 2683.150 ;
        RECT 380.575 2680.050 417.780 2680.550 ;
        RECT 3441.860 2680.050 3494.610 2683.150 ;
        RECT 380.575 2679.550 400.390 2680.050 ;
        RECT 380.575 2677.550 382.175 2679.550 ;
        RECT 384.575 2677.550 393.390 2678.550 ;
        RECT 3489.610 2676.280 3513.120 2677.880 ;
        RECT 3496.610 2658.780 3513.440 2660.380 ;
        RECT 3489.610 2641.280 3513.120 2642.880 ;
        RECT 3496.610 2623.780 3513.440 2625.380 ;
        RECT 3489.610 2606.280 3513.120 2607.880 ;
        RECT 376.880 2597.120 400.390 2598.720 ;
        RECT 388.390 2590.050 422.580 2593.150 ;
        RECT 3437.060 2590.050 3501.610 2593.150 ;
        RECT 376.560 2579.620 393.390 2581.220 ;
        RECT 376.880 2562.120 400.390 2563.720 ;
        RECT 376.560 2544.620 393.390 2546.220 ;
        RECT 376.880 2527.120 400.390 2528.720 ;
        RECT 3496.610 2526.450 3505.425 2527.450 ;
        RECT 3507.825 2525.450 3509.425 2527.450 ;
        RECT 3489.610 2524.450 3509.425 2525.450 ;
        RECT 376.560 2509.620 393.390 2511.220 ;
        RECT 395.390 2500.050 417.780 2503.150 ;
        RECT 3441.860 2500.050 3494.610 2503.150 ;
        RECT 3496.610 2474.140 3540.000 2483.640 ;
        RECT 3496.610 2460.990 3540.000 2471.240 ;
        RECT 3496.610 2449.140 3540.000 2459.390 ;
        RECT 3496.610 2435.610 3540.000 2445.860 ;
        RECT 3496.610 2423.760 3540.000 2434.010 ;
        RECT 3496.610 2413.150 3540.000 2420.860 ;
        RECT 388.390 2410.050 422.580 2413.150 ;
        RECT 3437.060 2411.360 3540.000 2413.150 ;
        RECT 3437.060 2410.050 3501.610 2411.360 ;
        RECT 350.000 2364.140 393.390 2373.640 ;
        RECT 350.000 2350.990 393.390 2361.240 ;
        RECT 350.000 2339.140 393.390 2349.390 ;
        RECT 350.000 2325.610 393.390 2335.860 ;
        RECT 350.000 2313.760 393.390 2324.010 ;
        RECT 3441.860 2320.050 3494.610 2323.150 ;
        RECT 350.000 2301.360 393.390 2310.860 ;
        RECT 3489.610 2259.140 3540.000 2268.640 ;
        RECT 3489.610 2245.990 3540.000 2256.240 ;
        RECT 3489.610 2234.140 3540.000 2244.390 ;
        RECT 388.390 2230.050 422.580 2233.150 ;
        RECT 3489.610 2220.610 3540.000 2230.860 ;
        RECT 3489.610 2208.760 3540.000 2219.010 ;
        RECT 3489.610 2196.360 3540.000 2205.860 ;
        RECT 350.000 2159.140 400.390 2168.640 ;
        RECT 350.000 2145.990 400.390 2156.240 ;
        RECT 350.000 2134.140 400.390 2144.390 ;
        RECT 3441.860 2140.050 3494.610 2143.150 ;
        RECT 350.000 2120.610 400.390 2130.860 ;
        RECT 350.000 2108.760 400.390 2119.010 ;
        RECT 350.000 2096.360 400.390 2105.860 ;
        RECT 380.575 2064.550 400.390 2065.550 ;
        RECT 380.575 2062.550 382.175 2064.550 ;
        RECT 384.575 2062.550 393.390 2063.550 ;
        RECT 388.390 2050.050 422.580 2053.150 ;
        RECT 3489.610 2044.140 3540.000 2053.640 ;
        RECT 3489.610 2030.990 3540.000 2041.240 ;
        RECT 3489.610 2019.140 3540.000 2029.390 ;
        RECT 3489.610 2005.610 3540.000 2015.860 ;
        RECT 3489.610 1993.760 3540.000 2004.010 ;
        RECT 376.880 1982.120 400.390 1983.720 ;
        RECT 3489.610 1981.360 3540.000 1990.860 ;
        RECT 376.560 1964.620 393.390 1966.220 ;
        RECT 395.390 1960.050 417.780 1963.150 ;
        RECT 3441.860 1960.050 3494.610 1963.150 ;
        RECT 376.880 1947.120 400.390 1948.720 ;
        RECT 376.560 1929.620 393.390 1931.220 ;
        RECT 376.880 1912.120 400.390 1913.720 ;
        RECT 376.560 1894.620 393.390 1896.220 ;
        RECT 388.390 1870.050 422.580 1873.150 ;
        RECT 3437.060 1870.050 3501.610 1873.150 ;
        RECT 380.575 1859.550 400.390 1860.550 ;
        RECT 380.575 1857.550 382.175 1859.550 ;
        RECT 384.575 1857.550 393.390 1858.550 ;
        RECT 3496.610 1833.780 3513.440 1835.380 ;
        RECT 3489.610 1816.280 3513.120 1817.880 ;
        RECT 3496.610 1798.780 3513.440 1800.380 ;
        RECT 395.390 1780.050 417.780 1783.150 ;
        RECT 3441.860 1782.880 3494.610 1783.150 ;
        RECT 3441.860 1781.280 3513.120 1782.880 ;
        RECT 3441.860 1780.050 3494.610 1781.280 ;
        RECT 376.880 1777.120 400.390 1778.720 ;
        RECT 3496.610 1763.780 3513.440 1765.380 ;
        RECT 376.560 1759.620 393.390 1761.220 ;
        RECT 3489.610 1746.280 3513.120 1747.880 ;
        RECT 376.880 1742.120 400.390 1743.720 ;
        RECT 376.560 1724.620 393.390 1726.220 ;
        RECT 376.880 1707.120 400.390 1708.720 ;
        RECT 388.390 1691.220 422.580 1693.150 ;
        RECT 376.560 1690.050 422.580 1691.220 ;
        RECT 3437.060 1690.050 3501.610 1693.150 ;
        RECT 376.560 1689.620 393.390 1690.050 ;
        RECT 3496.610 1666.450 3505.425 1667.450 ;
        RECT 3507.825 1665.450 3509.425 1667.450 ;
        RECT 3489.610 1664.450 3509.425 1665.450 ;
        RECT 380.575 1654.550 3494.610 1655.550 ;
        RECT 380.575 1652.550 382.175 1654.550 ;
        RECT 384.575 1652.550 393.390 1653.550 ;
        RECT 395.390 1650.550 3494.610 1654.550 ;
        RECT 388.390 1643.550 3501.610 1648.550 ;
        RECT 3496.610 1618.780 3513.440 1620.380 ;
        RECT 3489.610 1601.280 3513.120 1602.880 ;
        RECT 785.440 1591.185 808.420 1592.785 ;
        RECT 1891.420 1591.185 1914.400 1592.785 ;
        RECT 790.540 1587.690 808.420 1589.290 ;
        RECT 1891.420 1587.690 1909.300 1589.290 ;
        RECT 785.440 1584.195 808.420 1585.795 ;
        RECT 1891.420 1584.195 1914.400 1585.795 ;
        RECT 3496.610 1583.780 3513.440 1585.380 ;
        RECT 790.540 1580.700 808.420 1582.300 ;
        RECT 1891.420 1580.700 1909.300 1582.300 ;
        RECT 785.440 1577.205 808.420 1578.805 ;
        RECT 1891.420 1577.205 1914.400 1578.805 ;
        RECT 376.880 1572.120 400.390 1573.720 ;
        RECT 790.540 1573.710 808.420 1575.310 ;
        RECT 1891.420 1573.710 1909.300 1575.310 ;
        RECT 785.440 1570.215 808.420 1571.815 ;
        RECT 1891.420 1570.215 1914.400 1571.815 ;
        RECT 3489.610 1566.280 3513.120 1567.880 ;
        RECT 376.560 1554.620 393.390 1556.220 ;
        RECT 3496.610 1548.780 3513.440 1550.380 ;
        RECT 376.880 1537.120 400.390 1538.720 ;
        RECT 395.390 1532.880 3494.610 1536.280 ;
        RECT 395.390 1531.280 3513.120 1532.880 ;
        RECT 388.390 1524.280 3501.610 1529.280 ;
        RECT 376.560 1519.620 393.390 1521.220 ;
        RECT 376.880 1502.120 400.390 1503.720 ;
        RECT 376.560 1484.620 393.390 1486.220 ;
        RECT 3496.610 1451.450 3505.425 1452.450 ;
        RECT 380.575 1449.550 400.390 1450.550 ;
        RECT 3507.825 1450.450 3509.425 1452.450 ;
        RECT 380.575 1447.550 382.175 1449.550 ;
        RECT 3489.610 1449.450 3509.425 1450.450 ;
        RECT 384.575 1447.550 393.390 1448.550 ;
        RECT 3330.660 1418.735 3494.610 1420.335 ;
        RECT 395.390 1412.210 2959.200 1417.210 ;
        RECT 388.390 1405.210 2966.200 1410.210 ;
        RECT 3496.610 1403.780 3513.440 1405.380 ;
        RECT 3489.610 1386.280 3513.120 1387.880 ;
        RECT 3496.610 1368.780 3513.440 1370.380 ;
        RECT 376.880 1367.120 400.390 1368.720 ;
        RECT 3489.610 1351.280 3513.120 1352.880 ;
        RECT 376.560 1349.620 393.390 1351.220 ;
        RECT 388.390 1340.610 449.600 1342.210 ;
        RECT 2800.160 1340.610 2966.200 1342.210 ;
        RECT 3330.660 1342.145 3501.610 1343.745 ;
        RECT 3496.610 1333.780 3513.440 1335.380 ;
        RECT 376.880 1332.120 400.390 1333.720 ;
        RECT 3489.610 1316.280 3513.120 1317.880 ;
        RECT 376.560 1314.620 393.390 1316.220 ;
        RECT 376.880 1297.120 400.390 1298.720 ;
        RECT 376.560 1279.620 393.390 1281.220 ;
        RECT 395.390 1275.610 449.600 1277.210 ;
        RECT 2800.160 1275.610 2959.200 1277.210 ;
        RECT 3330.660 1265.555 3494.610 1267.155 ;
        RECT 380.575 1244.550 400.390 1245.550 ;
        RECT 380.575 1242.550 382.175 1244.550 ;
        RECT 384.575 1242.550 393.390 1243.550 ;
        RECT 3496.610 1236.450 3505.425 1237.450 ;
        RECT 3507.825 1235.450 3509.425 1237.450 ;
        RECT 3489.610 1234.450 3509.425 1235.450 ;
        RECT 388.390 1210.610 449.600 1212.210 ;
        RECT 2800.160 1210.610 2966.200 1212.210 ;
        RECT 3496.610 1188.780 3513.440 1190.380 ;
        RECT 3489.610 1171.280 3513.120 1172.880 ;
        RECT 376.880 1162.120 400.390 1163.720 ;
        RECT 3496.610 1153.780 3513.440 1155.380 ;
        RECT 376.560 1144.620 393.390 1146.220 ;
        RECT 395.390 1145.610 449.600 1147.210 ;
        RECT 2800.160 1145.610 2959.200 1147.210 ;
        RECT 3489.610 1136.280 3513.120 1137.880 ;
        RECT 376.880 1127.120 400.390 1128.720 ;
        RECT 3496.610 1118.780 3513.440 1120.380 ;
        RECT 3330.660 1112.375 3494.610 1113.975 ;
        RECT 376.560 1109.620 393.390 1111.220 ;
        RECT 3489.610 1101.280 3513.120 1102.880 ;
        RECT 376.880 1092.120 400.390 1093.720 ;
        RECT 388.390 1080.610 449.600 1082.210 ;
        RECT 2800.160 1080.610 2966.200 1082.210 ;
        RECT 376.560 1074.620 393.390 1076.220 ;
        RECT 380.575 1039.550 400.390 1040.550 ;
        RECT 380.575 1037.550 382.175 1039.550 ;
        RECT 384.575 1037.550 393.390 1038.550 ;
        RECT 3330.660 1035.785 3501.610 1037.385 ;
        RECT 3496.610 1021.450 3505.425 1022.450 ;
        RECT 3507.825 1020.450 3509.425 1022.450 ;
        RECT 3489.610 1019.450 3509.425 1020.450 ;
        RECT 395.390 1015.610 449.600 1017.210 ;
        RECT 2800.160 1015.610 2959.200 1017.210 ;
        RECT 3496.610 973.780 3513.440 975.380 ;
        RECT 3330.660 959.195 3494.610 960.795 ;
        RECT 376.880 957.120 400.390 958.720 ;
        RECT 3489.610 956.280 3513.120 957.880 ;
        RECT 388.390 950.610 449.600 952.210 ;
        RECT 2800.160 950.610 2966.200 952.210 ;
        RECT 376.560 939.620 393.390 941.220 ;
        RECT 3496.610 938.780 3513.440 940.380 ;
        RECT 376.880 922.120 400.390 923.720 ;
        RECT 3489.610 921.280 3513.120 922.880 ;
        RECT 376.560 904.620 393.390 906.220 ;
        RECT 3496.610 903.780 3513.440 905.380 ;
        RECT 376.880 887.210 400.390 888.720 ;
        RECT 376.880 887.120 449.600 887.210 ;
        RECT 395.390 885.610 449.600 887.120 ;
        RECT 2800.160 885.610 2959.200 887.210 ;
        RECT 3489.610 886.280 3513.120 887.880 ;
        RECT 3330.660 882.605 3501.610 884.205 ;
        RECT 376.560 869.620 393.390 871.220 ;
        RECT 388.390 820.610 449.600 822.210 ;
        RECT 2800.160 820.610 2966.200 822.210 ;
        RECT 3330.660 806.015 3494.610 807.615 ;
        RECT 3496.610 806.450 3505.425 807.450 ;
        RECT 3507.825 805.450 3509.425 807.450 ;
        RECT 3489.610 804.450 3509.425 805.450 ;
        RECT 3496.610 758.780 3513.440 760.380 ;
        RECT 395.390 755.610 449.600 757.210 ;
        RECT 2800.160 755.610 2959.200 757.210 ;
        RECT 3489.610 741.280 3513.120 742.880 ;
        RECT 350.000 724.140 393.390 733.640 ;
        RECT 3330.660 729.425 3501.610 731.025 ;
        RECT 3496.610 723.780 3513.440 725.380 ;
        RECT 350.000 710.990 393.390 721.240 ;
        RECT 350.000 699.140 393.390 709.390 ;
        RECT 3489.610 706.280 3513.120 707.880 ;
        RECT 350.000 685.610 393.390 695.860 ;
        RECT 2800.160 690.610 2966.200 692.210 ;
        RECT 3496.610 688.780 3513.440 690.380 ;
        RECT 350.000 673.760 393.390 684.010 ;
        RECT 3489.610 671.280 3513.120 672.880 ;
        RECT 350.000 661.360 393.390 670.860 ;
        RECT 3350.805 668.125 3501.610 669.725 ;
        RECT 3350.805 664.125 3494.610 665.725 ;
        RECT 395.390 625.610 449.600 627.210 ;
        RECT 2800.160 625.610 2959.200 627.210 ;
        RECT 2961.200 607.510 3103.110 609.110 ;
        RECT 2954.200 599.740 3103.110 601.340 ;
        RECT 2961.200 591.970 3103.110 593.570 ;
        RECT 3496.610 591.450 3505.425 592.450 ;
        RECT 3507.825 590.450 3509.425 592.450 ;
        RECT 3489.610 589.450 3509.425 590.450 ;
        RECT 2954.200 584.200 3103.110 585.800 ;
        RECT 2961.200 576.430 3103.110 578.030 ;
        RECT 2954.200 568.660 3103.110 570.260 ;
        RECT 2961.200 562.210 3103.110 562.490 ;
        RECT 388.390 560.610 449.600 562.210 ;
        RECT 2800.160 560.890 3103.110 562.210 ;
        RECT 2800.160 560.610 2966.200 560.890 ;
        RECT 3496.610 543.780 3513.440 545.380 ;
        RECT 350.000 519.140 393.390 528.640 ;
        RECT 3489.610 526.280 3513.120 527.880 ;
        RECT 350.000 505.990 393.390 516.240 ;
        RECT 3496.610 508.780 3513.440 510.380 ;
        RECT 350.000 494.140 393.390 504.390 ;
        RECT 3340.300 497.265 3340.580 497.545 ;
        RECT 3340.920 497.265 3341.200 497.545 ;
        RECT 3341.540 497.265 3341.820 497.545 ;
        RECT 3342.160 497.265 3342.440 497.545 ;
        RECT 3342.780 497.265 3343.060 497.545 ;
        RECT 3343.400 497.265 3343.680 497.545 ;
        RECT 3350.450 497.265 3350.730 497.545 ;
        RECT 3351.070 497.265 3351.350 497.545 ;
        RECT 3351.690 497.265 3351.970 497.545 ;
        RECT 3352.310 497.265 3352.590 497.545 ;
        RECT 3352.930 497.265 3353.210 497.545 ;
        RECT 3353.550 497.265 3353.830 497.545 ;
        RECT 395.390 495.610 449.600 497.210 ;
        RECT 2800.160 495.610 2959.200 497.210 ;
        RECT 3340.300 496.645 3340.580 496.925 ;
        RECT 3340.920 496.645 3341.200 496.925 ;
        RECT 3341.540 496.645 3341.820 496.925 ;
        RECT 3342.160 496.645 3342.440 496.925 ;
        RECT 3342.780 496.645 3343.060 496.925 ;
        RECT 3343.400 496.645 3343.680 496.925 ;
        RECT 3350.450 496.645 3350.730 496.925 ;
        RECT 3351.070 496.645 3351.350 496.925 ;
        RECT 3351.690 496.645 3351.970 496.925 ;
        RECT 3352.310 496.645 3352.590 496.925 ;
        RECT 3352.930 496.645 3353.210 496.925 ;
        RECT 3353.550 496.645 3353.830 496.925 ;
        RECT 3340.300 496.025 3340.580 496.305 ;
        RECT 3340.920 496.025 3341.200 496.305 ;
        RECT 3341.540 496.025 3341.820 496.305 ;
        RECT 3342.160 496.025 3342.440 496.305 ;
        RECT 3342.780 496.025 3343.060 496.305 ;
        RECT 3343.400 496.025 3343.680 496.305 ;
        RECT 3350.450 496.025 3350.730 496.305 ;
        RECT 3351.070 496.025 3351.350 496.305 ;
        RECT 3351.690 496.025 3351.970 496.305 ;
        RECT 3352.310 496.025 3352.590 496.305 ;
        RECT 3352.930 496.025 3353.210 496.305 ;
        RECT 3353.550 496.025 3353.830 496.305 ;
        RECT 3340.300 495.405 3340.580 495.685 ;
        RECT 3340.920 495.405 3341.200 495.685 ;
        RECT 3341.540 495.405 3341.820 495.685 ;
        RECT 3342.160 495.405 3342.440 495.685 ;
        RECT 3342.780 495.405 3343.060 495.685 ;
        RECT 3343.400 495.405 3343.680 495.685 ;
        RECT 3350.450 495.405 3350.730 495.685 ;
        RECT 3351.070 495.405 3351.350 495.685 ;
        RECT 3351.690 495.405 3351.970 495.685 ;
        RECT 3352.310 495.405 3352.590 495.685 ;
        RECT 3352.930 495.405 3353.210 495.685 ;
        RECT 3353.550 495.405 3353.830 495.685 ;
        RECT 3340.300 494.785 3340.580 495.065 ;
        RECT 3340.920 494.785 3341.200 495.065 ;
        RECT 3341.540 494.785 3341.820 495.065 ;
        RECT 3342.160 494.785 3342.440 495.065 ;
        RECT 3342.780 494.785 3343.060 495.065 ;
        RECT 3343.400 494.785 3343.680 495.065 ;
        RECT 3350.450 494.785 3350.730 495.065 ;
        RECT 3351.070 494.785 3351.350 495.065 ;
        RECT 3351.690 494.785 3351.970 495.065 ;
        RECT 3352.310 494.785 3352.590 495.065 ;
        RECT 3352.930 494.785 3353.210 495.065 ;
        RECT 3353.550 494.785 3353.830 495.065 ;
        RECT 3340.300 494.165 3340.580 494.445 ;
        RECT 3340.920 494.165 3341.200 494.445 ;
        RECT 3341.540 494.165 3341.820 494.445 ;
        RECT 3342.160 494.165 3342.440 494.445 ;
        RECT 3342.780 494.165 3343.060 494.445 ;
        RECT 3343.400 494.165 3343.680 494.445 ;
        RECT 3350.450 494.165 3350.730 494.445 ;
        RECT 3351.070 494.165 3351.350 494.445 ;
        RECT 3351.690 494.165 3351.970 494.445 ;
        RECT 3352.310 494.165 3352.590 494.445 ;
        RECT 3352.930 494.165 3353.210 494.445 ;
        RECT 3353.550 494.165 3353.830 494.445 ;
        RECT 3340.300 493.545 3340.580 493.825 ;
        RECT 3340.920 493.545 3341.200 493.825 ;
        RECT 3341.540 493.545 3341.820 493.825 ;
        RECT 3342.160 493.545 3342.440 493.825 ;
        RECT 3342.780 493.545 3343.060 493.825 ;
        RECT 3343.400 493.545 3343.680 493.825 ;
        RECT 3350.450 493.545 3350.730 493.825 ;
        RECT 3351.070 493.545 3351.350 493.825 ;
        RECT 3351.690 493.545 3351.970 493.825 ;
        RECT 3352.310 493.545 3352.590 493.825 ;
        RECT 3352.930 493.545 3353.210 493.825 ;
        RECT 3353.550 493.545 3353.830 493.825 ;
        RECT 3489.610 491.280 3513.120 492.880 ;
        RECT 350.000 480.610 393.390 490.860 ;
        RECT 350.000 468.760 393.390 479.010 ;
        RECT 3496.610 473.780 3513.440 475.380 ;
        RECT 350.000 456.360 393.390 465.860 ;
        RECT 3489.610 456.280 3513.120 457.880 ;
        RECT 388.390 430.610 449.600 432.210 ;
        RECT 2800.160 430.610 2966.200 432.210 ;
        RECT 395.390 395.390 3494.610 400.390 ;
        RECT 388.390 388.390 3501.610 393.390 ;
        RECT 3496.610 376.450 3505.425 377.450 ;
        RECT 3507.825 375.450 3509.425 377.450 ;
        RECT 3489.610 374.450 3509.425 375.450 ;
  END
END caravel_gf180_pdn
END LIBRARY

