VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO copyright_block
  CLASS BLOCK ;
  FOREIGN copyright_block ;
  ORIGIN 0.00 0.00 ;
  SIZE 93.495 BY 44.990 ;
  OBS
      LAYER Metal5 ;
        RECT 0.490 11.125 3.010 11.485 ;
        RECT 0.130 10.765 3.010 11.125 ;
        RECT -0.230 10.045 3.010 10.765 ;
        RECT -0.230 5.365 0.850 10.045 ;
        RECT 4.030 8.920 6.910 9.280 ;
        RECT 8.335 8.920 10.855 9.280 ;
        RECT 12.685 8.920 15.565 9.280 ;
        RECT 4.030 8.200 7.270 8.920 ;
        RECT 6.190 7.120 7.270 8.200 ;
        RECT 4.390 6.760 7.270 7.120 ;
        RECT 4.030 6.040 7.270 6.760 ;
        RECT -0.230 4.645 3.010 5.365 ;
        RECT 0.130 4.285 3.010 4.645 ;
        RECT 0.490 3.925 3.010 4.285 ;
        RECT 4.030 4.960 5.110 6.040 ;
        RECT 6.190 4.960 7.270 6.040 ;
        RECT 4.030 4.240 7.270 4.960 ;
        RECT 4.390 3.880 7.270 4.240 ;
        RECT 8.335 8.560 11.215 8.920 ;
        RECT 8.335 7.840 11.575 8.560 ;
        RECT 12.685 8.200 15.925 8.920 ;
        RECT 8.335 3.880 9.415 7.840 ;
        RECT 10.495 7.120 11.575 7.840 ;
        RECT 14.845 7.120 15.925 8.200 ;
        RECT 13.045 6.760 15.925 7.120 ;
        RECT 12.685 6.040 15.925 6.760 ;
        RECT 12.685 4.960 13.765 6.040 ;
        RECT 14.845 4.960 15.925 6.040 ;
        RECT 17.225 6.040 18.305 9.280 ;
        RECT 19.385 6.040 20.465 9.280 ;
        RECT 21.745 9.010 24.265 9.370 ;
        RECT 17.225 4.960 20.465 6.040 ;
        RECT 21.385 8.290 24.625 9.010 ;
        RECT 21.385 7.210 22.465 8.290 ;
        RECT 23.545 7.210 24.625 8.290 ;
        RECT 21.385 6.490 24.625 7.210 ;
        RECT 21.385 6.130 24.265 6.490 ;
        RECT 21.385 5.050 22.465 6.130 ;
        RECT 12.685 4.240 15.925 4.960 ;
        RECT 17.585 4.600 20.105 4.960 ;
        RECT 13.045 3.880 15.925 4.240 ;
        RECT 18.305 3.880 19.385 4.600 ;
        RECT 21.385 4.330 24.625 5.050 ;
        RECT 21.745 3.970 24.625 4.330 ;
        RECT 25.690 3.880 26.770 11.440 ;
        RECT 30.855 11.170 32.655 11.530 ;
        RECT 30.495 10.810 33.015 11.170 ;
        RECT 30.135 10.090 33.375 10.810 ;
        RECT 30.135 5.410 31.215 10.090 ;
        RECT 32.295 9.370 33.375 10.090 ;
        RECT 34.535 10.450 37.775 11.530 ;
        RECT 41.420 11.200 42.860 11.560 ;
        RECT 41.060 10.840 42.860 11.200 ;
        RECT 34.535 8.290 35.615 10.450 ;
        RECT 40.700 10.120 42.860 10.840 ;
        RECT 48.200 11.110 49.640 11.470 ;
        RECT 48.200 10.750 50.000 11.110 ;
        RECT 32.295 5.410 33.375 8.290 ;
        RECT 30.135 4.690 33.375 5.410 ;
        RECT 30.495 4.330 33.375 4.690 ;
        RECT 30.855 3.970 33.375 4.330 ;
        RECT 34.535 7.210 36.695 8.290 ;
        RECT 34.535 3.970 35.615 7.210 ;
        RECT 40.700 5.440 41.780 10.120 ;
        RECT 44.620 9.890 46.420 10.250 ;
        RECT 48.200 10.030 50.360 10.750 ;
        RECT 44.260 9.530 46.780 9.890 ;
        RECT 43.900 8.810 47.140 9.530 ;
        RECT 43.900 6.290 44.980 8.810 ;
        RECT 46.060 8.090 47.140 8.810 ;
        RECT 46.060 6.290 47.140 6.650 ;
        RECT 43.900 5.570 47.140 6.290 ;
        RECT 40.700 4.720 42.860 5.440 ;
        RECT 44.260 5.210 46.780 5.570 ;
        RECT 49.280 5.350 50.360 10.030 ;
        RECT 44.620 4.850 46.420 5.210 ;
        RECT 41.060 4.360 42.860 4.720 ;
        RECT 41.420 4.000 42.860 4.360 ;
        RECT 48.200 4.630 50.360 5.350 ;
        RECT 55.150 10.390 58.390 11.470 ;
        RECT 60.890 11.110 62.690 11.470 ;
        RECT 60.530 10.390 62.690 11.110 ;
        RECT 55.150 8.230 56.230 10.390 ;
        RECT 60.530 9.310 61.610 10.390 ;
        RECT 68.150 9.310 69.230 11.470 ;
        RECT 59.450 8.230 62.690 9.310 ;
        RECT 63.800 8.900 66.680 9.260 ;
        RECT 68.150 8.950 70.670 9.310 ;
        RECT 55.150 7.150 57.310 8.230 ;
        RECT 55.150 4.990 56.230 7.150 ;
        RECT 48.200 4.270 50.000 4.630 ;
        RECT 48.200 3.910 49.640 4.270 ;
        RECT 55.150 3.910 58.390 4.990 ;
        RECT 60.530 3.910 61.610 8.230 ;
        RECT 63.800 8.180 67.040 8.900 ;
        RECT 65.960 7.100 67.040 8.180 ;
        RECT 64.160 6.740 67.040 7.100 ;
        RECT 63.800 6.020 67.040 6.740 ;
        RECT 63.800 4.940 64.880 6.020 ;
        RECT 65.960 4.940 67.040 6.020 ;
        RECT 63.800 4.220 67.040 4.940 ;
        RECT 64.160 3.860 67.040 4.220 ;
        RECT 68.150 8.590 71.030 8.950 ;
        RECT 68.150 7.870 71.390 8.590 ;
        RECT 68.150 5.350 69.230 7.870 ;
        RECT 70.310 5.350 71.390 7.870 ;
        RECT 68.150 4.630 71.390 5.350 ;
        RECT 68.150 4.270 71.030 4.630 ;
        RECT 68.150 3.910 70.670 4.270 ;
        RECT 72.500 3.910 73.580 11.470 ;
        RECT 75.010 8.950 77.530 9.310 ;
        RECT 79.720 8.990 82.240 9.350 ;
        RECT 84.020 8.990 86.540 9.350 ;
        RECT 74.650 8.230 77.890 8.950 ;
        RECT 79.360 8.630 82.240 8.990 ;
        RECT 83.660 8.630 86.540 8.990 ;
        RECT 74.650 7.150 75.730 8.230 ;
        RECT 76.810 7.150 77.890 8.230 ;
        RECT 74.650 6.430 77.890 7.150 ;
        RECT 79.000 8.270 82.240 8.630 ;
        RECT 83.300 8.270 86.540 8.630 ;
        RECT 79.000 7.190 80.440 8.270 ;
        RECT 83.300 7.190 84.740 8.270 ;
        RECT 79.000 6.830 81.520 7.190 ;
        RECT 83.300 6.830 85.820 7.190 ;
        RECT 79.360 6.470 81.880 6.830 ;
        RECT 83.660 6.470 86.180 6.830 ;
        RECT 74.650 6.070 77.530 6.430 ;
        RECT 79.720 6.110 82.240 6.470 ;
        RECT 84.020 6.110 86.540 6.470 ;
        RECT 74.650 4.990 75.730 6.070 ;
        RECT 80.800 5.030 82.240 6.110 ;
        RECT 85.100 5.030 86.540 6.110 ;
        RECT 74.650 4.270 77.890 4.990 ;
        RECT 75.010 3.910 77.890 4.270 ;
        RECT 79.000 4.670 82.240 5.030 ;
        RECT 83.300 4.670 86.540 5.030 ;
        RECT 79.000 4.310 81.880 4.670 ;
        RECT 83.300 4.310 86.180 4.670 ;
        RECT 79.000 3.950 81.520 4.310 ;
        RECT 83.300 3.950 85.820 4.310 ;
        RECT 0.915 0.550 2.715 0.910 ;
        RECT 0.555 0.190 3.075 0.550 ;
        RECT 0.195 -0.530 3.435 0.190 ;
        RECT 0.195 -5.210 1.275 -0.530 ;
        RECT 2.355 -1.250 3.435 -0.530 ;
        RECT 5.115 -1.525 6.915 -1.165 ;
        RECT 4.755 -1.885 7.275 -1.525 ;
        RECT 9.370 -1.575 11.170 -1.215 ;
        RECT 2.355 -5.210 3.435 -2.330 ;
        RECT 0.195 -5.930 3.435 -5.210 ;
        RECT 4.395 -2.605 7.635 -1.885 ;
        RECT 9.010 -1.935 11.530 -1.575 ;
        RECT 13.765 -1.620 15.565 -1.260 ;
        RECT 4.395 -5.125 5.475 -2.605 ;
        RECT 6.555 -5.125 7.635 -2.605 ;
        RECT 4.395 -5.845 7.635 -5.125 ;
        RECT 8.650 -2.655 11.890 -1.935 ;
        RECT 13.405 -1.980 15.925 -1.620 ;
        RECT 8.650 -5.175 9.730 -2.655 ;
        RECT 10.810 -5.175 11.890 -2.655 ;
        RECT 0.555 -6.290 3.435 -5.930 ;
        RECT 4.755 -6.205 7.275 -5.845 ;
        RECT 8.650 -5.895 11.890 -5.175 ;
        RECT 13.045 -2.700 16.285 -1.980 ;
        RECT 13.045 -5.220 14.125 -2.700 ;
        RECT 15.205 -5.220 16.285 -2.700 ;
        RECT 0.915 -6.650 3.435 -6.290 ;
        RECT 5.115 -6.565 6.915 -6.205 ;
        RECT 9.010 -6.255 11.530 -5.895 ;
        RECT 13.045 -5.940 16.285 -5.220 ;
        RECT 9.370 -6.615 11.170 -6.255 ;
        RECT 13.405 -6.300 16.285 -5.940 ;
        RECT 13.765 -6.660 16.285 -6.300 ;
        RECT 14.845 -7.740 16.285 -6.660 ;
        RECT 17.390 -6.705 18.470 0.855 ;
        RECT 29.875 0.550 31.675 0.910 ;
        RECT 29.515 0.190 32.035 0.550 ;
        RECT 29.155 -0.530 32.395 0.190 ;
        RECT 19.950 -1.665 22.470 -1.305 ;
        RECT 19.590 -2.385 22.830 -1.665 ;
        RECT 19.590 -3.465 20.670 -2.385 ;
        RECT 21.750 -3.465 22.830 -2.385 ;
        RECT 19.590 -4.185 22.830 -3.465 ;
        RECT 23.840 -3.515 28.160 -2.435 ;
        RECT 19.590 -4.545 22.470 -4.185 ;
        RECT 19.590 -5.625 20.670 -4.545 ;
        RECT 29.155 -5.210 30.235 -0.530 ;
        RECT 31.315 -1.250 32.395 -0.530 ;
        RECT 31.315 -5.210 32.395 -2.330 ;
        RECT 19.590 -6.345 22.830 -5.625 ;
        RECT 29.155 -5.930 32.395 -5.210 ;
        RECT 29.515 -6.290 32.395 -5.930 ;
        RECT 19.950 -6.705 22.830 -6.345 ;
        RECT 29.875 -6.650 32.395 -6.290 ;
        RECT 33.455 -6.780 34.535 0.780 ;
        RECT 39.960 -1.335 41.040 0.825 ;
        RECT 36.375 -1.790 38.175 -1.430 ;
        RECT 39.960 -1.695 42.480 -1.335 ;
        RECT 44.265 -1.695 47.145 -1.335 ;
        RECT 36.015 -2.150 38.535 -1.790 ;
        RECT 39.960 -2.055 42.840 -1.695 ;
        RECT 35.655 -2.870 38.895 -2.150 ;
        RECT 35.655 -5.390 36.735 -2.870 ;
        RECT 37.815 -5.390 38.895 -2.870 ;
        RECT 35.655 -6.110 38.895 -5.390 ;
        RECT 39.960 -2.775 43.200 -2.055 ;
        RECT 44.265 -2.415 47.505 -1.695 ;
        RECT 39.960 -5.295 41.040 -2.775 ;
        RECT 42.120 -5.295 43.200 -2.775 ;
        RECT 46.425 -3.495 47.505 -2.415 ;
        RECT 44.625 -3.855 47.505 -3.495 ;
        RECT 39.960 -6.015 43.200 -5.295 ;
        RECT 44.265 -4.575 47.505 -3.855 ;
        RECT 44.265 -5.655 45.345 -4.575 ;
        RECT 46.425 -5.655 47.505 -4.575 ;
        RECT 36.015 -6.470 38.535 -6.110 ;
        RECT 39.960 -6.375 42.840 -6.015 ;
        RECT 44.265 -6.375 47.505 -5.655 ;
        RECT 36.375 -6.830 38.175 -6.470 ;
        RECT 39.960 -6.735 42.480 -6.375 ;
        RECT 44.625 -6.735 47.505 -6.375 ;
        RECT 48.615 -6.830 49.695 0.730 ;
        RECT 53.105 -0.395 56.345 0.685 ;
        RECT 53.105 -2.555 54.185 -0.395 ;
        RECT 72.435 -1.250 73.515 0.910 ;
        RECT 78.885 -1.250 81.045 0.910 ;
        RECT 58.085 -1.655 59.885 -1.295 ;
        RECT 57.725 -2.015 60.245 -1.655 ;
        RECT 53.105 -3.635 55.265 -2.555 ;
        RECT 57.365 -2.735 60.605 -2.015 ;
        RECT 53.105 -6.875 54.185 -3.635 ;
        RECT 57.365 -5.255 58.445 -2.735 ;
        RECT 59.525 -5.255 60.605 -2.735 ;
        RECT 57.365 -5.975 60.605 -5.255 ;
        RECT 61.670 -5.210 62.750 -1.250 ;
        RECT 63.830 -5.210 64.910 -1.250 ;
        RECT 61.670 -5.930 64.910 -5.210 ;
        RECT 57.725 -6.335 60.245 -5.975 ;
        RECT 62.030 -6.290 64.910 -5.930 ;
        RECT 58.085 -6.695 59.885 -6.335 ;
        RECT 62.390 -6.650 64.910 -6.290 ;
        RECT 65.880 -1.700 68.400 -1.340 ;
        RECT 70.995 -1.610 73.515 -1.250 ;
        RECT 65.880 -2.060 68.760 -1.700 ;
        RECT 70.635 -1.970 73.515 -1.610 ;
        RECT 65.880 -2.780 69.120 -2.060 ;
        RECT 65.880 -6.740 66.960 -2.780 ;
        RECT 68.040 -6.740 69.120 -2.780 ;
        RECT 70.275 -2.690 73.515 -1.970 ;
        RECT 70.275 -5.210 71.355 -2.690 ;
        RECT 72.435 -5.210 73.515 -2.690 ;
        RECT 70.275 -5.930 73.515 -5.210 ;
        RECT 70.635 -6.290 73.515 -5.930 ;
        RECT 70.995 -6.650 73.515 -6.290 ;
        RECT 74.580 -1.655 77.100 -1.295 ;
        RECT 82.520 -1.655 85.040 -1.295 ;
        RECT 87.230 -1.610 89.750 -1.250 ;
        RECT 74.580 -2.015 77.460 -1.655 ;
        RECT 74.580 -2.735 77.820 -2.015 ;
        RECT 74.580 -6.695 75.660 -2.735 ;
        RECT 76.740 -3.455 77.820 -2.735 ;
        RECT 78.885 -3.410 81.045 -2.330 ;
        RECT 79.965 -5.570 81.045 -3.410 ;
        RECT 78.885 -6.650 81.045 -5.570 ;
        RECT 82.160 -2.375 85.400 -1.655 ;
        RECT 86.870 -1.970 89.750 -1.610 ;
        RECT 82.160 -3.455 83.240 -2.375 ;
        RECT 84.320 -3.455 85.400 -2.375 ;
        RECT 82.160 -4.175 85.400 -3.455 ;
        RECT 86.510 -2.330 89.750 -1.970 ;
        RECT 86.510 -3.410 87.950 -2.330 ;
        RECT 86.510 -3.770 89.030 -3.410 ;
        RECT 86.870 -4.130 89.390 -3.770 ;
        RECT 82.160 -4.535 85.040 -4.175 ;
        RECT 87.230 -4.490 89.750 -4.130 ;
        RECT 82.160 -5.615 83.240 -4.535 ;
        RECT 88.310 -5.570 89.750 -4.490 ;
        RECT 82.160 -6.335 85.400 -5.615 ;
        RECT 82.520 -6.695 85.400 -6.335 ;
        RECT 86.510 -5.930 89.750 -5.570 ;
        RECT 86.510 -6.290 89.390 -5.930 ;
        RECT 86.510 -6.650 89.030 -6.290 ;
        RECT 13.045 -8.100 16.285 -7.740 ;
        RECT 13.045 -8.460 15.925 -8.100 ;
        RECT 13.045 -8.820 15.565 -8.460 ;
        RECT 20.920 -10.670 23.440 -10.310 ;
        RECT 20.920 -11.030 23.800 -10.670 ;
        RECT 25.225 -10.760 27.745 -10.400 ;
        RECT 20.920 -11.750 24.160 -11.030 ;
        RECT 0.445 -12.735 2.245 -12.375 ;
        RECT 4.750 -12.690 6.550 -12.330 ;
        RECT 0.085 -13.095 2.605 -12.735 ;
        RECT 4.390 -13.050 6.910 -12.690 ;
        RECT 8.740 -12.780 11.260 -12.420 ;
        RECT -0.275 -13.815 2.965 -13.095 ;
        RECT -0.275 -16.335 0.805 -13.815 ;
        RECT 1.885 -16.335 2.965 -13.815 ;
        RECT -0.275 -17.055 2.965 -16.335 ;
        RECT 4.030 -13.770 7.270 -13.050 ;
        RECT 4.030 -16.290 5.110 -13.770 ;
        RECT 6.190 -16.290 7.270 -13.770 ;
        RECT 4.030 -17.010 7.270 -16.290 ;
        RECT 8.380 -13.500 11.620 -12.780 ;
        RECT 8.380 -14.580 9.460 -13.500 ;
        RECT 10.540 -14.580 11.620 -13.500 ;
        RECT 8.380 -15.300 11.620 -14.580 ;
        RECT 12.640 -12.875 15.160 -12.515 ;
        RECT 12.640 -13.235 15.520 -12.875 ;
        RECT 12.640 -13.955 15.880 -13.235 ;
        RECT 8.380 -15.660 11.260 -15.300 ;
        RECT 8.380 -16.740 9.460 -15.660 ;
        RECT 0.085 -17.415 2.605 -17.055 ;
        RECT 4.030 -17.370 6.910 -17.010 ;
        RECT 0.445 -17.775 2.245 -17.415 ;
        RECT 4.030 -17.730 6.550 -17.370 ;
        RECT 8.380 -17.460 11.620 -16.740 ;
        RECT 4.030 -19.890 5.110 -17.730 ;
        RECT 8.740 -17.820 11.620 -17.460 ;
        RECT 12.640 -17.915 13.720 -13.955 ;
        RECT 14.800 -17.915 15.880 -13.955 ;
        RECT 20.920 -14.270 22.000 -11.750 ;
        RECT 23.080 -14.270 24.160 -11.750 ;
        RECT 20.920 -14.990 24.160 -14.270 ;
        RECT 25.225 -11.120 28.105 -10.760 ;
        RECT 25.225 -11.840 28.465 -11.120 ;
        RECT 20.920 -15.350 23.800 -14.990 ;
        RECT 20.920 -15.710 23.440 -15.350 ;
        RECT 20.920 -17.870 22.000 -15.710 ;
        RECT 25.225 -16.520 26.305 -11.840 ;
        RECT 27.385 -16.520 28.465 -11.840 ;
        RECT 25.225 -17.240 28.465 -16.520 ;
        RECT 29.525 -12.200 30.605 -10.400 ;
        RECT 31.685 -12.200 32.765 -10.400 ;
        RECT 29.525 -12.920 32.765 -12.200 ;
        RECT 29.525 -13.640 32.405 -12.920 ;
        RECT 29.525 -14.720 32.045 -13.640 ;
        RECT 29.525 -15.440 32.405 -14.720 ;
        RECT 29.525 -16.160 32.765 -15.440 ;
        RECT 25.225 -17.600 28.105 -17.240 ;
        RECT 25.225 -17.960 27.745 -17.600 ;
        RECT 29.525 -17.960 30.605 -16.160 ;
        RECT 31.685 -17.960 32.765 -16.160 ;
        RECT -0.790 -28.595 0.290 -27.875 ;
        RECT 1.370 -28.595 2.450 -22.475 ;
        RECT 20.265 -23.560 23.505 -22.480 ;
        RECT 22.425 -24.640 23.505 -23.560 ;
        RECT -0.790 -29.315 2.450 -28.595 ;
        RECT 3.515 -28.640 4.595 -24.680 ;
        RECT 5.675 -28.640 6.755 -24.680 ;
        RECT -0.430 -29.675 2.090 -29.315 ;
        RECT 3.515 -29.360 6.755 -28.640 ;
        RECT -0.070 -30.035 1.730 -29.675 ;
        RECT 3.875 -29.720 6.755 -29.360 ;
        RECT 4.235 -30.080 6.755 -29.720 ;
        RECT 7.820 -25.040 10.340 -24.680 ;
        RECT 12.485 -25.000 15.005 -24.640 ;
        RECT 7.820 -25.400 10.700 -25.040 ;
        RECT 7.820 -26.120 11.060 -25.400 ;
        RECT 7.820 -30.080 8.900 -26.120 ;
        RECT 9.980 -30.080 11.060 -26.120 ;
        RECT 12.125 -25.720 15.365 -25.000 ;
        RECT 12.125 -26.800 13.205 -25.720 ;
        RECT 14.285 -26.800 15.365 -25.720 ;
        RECT 12.125 -27.520 15.365 -26.800 ;
        RECT 20.265 -25.720 23.505 -24.640 ;
        RECT 24.615 -23.515 27.855 -22.435 ;
        RECT 12.125 -27.880 15.005 -27.520 ;
        RECT 12.125 -28.960 13.205 -27.880 ;
        RECT 20.265 -28.960 21.345 -25.720 ;
        RECT 24.615 -28.915 25.695 -23.515 ;
        RECT 26.775 -28.915 27.855 -23.515 ;
        RECT 29.015 -23.555 32.255 -22.475 ;
        RECT 33.455 -23.515 36.695 -22.435 ;
        RECT 31.175 -24.635 32.255 -23.555 ;
        RECT 35.615 -24.595 36.695 -23.515 ;
        RECT 12.125 -29.680 15.365 -28.960 ;
        RECT 12.485 -30.040 15.365 -29.680 ;
        RECT 20.265 -30.040 23.505 -28.960 ;
        RECT 24.615 -29.995 27.855 -28.915 ;
        RECT 29.015 -25.715 32.255 -24.635 ;
        RECT 33.455 -25.675 36.695 -24.595 ;
        RECT 29.015 -28.955 30.095 -25.715 ;
        RECT 33.455 -28.915 34.535 -25.675 ;
        RECT 29.015 -30.035 32.255 -28.955 ;
        RECT 33.455 -29.995 36.695 -28.915 ;
  END
END copyright_block
END LIBRARY

