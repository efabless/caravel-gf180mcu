magic
tech gf180mcuC
magscale 1 10
timestamp 1669928529
<< metal1 >>
rect 1494 1198 1569 1452
rect 1812 1238 1887 1462
rect 2838 1198 2913 1452
rect 3156 1238 3231 1462
rect 3958 1198 4033 1452
rect 4276 1238 4351 1462
rect 5302 1198 5377 1452
rect 5620 1238 5695 1462
rect 6422 1198 6497 1452
rect 6740 1238 6815 1462
rect 7766 1198 7841 1452
rect 8084 1238 8159 1462
rect 8886 1198 8961 1452
rect 9204 1238 9279 1462
rect 10230 1198 10305 1452
rect 10548 1238 10623 1462
rect 11350 1198 11425 1452
rect 11668 1238 11743 1462
rect 12694 1198 12769 1452
rect 13012 1238 13087 1462
rect 13814 1198 13889 1452
rect 14132 1238 14207 1462
rect 15158 1198 15233 1452
rect 15476 1238 15551 1462
rect 16278 1198 16353 1452
rect 16596 1238 16671 1462
rect 17622 1198 17697 1452
rect 17940 1238 18015 1462
rect 18742 1198 18817 1452
rect 19060 1238 19135 1462
rect 20086 1198 20161 1452
rect 20404 1238 20479 1462
rect 1364 1126 1569 1198
rect 2708 1126 2913 1198
rect 3828 1126 4033 1198
rect 5172 1126 5377 1198
rect 6292 1126 6497 1198
rect 7636 1126 7841 1198
rect 8756 1126 8961 1198
rect 10100 1126 10305 1198
rect 11220 1126 11425 1198
rect 12564 1126 12769 1198
rect 13684 1126 13889 1198
rect 15028 1126 15233 1198
rect 16148 1126 16353 1198
rect 17492 1126 17697 1198
rect 18612 1126 18817 1198
rect 19956 1126 20161 1198
rect 1364 1107 1436 1126
rect 2708 1107 2780 1126
rect 3828 1107 3900 1126
rect 5172 1107 5244 1126
rect 6292 1107 6364 1126
rect 7636 1107 7708 1126
rect 8756 1107 8828 1126
rect 10100 1107 10172 1126
rect 11220 1107 11292 1126
rect 12564 1107 12636 1126
rect 13684 1107 13756 1126
rect 15028 1107 15100 1126
rect 16148 1107 16220 1126
rect 17492 1107 17564 1126
rect 18612 1107 18684 1126
rect 19956 1107 20028 1126
rect 1364 442 1436 461
rect 2708 442 2780 461
rect 3828 442 3900 461
rect 5172 442 5244 461
rect 6292 442 6364 461
rect 7636 442 7708 461
rect 8756 442 8828 461
rect 10100 442 10172 461
rect 11220 442 11292 461
rect 12564 442 12636 461
rect 13684 442 13756 461
rect 15028 442 15100 461
rect 16148 442 16220 461
rect 16718 449 16778 461
rect 1364 370 1569 442
rect 2708 370 2913 442
rect 3828 370 4033 442
rect 5172 370 5377 442
rect 6292 370 6497 442
rect 7636 370 7841 442
rect 8756 370 8961 442
rect 10100 370 10305 442
rect 11220 370 11425 442
rect 12564 370 12769 442
rect 13684 370 13889 442
rect 15028 370 15233 442
rect 16148 370 16353 442
rect 16718 377 16778 389
rect 17492 442 17564 461
rect 18075 444 18135 456
rect 1494 116 1569 370
rect 1812 106 1887 330
rect 2838 116 2913 370
rect 3156 106 3231 330
rect 3958 116 4033 370
rect 4276 106 4351 330
rect 5302 116 5377 370
rect 5620 106 5695 330
rect 6422 116 6497 370
rect 6740 106 6815 330
rect 7766 116 7841 370
rect 8084 106 8159 330
rect 8886 116 8961 370
rect 9204 106 9279 330
rect 10230 116 10305 370
rect 10548 106 10623 330
rect 11350 116 11425 370
rect 11668 106 11743 330
rect 12694 116 12769 370
rect 13012 106 13087 330
rect 13814 116 13889 370
rect 14132 106 14207 330
rect 15158 116 15233 370
rect 15476 106 15551 330
rect 16278 116 16353 370
rect 16596 106 16671 330
rect 16722 201 16775 377
rect 17492 370 17697 442
rect 18075 372 18135 384
rect 18612 442 18684 461
rect 19190 449 19250 461
rect 16718 189 16778 201
rect 16718 117 16778 129
rect 17622 116 17697 370
rect 17940 106 18015 330
rect 18079 196 18132 372
rect 18612 370 18817 442
rect 19190 377 19250 389
rect 19956 442 20028 461
rect 20531 444 20591 456
rect 18075 184 18135 196
rect 18075 112 18135 124
rect 18742 116 18817 370
rect 19060 106 19135 330
rect 19194 201 19247 377
rect 19956 370 20161 442
rect 20531 372 20591 384
rect 19190 189 19250 201
rect 19190 117 19250 129
rect 20086 116 20161 370
rect 20404 106 20479 330
rect 20536 196 20589 372
rect 20531 184 20591 196
rect 20531 112 20591 124
rect 1716 57 2009 60
rect 2004 -57 2009 57
rect 1716 -60 2009 -57
<< via1 >>
rect 1714 1510 2007 1624
rect 10714 1510 11007 1624
rect 19714 1510 20007 1624
rect 1818 1258 1878 1318
rect 3162 1258 3222 1318
rect 4282 1258 4342 1318
rect 5626 1258 5686 1318
rect 6746 1258 6806 1318
rect 8090 1258 8150 1318
rect 9210 1258 9270 1318
rect 10554 1258 10614 1318
rect 11674 1258 11734 1318
rect 13018 1258 13078 1318
rect 14138 1258 14198 1318
rect 15482 1258 15542 1318
rect 16602 1258 16662 1318
rect 17946 1258 18006 1318
rect 19066 1258 19126 1318
rect 20410 1258 20470 1318
rect 6216 724 6506 844
rect 15216 724 15506 844
rect 16718 389 16778 449
rect 1818 250 1878 310
rect 3162 250 3222 310
rect 4282 250 4342 310
rect 5626 250 5686 310
rect 6746 250 6806 310
rect 8090 250 8150 310
rect 9210 250 9270 310
rect 10554 250 10614 310
rect 11674 250 11734 310
rect 13018 250 13078 310
rect 14138 250 14198 310
rect 15482 250 15542 310
rect 16602 250 16662 310
rect 18075 384 18135 444
rect 16718 129 16778 189
rect 17946 250 18006 310
rect 19190 389 19250 449
rect 18075 124 18135 184
rect 19066 250 19126 310
rect 20531 384 20591 444
rect 19190 129 19250 189
rect 20410 250 20470 310
rect 20531 124 20591 184
rect 1716 -57 2004 57
rect 10716 -57 11004 57
rect 19716 -57 20004 57
<< metal2 >>
rect 1701 1714 2021 1725
rect 1701 1507 1714 1714
rect 1703 1414 1714 1507
rect 2007 1414 2021 1714
rect 10703 1714 11021 1725
rect 10703 1628 10714 1714
rect 10701 1507 10714 1628
rect 1703 1405 2021 1414
rect 10703 1414 10714 1507
rect 11007 1414 11021 1714
rect 19703 1714 20021 1725
rect 19703 1628 19714 1714
rect 19701 1507 19714 1628
rect 10703 1405 11021 1414
rect 19703 1414 19714 1507
rect 20007 1414 20021 1714
rect 19703 1405 20021 1414
rect 1058 1256 1900 1320
rect 2345 1256 3244 1320
rect 3320 1256 4364 1320
rect 4747 1256 5708 1320
rect 6074 1256 6828 1320
rect 6972 1256 8172 1320
rect 8428 1256 9294 1320
rect 9772 1256 10634 1320
rect 11228 1256 11754 1320
rect 12572 1256 13098 1320
rect 13632 1256 14218 1320
rect 14985 1256 15560 1320
rect 16264 1256 16778 1320
rect 17609 1256 18133 1320
rect 18730 1256 19248 1320
rect 20073 1256 20589 1320
rect 1058 488 1114 1256
rect 28 432 1114 488
rect 28 -420 84 432
rect 700 248 1900 312
rect 700 -420 756 248
rect 2345 178 2401 1256
rect 1484 122 2401 178
rect 2549 248 3244 312
rect 1484 -420 1540 122
rect 1703 57 2020 60
rect 1703 -57 1716 57
rect 2004 -57 2020 57
rect 2549 38 2605 248
rect 3320 48 3376 1256
rect 3478 248 4364 312
rect 1703 -144 1726 -57
rect 2000 -144 2020 -57
rect 1703 -163 2020 -144
rect 2156 -18 2605 38
rect 2828 -8 3376 48
rect 2156 -420 2212 -18
rect 2828 -420 2884 -8
rect 3500 -420 3556 248
rect 4747 134 4803 1256
rect 4934 248 5708 312
rect 4172 78 4803 134
rect 4172 -420 4228 78
rect 4956 -420 5012 248
rect 6074 89 6130 1256
rect 6203 942 6520 957
rect 6203 652 6216 942
rect 6506 652 6520 942
rect 6203 637 6520 652
rect 5628 33 6130 89
rect 6300 248 6828 312
rect 5628 -420 5684 33
rect 6300 -420 6356 248
rect 6972 -420 7028 1256
rect 7756 248 8172 312
rect 7756 -420 7812 248
rect 8428 -420 8484 1256
rect 8873 248 9300 312
rect 9100 -420 9156 248
rect 9772 -420 9828 1256
rect 11228 606 11284 1256
rect 12572 632 12628 1256
rect 11223 545 11284 606
rect 12567 572 12628 632
rect 10217 248 10635 312
rect 10444 -420 10500 248
rect 11223 79 11279 545
rect 11337 248 11956 312
rect 10703 57 11020 60
rect 10703 -57 10716 57
rect 11004 -57 11020 57
rect 11223 23 11284 79
rect 10703 -144 10726 -57
rect 11000 -144 11020 -57
rect 10703 -163 11020 -144
rect 11228 -420 11284 23
rect 11900 -420 11956 248
rect 12567 15 12623 572
rect 12681 248 13300 312
rect 12567 -42 12628 15
rect 12572 -420 12628 -42
rect 13244 -420 13300 248
rect 13632 39 13688 1256
rect 13801 248 14756 312
rect 13632 -17 14084 39
rect 14028 -420 14084 -17
rect 14700 -420 14756 248
rect 14985 121 15041 1256
rect 15203 942 15520 957
rect 15203 652 15216 942
rect 15506 652 15520 942
rect 15203 637 15520 652
rect 16722 451 16778 1256
rect 16704 449 16797 451
rect 16704 389 16718 449
rect 16778 389 16797 449
rect 18077 446 18133 1256
rect 19192 451 19248 1256
rect 19178 449 19262 451
rect 16704 387 16797 389
rect 18063 444 18147 446
rect 18063 384 18075 444
rect 18135 384 18147 444
rect 19178 389 19190 449
rect 19250 389 19262 449
rect 20533 446 20589 1256
rect 19178 386 19262 389
rect 20519 444 20603 446
rect 18063 382 18147 384
rect 20519 384 20531 444
rect 20591 384 20603 444
rect 20519 382 20603 384
rect 15145 248 16100 312
rect 16265 248 17551 312
rect 17609 248 18407 312
rect 18727 248 19799 312
rect 20073 248 21700 312
rect 14985 65 15428 121
rect 15372 -420 15428 65
rect 16044 -420 16100 248
rect 16695 189 16797 191
rect 16695 129 16718 189
rect 16778 129 16797 189
rect 16716 127 16797 129
rect 16716 -420 16772 127
rect 17495 -8 17551 248
rect 18063 184 18228 186
rect 18063 124 18075 184
rect 18135 124 18228 184
rect 18063 122 18228 124
rect 17495 -103 17556 -8
rect 17500 -420 17556 -103
rect 18172 -420 18228 122
rect 18351 143 18407 248
rect 19178 189 19572 191
rect 18351 87 18900 143
rect 19178 129 19190 189
rect 19250 135 19572 189
rect 19250 129 19262 135
rect 19178 126 19262 129
rect 18844 -420 18900 87
rect 19516 -420 19572 135
rect 19743 179 19799 248
rect 20519 184 20603 186
rect 19743 123 20356 179
rect 19703 57 20020 60
rect 19703 -57 19716 57
rect 20004 -57 20020 57
rect 19703 -144 19726 -57
rect 20000 -144 20020 -57
rect 19703 -163 20020 -144
rect 20300 -420 20356 123
rect 20519 124 20531 184
rect 20591 181 20603 184
rect 20591 125 21028 181
rect 20591 124 20603 125
rect 20519 122 20603 124
rect 20972 -420 21028 125
rect 21644 -420 21700 248
<< via2 >>
rect 1714 1624 2007 1714
rect 1714 1510 2007 1624
rect 1714 1414 2007 1510
rect 10714 1624 11007 1714
rect 10714 1510 11007 1624
rect 10714 1414 11007 1510
rect 19714 1624 20007 1714
rect 19714 1510 20007 1624
rect 19714 1414 20007 1510
rect 1726 -57 2000 51
rect 1726 -144 2000 -57
rect 6216 844 6506 942
rect 6216 724 6506 844
rect 6216 652 6506 724
rect 10726 -57 11000 51
rect 10726 -144 11000 -57
rect 15216 844 15506 942
rect 15216 724 15506 844
rect 15216 652 15506 724
rect 19726 -57 20000 51
rect 19726 -144 20000 -57
<< metal3 >>
rect 1697 1714 2027 1732
rect 1697 1414 1714 1714
rect 2007 1414 2027 1714
rect 1697 51 2027 1414
rect 1697 -144 1726 51
rect 2000 -144 2027 51
rect 1697 -168 2027 -144
rect 6197 942 6527 1732
rect 6197 652 6216 942
rect 6506 652 6527 942
rect 6197 -168 6527 652
rect 10697 1714 11027 1732
rect 10697 1414 10714 1714
rect 11007 1414 11027 1714
rect 10697 51 11027 1414
rect 10697 -144 10726 51
rect 11000 -144 11027 51
rect 10697 -168 11027 -144
rect 15197 942 15527 1732
rect 15197 652 15216 942
rect 15506 652 15527 942
rect 15197 -168 15527 652
rect 19697 1714 20027 1732
rect 19697 1414 19714 1714
rect 20007 1414 20027 1714
rect 19697 51 20027 1414
rect 19697 -144 19726 51
rect 20000 -144 20027 51
rect 19697 -168 20027 -144
use gf180mcu_fd_sc_mcu7t5v0__endcap  ENDCAP_0 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_scmcu7t5v0/mag
timestamp 1669862171
transform 1 0 896 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  ENDCAP_1
timestamp 1669862171
transform 1 0 20608 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  ENDCAP_2
timestamp 1669862171
transform 1 0 20608 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  ENDCAP_3
timestamp 1669862171
transform 1 0 896 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_0 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_scmcu7t5v0/mag
timestamp 1669862171
transform 1 0 14336 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_1
timestamp 1669862171
transform 1 0 11872 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_2
timestamp 1669862171
transform 1 0 16800 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_3
timestamp 1669862171
transform 1 0 9408 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_4
timestamp 1669862171
transform 1 0 19264 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_5
timestamp 1669862171
transform 1 0 6944 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_6
timestamp 1669862171
transform 1 0 2016 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_7
timestamp 1669862171
transform 1 0 4480 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_8
timestamp 1669862171
transform 1 0 448 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_9
timestamp 1669862171
transform 1 0 448 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_10
timestamp 1669862171
transform 1 0 4480 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_11
timestamp 1669862171
transform 1 0 6944 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_12
timestamp 1669862171
transform 1 0 9408 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_13
timestamp 1669862171
transform 1 0 11872 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_14
timestamp 1669862171
transform 1 0 14336 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_15
timestamp 1669862171
transform 1 0 16800 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_16
timestamp 1669862171
transform 1 0 19264 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_17
timestamp 1669862171
transform 1 0 2016 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_18
timestamp 1669862171
transform 1 0 0 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_19
timestamp 1669862171
transform 1 0 0 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_20
timestamp 1669862171
transform 1 0 21280 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_21
timestamp 1669862171
transform 1 0 21280 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_22
timestamp 1669862171
transform 1 0 20832 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLCAP_4_23
timestamp 1669862171
transform 1 0 20832 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_0 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_scmcu7t5v0/mag
timestamp 1669862171
transform 1 0 13216 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_1
timestamp 1669862171
transform 1 0 15680 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_2
timestamp 1669862171
transform 1 0 18144 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_4
timestamp 1669862171
transform 1 0 10752 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_5
timestamp 1669862171
transform 1 0 8288 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_6
timestamp 1669862171
transform 1 0 5824 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_7
timestamp 1669862171
transform 1 0 3360 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_8
timestamp 1669862171
transform 1 0 3360 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_9
timestamp 1669862171
transform 1 0 5824 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_10
timestamp 1669862171
transform 1 0 8288 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_11
timestamp 1669862171
transform 1 0 10752 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_12
timestamp 1669862171
transform 1 0 13216 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_13
timestamp 1669862171
transform 1 0 15680 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLTIE_14
timestamp 1669862171
transform 1 0 18144 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[0] $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_scmcu7t5v0/mag
timestamp 1669862171
transform 1 0 1120 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[1]
timestamp 1669862171
transform 1 0 1120 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[2]
timestamp 1669862171
transform 1 0 2464 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[3]
timestamp 1669862171
transform 1 0 2464 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[4]
timestamp 1669862171
transform 1 0 3584 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[5]
timestamp 1669862171
transform 1 0 3584 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[6]
timestamp 1669862171
transform 1 0 4928 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[7]
timestamp 1669862171
transform 1 0 4928 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[8]
timestamp 1669862171
transform 1 0 6048 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[9]
timestamp 1669862171
transform 1 0 6048 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[10]
timestamp 1669862171
transform 1 0 7392 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[11]
timestamp 1669862171
transform 1 0 7392 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[12]
timestamp 1669862171
transform 1 0 8512 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[13]
timestamp 1669862171
transform 1 0 8512 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[14]
timestamp 1669862171
transform 1 0 9856 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[15]
timestamp 1669862171
transform 1 0 9856 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[16]
timestamp 1669862171
transform 1 0 10976 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[17]
timestamp 1669862171
transform 1 0 10976 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[18]
timestamp 1669862171
transform 1 0 12320 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[19]
timestamp 1669862171
transform 1 0 12320 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[20]
timestamp 1669862171
transform 1 0 13440 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[21]
timestamp 1669862171
transform 1 0 13440 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[22]
timestamp 1669862171
transform 1 0 14784 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[23]
timestamp 1669862171
transform 1 0 14784 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[24]
timestamp 1669862171
transform 1 0 15904 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[25]
timestamp 1669862171
transform 1 0 15904 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[26]
timestamp 1669862171
transform 1 0 17248 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[27]
timestamp 1669862171
transform 1 0 17248 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[28]
timestamp 1669862171
transform 1 0 18368 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[29]
timestamp 1669862171
transform 1 0 18368 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[30]
timestamp 1669862171
transform 1 0 19712 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  mask_rev_value_one[31]
timestamp 1669862171
transform 1 0 19712 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[0] $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_scmcu7t5v0/mag
timestamp 1669862171
transform 1 0 1568 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[1]
timestamp 1669862171
transform 1 0 1568 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[2]
timestamp 1669862171
transform 1 0 2912 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[3]
timestamp 1669862171
transform 1 0 2912 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[4]
timestamp 1669862171
transform 1 0 4032 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[5]
timestamp 1669862171
transform 1 0 4032 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[6]
timestamp 1669862171
transform 1 0 5376 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[7]
timestamp 1669862171
transform 1 0 5376 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[8]
timestamp 1669862171
transform 1 0 6496 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[9]
timestamp 1669862171
transform 1 0 6496 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[10]
timestamp 1669862171
transform 1 0 7840 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[11]
timestamp 1669862171
transform 1 0 7840 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[12]
timestamp 1669862171
transform 1 0 8960 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[13]
timestamp 1669862171
transform 1 0 8960 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[14]
timestamp 1669862171
transform 1 0 10304 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[15]
timestamp 1669862171
transform 1 0 10304 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[16]
timestamp 1669862171
transform 1 0 11424 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[17]
timestamp 1669862171
transform 1 0 11424 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[18]
timestamp 1669862171
transform 1 0 12768 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[19]
timestamp 1669862171
transform 1 0 12768 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[20]
timestamp 1669862171
transform 1 0 13888 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[21]
timestamp 1669862171
transform 1 0 13888 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[22]
timestamp 1669862171
transform 1 0 15232 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[23]
timestamp 1669862171
transform 1 0 15232 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[24]
timestamp 1669862171
transform 1 0 16352 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[25]
timestamp 1669862171
transform 1 0 16352 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[26]
timestamp 1669862171
transform 1 0 17696 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[27]
timestamp 1669862171
transform 1 0 17696 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[28]
timestamp 1669862171
transform 1 0 18816 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[29]
timestamp 1669862171
transform 1 0 18816 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[30]
timestamp 1669862171
transform 1 0 20160 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  mask_rev_value_zero[31]
timestamp 1669862171
transform 1 0 20160 0 1 0
box -86 -86 534 870
<< labels >>
flabel metal3 6197 -168 6527 162 0 FreeSans 1600 0 0 0 VDD
port 32 nsew
flabel metal3 10697 51 11027 1414 0 FreeSans 1600 0 0 0 VSS
port 33 nsew
flabel metal2 28 -420 84 -10 0 FreeSans 400 90 0 0 mask_rev[0]
port 0 nsew
flabel metal2 700 -420 756 -10 0 FreeSans 400 90 0 0 mask_rev[1]
port 11 nsew
flabel metal2 1484 -420 1540 -10 0 FreeSans 400 90 0 0 mask_rev[2]
port 22 nsew
flabel metal2 2156 -420 2212 -10 0 FreeSans 400 90 0 0 mask_rev[3]
port 25 nsew
flabel metal2 2828 -420 2884 -10 0 FreeSans 400 90 0 0 mask_rev[4]
port 26 nsew
flabel metal2 3500 -420 3556 -10 0 FreeSans 400 90 0 0 mask_rev[5]
port 27 nsew
flabel metal2 4172 -420 4228 -10 0 FreeSans 400 90 0 0 mask_rev[6]
port 28 nsew
flabel metal2 4956 -420 5012 -10 0 FreeSans 400 90 0 0 mask_rev[7]
port 29 nsew
flabel metal2 5628 -420 5684 -10 0 FreeSans 400 90 0 0 mask_rev[8]
port 30 nsew
flabel metal2 6300 -420 6356 -10 0 FreeSans 400 90 0 0 mask_rev[9]
port 31 nsew
flabel metal2 6972 -420 7028 -10 0 FreeSans 400 90 0 0 mask_rev[10]
port 1 nsew
flabel metal2 7756 -420 7812 -10 0 FreeSans 400 90 0 0 mask_rev[11]
port 2 nsew
flabel metal2 8428 -420 8484 -10 0 FreeSans 400 90 0 0 mask_rev[12]
port 3 nsew
flabel metal2 9100 -420 9156 -10 0 FreeSans 400 90 0 0 mask_rev[13]
port 4 nsew
flabel metal2 9772 -420 9828 -10 0 FreeSans 400 90 0 0 mask_rev[14]
port 5 nsew
flabel metal2 10444 -420 10500 -10 0 FreeSans 400 90 0 0 mask_rev[15]
port 6 nsew
flabel metal2 11228 -420 11284 -10 0 FreeSans 400 90 0 0 mask_rev[16]
port 7 nsew
flabel metal2 11900 -420 11956 -10 0 FreeSans 400 90 0 0 mask_rev[17]
port 8 nsew
flabel metal2 12572 -420 12628 -10 0 FreeSans 400 90 0 0 mask_rev[18]
port 9 nsew
flabel metal2 13244 -420 13300 -10 0 FreeSans 400 90 0 0 mask_rev[19]
port 10 nsew
flabel metal2 14028 -420 14084 -10 0 FreeSans 400 90 0 0 mask_rev[20]
port 12 nsew
flabel metal2 14700 -420 14756 -10 0 FreeSans 400 90 0 0 mask_rev[21]
port 13 nsew
flabel metal2 15372 -420 15428 -10 0 FreeSans 400 90 0 0 mask_rev[22]
port 14 nsew
flabel metal2 16044 -420 16100 -10 0 FreeSans 400 90 0 0 mask_rev[23]
port 15 nsew
flabel metal2 16716 -420 16772 -10 0 FreeSans 400 90 0 0 mask_rev[24]
port 16 nsew
flabel metal2 17500 -420 17556 -10 0 FreeSans 400 90 0 0 mask_rev[25]
port 17 nsew
flabel metal2 18172 -420 18228 -10 0 FreeSans 400 90 0 0 mask_rev[26]
port 18 nsew
flabel metal2 18844 -420 18900 -10 0 FreeSans 400 90 0 0 mask_rev[27]
port 19 nsew
flabel metal2 19516 -420 19572 -10 0 FreeSans 400 90 0 0 mask_rev[28]
port 20 nsew
flabel metal2 20300 -420 20356 -10 0 FreeSans 400 90 0 0 mask_rev[29]
port 21 nsew
flabel metal2 20972 -420 21028 -10 0 FreeSans 400 90 0 0 mask_rev[30]
port 23 nsew
flabel metal2 21644 -420 21700 -10 0 FreeSans 400 90 0 0 mask_rev[31]
port 24 nsew
<< end >>
