magic
tech gf180mcuC
magscale 1 10
timestamp 1655130296
<< metal1 >>
rect 1194 33910 1206 33962
rect 1258 33959 1270 33962
rect 2202 33959 2214 33962
rect 1258 33913 2214 33959
rect 1258 33910 1270 33913
rect 2202 33910 2214 33913
rect 2266 33959 2278 33962
rect 2986 33959 2998 33962
rect 2266 33913 2998 33959
rect 2266 33910 2278 33913
rect 2986 33910 2998 33913
rect 3050 33959 3062 33962
rect 4386 33959 4398 33962
rect 3050 33913 4398 33959
rect 3050 33910 3062 33913
rect 4386 33910 4398 33913
rect 4450 33959 4462 33962
rect 5002 33959 5014 33962
rect 4450 33913 5014 33959
rect 4450 33910 4462 33913
rect 5002 33910 5014 33913
rect 5066 33910 5078 33962
rect 336 33738 5696 33772
rect 336 33686 1406 33738
rect 1458 33686 1510 33738
rect 1562 33686 1614 33738
rect 1666 33686 3406 33738
rect 3458 33686 3510 33738
rect 3562 33686 3614 33738
rect 3666 33686 5406 33738
rect 5458 33686 5510 33738
rect 5562 33686 5614 33738
rect 5666 33686 5696 33738
rect 336 33652 5696 33686
rect 4174 33290 4226 33302
rect 4174 33226 4226 33238
rect 4398 33290 4450 33302
rect 4398 33226 4450 33238
rect 4622 33290 4674 33302
rect 4622 33226 4674 33238
rect 5182 33290 5234 33302
rect 5182 33226 5234 33238
rect 336 32954 5600 32988
rect 336 32902 406 32954
rect 458 32902 510 32954
rect 562 32902 614 32954
rect 666 32902 2406 32954
rect 2458 32902 2510 32954
rect 2562 32902 2614 32954
rect 2666 32902 4406 32954
rect 4458 32902 4510 32954
rect 4562 32902 4614 32954
rect 4666 32902 5600 32954
rect 336 32868 5600 32902
rect 3502 32618 3554 32630
rect 3502 32554 3554 32566
rect 5182 32618 5234 32630
rect 5182 32554 5234 32566
rect 4554 32454 4566 32506
rect 4618 32454 4630 32506
rect 3390 32394 3442 32406
rect 3390 32330 3442 32342
rect 3838 32394 3890 32406
rect 3838 32330 3890 32342
rect 3950 32394 4002 32406
rect 3950 32330 4002 32342
rect 4174 32394 4226 32406
rect 4174 32330 4226 32342
rect 4398 32394 4450 32406
rect 4398 32330 4450 32342
rect 4734 32394 4786 32406
rect 4734 32330 4786 32342
rect 336 32170 5696 32204
rect 336 32118 1406 32170
rect 1458 32118 1510 32170
rect 1562 32118 1614 32170
rect 1666 32118 3406 32170
rect 3458 32118 3510 32170
rect 3562 32118 3614 32170
rect 3666 32118 5406 32170
rect 5458 32118 5510 32170
rect 5562 32118 5614 32170
rect 5666 32118 5696 32170
rect 336 32084 5696 32118
rect 1318 31834 1370 31846
rect 1318 31770 1370 31782
rect 3658 31738 3670 31790
rect 3722 31738 3734 31790
rect 5114 31782 5126 31834
rect 5178 31782 5190 31834
rect 4106 31714 4118 31766
rect 4170 31714 4182 31766
rect 4510 31722 4562 31734
rect 4510 31658 4562 31670
rect 646 31610 698 31622
rect 646 31546 698 31558
rect 4790 31610 4842 31622
rect 4790 31546 4842 31558
rect 336 31386 5600 31420
rect 336 31334 406 31386
rect 458 31334 510 31386
rect 562 31334 614 31386
rect 666 31334 2406 31386
rect 2458 31334 2510 31386
rect 2562 31334 2614 31386
rect 2666 31334 4406 31386
rect 4458 31334 4510 31386
rect 4562 31334 4614 31386
rect 4666 31334 5600 31386
rect 336 31300 5600 31334
rect 646 31050 698 31062
rect 646 30986 698 30998
rect 3658 30954 3670 31006
rect 3722 30954 3734 31006
rect 1318 30938 1370 30950
rect 4106 30930 4118 30982
rect 4170 30930 4182 30982
rect 4734 30938 4786 30950
rect 4554 30886 4566 30938
rect 4618 30886 4630 30938
rect 1318 30874 1370 30886
rect 4734 30874 4786 30886
rect 4398 30826 4450 30838
rect 4398 30762 4450 30774
rect 5182 30826 5234 30838
rect 5182 30762 5234 30774
rect 336 30602 5696 30636
rect 336 30550 1406 30602
rect 1458 30550 1510 30602
rect 1562 30550 1614 30602
rect 1666 30550 3406 30602
rect 3458 30550 3510 30602
rect 3562 30550 3614 30602
rect 3666 30550 5406 30602
rect 5458 30550 5510 30602
rect 5562 30550 5614 30602
rect 5666 30550 5696 30602
rect 336 30516 5696 30550
rect 3546 30326 3558 30378
rect 3610 30326 3622 30378
rect 746 30146 758 30198
rect 810 30146 822 30198
rect 1194 30146 1206 30198
rect 1258 30146 1270 30198
rect 4622 30098 4674 30110
rect 4230 30042 4282 30054
rect 4622 30034 4674 30046
rect 4230 29978 4282 29990
rect 4846 29986 4898 29998
rect 5226 29990 5238 30042
rect 5290 29990 5302 30042
rect 4846 29922 4898 29934
rect 336 29818 5600 29852
rect 336 29766 406 29818
rect 458 29766 510 29818
rect 562 29766 614 29818
rect 666 29766 2406 29818
rect 2458 29766 2510 29818
rect 2562 29766 2614 29818
rect 2666 29766 4406 29818
rect 4458 29766 4510 29818
rect 4562 29766 4614 29818
rect 4666 29766 5600 29818
rect 336 29732 5600 29766
rect 1418 29365 1430 29417
rect 1482 29365 1494 29417
rect 1866 29386 1878 29438
rect 1930 29386 1942 29438
rect 4218 29362 4230 29414
rect 4282 29362 4294 29414
rect 4666 29362 4678 29414
rect 4730 29362 4742 29414
rect 646 29258 698 29270
rect 646 29194 698 29206
rect 5182 29258 5234 29270
rect 5182 29194 5234 29206
rect 336 29034 5696 29068
rect 336 28982 1406 29034
rect 1458 28982 1510 29034
rect 1562 28982 1614 29034
rect 1666 28982 3406 29034
rect 3458 28982 3510 29034
rect 3562 28982 3614 29034
rect 3666 28982 5406 29034
rect 5458 28982 5510 29034
rect 5562 28982 5614 29034
rect 5666 28982 5696 29034
rect 336 28948 5696 28982
rect 1082 28582 1094 28634
rect 1146 28582 1158 28634
rect 1586 28590 1598 28642
rect 1650 28590 1662 28642
rect 3994 28578 4006 28630
rect 4058 28578 4070 28630
rect 4554 28578 4566 28630
rect 4618 28578 4630 28630
rect 5238 28474 5290 28486
rect 5238 28410 5290 28422
rect 336 28250 5600 28284
rect 336 28198 406 28250
rect 458 28198 510 28250
rect 562 28198 614 28250
rect 666 28198 2406 28250
rect 2458 28198 2510 28250
rect 2562 28198 2614 28250
rect 2666 28198 4406 28250
rect 4458 28198 4510 28250
rect 4562 28198 4614 28250
rect 4666 28198 5600 28250
rect 336 28164 5600 28198
rect 802 27806 814 27858
rect 866 27806 878 27858
rect 1194 27818 1206 27870
rect 1258 27818 1270 27870
rect 3658 27818 3670 27870
rect 3722 27818 3734 27870
rect 3994 27818 4006 27870
rect 4058 27818 4070 27870
rect 4790 27690 4842 27702
rect 4790 27626 4842 27638
rect 5182 27690 5234 27702
rect 5182 27626 5234 27638
rect 336 27466 5696 27500
rect 336 27414 1406 27466
rect 1458 27414 1510 27466
rect 1562 27414 1614 27466
rect 1666 27414 3406 27466
rect 3458 27414 3510 27466
rect 3562 27414 3614 27466
rect 3666 27414 5406 27466
rect 5458 27414 5510 27466
rect 5562 27414 5614 27466
rect 5666 27414 5696 27466
rect 336 27380 5696 27414
rect 1306 27190 1318 27242
rect 1370 27190 1382 27242
rect 5070 27130 5122 27142
rect 3658 27034 3670 27086
rect 3722 27034 3734 27086
rect 5070 27066 5122 27078
rect 4106 27010 4118 27062
rect 4170 27010 4182 27062
rect 646 26906 698 26918
rect 4846 26906 4898 26918
rect 4442 26854 4454 26906
rect 4506 26854 4518 26906
rect 646 26842 698 26854
rect 4846 26842 4898 26854
rect 336 26682 5600 26716
rect 336 26630 406 26682
rect 458 26630 510 26682
rect 562 26630 614 26682
rect 666 26630 2406 26682
rect 2458 26630 2510 26682
rect 2562 26630 2614 26682
rect 2666 26630 4406 26682
rect 4458 26630 4510 26682
rect 4562 26630 4614 26682
rect 4666 26630 5600 26682
rect 336 26596 5600 26630
rect 3166 26346 3218 26358
rect 3166 26282 3218 26294
rect 4398 26346 4450 26358
rect 4398 26282 4450 26294
rect 4790 26346 4842 26358
rect 4790 26282 4842 26294
rect 5294 26346 5346 26358
rect 5294 26282 5346 26294
rect 4174 26178 4226 26190
rect 3446 26122 3498 26134
rect 3446 26058 3498 26070
rect 3782 26122 3834 26134
rect 4174 26114 4226 26126
rect 3782 26058 3834 26070
rect 336 25898 5696 25932
rect 336 25846 1406 25898
rect 1458 25846 1510 25898
rect 1562 25846 1614 25898
rect 1666 25846 3406 25898
rect 3458 25846 3510 25898
rect 3562 25846 3614 25898
rect 3666 25846 5406 25898
rect 5458 25846 5510 25898
rect 5562 25846 5614 25898
rect 5666 25846 5696 25898
rect 336 25812 5696 25846
rect 4174 25674 4226 25686
rect 4174 25610 4226 25622
rect 4510 25674 4562 25686
rect 4510 25610 4562 25622
rect 4790 25674 4842 25686
rect 4790 25610 4842 25622
rect 5126 25674 5178 25686
rect 5126 25610 5178 25622
rect 4062 25562 4114 25574
rect 4330 25510 4342 25562
rect 4394 25510 4406 25562
rect 4062 25498 4114 25510
rect 336 25114 5600 25148
rect 336 25062 406 25114
rect 458 25062 510 25114
rect 562 25062 614 25114
rect 666 25062 2406 25114
rect 2458 25062 2510 25114
rect 2562 25062 2614 25114
rect 2666 25062 4406 25114
rect 4458 25062 4510 25114
rect 4562 25062 4614 25114
rect 4666 25062 5600 25114
rect 336 25028 5600 25062
rect 4398 24778 4450 24790
rect 4398 24714 4450 24726
rect 5294 24778 5346 24790
rect 5294 24714 5346 24726
rect 4622 24554 4674 24566
rect 4622 24490 4674 24502
rect 336 24330 5696 24364
rect 336 24278 1406 24330
rect 1458 24278 1510 24330
rect 1562 24278 1614 24330
rect 1666 24278 3406 24330
rect 3458 24278 3510 24330
rect 3562 24278 3614 24330
rect 3666 24278 5406 24330
rect 5458 24278 5510 24330
rect 5562 24278 5614 24330
rect 5666 24278 5696 24330
rect 336 24244 5696 24278
rect 4958 24106 5010 24118
rect 3546 24054 3558 24106
rect 3610 24054 3622 24106
rect 4958 24042 5010 24054
rect 5182 24106 5234 24118
rect 5182 24042 5234 24054
rect 746 23898 758 23950
rect 810 23898 822 23950
rect 1194 23874 1206 23926
rect 1258 23874 1270 23926
rect 4398 23882 4450 23894
rect 4398 23818 4450 23830
rect 4622 23882 4674 23894
rect 4622 23818 4674 23830
rect 4230 23770 4282 23782
rect 4230 23706 4282 23718
rect 336 23546 5600 23580
rect 336 23494 406 23546
rect 458 23494 510 23546
rect 562 23494 614 23546
rect 666 23494 2406 23546
rect 2458 23494 2510 23546
rect 2562 23494 2614 23546
rect 2666 23494 4406 23546
rect 4458 23494 4510 23546
rect 4562 23494 4614 23546
rect 4666 23494 5600 23546
rect 336 23460 5600 23494
rect 646 23210 698 23222
rect 646 23146 698 23158
rect 5182 23210 5234 23222
rect 3714 23102 3726 23154
rect 3778 23102 3790 23154
rect 5182 23146 5234 23158
rect 4106 23090 4118 23142
rect 4170 23090 4182 23142
rect 4554 23046 4566 23098
rect 4618 23046 4630 23098
rect 4734 23042 4786 23054
rect 4398 22986 4450 22998
rect 1306 22934 1318 22986
rect 1370 22934 1382 22986
rect 4734 22978 4786 22990
rect 4398 22922 4450 22934
rect 336 22762 5696 22796
rect 336 22710 1406 22762
rect 1458 22710 1510 22762
rect 1562 22710 1614 22762
rect 1666 22710 3406 22762
rect 3458 22710 3510 22762
rect 3562 22710 3614 22762
rect 3666 22710 5406 22762
rect 5458 22710 5510 22762
rect 5562 22710 5614 22762
rect 5666 22710 5696 22762
rect 336 22676 5696 22710
rect 2382 22538 2434 22550
rect 2382 22474 2434 22486
rect 3446 22538 3498 22550
rect 3446 22474 3498 22486
rect 3726 22482 3778 22494
rect 2718 22426 2770 22438
rect 2538 22374 2550 22426
rect 2602 22374 2614 22426
rect 3726 22418 3778 22430
rect 4622 22482 4674 22494
rect 4622 22418 4674 22430
rect 2718 22362 2770 22374
rect 4846 22370 4898 22382
rect 1934 22314 1986 22326
rect 1934 22250 1986 22262
rect 2270 22314 2322 22326
rect 3098 22306 3110 22358
rect 3162 22306 3174 22358
rect 4846 22306 4898 22318
rect 2270 22250 2322 22262
rect 3950 22202 4002 22214
rect 4330 22150 4342 22202
rect 4394 22150 4406 22202
rect 5226 22150 5238 22202
rect 5290 22150 5302 22202
rect 3950 22138 4002 22150
rect 336 21978 5600 22012
rect 336 21926 406 21978
rect 458 21926 510 21978
rect 562 21926 614 21978
rect 666 21926 2406 21978
rect 2458 21926 2510 21978
rect 2562 21926 2614 21978
rect 2666 21926 4406 21978
rect 4458 21926 4510 21978
rect 4562 21926 4614 21978
rect 4666 21926 5600 21978
rect 336 21892 5600 21926
rect 1418 21525 1430 21577
rect 1482 21525 1494 21577
rect 1866 21546 1878 21598
rect 1930 21546 1942 21598
rect 4218 21546 4230 21598
rect 4282 21546 4294 21598
rect 4666 21522 4678 21574
rect 4730 21522 4742 21574
rect 646 21418 698 21430
rect 646 21354 698 21366
rect 5182 21418 5234 21430
rect 5182 21354 5234 21366
rect 336 21194 5696 21228
rect 336 21142 1406 21194
rect 1458 21142 1510 21194
rect 1562 21142 1614 21194
rect 1666 21142 3406 21194
rect 3458 21142 3510 21194
rect 3562 21142 3614 21194
rect 3666 21142 5406 21194
rect 5458 21142 5510 21194
rect 5562 21142 5614 21194
rect 5666 21142 5696 21194
rect 336 21108 5696 21142
rect 1082 20762 1094 20814
rect 1146 20762 1158 20814
rect 1586 20750 1598 20802
rect 1650 20750 1662 20802
rect 4106 20776 4118 20828
rect 4170 20776 4182 20828
rect 4554 20738 4566 20790
rect 4618 20738 4630 20790
rect 5238 20634 5290 20646
rect 5238 20570 5290 20582
rect 336 20410 5600 20444
rect 336 20358 406 20410
rect 458 20358 510 20410
rect 562 20358 614 20410
rect 666 20358 2406 20410
rect 2458 20358 2510 20410
rect 2562 20358 2614 20410
rect 2666 20358 4406 20410
rect 4458 20358 4510 20410
rect 4562 20358 4614 20410
rect 4666 20358 5600 20410
rect 336 20324 5600 20358
rect 3222 20186 3274 20198
rect 3222 20122 3274 20134
rect 5182 20074 5234 20086
rect 5182 20010 5234 20022
rect 4230 19962 4282 19974
rect 4554 19910 4566 19962
rect 4618 19910 4630 19962
rect 4230 19898 4282 19910
rect 2886 19850 2938 19862
rect 2886 19786 2938 19798
rect 336 19626 5696 19660
rect 336 19574 1406 19626
rect 1458 19574 1510 19626
rect 1562 19574 1614 19626
rect 1666 19574 3406 19626
rect 3458 19574 3510 19626
rect 3562 19574 3614 19626
rect 3666 19574 5406 19626
rect 5458 19574 5510 19626
rect 5562 19574 5614 19626
rect 5666 19574 5696 19626
rect 336 19540 5696 19574
rect 2270 19402 2322 19414
rect 2270 19338 2322 19350
rect 2606 19402 2658 19414
rect 2606 19338 2658 19350
rect 4790 19402 4842 19414
rect 4790 19338 4842 19350
rect 5126 19402 5178 19414
rect 5126 19338 5178 19350
rect 2718 19066 2770 19078
rect 2718 19002 2770 19014
rect 336 18842 5600 18876
rect 336 18790 406 18842
rect 458 18790 510 18842
rect 562 18790 614 18842
rect 666 18790 2406 18842
rect 2458 18790 2510 18842
rect 2562 18790 2614 18842
rect 2666 18790 4406 18842
rect 4458 18790 4510 18842
rect 4562 18790 4614 18842
rect 4666 18790 5600 18842
rect 336 18756 5600 18790
rect 3950 18394 4002 18406
rect 3950 18330 4002 18342
rect 4174 18282 4226 18294
rect 4174 18218 4226 18230
rect 4286 18282 4338 18294
rect 5182 18282 5234 18294
rect 4286 18218 4338 18230
rect 4734 18226 4786 18238
rect 5182 18218 5234 18230
rect 4734 18162 4786 18174
rect 336 18058 5696 18092
rect 336 18006 1406 18058
rect 1458 18006 1510 18058
rect 1562 18006 1614 18058
rect 1666 18006 3406 18058
rect 3458 18006 3510 18058
rect 3562 18006 3614 18058
rect 3666 18006 5406 18058
rect 5458 18006 5510 18058
rect 5562 18006 5614 18058
rect 5666 18006 5696 18058
rect 336 17972 5696 18006
rect 2886 17834 2938 17846
rect 2886 17770 2938 17782
rect 4678 17722 4730 17734
rect 5002 17730 5014 17782
rect 5066 17730 5078 17782
rect 4678 17658 4730 17670
rect 2550 17498 2602 17510
rect 3950 17498 4002 17510
rect 2550 17434 2602 17446
rect 3502 17442 3554 17454
rect 3950 17434 4002 17446
rect 4286 17498 4338 17510
rect 4286 17434 4338 17446
rect 3502 17378 3554 17390
rect 336 17274 5600 17308
rect 336 17222 406 17274
rect 458 17222 510 17274
rect 562 17222 614 17274
rect 666 17222 2406 17274
rect 2458 17222 2510 17274
rect 2562 17222 2614 17274
rect 2666 17222 4406 17274
rect 4458 17222 4510 17274
rect 4562 17222 4614 17274
rect 4666 17222 5600 17274
rect 336 17188 5600 17222
rect 2270 17050 2322 17062
rect 4162 16998 4174 17050
rect 4226 16998 4238 17050
rect 2270 16986 2322 16998
rect 3838 16938 3890 16950
rect 3838 16874 3890 16886
rect 5294 16938 5346 16950
rect 5294 16874 5346 16886
rect 2942 16826 2994 16838
rect 2762 16774 2774 16826
rect 2826 16774 2838 16826
rect 4498 16774 4510 16826
rect 4562 16774 4574 16826
rect 4722 16774 4734 16826
rect 4786 16774 4798 16826
rect 2942 16762 2994 16774
rect 2382 16714 2434 16726
rect 2382 16650 2434 16662
rect 2606 16714 2658 16726
rect 2606 16650 2658 16662
rect 3222 16714 3274 16726
rect 3222 16650 3274 16662
rect 3558 16714 3610 16726
rect 3558 16650 3610 16662
rect 336 16490 5696 16524
rect 336 16438 1406 16490
rect 1458 16438 1510 16490
rect 1562 16438 1614 16490
rect 1666 16438 3406 16490
rect 3458 16438 3510 16490
rect 3562 16438 3614 16490
rect 3666 16438 5406 16490
rect 5458 16438 5510 16490
rect 5562 16438 5614 16490
rect 5666 16438 5696 16490
rect 336 16404 5696 16438
rect 1934 16266 1986 16278
rect 1934 16202 1986 16214
rect 2998 16266 3050 16278
rect 2998 16202 3050 16214
rect 3950 16266 4002 16278
rect 3950 16202 4002 16214
rect 4062 16266 4114 16278
rect 4062 16202 4114 16214
rect 2090 16124 2102 16176
rect 2154 16124 2166 16176
rect 2382 16154 2434 16166
rect 2538 16102 2550 16154
rect 2602 16102 2614 16154
rect 2382 16090 2434 16102
rect 2718 16098 2770 16110
rect 1710 16042 1762 16054
rect 2090 15990 2102 16042
rect 2154 15990 2166 16042
rect 2718 16034 2770 16046
rect 3390 16098 3442 16110
rect 4666 16075 4678 16127
rect 4730 16075 4742 16127
rect 4846 16098 4898 16110
rect 3390 16034 3442 16046
rect 5070 16098 5122 16110
rect 4846 16034 4898 16046
rect 4958 16042 5010 16054
rect 1710 15978 1762 15990
rect 3614 15986 3666 15998
rect 5070 16034 5122 16046
rect 4958 15978 5010 15990
rect 3614 15922 3666 15934
rect 4398 15930 4450 15942
rect 4398 15866 4450 15878
rect 336 15706 5600 15740
rect 336 15654 406 15706
rect 458 15654 510 15706
rect 562 15654 614 15706
rect 666 15654 2406 15706
rect 2458 15654 2510 15706
rect 2562 15654 2614 15706
rect 2666 15654 4406 15706
rect 4458 15654 4510 15706
rect 4562 15654 4614 15706
rect 4666 15654 5600 15706
rect 336 15620 5600 15654
rect 1418 15274 1430 15326
rect 1482 15274 1494 15326
rect 1866 15274 1878 15326
rect 1930 15274 1942 15326
rect 4218 15250 4230 15302
rect 4282 15250 4294 15302
rect 4666 15270 4678 15322
rect 4730 15270 4742 15322
rect 5294 15258 5346 15270
rect 5294 15194 5346 15206
rect 646 15146 698 15158
rect 646 15082 698 15094
rect 336 14922 5696 14956
rect 336 14870 1406 14922
rect 1458 14870 1510 14922
rect 1562 14870 1614 14922
rect 1666 14870 3406 14922
rect 3458 14870 3510 14922
rect 3562 14870 3614 14922
rect 3666 14870 5406 14922
rect 5458 14870 5510 14922
rect 5562 14870 5614 14922
rect 5666 14870 5696 14922
rect 336 14836 5696 14870
rect 2158 14698 2210 14710
rect 2158 14634 2210 14646
rect 2494 14698 2546 14710
rect 4958 14698 5010 14710
rect 2494 14634 2546 14646
rect 3390 14642 3442 14654
rect 4386 14646 4398 14698
rect 4450 14646 4462 14698
rect 4958 14634 5010 14646
rect 3390 14578 3442 14590
rect 4846 14586 4898 14598
rect 4846 14522 4898 14534
rect 5114 14486 5126 14538
rect 5178 14486 5190 14538
rect 2886 14362 2938 14374
rect 2886 14298 2938 14310
rect 336 14138 5600 14172
rect 336 14086 406 14138
rect 458 14086 510 14138
rect 562 14086 614 14138
rect 666 14086 2406 14138
rect 2458 14086 2510 14138
rect 2562 14086 2614 14138
rect 2666 14086 4406 14138
rect 4458 14086 4510 14138
rect 4562 14086 4614 14138
rect 4666 14086 5600 14138
rect 336 14052 5600 14086
rect 4790 13914 4842 13926
rect 4790 13850 4842 13862
rect 2830 13802 2882 13814
rect 5182 13802 5234 13814
rect 2830 13738 2882 13750
rect 3054 13746 3106 13758
rect 5182 13738 5234 13750
rect 2314 13638 2326 13690
rect 2378 13638 2390 13690
rect 3054 13682 3106 13694
rect 2046 13578 2098 13590
rect 2046 13514 2098 13526
rect 2158 13578 2210 13590
rect 2158 13514 2210 13526
rect 2494 13578 2546 13590
rect 2494 13514 2546 13526
rect 3446 13578 3498 13590
rect 3446 13514 3498 13526
rect 3670 13578 3722 13590
rect 3670 13514 3722 13526
rect 4006 13578 4058 13590
rect 4006 13514 4058 13526
rect 4454 13578 4506 13590
rect 4454 13514 4506 13526
rect 336 13354 5696 13388
rect 336 13302 1406 13354
rect 1458 13302 1510 13354
rect 1562 13302 1614 13354
rect 1666 13302 3406 13354
rect 3458 13302 3510 13354
rect 3562 13302 3614 13354
rect 3666 13302 5406 13354
rect 5458 13302 5510 13354
rect 5562 13302 5614 13354
rect 5666 13302 5696 13354
rect 336 13268 5696 13302
rect 4622 13130 4674 13142
rect 2046 13074 2098 13086
rect 3042 13078 3054 13130
rect 3106 13078 3118 13130
rect 4622 13066 4674 13078
rect 5238 13130 5290 13142
rect 5238 13066 5290 13078
rect 2046 13010 2098 13022
rect 4890 12966 4902 13018
rect 4954 12966 4966 13018
rect 3390 12906 3442 12918
rect 3390 12842 3442 12854
rect 4286 12850 4338 12862
rect 3658 12742 3670 12794
rect 3722 12742 3734 12794
rect 4286 12786 4338 12798
rect 4062 12738 4114 12750
rect 4062 12674 4114 12686
rect 336 12570 5600 12604
rect 336 12518 406 12570
rect 458 12518 510 12570
rect 562 12518 614 12570
rect 666 12518 2406 12570
rect 2458 12518 2510 12570
rect 2562 12518 2614 12570
rect 2666 12518 4406 12570
rect 4458 12518 4510 12570
rect 4562 12518 4614 12570
rect 4666 12518 5600 12570
rect 336 12484 5600 12518
rect 646 12346 698 12358
rect 646 12282 698 12294
rect 5182 12234 5234 12246
rect 1418 12138 1430 12190
rect 1482 12138 1494 12190
rect 1866 12138 1878 12190
rect 1930 12138 1942 12190
rect 5182 12170 5234 12182
rect 4218 12114 4230 12166
rect 4282 12114 4294 12166
rect 4666 12114 4678 12166
rect 4730 12114 4742 12166
rect 336 11786 5696 11820
rect 336 11734 1406 11786
rect 1458 11734 1510 11786
rect 1562 11734 1614 11786
rect 1666 11734 3406 11786
rect 3458 11734 3510 11786
rect 3562 11734 3614 11786
rect 3666 11734 5406 11786
rect 5458 11734 5510 11786
rect 5562 11734 5614 11786
rect 5666 11734 5696 11786
rect 336 11700 5696 11734
rect 4790 11562 4842 11574
rect 4790 11498 4842 11510
rect 5182 11562 5234 11574
rect 5182 11498 5234 11510
rect 746 11334 758 11386
rect 810 11334 822 11386
rect 1194 11330 1206 11382
rect 1258 11330 1270 11382
rect 3658 11330 3670 11382
rect 3722 11330 3734 11382
rect 4106 11330 4118 11382
rect 4170 11330 4182 11382
rect 4958 11338 5010 11350
rect 4958 11274 5010 11286
rect 336 11002 5600 11036
rect 336 10950 406 11002
rect 458 10950 510 11002
rect 562 10950 614 11002
rect 666 10950 2406 11002
rect 2458 10950 2510 11002
rect 2562 10950 2614 11002
rect 2666 10950 4406 11002
rect 4458 10950 4510 11002
rect 4562 10950 4614 11002
rect 4666 10950 5600 11002
rect 336 10916 5600 10950
rect 4230 10778 4282 10790
rect 4230 10714 4282 10726
rect 4622 10778 4674 10790
rect 4622 10714 4674 10726
rect 5182 10666 5234 10678
rect 4734 10610 4786 10622
rect 5182 10602 5234 10614
rect 3882 10502 3894 10554
rect 3946 10502 3958 10554
rect 4554 10502 4566 10554
rect 4618 10502 4630 10554
rect 4734 10546 4786 10558
rect 3110 10442 3162 10454
rect 3110 10378 3162 10390
rect 3446 10442 3498 10454
rect 3446 10378 3498 10390
rect 336 10218 5696 10252
rect 336 10166 1406 10218
rect 1458 10166 1510 10218
rect 1562 10166 1614 10218
rect 1666 10166 3406 10218
rect 3458 10166 3510 10218
rect 3562 10166 3614 10218
rect 3666 10166 5406 10218
rect 5458 10166 5510 10218
rect 5562 10166 5614 10218
rect 5666 10166 5696 10218
rect 336 10132 5696 10166
rect 646 9994 698 10006
rect 646 9930 698 9942
rect 5070 9994 5122 10006
rect 5070 9930 5122 9942
rect 5182 9994 5234 10006
rect 5182 9930 5234 9942
rect 1418 9783 1430 9835
rect 1482 9783 1494 9835
rect 1866 9762 1878 9814
rect 1930 9762 1942 9814
rect 4218 9762 4230 9814
rect 4282 9762 4294 9814
rect 4834 9774 4846 9826
rect 4898 9774 4910 9826
rect 336 9434 5600 9468
rect 336 9382 406 9434
rect 458 9382 510 9434
rect 562 9382 614 9434
rect 666 9382 2406 9434
rect 2458 9382 2510 9434
rect 2562 9382 2614 9434
rect 2666 9382 4406 9434
rect 4458 9382 4510 9434
rect 4562 9382 4614 9434
rect 4666 9382 5600 9434
rect 336 9348 5600 9382
rect 2718 9210 2770 9222
rect 2718 9146 2770 9158
rect 3390 9210 3442 9222
rect 3994 9158 4006 9210
rect 4058 9158 4070 9210
rect 3390 9146 3442 9158
rect 3166 9098 3218 9110
rect 4622 9098 4674 9110
rect 3166 9034 3218 9046
rect 4398 9042 4450 9054
rect 4622 9034 4674 9046
rect 5182 9098 5234 9110
rect 5182 9034 5234 9046
rect 2650 8934 2662 8986
rect 2714 8934 2726 8986
rect 4398 8978 4450 8990
rect 2382 8874 2434 8886
rect 2382 8810 2434 8822
rect 2830 8874 2882 8886
rect 2830 8810 2882 8822
rect 3782 8874 3834 8886
rect 3782 8810 3834 8822
rect 336 8650 5696 8684
rect 336 8598 1406 8650
rect 1458 8598 1510 8650
rect 1562 8598 1614 8650
rect 1666 8598 3406 8650
rect 3458 8598 3510 8650
rect 3562 8598 3614 8650
rect 3666 8598 5406 8650
rect 5458 8598 5510 8650
rect 5562 8598 5614 8650
rect 5666 8598 5696 8650
rect 336 8564 5696 8598
rect 5238 8426 5290 8438
rect 5238 8362 5290 8374
rect 1082 8198 1094 8250
rect 1146 8198 1158 8250
rect 1698 8206 1710 8258
rect 1762 8206 1774 8258
rect 3994 8194 4006 8246
rect 4058 8194 4070 8246
rect 4554 8194 4566 8246
rect 4618 8194 4630 8246
rect 336 7866 5600 7900
rect 336 7814 406 7866
rect 458 7814 510 7866
rect 562 7814 614 7866
rect 666 7814 2406 7866
rect 2458 7814 2510 7866
rect 2562 7814 2614 7866
rect 2666 7814 4406 7866
rect 4458 7814 4510 7866
rect 4562 7814 4614 7866
rect 4666 7814 5600 7866
rect 336 7780 5600 7814
rect 4790 7642 4842 7654
rect 4790 7578 4842 7590
rect 5294 7530 5346 7542
rect 3994 7478 4006 7530
rect 4058 7478 4070 7530
rect 5294 7466 5346 7478
rect 3994 7344 4006 7396
rect 4058 7344 4070 7396
rect 4442 7366 4454 7418
rect 4506 7366 4518 7418
rect 3502 7306 3554 7318
rect 3502 7242 3554 7254
rect 3838 7306 3890 7318
rect 3838 7242 3890 7254
rect 336 7082 5696 7116
rect 336 7030 1406 7082
rect 1458 7030 1510 7082
rect 1562 7030 1614 7082
rect 1666 7030 3406 7082
rect 3458 7030 3510 7082
rect 3562 7030 3614 7082
rect 3666 7030 5406 7082
rect 5458 7030 5510 7082
rect 5562 7030 5614 7082
rect 5666 7030 5696 7082
rect 336 6996 5696 7030
rect 5182 6634 5234 6646
rect 5182 6570 5234 6582
rect 336 6298 5600 6332
rect 336 6246 406 6298
rect 458 6246 510 6298
rect 562 6246 614 6298
rect 666 6246 2406 6298
rect 2458 6246 2510 6298
rect 2562 6246 2614 6298
rect 2666 6246 4406 6298
rect 4458 6246 4510 6298
rect 4562 6246 4614 6298
rect 4666 6246 5600 6298
rect 336 6212 5600 6246
rect 4622 5962 4674 5974
rect 746 5842 758 5894
rect 810 5842 822 5894
rect 1138 5854 1150 5906
rect 1202 5854 1214 5906
rect 4622 5898 4674 5910
rect 3558 5850 3610 5862
rect 3558 5786 3610 5798
rect 4398 5738 4450 5750
rect 4230 5682 4282 5694
rect 4398 5674 4450 5686
rect 4230 5618 4282 5630
rect 336 5514 5696 5548
rect 336 5462 1406 5514
rect 1458 5462 1510 5514
rect 1562 5462 1614 5514
rect 1666 5462 3406 5514
rect 3458 5462 3510 5514
rect 3562 5462 3614 5514
rect 3666 5462 5406 5514
rect 5458 5462 5510 5514
rect 5562 5462 5614 5514
rect 5666 5462 5696 5514
rect 336 5428 5696 5462
rect 4398 5290 4450 5302
rect 4398 5226 4450 5238
rect 4622 5290 4674 5302
rect 4622 5226 4674 5238
rect 1318 5178 1370 5190
rect 1318 5114 1370 5126
rect 646 5066 698 5078
rect 3714 5070 3726 5122
rect 3778 5070 3790 5122
rect 4218 5082 4230 5134
rect 4282 5082 4294 5134
rect 646 5002 698 5014
rect 336 4730 5600 4764
rect 336 4678 406 4730
rect 458 4678 510 4730
rect 562 4678 614 4730
rect 666 4678 2406 4730
rect 2458 4678 2510 4730
rect 2562 4678 2614 4730
rect 2666 4678 4406 4730
rect 4458 4678 4510 4730
rect 4562 4678 4614 4730
rect 4666 4678 5600 4730
rect 336 4644 5600 4678
rect 4398 4394 4450 4406
rect 746 4298 758 4350
rect 810 4298 822 4350
rect 1194 4298 1206 4350
rect 1258 4298 1270 4350
rect 4398 4330 4450 4342
rect 4622 4394 4674 4406
rect 4622 4330 4674 4342
rect 3558 4282 3610 4294
rect 3558 4218 3610 4230
rect 4230 4114 4282 4126
rect 4230 4050 4282 4062
rect 336 3946 5696 3980
rect 336 3894 1406 3946
rect 1458 3894 1510 3946
rect 1562 3894 1614 3946
rect 1666 3894 3406 3946
rect 3458 3894 3510 3946
rect 3562 3894 3614 3946
rect 3666 3894 5406 3946
rect 5458 3894 5510 3946
rect 5562 3894 5614 3946
rect 5666 3894 5696 3946
rect 336 3860 5696 3894
rect 4790 3722 4842 3734
rect 1306 3670 1318 3722
rect 1370 3670 1382 3722
rect 4790 3658 4842 3670
rect 5070 3610 5122 3622
rect 646 3498 698 3510
rect 3714 3502 3726 3554
rect 3778 3502 3790 3554
rect 4218 3514 4230 3566
rect 4282 3514 4294 3566
rect 5070 3546 5122 3558
rect 646 3434 698 3446
rect 4454 3498 4506 3510
rect 4454 3434 4506 3446
rect 336 3162 5600 3196
rect 336 3110 406 3162
rect 458 3110 510 3162
rect 562 3110 614 3162
rect 666 3110 2406 3162
rect 2458 3110 2510 3162
rect 2562 3110 2614 3162
rect 2666 3110 4406 3162
rect 4458 3110 4510 3162
rect 4562 3110 4614 3162
rect 4666 3110 5600 3162
rect 336 3076 5600 3110
rect 2942 2826 2994 2838
rect 2942 2762 2994 2774
rect 4398 2826 4450 2838
rect 4398 2762 4450 2774
rect 4734 2826 4786 2838
rect 4734 2762 4786 2774
rect 3334 2714 3386 2726
rect 1306 2662 1318 2714
rect 1370 2662 1382 2714
rect 1754 2662 1766 2714
rect 1818 2662 1830 2714
rect 2426 2662 2438 2714
rect 2490 2662 2502 2714
rect 3658 2662 3670 2714
rect 3722 2662 3734 2714
rect 3334 2650 3386 2662
rect 982 2602 1034 2614
rect 982 2538 1034 2550
rect 2102 2602 2154 2614
rect 2102 2538 2154 2550
rect 2774 2602 2826 2614
rect 2774 2538 2826 2550
rect 336 2378 5696 2412
rect 336 2326 1406 2378
rect 1458 2326 1510 2378
rect 1562 2326 1614 2378
rect 1666 2326 3406 2378
rect 3458 2326 3510 2378
rect 3562 2326 3614 2378
rect 3666 2326 5406 2378
rect 5458 2326 5510 2378
rect 5562 2326 5614 2378
rect 5666 2326 5696 2378
rect 336 2292 5696 2326
rect 1766 2154 1818 2166
rect 1766 2090 1818 2102
rect 2382 2154 2434 2166
rect 2382 2090 2434 2102
rect 1430 1818 1482 1830
rect 1430 1754 1482 1766
rect 336 1594 5600 1628
rect 336 1542 406 1594
rect 458 1542 510 1594
rect 562 1542 614 1594
rect 666 1542 2406 1594
rect 2458 1542 2510 1594
rect 2562 1542 2614 1594
rect 2666 1542 4406 1594
rect 4458 1542 4510 1594
rect 4562 1542 4614 1594
rect 4666 1542 5600 1594
rect 336 1508 5600 1542
rect 336 810 5696 844
rect 336 758 1406 810
rect 1458 758 1510 810
rect 1562 758 1614 810
rect 1666 758 3406 810
rect 3458 758 3510 810
rect 3562 758 3614 810
rect 3666 758 5406 810
rect 5458 758 5510 810
rect 5562 758 5614 810
rect 5666 758 5696 810
rect 336 724 5696 758
<< via1 >>
rect 1206 33910 1258 33962
rect 2214 33910 2266 33962
rect 2998 33910 3050 33962
rect 4398 33910 4450 33962
rect 5014 33910 5066 33962
rect 1406 33686 1458 33738
rect 1510 33686 1562 33738
rect 1614 33686 1666 33738
rect 3406 33686 3458 33738
rect 3510 33686 3562 33738
rect 3614 33686 3666 33738
rect 5406 33686 5458 33738
rect 5510 33686 5562 33738
rect 5614 33686 5666 33738
rect 4174 33238 4226 33290
rect 4398 33238 4450 33290
rect 4622 33238 4674 33290
rect 5182 33238 5234 33290
rect 406 32902 458 32954
rect 510 32902 562 32954
rect 614 32902 666 32954
rect 2406 32902 2458 32954
rect 2510 32902 2562 32954
rect 2614 32902 2666 32954
rect 4406 32902 4458 32954
rect 4510 32902 4562 32954
rect 4614 32902 4666 32954
rect 3502 32566 3554 32618
rect 5182 32566 5234 32618
rect 4566 32454 4618 32506
rect 3390 32342 3442 32394
rect 3838 32342 3890 32394
rect 3950 32342 4002 32394
rect 4174 32342 4226 32394
rect 4398 32342 4450 32394
rect 4734 32342 4786 32394
rect 1406 32118 1458 32170
rect 1510 32118 1562 32170
rect 1614 32118 1666 32170
rect 3406 32118 3458 32170
rect 3510 32118 3562 32170
rect 3614 32118 3666 32170
rect 5406 32118 5458 32170
rect 5510 32118 5562 32170
rect 5614 32118 5666 32170
rect 1318 31782 1370 31834
rect 3670 31738 3722 31790
rect 5126 31782 5178 31834
rect 4118 31714 4170 31766
rect 4510 31670 4562 31722
rect 646 31558 698 31610
rect 4790 31558 4842 31610
rect 406 31334 458 31386
rect 510 31334 562 31386
rect 614 31334 666 31386
rect 2406 31334 2458 31386
rect 2510 31334 2562 31386
rect 2614 31334 2666 31386
rect 4406 31334 4458 31386
rect 4510 31334 4562 31386
rect 4614 31334 4666 31386
rect 646 30998 698 31050
rect 3670 30954 3722 31006
rect 1318 30886 1370 30938
rect 4118 30930 4170 30982
rect 4566 30886 4618 30938
rect 4734 30886 4786 30938
rect 4398 30774 4450 30826
rect 5182 30774 5234 30826
rect 1406 30550 1458 30602
rect 1510 30550 1562 30602
rect 1614 30550 1666 30602
rect 3406 30550 3458 30602
rect 3510 30550 3562 30602
rect 3614 30550 3666 30602
rect 5406 30550 5458 30602
rect 5510 30550 5562 30602
rect 5614 30550 5666 30602
rect 3558 30326 3610 30378
rect 758 30146 810 30198
rect 1206 30146 1258 30198
rect 4230 29990 4282 30042
rect 4622 30046 4674 30098
rect 5238 29990 5290 30042
rect 4846 29934 4898 29986
rect 406 29766 458 29818
rect 510 29766 562 29818
rect 614 29766 666 29818
rect 2406 29766 2458 29818
rect 2510 29766 2562 29818
rect 2614 29766 2666 29818
rect 4406 29766 4458 29818
rect 4510 29766 4562 29818
rect 4614 29766 4666 29818
rect 1430 29365 1482 29417
rect 1878 29386 1930 29438
rect 4230 29362 4282 29414
rect 4678 29362 4730 29414
rect 646 29206 698 29258
rect 5182 29206 5234 29258
rect 1406 28982 1458 29034
rect 1510 28982 1562 29034
rect 1614 28982 1666 29034
rect 3406 28982 3458 29034
rect 3510 28982 3562 29034
rect 3614 28982 3666 29034
rect 5406 28982 5458 29034
rect 5510 28982 5562 29034
rect 5614 28982 5666 29034
rect 1094 28582 1146 28634
rect 1598 28590 1650 28642
rect 4006 28578 4058 28630
rect 4566 28578 4618 28630
rect 5238 28422 5290 28474
rect 406 28198 458 28250
rect 510 28198 562 28250
rect 614 28198 666 28250
rect 2406 28198 2458 28250
rect 2510 28198 2562 28250
rect 2614 28198 2666 28250
rect 4406 28198 4458 28250
rect 4510 28198 4562 28250
rect 4614 28198 4666 28250
rect 814 27806 866 27858
rect 1206 27818 1258 27870
rect 3670 27818 3722 27870
rect 4006 27818 4058 27870
rect 4790 27638 4842 27690
rect 5182 27638 5234 27690
rect 1406 27414 1458 27466
rect 1510 27414 1562 27466
rect 1614 27414 1666 27466
rect 3406 27414 3458 27466
rect 3510 27414 3562 27466
rect 3614 27414 3666 27466
rect 5406 27414 5458 27466
rect 5510 27414 5562 27466
rect 5614 27414 5666 27466
rect 1318 27190 1370 27242
rect 3670 27034 3722 27086
rect 5070 27078 5122 27130
rect 4118 27010 4170 27062
rect 646 26854 698 26906
rect 4454 26854 4506 26906
rect 4846 26854 4898 26906
rect 406 26630 458 26682
rect 510 26630 562 26682
rect 614 26630 666 26682
rect 2406 26630 2458 26682
rect 2510 26630 2562 26682
rect 2614 26630 2666 26682
rect 4406 26630 4458 26682
rect 4510 26630 4562 26682
rect 4614 26630 4666 26682
rect 3166 26294 3218 26346
rect 4398 26294 4450 26346
rect 4790 26294 4842 26346
rect 5294 26294 5346 26346
rect 3446 26070 3498 26122
rect 3782 26070 3834 26122
rect 4174 26126 4226 26178
rect 1406 25846 1458 25898
rect 1510 25846 1562 25898
rect 1614 25846 1666 25898
rect 3406 25846 3458 25898
rect 3510 25846 3562 25898
rect 3614 25846 3666 25898
rect 5406 25846 5458 25898
rect 5510 25846 5562 25898
rect 5614 25846 5666 25898
rect 4174 25622 4226 25674
rect 4510 25622 4562 25674
rect 4790 25622 4842 25674
rect 5126 25622 5178 25674
rect 4062 25510 4114 25562
rect 4342 25510 4394 25562
rect 406 25062 458 25114
rect 510 25062 562 25114
rect 614 25062 666 25114
rect 2406 25062 2458 25114
rect 2510 25062 2562 25114
rect 2614 25062 2666 25114
rect 4406 25062 4458 25114
rect 4510 25062 4562 25114
rect 4614 25062 4666 25114
rect 4398 24726 4450 24778
rect 5294 24726 5346 24778
rect 4622 24502 4674 24554
rect 1406 24278 1458 24330
rect 1510 24278 1562 24330
rect 1614 24278 1666 24330
rect 3406 24278 3458 24330
rect 3510 24278 3562 24330
rect 3614 24278 3666 24330
rect 5406 24278 5458 24330
rect 5510 24278 5562 24330
rect 5614 24278 5666 24330
rect 3558 24054 3610 24106
rect 4958 24054 5010 24106
rect 5182 24054 5234 24106
rect 758 23898 810 23950
rect 1206 23874 1258 23926
rect 4398 23830 4450 23882
rect 4622 23830 4674 23882
rect 4230 23718 4282 23770
rect 406 23494 458 23546
rect 510 23494 562 23546
rect 614 23494 666 23546
rect 2406 23494 2458 23546
rect 2510 23494 2562 23546
rect 2614 23494 2666 23546
rect 4406 23494 4458 23546
rect 4510 23494 4562 23546
rect 4614 23494 4666 23546
rect 646 23158 698 23210
rect 5182 23158 5234 23210
rect 3726 23102 3778 23154
rect 4118 23090 4170 23142
rect 4566 23046 4618 23098
rect 1318 22934 1370 22986
rect 4398 22934 4450 22986
rect 4734 22990 4786 23042
rect 1406 22710 1458 22762
rect 1510 22710 1562 22762
rect 1614 22710 1666 22762
rect 3406 22710 3458 22762
rect 3510 22710 3562 22762
rect 3614 22710 3666 22762
rect 5406 22710 5458 22762
rect 5510 22710 5562 22762
rect 5614 22710 5666 22762
rect 2382 22486 2434 22538
rect 3446 22486 3498 22538
rect 2550 22374 2602 22426
rect 2718 22374 2770 22426
rect 3726 22430 3778 22482
rect 4622 22430 4674 22482
rect 1934 22262 1986 22314
rect 2270 22262 2322 22314
rect 3110 22306 3162 22358
rect 4846 22318 4898 22370
rect 3950 22150 4002 22202
rect 4342 22150 4394 22202
rect 5238 22150 5290 22202
rect 406 21926 458 21978
rect 510 21926 562 21978
rect 614 21926 666 21978
rect 2406 21926 2458 21978
rect 2510 21926 2562 21978
rect 2614 21926 2666 21978
rect 4406 21926 4458 21978
rect 4510 21926 4562 21978
rect 4614 21926 4666 21978
rect 1430 21525 1482 21577
rect 1878 21546 1930 21598
rect 4230 21546 4282 21598
rect 4678 21522 4730 21574
rect 646 21366 698 21418
rect 5182 21366 5234 21418
rect 1406 21142 1458 21194
rect 1510 21142 1562 21194
rect 1614 21142 1666 21194
rect 3406 21142 3458 21194
rect 3510 21142 3562 21194
rect 3614 21142 3666 21194
rect 5406 21142 5458 21194
rect 5510 21142 5562 21194
rect 5614 21142 5666 21194
rect 1094 20762 1146 20814
rect 1598 20750 1650 20802
rect 4118 20776 4170 20828
rect 4566 20738 4618 20790
rect 5238 20582 5290 20634
rect 406 20358 458 20410
rect 510 20358 562 20410
rect 614 20358 666 20410
rect 2406 20358 2458 20410
rect 2510 20358 2562 20410
rect 2614 20358 2666 20410
rect 4406 20358 4458 20410
rect 4510 20358 4562 20410
rect 4614 20358 4666 20410
rect 3222 20134 3274 20186
rect 5182 20022 5234 20074
rect 4230 19910 4282 19962
rect 4566 19910 4618 19962
rect 2886 19798 2938 19850
rect 1406 19574 1458 19626
rect 1510 19574 1562 19626
rect 1614 19574 1666 19626
rect 3406 19574 3458 19626
rect 3510 19574 3562 19626
rect 3614 19574 3666 19626
rect 5406 19574 5458 19626
rect 5510 19574 5562 19626
rect 5614 19574 5666 19626
rect 2270 19350 2322 19402
rect 2606 19350 2658 19402
rect 4790 19350 4842 19402
rect 5126 19350 5178 19402
rect 2718 19014 2770 19066
rect 406 18790 458 18842
rect 510 18790 562 18842
rect 614 18790 666 18842
rect 2406 18790 2458 18842
rect 2510 18790 2562 18842
rect 2614 18790 2666 18842
rect 4406 18790 4458 18842
rect 4510 18790 4562 18842
rect 4614 18790 4666 18842
rect 3950 18342 4002 18394
rect 4174 18230 4226 18282
rect 4286 18230 4338 18282
rect 4734 18174 4786 18226
rect 5182 18230 5234 18282
rect 1406 18006 1458 18058
rect 1510 18006 1562 18058
rect 1614 18006 1666 18058
rect 3406 18006 3458 18058
rect 3510 18006 3562 18058
rect 3614 18006 3666 18058
rect 5406 18006 5458 18058
rect 5510 18006 5562 18058
rect 5614 18006 5666 18058
rect 2886 17782 2938 17834
rect 5014 17730 5066 17782
rect 4678 17670 4730 17722
rect 2550 17446 2602 17498
rect 3502 17390 3554 17442
rect 3950 17446 4002 17498
rect 4286 17446 4338 17498
rect 406 17222 458 17274
rect 510 17222 562 17274
rect 614 17222 666 17274
rect 2406 17222 2458 17274
rect 2510 17222 2562 17274
rect 2614 17222 2666 17274
rect 4406 17222 4458 17274
rect 4510 17222 4562 17274
rect 4614 17222 4666 17274
rect 2270 16998 2322 17050
rect 4174 16998 4226 17050
rect 3838 16886 3890 16938
rect 5294 16886 5346 16938
rect 2774 16774 2826 16826
rect 2942 16774 2994 16826
rect 4510 16774 4562 16826
rect 4734 16774 4786 16826
rect 2382 16662 2434 16714
rect 2606 16662 2658 16714
rect 3222 16662 3274 16714
rect 3558 16662 3610 16714
rect 1406 16438 1458 16490
rect 1510 16438 1562 16490
rect 1614 16438 1666 16490
rect 3406 16438 3458 16490
rect 3510 16438 3562 16490
rect 3614 16438 3666 16490
rect 5406 16438 5458 16490
rect 5510 16438 5562 16490
rect 5614 16438 5666 16490
rect 1934 16214 1986 16266
rect 2998 16214 3050 16266
rect 3950 16214 4002 16266
rect 4062 16214 4114 16266
rect 2102 16124 2154 16176
rect 2382 16102 2434 16154
rect 2550 16102 2602 16154
rect 2718 16046 2770 16098
rect 1710 15990 1762 16042
rect 2102 15990 2154 16042
rect 3390 16046 3442 16098
rect 4678 16075 4730 16127
rect 4846 16046 4898 16098
rect 3614 15934 3666 15986
rect 4958 15990 5010 16042
rect 5070 16046 5122 16098
rect 4398 15878 4450 15930
rect 406 15654 458 15706
rect 510 15654 562 15706
rect 614 15654 666 15706
rect 2406 15654 2458 15706
rect 2510 15654 2562 15706
rect 2614 15654 2666 15706
rect 4406 15654 4458 15706
rect 4510 15654 4562 15706
rect 4614 15654 4666 15706
rect 1430 15274 1482 15326
rect 1878 15274 1930 15326
rect 4230 15250 4282 15302
rect 4678 15270 4730 15322
rect 5294 15206 5346 15258
rect 646 15094 698 15146
rect 1406 14870 1458 14922
rect 1510 14870 1562 14922
rect 1614 14870 1666 14922
rect 3406 14870 3458 14922
rect 3510 14870 3562 14922
rect 3614 14870 3666 14922
rect 5406 14870 5458 14922
rect 5510 14870 5562 14922
rect 5614 14870 5666 14922
rect 2158 14646 2210 14698
rect 2494 14646 2546 14698
rect 4398 14646 4450 14698
rect 4958 14646 5010 14698
rect 3390 14590 3442 14642
rect 4846 14534 4898 14586
rect 5126 14486 5178 14538
rect 2886 14310 2938 14362
rect 406 14086 458 14138
rect 510 14086 562 14138
rect 614 14086 666 14138
rect 2406 14086 2458 14138
rect 2510 14086 2562 14138
rect 2614 14086 2666 14138
rect 4406 14086 4458 14138
rect 4510 14086 4562 14138
rect 4614 14086 4666 14138
rect 4790 13862 4842 13914
rect 2830 13750 2882 13802
rect 3054 13694 3106 13746
rect 5182 13750 5234 13802
rect 2326 13638 2378 13690
rect 2046 13526 2098 13578
rect 2158 13526 2210 13578
rect 2494 13526 2546 13578
rect 3446 13526 3498 13578
rect 3670 13526 3722 13578
rect 4006 13526 4058 13578
rect 4454 13526 4506 13578
rect 1406 13302 1458 13354
rect 1510 13302 1562 13354
rect 1614 13302 1666 13354
rect 3406 13302 3458 13354
rect 3510 13302 3562 13354
rect 3614 13302 3666 13354
rect 5406 13302 5458 13354
rect 5510 13302 5562 13354
rect 5614 13302 5666 13354
rect 3054 13078 3106 13130
rect 4622 13078 4674 13130
rect 2046 13022 2098 13074
rect 5238 13078 5290 13130
rect 4902 12966 4954 13018
rect 3390 12854 3442 12906
rect 4286 12798 4338 12850
rect 3670 12742 3722 12794
rect 4062 12686 4114 12738
rect 406 12518 458 12570
rect 510 12518 562 12570
rect 614 12518 666 12570
rect 2406 12518 2458 12570
rect 2510 12518 2562 12570
rect 2614 12518 2666 12570
rect 4406 12518 4458 12570
rect 4510 12518 4562 12570
rect 4614 12518 4666 12570
rect 646 12294 698 12346
rect 1430 12138 1482 12190
rect 1878 12138 1930 12190
rect 5182 12182 5234 12234
rect 4230 12114 4282 12166
rect 4678 12114 4730 12166
rect 1406 11734 1458 11786
rect 1510 11734 1562 11786
rect 1614 11734 1666 11786
rect 3406 11734 3458 11786
rect 3510 11734 3562 11786
rect 3614 11734 3666 11786
rect 5406 11734 5458 11786
rect 5510 11734 5562 11786
rect 5614 11734 5666 11786
rect 4790 11510 4842 11562
rect 5182 11510 5234 11562
rect 758 11334 810 11386
rect 1206 11330 1258 11382
rect 3670 11330 3722 11382
rect 4118 11330 4170 11382
rect 4958 11286 5010 11338
rect 406 10950 458 11002
rect 510 10950 562 11002
rect 614 10950 666 11002
rect 2406 10950 2458 11002
rect 2510 10950 2562 11002
rect 2614 10950 2666 11002
rect 4406 10950 4458 11002
rect 4510 10950 4562 11002
rect 4614 10950 4666 11002
rect 4230 10726 4282 10778
rect 4622 10726 4674 10778
rect 4734 10558 4786 10610
rect 5182 10614 5234 10666
rect 3894 10502 3946 10554
rect 4566 10502 4618 10554
rect 3110 10390 3162 10442
rect 3446 10390 3498 10442
rect 1406 10166 1458 10218
rect 1510 10166 1562 10218
rect 1614 10166 1666 10218
rect 3406 10166 3458 10218
rect 3510 10166 3562 10218
rect 3614 10166 3666 10218
rect 5406 10166 5458 10218
rect 5510 10166 5562 10218
rect 5614 10166 5666 10218
rect 646 9942 698 9994
rect 5070 9942 5122 9994
rect 5182 9942 5234 9994
rect 1430 9783 1482 9835
rect 1878 9762 1930 9814
rect 4230 9762 4282 9814
rect 4846 9774 4898 9826
rect 406 9382 458 9434
rect 510 9382 562 9434
rect 614 9382 666 9434
rect 2406 9382 2458 9434
rect 2510 9382 2562 9434
rect 2614 9382 2666 9434
rect 4406 9382 4458 9434
rect 4510 9382 4562 9434
rect 4614 9382 4666 9434
rect 2718 9158 2770 9210
rect 3390 9158 3442 9210
rect 4006 9158 4058 9210
rect 3166 9046 3218 9098
rect 4398 8990 4450 9042
rect 4622 9046 4674 9098
rect 5182 9046 5234 9098
rect 2662 8934 2714 8986
rect 2382 8822 2434 8874
rect 2830 8822 2882 8874
rect 3782 8822 3834 8874
rect 1406 8598 1458 8650
rect 1510 8598 1562 8650
rect 1614 8598 1666 8650
rect 3406 8598 3458 8650
rect 3510 8598 3562 8650
rect 3614 8598 3666 8650
rect 5406 8598 5458 8650
rect 5510 8598 5562 8650
rect 5614 8598 5666 8650
rect 5238 8374 5290 8426
rect 1094 8198 1146 8250
rect 1710 8206 1762 8258
rect 4006 8194 4058 8246
rect 4566 8194 4618 8246
rect 406 7814 458 7866
rect 510 7814 562 7866
rect 614 7814 666 7866
rect 2406 7814 2458 7866
rect 2510 7814 2562 7866
rect 2614 7814 2666 7866
rect 4406 7814 4458 7866
rect 4510 7814 4562 7866
rect 4614 7814 4666 7866
rect 4790 7590 4842 7642
rect 4006 7478 4058 7530
rect 5294 7478 5346 7530
rect 4006 7344 4058 7396
rect 4454 7366 4506 7418
rect 3502 7254 3554 7306
rect 3838 7254 3890 7306
rect 1406 7030 1458 7082
rect 1510 7030 1562 7082
rect 1614 7030 1666 7082
rect 3406 7030 3458 7082
rect 3510 7030 3562 7082
rect 3614 7030 3666 7082
rect 5406 7030 5458 7082
rect 5510 7030 5562 7082
rect 5614 7030 5666 7082
rect 5182 6582 5234 6634
rect 406 6246 458 6298
rect 510 6246 562 6298
rect 614 6246 666 6298
rect 2406 6246 2458 6298
rect 2510 6246 2562 6298
rect 2614 6246 2666 6298
rect 4406 6246 4458 6298
rect 4510 6246 4562 6298
rect 4614 6246 4666 6298
rect 4622 5910 4674 5962
rect 758 5842 810 5894
rect 1150 5854 1202 5906
rect 3558 5798 3610 5850
rect 4230 5630 4282 5682
rect 4398 5686 4450 5738
rect 1406 5462 1458 5514
rect 1510 5462 1562 5514
rect 1614 5462 1666 5514
rect 3406 5462 3458 5514
rect 3510 5462 3562 5514
rect 3614 5462 3666 5514
rect 5406 5462 5458 5514
rect 5510 5462 5562 5514
rect 5614 5462 5666 5514
rect 4398 5238 4450 5290
rect 4622 5238 4674 5290
rect 1318 5126 1370 5178
rect 3726 5070 3778 5122
rect 4230 5082 4282 5134
rect 646 5014 698 5066
rect 406 4678 458 4730
rect 510 4678 562 4730
rect 614 4678 666 4730
rect 2406 4678 2458 4730
rect 2510 4678 2562 4730
rect 2614 4678 2666 4730
rect 4406 4678 4458 4730
rect 4510 4678 4562 4730
rect 4614 4678 4666 4730
rect 758 4298 810 4350
rect 1206 4298 1258 4350
rect 4398 4342 4450 4394
rect 4622 4342 4674 4394
rect 3558 4230 3610 4282
rect 4230 4062 4282 4114
rect 1406 3894 1458 3946
rect 1510 3894 1562 3946
rect 1614 3894 1666 3946
rect 3406 3894 3458 3946
rect 3510 3894 3562 3946
rect 3614 3894 3666 3946
rect 5406 3894 5458 3946
rect 5510 3894 5562 3946
rect 5614 3894 5666 3946
rect 1318 3670 1370 3722
rect 4790 3670 4842 3722
rect 3726 3502 3778 3554
rect 4230 3514 4282 3566
rect 5070 3558 5122 3610
rect 646 3446 698 3498
rect 4454 3446 4506 3498
rect 406 3110 458 3162
rect 510 3110 562 3162
rect 614 3110 666 3162
rect 2406 3110 2458 3162
rect 2510 3110 2562 3162
rect 2614 3110 2666 3162
rect 4406 3110 4458 3162
rect 4510 3110 4562 3162
rect 4614 3110 4666 3162
rect 2942 2774 2994 2826
rect 4398 2774 4450 2826
rect 4734 2774 4786 2826
rect 1318 2662 1370 2714
rect 1766 2662 1818 2714
rect 2438 2662 2490 2714
rect 3334 2662 3386 2714
rect 3670 2662 3722 2714
rect 982 2550 1034 2602
rect 2102 2550 2154 2602
rect 2774 2550 2826 2602
rect 1406 2326 1458 2378
rect 1510 2326 1562 2378
rect 1614 2326 1666 2378
rect 3406 2326 3458 2378
rect 3510 2326 3562 2378
rect 3614 2326 3666 2378
rect 5406 2326 5458 2378
rect 5510 2326 5562 2378
rect 5614 2326 5666 2378
rect 1766 2102 1818 2154
rect 2382 2102 2434 2154
rect 1430 1766 1482 1818
rect 406 1542 458 1594
rect 510 1542 562 1594
rect 614 1542 666 1594
rect 2406 1542 2458 1594
rect 2510 1542 2562 1594
rect 2614 1542 2666 1594
rect 4406 1542 4458 1594
rect 4510 1542 4562 1594
rect 4614 1542 4666 1594
rect 1406 758 1458 810
rect 1510 758 1562 810
rect 1614 758 1666 810
rect 3406 758 3458 810
rect 3510 758 3562 810
rect 3614 758 3666 810
rect 5406 758 5458 810
rect 5510 758 5562 810
rect 5614 758 5666 810
<< metal2 >>
rect 1204 33962 1260 33974
rect 1204 33910 1206 33962
rect 1258 33910 1260 33962
rect 404 32956 668 32966
rect 460 32900 508 32956
rect 564 32900 612 32956
rect 404 32890 668 32900
rect 1204 31948 1260 33910
rect 2212 33962 2268 35200
rect 2212 33910 2214 33962
rect 2266 33910 2268 33962
rect 2212 33898 2268 33910
rect 1404 33740 1668 33750
rect 1460 33684 1508 33740
rect 1564 33684 1612 33740
rect 1404 33674 1668 33684
rect 2660 33180 2716 35200
rect 2996 33962 3052 33974
rect 2996 33910 2998 33962
rect 3050 33910 3052 33962
rect 2660 33124 2828 33180
rect 2404 32956 2668 32966
rect 2460 32900 2508 32956
rect 2564 32900 2612 32956
rect 2404 32890 2668 32900
rect 1404 32172 1668 32182
rect 1460 32116 1508 32172
rect 1564 32116 1612 32172
rect 1404 32106 1668 32116
rect 2772 31948 2828 33124
rect 1204 31892 1372 31948
rect 1316 31834 1372 31892
rect 2996 31948 3052 33910
rect 3108 32620 3164 35200
rect 3556 34524 3612 35200
rect 4900 34944 6100 35000
rect 3668 34692 4172 34748
rect 3668 34524 3724 34692
rect 3556 34468 3724 34524
rect 3404 33740 3668 33750
rect 3460 33684 3508 33740
rect 3564 33684 3612 33740
rect 3404 33674 3668 33684
rect 4116 33302 4172 34692
rect 4396 33962 4452 33974
rect 4396 33910 4398 33962
rect 4450 33910 4452 33962
rect 4004 33292 4060 33302
rect 4116 33292 4228 33302
rect 4116 33290 4284 33292
rect 4116 33238 4174 33290
rect 4226 33238 4284 33290
rect 4116 33236 4284 33238
rect 3500 32620 3556 32630
rect 4004 32620 4060 33236
rect 4172 33226 4284 33236
rect 4396 33290 4452 33910
rect 4396 33238 4398 33290
rect 4450 33238 4452 33290
rect 4396 33226 4452 33238
rect 4620 33292 4676 33302
rect 4228 32620 4284 33226
rect 4620 33198 4676 33236
rect 4404 32956 4668 32966
rect 4460 32900 4508 32956
rect 4564 32900 4612 32956
rect 4404 32890 4668 32900
rect 3108 32618 4172 32620
rect 3108 32566 3502 32618
rect 3554 32566 4172 32618
rect 3108 32564 4172 32566
rect 4228 32564 4340 32620
rect 3500 32554 3556 32564
rect 3388 32396 3444 32434
rect 4116 32406 4172 32564
rect 3836 32396 3892 32406
rect 3388 32330 3444 32340
rect 3780 32394 3892 32396
rect 3780 32342 3838 32394
rect 3890 32342 3892 32394
rect 3780 32330 3892 32342
rect 3948 32394 4004 32406
rect 3948 32342 3950 32394
rect 4002 32342 4004 32394
rect 3404 32172 3668 32182
rect 3460 32116 3508 32172
rect 3564 32116 3612 32172
rect 3404 32106 3668 32116
rect 3220 32060 3276 32070
rect 3220 31948 3276 32004
rect 2996 31892 3276 31948
rect 2772 31882 2828 31892
rect 1316 31782 1318 31834
rect 1370 31782 1372 31834
rect 644 31612 700 31622
rect 308 31610 812 31612
rect 308 31558 646 31610
rect 698 31558 812 31610
rect 308 31556 812 31558
rect 308 31500 364 31556
rect 644 31546 700 31556
rect 196 31444 364 31500
rect 196 28476 252 31444
rect 404 31388 668 31398
rect 460 31332 508 31388
rect 564 31332 612 31388
rect 404 31322 668 31332
rect 756 31164 812 31556
rect 756 31098 812 31108
rect 644 31050 700 31062
rect 644 30998 646 31050
rect 698 30998 700 31050
rect 644 30940 700 30998
rect 644 30884 1260 30940
rect 756 30198 812 30210
rect 756 30156 758 30198
rect 810 30156 812 30198
rect 756 30090 812 30100
rect 1204 30198 1260 30884
rect 1316 30938 1372 31782
rect 2404 31388 2668 31398
rect 2460 31332 2508 31388
rect 2564 31332 2612 31388
rect 2404 31322 2668 31332
rect 1316 30886 1318 30938
rect 1370 30886 1372 30938
rect 1316 30874 1372 30886
rect 1404 30604 1668 30614
rect 1460 30548 1508 30604
rect 1564 30548 1612 30604
rect 1404 30538 1668 30548
rect 1204 30146 1206 30198
rect 1258 30146 1260 30198
rect 404 29820 668 29830
rect 460 29764 508 29820
rect 564 29764 612 29820
rect 404 29754 668 29764
rect 644 29260 700 29270
rect 1092 29260 1148 29270
rect 644 29258 812 29260
rect 644 29206 646 29258
rect 698 29206 812 29258
rect 644 29204 812 29206
rect 644 29194 700 29204
rect 196 28410 252 28420
rect 404 28252 668 28262
rect 460 28196 508 28252
rect 564 28196 612 28252
rect 404 28186 668 28196
rect 756 28028 812 29204
rect 644 27972 812 28028
rect 1092 28634 1148 29204
rect 1204 28700 1260 30146
rect 3220 30380 3276 31892
rect 3668 31836 3724 31846
rect 3668 31738 3670 31780
rect 3722 31738 3724 31780
rect 3668 31726 3724 31738
rect 3668 31164 3724 31174
rect 3668 31006 3724 31108
rect 3668 30954 3670 31006
rect 3722 30954 3724 31006
rect 3668 30942 3724 30954
rect 3780 30940 3836 32330
rect 3948 32060 4004 32342
rect 3948 31994 4004 32004
rect 4116 32394 4228 32406
rect 4116 32342 4174 32394
rect 4226 32342 4228 32394
rect 4116 32330 4228 32342
rect 4116 31766 4172 32330
rect 4284 32172 4340 32564
rect 4564 32506 4620 32518
rect 4564 32454 4566 32506
rect 4618 32454 4620 32506
rect 4396 32396 4452 32406
rect 4396 32394 4508 32396
rect 4396 32342 4398 32394
rect 4450 32342 4508 32394
rect 4396 32330 4508 32342
rect 4228 32116 4340 32172
rect 4228 31836 4284 32116
rect 4452 31948 4508 32330
rect 4228 31770 4284 31780
rect 4340 31892 4508 31948
rect 4564 31948 4620 32454
rect 4732 32396 4788 32406
rect 4900 32396 4956 34944
rect 5012 33962 5068 33974
rect 5012 33910 5014 33962
rect 5066 33910 5068 33962
rect 5012 32620 5068 33910
rect 5404 33740 5668 33750
rect 5460 33684 5508 33740
rect 5564 33684 5612 33740
rect 5404 33674 5668 33684
rect 5348 33488 6100 33544
rect 5180 33292 5236 33302
rect 5348 33292 5404 33488
rect 5180 33290 5404 33292
rect 5180 33238 5182 33290
rect 5234 33238 5404 33290
rect 5180 33236 5404 33238
rect 5180 33226 5236 33236
rect 5180 32620 5236 32630
rect 5012 32618 5236 32620
rect 5012 32566 5182 32618
rect 5234 32566 5236 32618
rect 5012 32564 5236 32566
rect 5180 32554 5236 32564
rect 5348 32396 5404 33236
rect 4732 32394 4956 32396
rect 4732 32342 4734 32394
rect 4786 32342 4956 32394
rect 4732 32340 4956 32342
rect 5236 32340 5404 32396
rect 4732 32172 4788 32340
rect 4732 32106 4788 32116
rect 5236 31982 5292 32340
rect 5404 32172 5668 32182
rect 5460 32116 5508 32172
rect 5564 32116 5612 32172
rect 5404 32106 5668 32116
rect 4564 31892 4956 31948
rect 5236 31926 5404 31982
rect 4004 31724 4060 31734
rect 3780 30874 3836 30884
rect 3892 31612 3948 31622
rect 3404 30604 3668 30614
rect 3460 30548 3508 30604
rect 3564 30548 3612 30604
rect 3404 30538 3668 30548
rect 3556 30380 3612 30390
rect 3220 30378 3612 30380
rect 3220 30326 3558 30378
rect 3610 30326 3612 30378
rect 3220 30324 3612 30326
rect 1876 30044 1932 30054
rect 1876 29438 1932 29988
rect 2404 29820 2668 29830
rect 2460 29764 2508 29820
rect 2564 29764 2612 29820
rect 2404 29754 2668 29764
rect 1428 29417 1484 29429
rect 1428 29372 1430 29417
rect 1482 29372 1484 29417
rect 1876 29386 1878 29438
rect 1930 29386 1932 29438
rect 1876 29374 1932 29386
rect 1428 29306 1484 29316
rect 1404 29036 1668 29046
rect 1460 28980 1508 29036
rect 1564 28980 1612 29036
rect 1404 28970 1668 28980
rect 1204 28644 1652 28700
rect 1092 28582 1094 28634
rect 1146 28582 1148 28634
rect 644 27132 700 27972
rect 812 27860 868 27870
rect 1092 27860 1148 28582
rect 1596 28642 1652 28644
rect 1596 28590 1598 28642
rect 1650 28590 1652 28642
rect 1596 28578 1652 28590
rect 3220 28588 3276 30324
rect 3556 30314 3612 30324
rect 3780 29372 3836 29382
rect 3404 29036 3668 29046
rect 3460 28980 3508 29036
rect 3564 28980 3612 29036
rect 3404 28970 3668 28980
rect 3668 28812 3724 28822
rect 3220 28532 3500 28588
rect 812 27858 1148 27860
rect 812 27806 814 27858
rect 866 27806 1148 27858
rect 1204 28476 1260 28486
rect 1204 27870 1260 28420
rect 2404 28252 2668 28262
rect 2460 28196 2508 28252
rect 2564 28196 2612 28252
rect 2404 28186 2668 28196
rect 1204 27818 1206 27870
rect 1258 27818 1260 27870
rect 1204 27806 1260 27818
rect 812 27804 1148 27806
rect 812 27794 868 27804
rect 644 27076 1036 27132
rect 644 26908 700 26918
rect 644 26906 812 26908
rect 644 26854 646 26906
rect 698 26854 812 26906
rect 644 26852 812 26854
rect 644 26842 700 26852
rect 756 26796 812 26852
rect 756 26730 812 26740
rect 404 26684 668 26694
rect 460 26628 508 26684
rect 564 26628 612 26684
rect 404 26618 668 26628
rect 404 25116 668 25126
rect 460 25060 508 25116
rect 564 25060 612 25116
rect 404 25050 668 25060
rect 756 23996 812 24006
rect 756 23898 758 23940
rect 810 23898 812 23940
rect 756 23886 812 23898
rect 404 23548 668 23558
rect 460 23492 508 23548
rect 564 23492 612 23548
rect 404 23482 668 23492
rect 644 23212 700 23222
rect 644 23210 812 23212
rect 644 23158 646 23210
rect 698 23158 812 23210
rect 644 23156 812 23158
rect 644 23146 700 23156
rect 404 21980 668 21990
rect 460 21924 508 21980
rect 564 21924 612 21980
rect 404 21914 668 21924
rect 756 21644 812 23156
rect 756 21578 812 21588
rect 644 21420 700 21430
rect 644 21418 924 21420
rect 644 21366 646 21418
rect 698 21366 924 21418
rect 644 21364 924 21366
rect 644 21354 700 21364
rect 404 20412 668 20422
rect 460 20356 508 20412
rect 564 20356 612 20412
rect 404 20346 668 20356
rect 404 18844 668 18854
rect 460 18788 508 18844
rect 564 18788 612 18844
rect 404 18778 668 18788
rect 404 17276 668 17286
rect 460 17220 508 17276
rect 564 17220 612 17276
rect 404 17210 668 17220
rect 404 15708 668 15718
rect 460 15652 508 15708
rect 564 15652 612 15708
rect 404 15642 668 15652
rect 644 15146 700 15158
rect 644 15094 646 15146
rect 698 15094 700 15146
rect -100 14308 100 14328
rect 644 14308 700 15094
rect -100 14252 700 14308
rect 404 14140 668 14150
rect 460 14084 508 14140
rect 564 14084 612 14140
rect 404 14074 668 14084
rect 196 14028 252 14038
rect -100 13804 100 13807
rect 196 13804 252 13972
rect -100 13748 252 13804
rect -100 13731 100 13748
rect -100 13568 100 13578
rect -100 13512 812 13568
rect -100 13502 100 13512
rect -100 13426 100 13436
rect -100 13370 252 13426
rect -100 13360 100 13370
rect 196 13132 252 13370
rect 196 13066 252 13076
rect -100 12924 100 12934
rect -100 12868 252 12924
rect -100 12858 100 12868
rect -100 12713 100 12723
rect -100 12647 140 12713
rect 84 12460 140 12647
rect 84 12394 140 12404
rect 196 9996 252 12868
rect 404 12572 668 12582
rect 460 12516 508 12572
rect 564 12516 612 12572
rect 404 12506 668 12516
rect 644 12348 700 12358
rect 756 12348 812 13512
rect 644 12346 812 12348
rect 644 12294 646 12346
rect 698 12294 812 12346
rect 644 12292 812 12294
rect 644 12282 700 12292
rect 756 11386 812 11398
rect 756 11334 758 11386
rect 810 11334 812 11386
rect 404 11004 668 11014
rect 460 10948 508 11004
rect 564 10948 612 11004
rect 404 10938 668 10948
rect 196 9930 252 9940
rect 644 9996 700 10006
rect 644 9902 700 9940
rect 196 9772 252 9782
rect -100 1260 100 1266
rect 196 1260 252 9716
rect 756 9548 812 11334
rect 868 9772 924 21364
rect 980 12460 1036 27076
rect 1092 21532 1148 27804
rect 1764 27804 1820 27814
rect 1404 27468 1668 27478
rect 1460 27412 1508 27468
rect 1564 27412 1612 27468
rect 1404 27402 1668 27412
rect 1316 27244 1372 27254
rect 1764 27244 1820 27748
rect 3444 27804 3500 28532
rect 3668 27870 3724 28756
rect 3668 27818 3670 27870
rect 3722 27818 3724 27870
rect 3668 27806 3724 27818
rect 3444 27738 3500 27748
rect 3404 27468 3668 27478
rect 3460 27412 3508 27468
rect 3564 27412 3612 27468
rect 3404 27402 3668 27412
rect 1316 27242 1820 27244
rect 1316 27190 1318 27242
rect 1370 27190 1820 27242
rect 1316 27188 1820 27190
rect 3668 27244 3724 27254
rect 1316 27178 1372 27188
rect 3668 27086 3724 27188
rect 3668 27034 3670 27086
rect 3722 27034 3724 27086
rect 3668 27022 3724 27034
rect 3780 26908 3836 29316
rect 3892 28476 3948 31556
rect 4004 28812 4060 31668
rect 4004 28746 4060 28756
rect 4116 31714 4118 31766
rect 4170 31714 4172 31766
rect 4116 30982 4172 31714
rect 4340 31724 4396 31892
rect 4340 31658 4396 31668
rect 4508 31724 4564 31734
rect 4508 31630 4564 31668
rect 4788 31612 4844 31622
rect 4788 31518 4844 31556
rect 4404 31388 4668 31398
rect 4460 31332 4508 31388
rect 4564 31332 4612 31388
rect 4404 31322 4668 31332
rect 4900 31164 4956 31892
rect 5124 31836 5180 31846
rect 5124 31742 5180 31780
rect 4116 30930 4118 30982
rect 4170 30930 4172 30982
rect 4116 30156 4172 30930
rect 4564 31108 4956 31164
rect 5236 31724 5292 31734
rect 4564 30938 4620 31108
rect 4564 30886 4566 30938
rect 4618 30886 4620 30938
rect 4396 30828 4452 30838
rect 3892 28410 3948 28420
rect 4004 28630 4060 28642
rect 4004 28578 4006 28630
rect 4058 28578 4060 28630
rect 4004 28252 4060 28578
rect 3444 26852 3836 26908
rect 3892 28196 4060 28252
rect 3892 26908 3948 28196
rect 4004 28028 4060 28038
rect 4004 27870 4060 27972
rect 4004 27818 4006 27870
rect 4058 27818 4060 27870
rect 4004 27806 4060 27818
rect 4116 27062 4172 30100
rect 4340 30826 4452 30828
rect 4340 30774 4398 30826
rect 4450 30774 4452 30826
rect 4340 30762 4452 30774
rect 4228 30042 4284 30054
rect 4228 29990 4230 30042
rect 4282 29990 4284 30042
rect 4228 29414 4284 29990
rect 4340 30044 4396 30762
rect 4564 30380 4620 30886
rect 4732 30940 4788 30950
rect 4732 30846 4788 30884
rect 4900 30940 4956 30950
rect 4564 30314 4620 30324
rect 4340 29978 4396 29988
rect 4620 30098 4676 30110
rect 4620 30046 4622 30098
rect 4674 30046 4676 30098
rect 4620 30044 4676 30046
rect 4900 29998 4956 30884
rect 5236 30838 5292 31668
rect 5348 30940 5404 31926
rect 5460 31926 6100 31982
rect 5460 31052 5516 31926
rect 5460 30986 5516 30996
rect 5348 30874 5404 30884
rect 5180 30826 5292 30838
rect 5180 30774 5182 30826
rect 5234 30774 5292 30826
rect 5180 30772 5292 30774
rect 5180 30268 5236 30772
rect 5404 30604 5668 30614
rect 5460 30548 5508 30604
rect 5564 30548 5612 30604
rect 5404 30538 5668 30548
rect 4620 29978 4676 29988
rect 4844 29986 4956 29998
rect 4844 29934 4846 29986
rect 4898 29934 4956 29986
rect 4844 29876 4956 29934
rect 4404 29820 4668 29830
rect 4460 29764 4508 29820
rect 4564 29764 4612 29820
rect 4404 29754 4668 29764
rect 4900 29708 4956 29876
rect 4900 29642 4956 29652
rect 5012 30212 5236 30268
rect 5796 30470 6100 30526
rect 4228 29362 4230 29414
rect 4282 29362 4284 29414
rect 4228 27244 4284 29362
rect 4676 29414 4732 29426
rect 4676 29362 4678 29414
rect 4730 29362 4732 29414
rect 4676 29260 4732 29362
rect 4676 29194 4732 29204
rect 5012 29260 5068 30212
rect 5236 30044 5292 30054
rect 5236 30042 5404 30044
rect 5236 29990 5238 30042
rect 5290 29990 5404 30042
rect 5236 29988 5404 29990
rect 5236 29978 5292 29988
rect 5012 29194 5068 29204
rect 5180 29260 5236 29270
rect 5348 29260 5404 29988
rect 5180 29166 5236 29204
rect 5292 29204 5404 29260
rect 5292 29036 5348 29204
rect 5796 29148 5852 30470
rect 5796 29082 5852 29092
rect 5236 28980 5348 29036
rect 5404 29036 5668 29046
rect 5460 28980 5508 29036
rect 5564 28980 5612 29036
rect 4564 28630 4620 28642
rect 4564 28578 4566 28630
rect 4618 28578 4620 28630
rect 4564 28476 4620 28578
rect 5236 28632 5292 28980
rect 5404 28970 5668 28980
rect 5796 28906 6100 28962
rect 5236 28576 5404 28632
rect 4564 28420 4844 28476
rect 4404 28252 4668 28262
rect 4460 28196 4508 28252
rect 4564 28196 4612 28252
rect 4404 28186 4668 28196
rect 4788 27916 4844 28420
rect 4228 27178 4284 27188
rect 4676 27860 4844 27916
rect 5236 28474 5292 28486
rect 5236 28422 5238 28474
rect 5290 28422 5292 28474
rect 5236 27916 5292 28422
rect 4116 27010 4118 27062
rect 4170 27010 4172 27062
rect 3892 26852 4060 26908
rect 1092 20814 1148 21476
rect 1092 20762 1094 20814
rect 1146 20762 1148 20814
rect 1204 26796 1260 26806
rect 1204 23926 1260 26740
rect 2404 26684 2668 26694
rect 2460 26628 2508 26684
rect 2564 26628 2612 26684
rect 2404 26618 2668 26628
rect 3164 26348 3220 26358
rect 3332 26348 3388 26358
rect 3164 26346 3332 26348
rect 3164 26294 3166 26346
rect 3218 26294 3332 26346
rect 3164 26292 3332 26294
rect 3164 26282 3220 26292
rect 3332 26282 3388 26292
rect 3444 26122 3500 26852
rect 3780 26684 3836 26694
rect 3780 26348 3836 26628
rect 3836 26292 3948 26348
rect 3780 26282 3836 26292
rect 3444 26070 3446 26122
rect 3498 26070 3500 26122
rect 3444 26058 3500 26070
rect 3780 26124 3836 26134
rect 3780 26030 3836 26068
rect 1404 25900 1668 25910
rect 1460 25844 1508 25900
rect 1564 25844 1612 25900
rect 1404 25834 1668 25844
rect 3404 25900 3668 25910
rect 3460 25844 3508 25900
rect 3564 25844 3612 25900
rect 3404 25834 3668 25844
rect 2404 25116 2668 25126
rect 2460 25060 2508 25116
rect 2564 25060 2612 25116
rect 2404 25050 2668 25060
rect 3780 25116 3836 25126
rect 1404 24332 1668 24342
rect 1460 24276 1508 24332
rect 1564 24276 1612 24332
rect 1404 24266 1668 24276
rect 3404 24332 3668 24342
rect 3460 24276 3508 24332
rect 3564 24276 3612 24332
rect 3404 24266 3668 24276
rect 3556 24108 3612 24118
rect 3780 24108 3836 25060
rect 1204 23874 1206 23926
rect 1258 23874 1260 23926
rect 1204 20860 1260 23874
rect 3108 24106 3836 24108
rect 3108 24054 3558 24106
rect 3610 24054 3836 24106
rect 3108 24052 3836 24054
rect 2404 23548 2668 23558
rect 2460 23492 2508 23548
rect 2564 23492 2612 23548
rect 2404 23482 2668 23492
rect 2884 23324 2940 23334
rect 1316 22988 1372 22998
rect 1316 22986 1820 22988
rect 1316 22934 1318 22986
rect 1370 22934 1820 22986
rect 1316 22932 1820 22934
rect 1316 22922 1372 22932
rect 1404 22764 1668 22774
rect 1460 22708 1508 22764
rect 1564 22708 1612 22764
rect 1404 22698 1668 22708
rect 1764 22092 1820 22932
rect 2380 22540 2436 22550
rect 2100 22538 2436 22540
rect 2100 22486 2382 22538
rect 2434 22486 2436 22538
rect 2100 22484 2436 22486
rect 1932 22314 1988 22326
rect 1932 22262 1934 22314
rect 1986 22262 1988 22314
rect 1932 22204 1988 22262
rect 1932 22092 1988 22148
rect 1764 22036 1988 22092
rect 1428 21577 1484 21589
rect 1428 21525 1430 21577
rect 1482 21525 1484 21577
rect 1428 21420 1484 21525
rect 1428 21354 1484 21364
rect 1404 21196 1668 21206
rect 1460 21140 1508 21196
rect 1564 21140 1612 21196
rect 1404 21130 1668 21140
rect 1204 20804 1652 20860
rect 1092 20750 1148 20762
rect 1596 20802 1652 20804
rect 1596 20750 1598 20802
rect 1650 20750 1652 20802
rect 1596 20738 1652 20750
rect 1404 19628 1668 19638
rect 1460 19572 1508 19628
rect 1564 19572 1612 19628
rect 1404 19562 1668 19572
rect 1764 19404 1820 22036
rect 2100 21980 2156 22484
rect 2380 22474 2436 22484
rect 2548 22426 2604 22438
rect 2548 22374 2550 22426
rect 2602 22374 2604 22426
rect 2268 22316 2324 22326
rect 2268 22222 2324 22260
rect 2548 22204 2604 22374
rect 2716 22428 2772 22438
rect 2716 22334 2772 22372
rect 2884 22204 2940 23268
rect 2548 22148 2940 22204
rect 1876 21924 2156 21980
rect 2404 21980 2668 21990
rect 2460 21924 2508 21980
rect 2564 21924 2612 21980
rect 1876 21598 1932 21924
rect 2404 21914 2668 21924
rect 2884 21868 2940 22148
rect 3108 22358 3164 24052
rect 3556 24042 3612 24052
rect 3892 23996 3948 26292
rect 4004 25788 4060 26852
rect 4116 26684 4172 27010
rect 4452 26908 4508 26918
rect 4116 26618 4172 26628
rect 4228 26906 4508 26908
rect 4228 26854 4454 26906
rect 4506 26854 4508 26906
rect 4228 26852 4508 26854
rect 4676 26908 4732 27860
rect 5236 27850 5292 27860
rect 5124 27804 5180 27814
rect 5124 27702 5180 27748
rect 4788 27690 4844 27702
rect 4788 27638 4790 27690
rect 4842 27638 4844 27690
rect 4788 27132 4844 27638
rect 5124 27690 5236 27702
rect 5348 27692 5404 28576
rect 5124 27638 5182 27690
rect 5234 27638 5236 27690
rect 5124 27636 5236 27638
rect 5180 27626 5236 27636
rect 5292 27636 5404 27692
rect 5796 27692 5852 28906
rect 5292 27506 5348 27636
rect 5796 27626 5852 27636
rect 5236 27450 5348 27506
rect 5404 27468 5668 27478
rect 4788 27066 4844 27076
rect 4900 27244 4956 27254
rect 4900 26918 4956 27188
rect 5068 27132 5180 27142
rect 5068 27130 5124 27132
rect 5068 27078 5070 27130
rect 5122 27078 5124 27130
rect 5068 27076 5124 27078
rect 5068 27066 5180 27076
rect 4844 26908 4956 26918
rect 5236 26908 5292 27450
rect 5460 27412 5508 27468
rect 5564 27412 5612 27468
rect 5404 27402 5668 27412
rect 5796 27450 6100 27506
rect 4676 26852 4788 26908
rect 4228 26460 4284 26852
rect 4452 26842 4508 26852
rect 4404 26684 4668 26694
rect 4460 26628 4508 26684
rect 4564 26628 4612 26684
rect 4732 26684 4788 26852
rect 4844 26906 4900 26908
rect 4844 26854 4846 26906
rect 4898 26854 4900 26906
rect 4844 26852 4900 26854
rect 4844 26842 4956 26852
rect 5124 26852 5292 26908
rect 4732 26628 4956 26684
rect 4404 26618 4668 26628
rect 4676 26460 4732 26470
rect 4228 26404 4340 26460
rect 4172 26178 4228 26190
rect 4172 26126 4174 26178
rect 4226 26126 4228 26178
rect 4172 26012 4228 26126
rect 4284 26134 4340 26404
rect 4396 26348 4452 26386
rect 4396 26282 4452 26292
rect 4508 26236 4564 26246
rect 4284 26124 4396 26134
rect 4284 26068 4340 26124
rect 4340 26058 4396 26068
rect 4172 25946 4228 25956
rect 4340 25900 4396 25910
rect 4004 25732 4228 25788
rect 4172 25674 4228 25732
rect 4172 25622 4174 25674
rect 4226 25622 4228 25674
rect 4172 25610 4228 25622
rect 4060 25564 4116 25574
rect 4060 25470 4116 25508
rect 4340 25562 4396 25844
rect 4340 25510 4342 25562
rect 4394 25510 4396 25562
rect 4340 25340 4396 25510
rect 4508 25674 4564 26180
rect 4508 25622 4510 25674
rect 4562 25622 4564 25674
rect 4508 25564 4564 25622
rect 4508 25498 4564 25508
rect 4116 25284 4396 25340
rect 4676 25340 4732 26404
rect 4788 26348 4844 26358
rect 4788 26254 4844 26292
rect 4788 25676 4844 25686
rect 4900 25676 4956 26628
rect 4788 25674 4956 25676
rect 4788 25622 4790 25674
rect 4842 25622 4956 25674
rect 4788 25620 4956 25622
rect 5012 26124 5068 26134
rect 4788 25610 4844 25620
rect 4676 25284 4844 25340
rect 4116 24108 4172 25284
rect 4228 25116 4284 25126
rect 4228 24780 4284 25060
rect 4404 25116 4668 25126
rect 4460 25060 4508 25116
rect 4564 25060 4612 25116
rect 4404 25050 4668 25060
rect 4396 24780 4452 24790
rect 4228 24778 4452 24780
rect 4228 24726 4398 24778
rect 4450 24726 4452 24778
rect 4228 24724 4452 24726
rect 3892 23930 3948 23940
rect 4004 24052 4172 24108
rect 3724 23154 3780 23166
rect 3724 23102 3726 23154
rect 3778 23102 3780 23154
rect 3724 23100 3780 23102
rect 4004 23100 4060 24052
rect 3724 23044 3948 23100
rect 3404 22764 3668 22774
rect 3460 22708 3508 22764
rect 3564 22708 3612 22764
rect 3404 22698 3668 22708
rect 3444 22540 3500 22550
rect 3724 22540 3780 22550
rect 3444 22538 3724 22540
rect 3444 22486 3446 22538
rect 3498 22486 3724 22538
rect 3444 22484 3724 22486
rect 3444 22474 3500 22484
rect 3724 22482 3780 22484
rect 3724 22430 3726 22482
rect 3778 22430 3780 22482
rect 3724 22418 3780 22430
rect 3892 22428 3948 23044
rect 4004 23034 4060 23044
rect 4116 23884 4172 23894
rect 4116 23142 4172 23828
rect 4396 23882 4452 24724
rect 4396 23830 4398 23882
rect 4450 23830 4452 23882
rect 4396 23818 4452 23830
rect 4620 24554 4676 24566
rect 4620 24502 4622 24554
rect 4674 24502 4676 24554
rect 4620 23884 4676 24502
rect 4620 23790 4676 23828
rect 4116 23090 4118 23142
rect 4170 23090 4172 23142
rect 3892 22362 3948 22372
rect 4004 22764 4060 22774
rect 3108 22306 3110 22358
rect 3162 22306 3164 22358
rect 3108 22204 3164 22306
rect 4004 22214 4060 22708
rect 3108 22138 3164 22148
rect 3948 22202 4060 22214
rect 3948 22150 3950 22202
rect 4002 22150 4060 22202
rect 3948 22148 4060 22150
rect 3948 22138 4004 22148
rect 4116 21980 4172 23090
rect 4228 23770 4284 23782
rect 4228 23718 4230 23770
rect 4282 23718 4284 23770
rect 4228 22428 4284 23718
rect 4404 23548 4668 23558
rect 4460 23492 4508 23548
rect 4564 23492 4612 23548
rect 4788 23548 4844 25284
rect 5012 24118 5068 26068
rect 5124 25674 5180 26852
rect 5460 26796 5516 26806
rect 5348 26572 5404 26582
rect 5348 26358 5404 26516
rect 5292 26346 5404 26358
rect 5292 26294 5294 26346
rect 5346 26294 5404 26346
rect 5292 26292 5404 26294
rect 5292 26282 5348 26292
rect 5460 26124 5516 26740
rect 5124 25622 5126 25674
rect 5178 25622 5180 25674
rect 5124 25610 5180 25622
rect 5236 26068 5516 26124
rect 5796 26124 5852 27450
rect 5236 24790 5292 26068
rect 5796 26058 5852 26068
rect 5404 25900 5668 25910
rect 5460 25844 5508 25900
rect 5564 25844 5612 25900
rect 5404 25834 5668 25844
rect 5796 25886 6100 25942
rect 5796 25676 5852 25886
rect 5684 25620 5852 25676
rect 5236 24778 5348 24790
rect 5236 24726 5294 24778
rect 5346 24726 5348 24778
rect 5236 24724 5348 24726
rect 5292 24714 5348 24724
rect 5684 24486 5740 25620
rect 5292 24430 5740 24486
rect 5796 24430 6100 24486
rect 4956 24108 5068 24118
rect 5180 24108 5236 24118
rect 4956 24106 5236 24108
rect 4956 24054 4958 24106
rect 5010 24054 5182 24106
rect 5234 24054 5236 24106
rect 4956 24052 5236 24054
rect 5292 24108 5348 24430
rect 5404 24332 5668 24342
rect 5460 24276 5508 24332
rect 5564 24276 5612 24332
rect 5404 24266 5668 24276
rect 5292 24052 5404 24108
rect 4788 23492 4900 23548
rect 4404 23482 4668 23492
rect 4676 23324 4732 23334
rect 4564 23100 4620 23138
rect 4676 23100 4732 23268
rect 4844 23212 4900 23492
rect 4956 23436 5012 24052
rect 5180 24042 5236 24052
rect 4956 23370 5012 23380
rect 5236 23884 5292 23894
rect 5236 23222 5292 23828
rect 4844 23156 5068 23212
rect 4676 23044 4788 23100
rect 4564 23034 4620 23044
rect 4732 23042 4788 23044
rect 4396 22988 4452 22998
rect 4732 22990 4734 23042
rect 4786 22990 4788 23042
rect 4396 22986 4508 22988
rect 4396 22934 4398 22986
rect 4450 22934 4508 22986
rect 4396 22922 4508 22934
rect 4228 22362 4284 22372
rect 4340 22204 4396 22214
rect 3780 21924 4172 21980
rect 4228 22202 4396 22204
rect 4228 22150 4342 22202
rect 4394 22150 4396 22202
rect 4228 22148 4396 22150
rect 2884 21812 3276 21868
rect 1876 21546 1878 21598
rect 1930 21546 1932 21598
rect 1876 21534 1932 21546
rect 1764 19338 1820 19348
rect 2100 20636 2156 20646
rect 1404 18060 1668 18070
rect 1460 18004 1508 18060
rect 1564 18004 1612 18060
rect 1404 17994 1668 18004
rect 2100 17052 2156 20580
rect 2404 20412 2668 20422
rect 2460 20356 2508 20412
rect 2564 20356 2612 20412
rect 2404 20346 2668 20356
rect 3220 20186 3276 21812
rect 3404 21196 3668 21206
rect 3460 21140 3508 21196
rect 3564 21140 3612 21196
rect 3404 21130 3668 21140
rect 3220 20134 3222 20186
rect 3274 20134 3276 20186
rect 3220 20122 3276 20134
rect 2884 19850 2940 19862
rect 2884 19798 2886 19850
rect 2938 19798 2940 19850
rect 2268 19404 2324 19414
rect 2268 19310 2324 19348
rect 2604 19404 2660 19414
rect 2604 19310 2660 19348
rect 2716 19068 2772 19078
rect 2884 19068 2940 19798
rect 3404 19628 3668 19638
rect 3460 19572 3508 19628
rect 3564 19572 3612 19628
rect 3404 19562 3668 19572
rect 2716 19066 2940 19068
rect 2716 19014 2718 19066
rect 2770 19014 2940 19066
rect 2716 19012 2940 19014
rect 2716 19002 2828 19012
rect 2404 18844 2668 18854
rect 2460 18788 2508 18844
rect 2564 18788 2612 18844
rect 2404 18778 2668 18788
rect 2772 17836 2828 19002
rect 3404 18060 3668 18070
rect 3460 18004 3508 18060
rect 3564 18004 3612 18060
rect 3404 17994 3668 18004
rect 3780 18060 3836 21924
rect 3892 21756 3948 21766
rect 4228 21756 4284 22148
rect 4340 22138 4396 22148
rect 4452 22204 4508 22922
rect 4620 22876 4676 22886
rect 4620 22540 4676 22820
rect 4732 22652 4788 22990
rect 4732 22596 4900 22652
rect 4620 22482 4676 22484
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22408 4676 22430
rect 4844 22370 4900 22596
rect 4844 22318 4846 22370
rect 4898 22318 4900 22370
rect 4844 22306 4900 22318
rect 4452 22138 4508 22148
rect 4404 21980 4668 21990
rect 4460 21924 4508 21980
rect 4564 21924 4612 21980
rect 4404 21914 4668 21924
rect 5012 21868 5068 23156
rect 5180 23210 5292 23222
rect 5180 23158 5182 23210
rect 5234 23158 5292 23210
rect 5180 23156 5292 23158
rect 5180 22988 5236 23156
rect 5180 22922 5236 22932
rect 5348 22922 5404 24052
rect 5796 23100 5852 24430
rect 5796 23034 5852 23044
rect 5292 22866 5404 22922
rect 5460 22922 5516 22932
rect 5516 22866 6100 22922
rect 5292 22764 5348 22866
rect 5460 22856 5516 22866
rect 4900 21812 5068 21868
rect 5124 22708 5348 22764
rect 5404 22764 5668 22774
rect 5460 22708 5508 22764
rect 5564 22708 5612 22764
rect 5124 21868 5180 22708
rect 5404 22698 5668 22708
rect 5236 22204 5292 22214
rect 5236 22202 5404 22204
rect 5236 22150 5238 22202
rect 5290 22150 5404 22202
rect 5236 22148 5404 22150
rect 5236 22138 5292 22148
rect 4452 21756 4508 21766
rect 3948 21700 4060 21756
rect 4228 21700 4396 21756
rect 3892 21690 3948 21700
rect 4004 21644 4060 21700
rect 4004 21598 4284 21644
rect 4004 21588 4230 21598
rect 4228 21546 4230 21588
rect 4282 21546 4284 21598
rect 4228 21534 4284 21546
rect 4340 21466 4396 21700
rect 4004 21420 4060 21430
rect 4004 19964 4060 21364
rect 4228 21410 4396 21466
rect 4116 21308 4172 21318
rect 4116 20828 4172 21252
rect 4116 20776 4118 20828
rect 4170 20776 4172 20828
rect 4116 20764 4172 20776
rect 4228 20188 4284 21410
rect 4452 21308 4508 21700
rect 4676 21574 4732 21586
rect 4676 21532 4678 21574
rect 4730 21532 4732 21574
rect 4676 21466 4732 21476
rect 4452 21242 4508 21252
rect 4564 20790 4620 20802
rect 4564 20738 4566 20790
rect 4618 20738 4620 20790
rect 4564 20636 4620 20738
rect 4564 20580 4844 20636
rect 4404 20412 4668 20422
rect 4460 20356 4508 20412
rect 4564 20356 4612 20412
rect 4404 20346 4668 20356
rect 4228 20132 4396 20188
rect 4228 19964 4284 19974
rect 4004 19962 4284 19964
rect 4004 19910 4230 19962
rect 4282 19910 4284 19962
rect 4004 19908 4284 19910
rect 4340 19964 4396 20132
rect 4564 19964 4620 19974
rect 4340 19962 4620 19964
rect 4340 19910 4566 19962
rect 4618 19910 4620 19962
rect 4340 19908 4620 19910
rect 4228 19898 4284 19908
rect 4564 19898 4620 19908
rect 4788 19402 4844 20580
rect 4788 19350 4790 19402
rect 4842 19350 4844 19402
rect 4788 19338 4844 19350
rect 4404 18844 4668 18854
rect 4460 18788 4508 18844
rect 4564 18788 4612 18844
rect 4404 18778 4668 18788
rect 3948 18396 4004 18406
rect 3948 18302 4004 18340
rect 4172 18284 4228 18294
rect 4172 18190 4228 18228
rect 4284 18282 4340 18294
rect 4284 18230 4286 18282
rect 4338 18230 4340 18282
rect 3780 17994 3836 18004
rect 2884 17836 2940 17846
rect 2772 17834 2940 17836
rect 2772 17782 2886 17834
rect 2938 17782 2940 17834
rect 2772 17780 2940 17782
rect 2884 17770 2940 17780
rect 4284 17724 4340 18230
rect 4732 18226 4788 18238
rect 4732 18174 4734 18226
rect 4786 18174 4788 18226
rect 4732 17948 4788 18174
rect 4732 17892 4844 17948
rect 4564 17836 4620 17846
rect 4564 17724 4620 17780
rect 4676 17724 4732 17734
rect 4564 17722 4732 17724
rect 4564 17670 4678 17722
rect 4730 17670 4732 17722
rect 4564 17668 4732 17670
rect 4284 17658 4340 17668
rect 4676 17658 4732 17668
rect 2772 17612 2828 17622
rect 2548 17500 2604 17538
rect 2548 17434 2604 17444
rect 2404 17276 2668 17286
rect 2460 17220 2508 17276
rect 2564 17220 2612 17276
rect 2404 17210 2668 17220
rect 2268 17052 2324 17062
rect 2100 17050 2324 17052
rect 2100 16998 2270 17050
rect 2322 16998 2324 17050
rect 2100 16996 2324 16998
rect 2268 16986 2324 16996
rect 2772 16826 2828 17556
rect 3780 17612 3836 17622
rect 3500 17442 3556 17454
rect 3500 17390 3502 17442
rect 3554 17390 3556 17442
rect 3500 16940 3556 17390
rect 3500 16874 3556 16884
rect 3780 16950 3836 17556
rect 3948 17498 4004 17510
rect 3948 17446 3950 17498
rect 4002 17446 4004 17498
rect 3948 17052 4004 17446
rect 4284 17500 4340 17510
rect 4284 17406 4340 17444
rect 4404 17276 4668 17286
rect 4460 17220 4508 17276
rect 4564 17220 4612 17276
rect 4404 17210 4668 17220
rect 4788 17164 4844 17892
rect 4788 17098 4844 17108
rect 3948 16986 4004 16996
rect 4172 17052 4228 17062
rect 4172 16958 4228 16996
rect 3780 16938 3892 16950
rect 3780 16886 3838 16938
rect 3890 16886 3892 16938
rect 3780 16874 3892 16886
rect 4732 16940 4788 16950
rect 2772 16774 2774 16826
rect 2826 16774 2828 16826
rect 2772 16762 2828 16774
rect 2940 16828 2996 16838
rect 2940 16734 2996 16772
rect 3780 16828 3836 16874
rect 3780 16762 3836 16772
rect 4060 16828 4116 16838
rect 4508 16828 4564 16838
rect 1932 16716 1988 16726
rect 1404 16492 1668 16502
rect 1460 16436 1508 16492
rect 1564 16436 1612 16492
rect 1404 16426 1668 16436
rect 1932 16266 1988 16660
rect 2380 16714 2436 16726
rect 2380 16662 2382 16714
rect 2434 16662 2436 16714
rect 2380 16380 2436 16662
rect 2548 16716 2660 16726
rect 2604 16714 2660 16716
rect 2604 16662 2606 16714
rect 2658 16662 2660 16714
rect 2604 16660 2660 16662
rect 2548 16650 2660 16660
rect 3108 16716 3164 16726
rect 2380 16314 2436 16324
rect 1932 16214 1934 16266
rect 1986 16214 1988 16266
rect 1932 16202 1988 16214
rect 2100 16268 2156 16278
rect 2100 16176 2156 16212
rect 2996 16268 3052 16278
rect 3108 16268 3164 16660
rect 2996 16266 3164 16268
rect 2996 16214 2998 16266
rect 3050 16214 3164 16266
rect 2996 16212 3164 16214
rect 3220 16714 3276 16726
rect 3220 16662 3222 16714
rect 3274 16662 3276 16714
rect 2996 16202 3052 16212
rect 2100 16124 2102 16176
rect 2154 16124 2156 16176
rect 2380 16156 2436 16166
rect 2100 16112 2156 16124
rect 2212 16154 2436 16156
rect 2212 16102 2382 16154
rect 2434 16102 2436 16154
rect 2212 16100 2436 16102
rect 1708 16042 1764 16054
rect 1708 15990 1710 16042
rect 1762 15990 1764 16042
rect 1708 15932 1764 15990
rect 2100 16044 2156 16054
rect 2100 15950 2156 15988
rect 1708 15866 1764 15876
rect 2212 15708 2268 16100
rect 2380 16090 2436 16100
rect 2548 16156 2604 16166
rect 2548 16062 2604 16100
rect 2716 16098 2772 16110
rect 2716 16046 2718 16098
rect 2770 16046 2772 16098
rect 2716 15932 2772 16046
rect 2716 15866 2772 15876
rect 1876 15652 2268 15708
rect 2404 15708 2668 15718
rect 2460 15652 2508 15708
rect 2564 15652 2612 15708
rect 1428 15372 1484 15382
rect 1428 15274 1430 15316
rect 1482 15274 1484 15316
rect 1428 15262 1484 15274
rect 1876 15326 1932 15652
rect 2404 15642 2668 15652
rect 1876 15274 1878 15326
rect 1930 15274 1932 15326
rect 3220 15372 3276 16662
rect 3556 16716 3612 16754
rect 3556 16650 3612 16660
rect 3404 16492 3668 16502
rect 3460 16436 3508 16492
rect 3564 16436 3612 16492
rect 3404 16426 3668 16436
rect 3948 16268 4004 16278
rect 3948 16174 4004 16212
rect 4060 16266 4116 16772
rect 4060 16214 4062 16266
rect 4114 16214 4116 16266
rect 4060 16202 4116 16214
rect 4340 16826 4564 16828
rect 4340 16774 4510 16826
rect 4562 16774 4564 16826
rect 4340 16772 4564 16774
rect 3388 16156 3444 16166
rect 4340 16156 4396 16772
rect 4508 16762 4564 16772
rect 4732 16826 4788 16884
rect 4732 16774 4734 16826
rect 4786 16774 4788 16826
rect 4732 16716 4788 16774
rect 4900 16828 4956 21812
rect 5124 21802 5180 21812
rect 5348 21644 5404 22148
rect 5012 21588 5404 21644
rect 5012 19404 5068 21588
rect 5180 21420 5236 21430
rect 5124 21364 5180 21420
rect 5124 21326 5236 21364
rect 5796 21410 6100 21466
rect 5124 20086 5180 21326
rect 5404 21196 5668 21206
rect 5460 21140 5508 21196
rect 5564 21140 5612 21196
rect 5404 21130 5668 21140
rect 5236 20636 5292 20646
rect 5236 20542 5292 20580
rect 5124 20074 5236 20086
rect 5124 20022 5182 20074
rect 5234 20022 5236 20074
rect 5124 20020 5236 20022
rect 5180 20010 5236 20020
rect 5796 19740 5852 21410
rect 5796 19674 5852 19684
rect 5404 19628 5668 19638
rect 5460 19572 5508 19628
rect 5564 19572 5612 19628
rect 5404 19562 5668 19572
rect 5124 19404 5180 19414
rect 5012 19402 5180 19404
rect 5012 19350 5126 19402
rect 5178 19350 5180 19402
rect 5012 19348 5180 19350
rect 5124 19338 5180 19348
rect 5012 18956 5068 18966
rect 5012 18396 5068 18900
rect 5012 17782 5068 18340
rect 5348 18508 5404 18518
rect 5180 18284 5236 18294
rect 5348 18284 5404 18452
rect 5180 18190 5236 18228
rect 5292 18228 5404 18284
rect 5012 17730 5014 17782
rect 5066 17730 5068 17782
rect 5292 17836 5348 18228
rect 5404 18060 5668 18070
rect 5460 18004 5508 18060
rect 5564 18004 5612 18060
rect 5404 17994 5668 18004
rect 5292 17780 5404 17836
rect 5012 17718 5068 17730
rect 5124 17724 5180 17734
rect 4900 16762 4956 16772
rect 4732 16650 4788 16660
rect 3388 16098 3444 16100
rect 3388 16046 3390 16098
rect 3442 16046 3444 16098
rect 3388 15932 3444 16046
rect 4228 16100 4396 16156
rect 4452 16380 4508 16390
rect 5124 16380 5180 17668
rect 5348 17500 5404 17780
rect 5348 16950 5404 17444
rect 5684 17052 5740 17062
rect 5740 16996 5964 17052
rect 5684 16986 5740 16996
rect 5292 16938 5404 16950
rect 5292 16886 5294 16938
rect 5346 16886 5404 16938
rect 5292 16884 5404 16886
rect 5292 16874 5348 16884
rect 5404 16492 5668 16502
rect 5460 16436 5508 16492
rect 5564 16436 5612 16492
rect 5404 16426 5668 16436
rect 5124 16324 5292 16380
rect 3388 15866 3444 15876
rect 3612 15986 3668 15998
rect 3612 15934 3614 15986
rect 3666 15934 3668 15986
rect 3612 15372 3668 15934
rect 4228 15484 4284 16100
rect 4452 15942 4508 16324
rect 4676 16268 4732 16278
rect 4676 16127 4732 16212
rect 4676 16075 4678 16127
rect 4730 16075 4732 16127
rect 4676 16063 4732 16075
rect 4844 16098 4900 16110
rect 4844 16054 4846 16098
rect 4788 16046 4846 16054
rect 4898 16046 4900 16098
rect 5068 16098 5124 16110
rect 4788 16044 4900 16046
rect 4844 15988 4900 16044
rect 4956 16044 5012 16054
rect 4788 15978 4844 15988
rect 4956 15950 5012 15988
rect 5068 16046 5070 16098
rect 5122 16046 5124 16098
rect 4396 15930 4508 15942
rect 4396 15878 4398 15930
rect 4450 15878 4508 15930
rect 4396 15876 4508 15878
rect 4396 15866 4452 15876
rect 4404 15708 4668 15718
rect 4460 15652 4508 15708
rect 4564 15652 4612 15708
rect 4404 15642 4668 15652
rect 5068 15596 5124 16046
rect 5012 15540 5124 15596
rect 4228 15428 4396 15484
rect 3612 15316 3836 15372
rect 3220 15306 3276 15316
rect 1876 15262 1932 15274
rect 1404 14924 1668 14934
rect 1460 14868 1508 14924
rect 1564 14868 1612 14924
rect 1404 14858 1668 14868
rect 3404 14924 3668 14934
rect 3460 14868 3508 14924
rect 3564 14868 3612 14924
rect 3404 14858 3668 14868
rect 2156 14700 2212 14710
rect 2156 14606 2212 14644
rect 2436 14700 2548 14710
rect 2492 14698 2548 14700
rect 2492 14646 2494 14698
rect 2546 14646 2548 14698
rect 2492 14644 2548 14646
rect 2436 14634 2548 14644
rect 3388 14642 3444 14654
rect 3388 14590 3390 14642
rect 3442 14590 3444 14642
rect 3388 14588 3444 14590
rect 3220 14532 3444 14588
rect 2884 14364 2940 14374
rect 2828 14362 2940 14364
rect 2828 14310 2886 14362
rect 2938 14310 2940 14362
rect 2828 14298 2940 14310
rect 2404 14140 2668 14150
rect 2460 14084 2508 14140
rect 2564 14084 2612 14140
rect 2404 14074 2668 14084
rect 2660 13916 2716 13926
rect 2324 13692 2380 13702
rect 2044 13580 2100 13618
rect 2324 13598 2380 13636
rect 2044 13514 2100 13524
rect 2156 13578 2212 13590
rect 2156 13526 2158 13578
rect 2210 13526 2212 13578
rect 980 12394 1036 12404
rect 1092 13468 1148 13478
rect 2156 13426 2212 13526
rect 868 9706 924 9716
rect 756 9492 924 9548
rect 404 9436 668 9446
rect 460 9380 508 9436
rect 564 9380 612 9436
rect 404 9370 668 9380
rect 756 9100 812 9110
rect 404 7868 668 7878
rect 460 7812 508 7868
rect 564 7812 612 7868
rect 404 7802 668 7812
rect 404 6300 668 6310
rect 460 6244 508 6300
rect 564 6244 612 6300
rect 404 6234 668 6244
rect 756 6076 812 9044
rect 868 8316 924 9492
rect 1092 8428 1148 13412
rect 1876 13370 2212 13426
rect 2492 13578 2548 13590
rect 2492 13526 2494 13578
rect 2546 13526 2548 13578
rect 1404 13356 1668 13366
rect 1460 13300 1508 13356
rect 1564 13300 1612 13356
rect 1404 13290 1668 13300
rect 1428 13020 1484 13030
rect 1428 12190 1484 12964
rect 1428 12138 1430 12190
rect 1482 12138 1484 12190
rect 1428 12126 1484 12138
rect 1876 12190 1932 13370
rect 2492 13356 2548 13526
rect 2492 13290 2548 13300
rect 2044 13074 2100 13086
rect 2044 13022 2046 13074
rect 2098 13022 2100 13074
rect 2044 13020 2100 13022
rect 1876 12138 1878 12190
rect 1930 12138 1932 12190
rect 1876 12126 1932 12138
rect 1988 12964 2100 13020
rect 1404 11788 1668 11798
rect 1460 11732 1508 11788
rect 1564 11732 1612 11788
rect 1404 11722 1668 11732
rect 1204 11382 1260 11394
rect 1204 11330 1206 11382
rect 1258 11330 1260 11382
rect 1204 9100 1260 11330
rect 1404 10220 1668 10230
rect 1460 10164 1508 10220
rect 1564 10164 1612 10220
rect 1404 10154 1668 10164
rect 1428 9884 1484 9894
rect 1428 9783 1430 9828
rect 1482 9783 1484 9828
rect 1428 9771 1484 9783
rect 1876 9814 1932 9826
rect 1876 9762 1878 9814
rect 1930 9762 1932 9814
rect 1876 9212 1932 9762
rect 1876 9146 1932 9156
rect 1204 9034 1260 9044
rect 1404 8652 1668 8662
rect 1460 8596 1508 8652
rect 1564 8596 1612 8652
rect 1404 8586 1668 8596
rect 1092 8372 1260 8428
rect 868 8260 1148 8316
rect 1092 8250 1148 8260
rect 1092 8204 1094 8250
rect 1146 8204 1148 8250
rect 1092 8138 1148 8148
rect 644 6020 812 6076
rect 980 6748 1036 6758
rect 1204 6748 1260 8372
rect 1988 8316 2044 12964
rect 2660 12924 2716 13860
rect 2828 13804 2884 14298
rect 2828 13710 2884 13748
rect 3052 13746 3108 13758
rect 3052 13694 3054 13746
rect 3106 13694 3108 13746
rect 3052 13356 3108 13694
rect 3052 13290 3108 13300
rect 3052 13132 3108 13142
rect 3220 13132 3276 14532
rect 3780 13804 3836 15316
rect 4228 15302 4284 15314
rect 4228 15260 4230 15302
rect 4282 15260 4284 15302
rect 4228 15194 4284 15204
rect 4340 14710 4396 15428
rect 4676 15372 4732 15382
rect 4676 15270 4678 15316
rect 4730 15270 4732 15316
rect 4340 14698 4452 14710
rect 4340 14646 4398 14698
rect 4450 14646 4452 14698
rect 4340 14644 4452 14646
rect 4396 14634 4452 14644
rect 4676 14364 4732 15270
rect 5012 14710 5068 15540
rect 5236 15484 5292 16324
rect 4956 14698 5068 14710
rect 4956 14646 4958 14698
rect 5010 14646 5068 14698
rect 4956 14644 5068 14646
rect 5124 15428 5292 15484
rect 5348 16156 5404 16166
rect 4956 14634 5012 14644
rect 4844 14588 4900 14598
rect 4844 14494 4900 14532
rect 5124 14538 5180 15428
rect 5348 15270 5404 16100
rect 5292 15258 5404 15270
rect 5292 15206 5294 15258
rect 5346 15206 5404 15258
rect 5292 15204 5404 15206
rect 5292 15194 5348 15204
rect 5796 15148 5852 15158
rect 5404 14924 5668 14934
rect 5460 14868 5508 14924
rect 5564 14868 5612 14924
rect 5404 14858 5668 14868
rect 5124 14486 5126 14538
rect 5178 14486 5180 14538
rect 5124 14474 5180 14486
rect 4676 14298 4732 14308
rect 5180 14364 5236 14374
rect 4404 14140 4668 14150
rect 4460 14084 4508 14140
rect 4564 14084 4612 14140
rect 4404 14074 4668 14084
rect 4564 13916 4620 13926
rect 4788 13916 4844 13926
rect 4620 13860 4732 13916
rect 4564 13850 4620 13860
rect 3780 13738 3836 13748
rect 3444 13580 3500 13618
rect 3444 13514 3500 13524
rect 3668 13580 3724 13590
rect 4004 13580 4060 13590
rect 3668 13578 3836 13580
rect 3668 13526 3670 13578
rect 3722 13526 3836 13578
rect 3668 13524 3836 13526
rect 3668 13514 3724 13524
rect 3404 13356 3668 13366
rect 3460 13300 3508 13356
rect 3564 13300 3612 13356
rect 3404 13290 3668 13300
rect 3052 13130 3276 13132
rect 3052 13078 3054 13130
rect 3106 13078 3276 13130
rect 3052 13076 3276 13078
rect 3052 13066 3108 13076
rect 3780 13020 3836 13524
rect 4004 13486 4060 13524
rect 4452 13580 4508 13590
rect 4452 13486 4508 13524
rect 4676 13468 4732 13860
rect 4788 13822 4844 13860
rect 5180 13802 5236 14308
rect 5180 13750 5182 13802
rect 5234 13750 5236 13802
rect 4900 13580 4956 13590
rect 4676 13412 4844 13468
rect 4620 13244 4676 13254
rect 4620 13130 4676 13188
rect 4620 13078 4622 13130
rect 4674 13078 4676 13130
rect 4620 13066 4676 13078
rect 3780 12954 3836 12964
rect 2660 12868 3052 12924
rect 2404 12572 2668 12582
rect 2460 12516 2508 12572
rect 2564 12516 2612 12572
rect 2404 12506 2668 12516
rect 2404 11004 2668 11014
rect 2460 10948 2508 11004
rect 2564 10948 2612 11004
rect 2404 10938 2668 10948
rect 2404 9436 2668 9446
rect 2460 9380 2508 9436
rect 2564 9380 2612 9436
rect 2404 9370 2668 9380
rect 2660 9212 2772 9222
rect 2716 9210 2772 9212
rect 2716 9158 2718 9210
rect 2770 9158 2772 9210
rect 2716 9156 2772 9158
rect 2660 9146 2772 9156
rect 2660 8988 2716 8998
rect 2660 8894 2716 8932
rect 2380 8876 2436 8886
rect 2380 8782 2436 8820
rect 2828 8876 2884 8886
rect 2828 8782 2884 8820
rect 1708 8260 2044 8316
rect 1708 8258 1820 8260
rect 1708 8206 1710 8258
rect 1762 8206 1820 8258
rect 1708 8194 1820 8206
rect 1404 7084 1668 7094
rect 1460 7028 1508 7084
rect 1564 7028 1612 7084
rect 1404 7018 1668 7028
rect 644 5066 700 6020
rect 644 5014 646 5066
rect 698 5014 700 5066
rect 644 4956 700 5014
rect 644 4890 700 4900
rect 756 5894 812 5906
rect 756 5842 758 5894
rect 810 5842 812 5894
rect 756 5068 812 5842
rect 404 4732 668 4742
rect 460 4676 508 4732
rect 564 4676 612 4732
rect 404 4666 668 4676
rect 756 4350 812 5012
rect 756 4298 758 4350
rect 810 4298 812 4350
rect 756 4286 812 4298
rect 644 3612 700 3622
rect 644 3498 700 3556
rect 644 3446 646 3498
rect 698 3446 700 3498
rect 644 3434 700 3446
rect 980 3500 1036 6692
rect 1092 6692 1260 6748
rect 1092 5964 1148 6692
rect 1092 5908 1204 5964
rect 1148 5906 1204 5908
rect 1148 5854 1150 5906
rect 1202 5854 1204 5906
rect 1148 5842 1204 5854
rect 1404 5516 1668 5526
rect 1460 5460 1508 5516
rect 1564 5460 1612 5516
rect 1404 5450 1668 5460
rect 1316 5178 1372 5190
rect 1316 5126 1318 5178
rect 1370 5126 1372 5178
rect 1204 4956 1260 4966
rect 980 3434 1036 3444
rect 1092 4844 1148 4854
rect 404 3164 668 3174
rect 460 3108 508 3164
rect 564 3108 612 3164
rect 404 3098 668 3108
rect 980 2604 1036 2614
rect 756 2602 1036 2604
rect 756 2550 982 2602
rect 1034 2550 1036 2602
rect 756 2548 1036 2550
rect 404 1596 668 1606
rect 460 1540 508 1596
rect 564 1540 612 1596
rect 404 1530 668 1540
rect -100 1204 252 1260
rect -100 1190 100 1204
rect -100 1110 100 1120
rect 756 1110 812 2548
rect 980 2538 1036 2548
rect -100 1054 812 1110
rect 868 1820 924 1830
rect -100 1044 100 1054
rect -100 964 100 974
rect 868 964 924 1764
rect -100 908 924 964
rect -100 898 100 908
rect -100 812 100 828
rect 1092 812 1148 4788
rect 1204 4350 1260 4900
rect 1204 4298 1206 4350
rect 1258 4298 1260 4350
rect 1204 4286 1260 4298
rect 1316 4172 1372 5126
rect 1204 4116 1372 4172
rect 1204 3724 1260 4116
rect 1404 3948 1668 3958
rect 1460 3892 1508 3948
rect 1564 3892 1612 3948
rect 1404 3882 1668 3892
rect 1316 3724 1372 3734
rect 1204 3722 1484 3724
rect 1204 3670 1318 3722
rect 1370 3670 1484 3722
rect 1204 3668 1484 3670
rect 1316 3658 1372 3668
rect 1316 3500 1372 3510
rect 1316 2714 1372 3444
rect 1428 2828 1484 3668
rect 1764 3612 1820 8194
rect 2404 7868 2668 7878
rect 2460 7812 2508 7868
rect 2564 7812 2612 7868
rect 2404 7802 2668 7812
rect 2404 6300 2668 6310
rect 2460 6244 2508 6300
rect 2564 6244 2612 6300
rect 2404 6234 2668 6244
rect 2996 5852 3052 12868
rect 3388 12908 3444 12918
rect 3388 12814 3444 12852
rect 4284 12850 4340 12862
rect 3668 12796 3724 12806
rect 4284 12798 4286 12850
rect 4338 12798 4340 12850
rect 4284 12796 4340 12798
rect 3668 12794 3948 12796
rect 3668 12742 3670 12794
rect 3722 12742 3948 12794
rect 3668 12740 3948 12742
rect 3668 12730 3724 12740
rect 3404 11788 3668 11798
rect 3460 11732 3508 11788
rect 3564 11732 3612 11788
rect 3404 11722 3668 11732
rect 3668 11382 3724 11394
rect 3668 11330 3670 11382
rect 3722 11330 3724 11382
rect 3668 10780 3724 11330
rect 3668 10714 3724 10724
rect 3892 10554 3948 12740
rect 4060 12738 4116 12750
rect 4060 12686 4062 12738
rect 4114 12686 4116 12738
rect 4284 12730 4340 12740
rect 4060 12236 4116 12686
rect 4404 12572 4668 12582
rect 4460 12516 4508 12572
rect 4564 12516 4612 12572
rect 4404 12506 4668 12516
rect 4060 12170 4116 12180
rect 4564 12236 4620 12246
rect 4228 12166 4284 12178
rect 4228 12114 4230 12166
rect 4282 12114 4284 12166
rect 4116 11382 4172 11394
rect 4116 11330 4118 11382
rect 4170 11330 4172 11382
rect 4116 10780 4172 11330
rect 4228 11004 4284 12114
rect 4564 11228 4620 12180
rect 4676 12166 4732 12178
rect 4676 12124 4678 12166
rect 4730 12124 4732 12166
rect 4676 12058 4732 12068
rect 4788 11562 4844 13412
rect 4788 11510 4790 11562
rect 4842 11510 4844 11562
rect 4788 11498 4844 11510
rect 4900 13018 4956 13524
rect 5180 13468 5236 13750
rect 4900 12966 4902 13018
rect 4954 12966 4956 13018
rect 4900 12908 4956 12966
rect 4900 11350 4956 12852
rect 5012 13412 5236 13468
rect 5012 12124 5068 13412
rect 5404 13356 5668 13366
rect 5460 13300 5508 13356
rect 5564 13300 5612 13356
rect 5404 13290 5668 13300
rect 5236 13132 5292 13142
rect 5236 13038 5292 13076
rect 5180 12236 5236 12246
rect 5180 12142 5236 12180
rect 5796 12236 5852 15092
rect 5796 12170 5852 12180
rect 5012 11676 5068 12068
rect 5404 11788 5668 11798
rect 5460 11732 5508 11788
rect 5564 11732 5612 11788
rect 5404 11722 5668 11732
rect 5012 11620 5236 11676
rect 5180 11562 5236 11620
rect 5180 11510 5182 11562
rect 5234 11510 5236 11562
rect 4900 11340 5012 11350
rect 4900 11284 4956 11340
rect 4956 11246 5012 11284
rect 4564 11172 4788 11228
rect 4228 10938 4284 10948
rect 4404 11004 4668 11014
rect 4460 10948 4508 11004
rect 4564 10948 4612 11004
rect 4404 10938 4668 10948
rect 4228 10780 4284 10790
rect 4116 10778 4284 10780
rect 4116 10726 4230 10778
rect 4282 10726 4284 10778
rect 4116 10724 4284 10726
rect 4228 10714 4284 10724
rect 4564 10780 4676 10790
rect 4620 10778 4676 10780
rect 4620 10726 4622 10778
rect 4674 10726 4676 10778
rect 4620 10724 4676 10726
rect 4564 10714 4676 10724
rect 4732 10610 4788 11172
rect 3892 10502 3894 10554
rect 3946 10502 3948 10554
rect 3892 10490 3948 10502
rect 4564 10556 4620 10566
rect 3108 10442 3164 10454
rect 3108 10390 3110 10442
rect 3162 10390 3164 10442
rect 3108 9884 3164 10390
rect 3444 10444 3500 10482
rect 4564 10462 4620 10500
rect 4732 10558 4734 10610
rect 4786 10558 4788 10610
rect 3444 10378 3500 10388
rect 4004 10444 4060 10454
rect 3404 10220 3668 10230
rect 3460 10164 3508 10220
rect 3564 10164 3612 10220
rect 3404 10154 3668 10164
rect 3108 9818 3164 9828
rect 3388 9212 3444 9222
rect 3388 9118 3444 9156
rect 3892 9212 3948 9222
rect 3164 9100 3220 9110
rect 3164 9006 3220 9044
rect 3780 8874 3836 8886
rect 3780 8822 3782 8874
rect 3834 8822 3836 8874
rect 3404 8652 3668 8662
rect 3460 8596 3508 8652
rect 3564 8596 3612 8652
rect 3404 8586 3668 8596
rect 3780 7532 3836 8822
rect 3780 7466 3836 7476
rect 3892 7318 3948 9156
rect 4004 9210 4060 10388
rect 4732 9996 4788 10558
rect 5180 10666 5236 11510
rect 5180 10614 5182 10666
rect 5234 10614 5236 10666
rect 5068 9996 5124 10006
rect 4732 9994 5124 9996
rect 4732 9942 5070 9994
rect 5122 9942 5124 9994
rect 4732 9940 5124 9942
rect 5068 9930 5124 9940
rect 5180 9994 5236 10614
rect 5796 11340 5852 11350
rect 5404 10220 5668 10230
rect 5460 10164 5508 10220
rect 5564 10164 5612 10220
rect 5404 10154 5668 10164
rect 5180 9942 5182 9994
rect 5234 9942 5236 9994
rect 4844 9826 4900 9838
rect 4004 9158 4006 9210
rect 4058 9158 4060 9210
rect 4004 9146 4060 9158
rect 4228 9814 4284 9826
rect 4228 9762 4230 9814
rect 4282 9762 4284 9814
rect 4228 8316 4284 9762
rect 4844 9774 4846 9826
rect 4898 9774 4900 9826
rect 4844 9772 4900 9774
rect 5180 9772 5236 9942
rect 4844 9716 5236 9772
rect 4404 9436 4668 9446
rect 4460 9380 4508 9436
rect 4564 9380 4612 9436
rect 4404 9370 4668 9380
rect 4620 9100 4676 9110
rect 4396 9042 4452 9054
rect 4396 8990 4398 9042
rect 4450 8990 4452 9042
rect 4620 9006 4676 9044
rect 4396 8988 4452 8990
rect 4452 8932 4508 8988
rect 4396 8922 4508 8932
rect 4004 8246 4060 8258
rect 4228 8250 4284 8260
rect 4004 8194 4006 8246
rect 4058 8194 4060 8246
rect 4004 7530 4060 8194
rect 4452 8092 4508 8922
rect 4900 8316 4956 8326
rect 4564 8246 4620 8258
rect 4564 8194 4566 8246
rect 4618 8194 4620 8246
rect 4564 8092 4620 8194
rect 4564 8036 4844 8092
rect 4452 8026 4508 8036
rect 4404 7868 4668 7878
rect 4460 7812 4508 7868
rect 4564 7812 4612 7868
rect 4404 7802 4668 7812
rect 4788 7642 4844 8036
rect 4788 7590 4790 7642
rect 4842 7590 4844 7642
rect 4788 7578 4844 7590
rect 4004 7478 4006 7530
rect 4058 7478 4060 7530
rect 4004 7466 4060 7478
rect 4452 7532 4508 7542
rect 4452 7418 4508 7476
rect 3500 7308 3556 7318
rect 3836 7308 3948 7318
rect 3500 7306 3948 7308
rect 3500 7254 3502 7306
rect 3554 7254 3838 7306
rect 3890 7254 3948 7306
rect 3500 7252 3948 7254
rect 4004 7396 4060 7408
rect 4004 7344 4006 7396
rect 4058 7344 4060 7396
rect 4452 7366 4454 7418
rect 4506 7366 4508 7418
rect 4452 7354 4508 7366
rect 4004 7308 4060 7344
rect 3500 7242 3556 7252
rect 3836 7242 3892 7252
rect 4004 7242 4060 7252
rect 3404 7084 3668 7094
rect 3460 7028 3508 7084
rect 3564 7028 3612 7084
rect 3404 7018 3668 7028
rect 4228 6748 4284 6758
rect 4228 6076 4284 6692
rect 4404 6300 4668 6310
rect 4460 6244 4508 6300
rect 4564 6244 4612 6300
rect 4404 6234 4668 6244
rect 4228 6020 4676 6076
rect 4620 5962 4676 6020
rect 4620 5910 4622 5962
rect 4674 5910 4676 5962
rect 2996 5786 3052 5796
rect 3556 5852 3612 5862
rect 3556 5758 3612 5796
rect 3780 5852 3836 5862
rect 3404 5516 3668 5526
rect 3460 5460 3508 5516
rect 3564 5460 3612 5516
rect 3404 5450 3668 5460
rect 3780 5180 3836 5796
rect 4228 5852 4284 5862
rect 4228 5682 4284 5796
rect 4228 5630 4230 5682
rect 4282 5630 4284 5682
rect 4228 5618 4284 5630
rect 4396 5740 4452 5750
rect 4396 5292 4452 5684
rect 4340 5290 4452 5292
rect 4340 5238 4398 5290
rect 4450 5238 4452 5290
rect 4340 5226 4452 5238
rect 4620 5290 4676 5910
rect 4900 5852 4956 8260
rect 5012 8204 5068 9716
rect 5180 9100 5236 9110
rect 5180 9006 5236 9044
rect 5404 8652 5668 8662
rect 5460 8596 5508 8652
rect 5564 8596 5612 8652
rect 5404 8586 5668 8596
rect 5236 8428 5292 8438
rect 5236 8334 5292 8372
rect 5012 7308 5068 8148
rect 5292 8092 5348 8102
rect 5292 7530 5348 8036
rect 5292 7478 5294 7530
rect 5346 7478 5348 7530
rect 5292 7466 5348 7478
rect 5012 7252 5292 7308
rect 4900 5786 4956 5796
rect 5012 6748 5068 6758
rect 4620 5238 4622 5290
rect 4674 5238 4676 5290
rect 3724 5124 3836 5180
rect 4228 5180 4284 5190
rect 3724 5122 3780 5124
rect 3724 5070 3726 5122
rect 3778 5070 3780 5122
rect 4228 5082 4230 5124
rect 4282 5082 4284 5124
rect 4228 5070 4284 5082
rect 3724 5058 3780 5070
rect 4340 4956 4396 5226
rect 4228 4900 4396 4956
rect 4620 5180 4676 5238
rect 4620 4956 4676 5124
rect 4620 4900 4844 4956
rect 2404 4732 2668 4742
rect 2460 4676 2508 4732
rect 2564 4676 2612 4732
rect 2404 4666 2668 4676
rect 4228 4620 4284 4900
rect 4404 4732 4668 4742
rect 4460 4676 4508 4732
rect 4564 4676 4612 4732
rect 4404 4666 4668 4676
rect 4228 4564 4340 4620
rect 4284 4508 4340 4564
rect 4284 4452 4452 4508
rect 3556 4396 3612 4406
rect 3556 4282 3612 4340
rect 4396 4396 4452 4452
rect 3556 4230 3558 4282
rect 3610 4230 3612 4282
rect 3556 4218 3612 4230
rect 4004 4284 4060 4294
rect 4396 4264 4452 4340
rect 4620 4396 4676 4406
rect 4788 4396 4844 4900
rect 4620 4394 4844 4396
rect 4620 4342 4622 4394
rect 4674 4342 4844 4394
rect 4620 4340 4844 4342
rect 4620 4330 4676 4340
rect 3780 4172 3836 4182
rect 3404 3948 3668 3958
rect 3460 3892 3508 3948
rect 3564 3892 3612 3948
rect 3404 3882 3668 3892
rect 3780 3566 3836 4116
rect 1764 3546 1820 3556
rect 3724 3554 3836 3566
rect 3332 3500 3388 3510
rect 3724 3502 3726 3554
rect 3778 3502 3836 3554
rect 3724 3500 3836 3502
rect 3724 3490 3780 3500
rect 3332 3388 3388 3444
rect 3108 3332 3388 3388
rect 2404 3164 2668 3174
rect 2460 3108 2508 3164
rect 2564 3108 2612 3164
rect 2404 3098 2668 3108
rect 2940 2940 2996 2950
rect 1428 2762 1484 2772
rect 1764 2828 1820 2838
rect 1316 2662 1318 2714
rect 1370 2662 1372 2714
rect 1316 2650 1372 2662
rect 1764 2714 1820 2772
rect 1764 2662 1766 2714
rect 1818 2662 1820 2714
rect 1764 2650 1820 2662
rect 2324 2828 2380 2838
rect 2940 2828 2996 2884
rect 2100 2604 2156 2614
rect 2100 2602 2268 2604
rect 2100 2550 2102 2602
rect 2154 2550 2268 2602
rect 2100 2548 2268 2550
rect 2100 2538 2156 2548
rect 1404 2380 1668 2390
rect 1460 2324 1508 2380
rect 1564 2324 1612 2380
rect 1404 2314 1668 2324
rect 1764 2156 1820 2166
rect 1764 2062 1820 2100
rect 1428 1820 1484 1830
rect 1428 1726 1484 1764
rect -100 756 1148 812
rect 1404 812 1668 822
rect 1460 756 1508 812
rect 1564 756 1612 812
rect -100 752 100 756
rect 1404 746 1668 756
rect 2212 -200 2268 2548
rect 2324 2166 2380 2772
rect 2436 2826 2996 2828
rect 2436 2774 2942 2826
rect 2994 2774 2996 2826
rect 2436 2772 2996 2774
rect 2436 2714 2492 2772
rect 2940 2762 2996 2772
rect 2436 2662 2438 2714
rect 2490 2662 2492 2714
rect 2436 2650 2492 2662
rect 2548 2604 2604 2614
rect 2324 2154 2436 2166
rect 2324 2102 2382 2154
rect 2434 2102 2436 2154
rect 2324 2100 2436 2102
rect 2380 2090 2436 2100
rect 2548 1820 2604 2548
rect 2772 2604 2828 2614
rect 2772 2510 2828 2548
rect 2548 1764 2828 1820
rect 2404 1596 2668 1606
rect 2460 1540 2508 1596
rect 2564 1540 2612 1596
rect 2404 1530 2668 1540
rect 2772 1372 2828 1764
rect 2660 1316 2828 1372
rect 2660 -200 2716 1316
rect 3108 -200 3164 3332
rect 4004 2940 4060 4228
rect 4228 4172 4284 4182
rect 4228 4114 4284 4116
rect 4228 4062 4230 4114
rect 4282 4062 4284 4114
rect 4228 4050 4284 4062
rect 4788 3724 4844 4340
rect 5012 4060 5068 6692
rect 5236 6646 5292 7252
rect 5404 7084 5668 7094
rect 5460 7028 5508 7084
rect 5564 7028 5612 7084
rect 5404 7018 5668 7028
rect 5180 6634 5292 6646
rect 5180 6582 5182 6634
rect 5234 6582 5292 6634
rect 5180 6580 5292 6582
rect 5180 6300 5236 6580
rect 5124 6244 5236 6300
rect 5124 4284 5180 6244
rect 5404 5516 5668 5526
rect 5460 5460 5508 5516
rect 5564 5460 5612 5516
rect 5404 5450 5668 5460
rect 5796 4844 5852 11284
rect 5796 4778 5852 4788
rect 5124 4218 5180 4228
rect 5012 4004 5292 4060
rect 4228 3722 4844 3724
rect 4228 3670 4790 3722
rect 4842 3670 4844 3722
rect 4228 3668 4844 3670
rect 4228 3566 4284 3668
rect 4228 3514 4230 3566
rect 4282 3514 4284 3566
rect 4228 3502 4284 3514
rect 4788 3612 4844 3668
rect 5068 3612 5124 3622
rect 4788 3610 5124 3612
rect 4788 3558 5070 3610
rect 5122 3558 5124 3610
rect 4788 3556 5124 3558
rect 4452 3500 4508 3510
rect 4452 3406 4508 3444
rect 4404 3164 4668 3174
rect 4460 3108 4508 3164
rect 4564 3108 4612 3164
rect 4404 3098 4668 3108
rect 4004 2874 4060 2884
rect 4788 2838 4844 3556
rect 5068 3546 5124 3556
rect 4396 2828 4452 2838
rect 3332 2716 3388 2754
rect 4396 2734 4452 2772
rect 4732 2826 4844 2838
rect 4732 2774 4734 2826
rect 4786 2774 4844 2826
rect 4732 2772 4844 2774
rect 4732 2762 4788 2772
rect 3332 2650 3388 2660
rect 3668 2716 3724 2726
rect 3668 2622 3724 2660
rect 3780 2604 3836 2614
rect 3404 2380 3668 2390
rect 3460 2324 3508 2380
rect 3564 2324 3612 2380
rect 3404 2314 3668 2324
rect 3404 812 3668 822
rect 3460 756 3508 812
rect 3564 756 3612 812
rect 3404 746 3668 756
rect 3780 588 3836 2548
rect 5236 2156 5292 4004
rect 5404 3948 5668 3958
rect 5460 3892 5508 3948
rect 5564 3892 5612 3948
rect 5404 3882 5668 3892
rect 5908 2716 5964 16996
rect 5908 2650 5964 2660
rect 5404 2380 5668 2390
rect 5460 2324 5508 2380
rect 5564 2324 5612 2380
rect 5404 2314 5668 2324
rect 5236 2090 5292 2100
rect 4404 1596 4668 1606
rect 4460 1540 4508 1596
rect 4564 1540 4612 1596
rect 4404 1530 4668 1540
rect 5404 812 5668 822
rect 5460 756 5508 812
rect 5564 756 5612 812
rect 5404 746 5668 756
rect 3556 532 3836 588
rect 3556 -200 3612 532
<< via2 >>
rect 404 32954 460 32956
rect 404 32902 406 32954
rect 406 32902 458 32954
rect 458 32902 460 32954
rect 404 32900 460 32902
rect 508 32954 564 32956
rect 508 32902 510 32954
rect 510 32902 562 32954
rect 562 32902 564 32954
rect 508 32900 564 32902
rect 612 32954 668 32956
rect 612 32902 614 32954
rect 614 32902 666 32954
rect 666 32902 668 32954
rect 612 32900 668 32902
rect 1404 33738 1460 33740
rect 1404 33686 1406 33738
rect 1406 33686 1458 33738
rect 1458 33686 1460 33738
rect 1404 33684 1460 33686
rect 1508 33738 1564 33740
rect 1508 33686 1510 33738
rect 1510 33686 1562 33738
rect 1562 33686 1564 33738
rect 1508 33684 1564 33686
rect 1612 33738 1668 33740
rect 1612 33686 1614 33738
rect 1614 33686 1666 33738
rect 1666 33686 1668 33738
rect 1612 33684 1668 33686
rect 2404 32954 2460 32956
rect 2404 32902 2406 32954
rect 2406 32902 2458 32954
rect 2458 32902 2460 32954
rect 2404 32900 2460 32902
rect 2508 32954 2564 32956
rect 2508 32902 2510 32954
rect 2510 32902 2562 32954
rect 2562 32902 2564 32954
rect 2508 32900 2564 32902
rect 2612 32954 2668 32956
rect 2612 32902 2614 32954
rect 2614 32902 2666 32954
rect 2666 32902 2668 32954
rect 2612 32900 2668 32902
rect 1404 32170 1460 32172
rect 1404 32118 1406 32170
rect 1406 32118 1458 32170
rect 1458 32118 1460 32170
rect 1404 32116 1460 32118
rect 1508 32170 1564 32172
rect 1508 32118 1510 32170
rect 1510 32118 1562 32170
rect 1562 32118 1564 32170
rect 1508 32116 1564 32118
rect 1612 32170 1668 32172
rect 1612 32118 1614 32170
rect 1614 32118 1666 32170
rect 1666 32118 1668 32170
rect 1612 32116 1668 32118
rect 2772 31892 2828 31948
rect 3404 33738 3460 33740
rect 3404 33686 3406 33738
rect 3406 33686 3458 33738
rect 3458 33686 3460 33738
rect 3404 33684 3460 33686
rect 3508 33738 3564 33740
rect 3508 33686 3510 33738
rect 3510 33686 3562 33738
rect 3562 33686 3564 33738
rect 3508 33684 3564 33686
rect 3612 33738 3668 33740
rect 3612 33686 3614 33738
rect 3614 33686 3666 33738
rect 3666 33686 3668 33738
rect 3612 33684 3668 33686
rect 4004 33236 4060 33292
rect 4620 33290 4676 33292
rect 4620 33238 4622 33290
rect 4622 33238 4674 33290
rect 4674 33238 4676 33290
rect 4620 33236 4676 33238
rect 4404 32954 4460 32956
rect 4404 32902 4406 32954
rect 4406 32902 4458 32954
rect 4458 32902 4460 32954
rect 4404 32900 4460 32902
rect 4508 32954 4564 32956
rect 4508 32902 4510 32954
rect 4510 32902 4562 32954
rect 4562 32902 4564 32954
rect 4508 32900 4564 32902
rect 4612 32954 4668 32956
rect 4612 32902 4614 32954
rect 4614 32902 4666 32954
rect 4666 32902 4668 32954
rect 4612 32900 4668 32902
rect 3388 32394 3444 32396
rect 3388 32342 3390 32394
rect 3390 32342 3442 32394
rect 3442 32342 3444 32394
rect 3388 32340 3444 32342
rect 3404 32170 3460 32172
rect 3404 32118 3406 32170
rect 3406 32118 3458 32170
rect 3458 32118 3460 32170
rect 3404 32116 3460 32118
rect 3508 32170 3564 32172
rect 3508 32118 3510 32170
rect 3510 32118 3562 32170
rect 3562 32118 3564 32170
rect 3508 32116 3564 32118
rect 3612 32170 3668 32172
rect 3612 32118 3614 32170
rect 3614 32118 3666 32170
rect 3666 32118 3668 32170
rect 3612 32116 3668 32118
rect 3220 32004 3276 32060
rect 404 31386 460 31388
rect 404 31334 406 31386
rect 406 31334 458 31386
rect 458 31334 460 31386
rect 404 31332 460 31334
rect 508 31386 564 31388
rect 508 31334 510 31386
rect 510 31334 562 31386
rect 562 31334 564 31386
rect 508 31332 564 31334
rect 612 31386 668 31388
rect 612 31334 614 31386
rect 614 31334 666 31386
rect 666 31334 668 31386
rect 612 31332 668 31334
rect 756 31108 812 31164
rect 756 30146 758 30156
rect 758 30146 810 30156
rect 810 30146 812 30156
rect 756 30100 812 30146
rect 2404 31386 2460 31388
rect 2404 31334 2406 31386
rect 2406 31334 2458 31386
rect 2458 31334 2460 31386
rect 2404 31332 2460 31334
rect 2508 31386 2564 31388
rect 2508 31334 2510 31386
rect 2510 31334 2562 31386
rect 2562 31334 2564 31386
rect 2508 31332 2564 31334
rect 2612 31386 2668 31388
rect 2612 31334 2614 31386
rect 2614 31334 2666 31386
rect 2666 31334 2668 31386
rect 2612 31332 2668 31334
rect 1404 30602 1460 30604
rect 1404 30550 1406 30602
rect 1406 30550 1458 30602
rect 1458 30550 1460 30602
rect 1404 30548 1460 30550
rect 1508 30602 1564 30604
rect 1508 30550 1510 30602
rect 1510 30550 1562 30602
rect 1562 30550 1564 30602
rect 1508 30548 1564 30550
rect 1612 30602 1668 30604
rect 1612 30550 1614 30602
rect 1614 30550 1666 30602
rect 1666 30550 1668 30602
rect 1612 30548 1668 30550
rect 404 29818 460 29820
rect 404 29766 406 29818
rect 406 29766 458 29818
rect 458 29766 460 29818
rect 404 29764 460 29766
rect 508 29818 564 29820
rect 508 29766 510 29818
rect 510 29766 562 29818
rect 562 29766 564 29818
rect 508 29764 564 29766
rect 612 29818 668 29820
rect 612 29766 614 29818
rect 614 29766 666 29818
rect 666 29766 668 29818
rect 612 29764 668 29766
rect 196 28420 252 28476
rect 404 28250 460 28252
rect 404 28198 406 28250
rect 406 28198 458 28250
rect 458 28198 460 28250
rect 404 28196 460 28198
rect 508 28250 564 28252
rect 508 28198 510 28250
rect 510 28198 562 28250
rect 562 28198 564 28250
rect 508 28196 564 28198
rect 612 28250 668 28252
rect 612 28198 614 28250
rect 614 28198 666 28250
rect 666 28198 668 28250
rect 612 28196 668 28198
rect 1092 29204 1148 29260
rect 3668 31790 3724 31836
rect 3668 31780 3670 31790
rect 3670 31780 3722 31790
rect 3722 31780 3724 31790
rect 3668 31108 3724 31164
rect 3948 32004 4004 32060
rect 4228 31780 4284 31836
rect 5404 33738 5460 33740
rect 5404 33686 5406 33738
rect 5406 33686 5458 33738
rect 5458 33686 5460 33738
rect 5404 33684 5460 33686
rect 5508 33738 5564 33740
rect 5508 33686 5510 33738
rect 5510 33686 5562 33738
rect 5562 33686 5564 33738
rect 5508 33684 5564 33686
rect 5612 33738 5668 33740
rect 5612 33686 5614 33738
rect 5614 33686 5666 33738
rect 5666 33686 5668 33738
rect 5612 33684 5668 33686
rect 4732 32116 4788 32172
rect 5404 32170 5460 32172
rect 5404 32118 5406 32170
rect 5406 32118 5458 32170
rect 5458 32118 5460 32170
rect 5404 32116 5460 32118
rect 5508 32170 5564 32172
rect 5508 32118 5510 32170
rect 5510 32118 5562 32170
rect 5562 32118 5564 32170
rect 5508 32116 5564 32118
rect 5612 32170 5668 32172
rect 5612 32118 5614 32170
rect 5614 32118 5666 32170
rect 5666 32118 5668 32170
rect 5612 32116 5668 32118
rect 4004 31668 4060 31724
rect 3780 30884 3836 30940
rect 3892 31556 3948 31612
rect 3404 30602 3460 30604
rect 3404 30550 3406 30602
rect 3406 30550 3458 30602
rect 3458 30550 3460 30602
rect 3404 30548 3460 30550
rect 3508 30602 3564 30604
rect 3508 30550 3510 30602
rect 3510 30550 3562 30602
rect 3562 30550 3564 30602
rect 3508 30548 3564 30550
rect 3612 30602 3668 30604
rect 3612 30550 3614 30602
rect 3614 30550 3666 30602
rect 3666 30550 3668 30602
rect 3612 30548 3668 30550
rect 1876 29988 1932 30044
rect 2404 29818 2460 29820
rect 2404 29766 2406 29818
rect 2406 29766 2458 29818
rect 2458 29766 2460 29818
rect 2404 29764 2460 29766
rect 2508 29818 2564 29820
rect 2508 29766 2510 29818
rect 2510 29766 2562 29818
rect 2562 29766 2564 29818
rect 2508 29764 2564 29766
rect 2612 29818 2668 29820
rect 2612 29766 2614 29818
rect 2614 29766 2666 29818
rect 2666 29766 2668 29818
rect 2612 29764 2668 29766
rect 1428 29365 1430 29372
rect 1430 29365 1482 29372
rect 1482 29365 1484 29372
rect 1428 29316 1484 29365
rect 1404 29034 1460 29036
rect 1404 28982 1406 29034
rect 1406 28982 1458 29034
rect 1458 28982 1460 29034
rect 1404 28980 1460 28982
rect 1508 29034 1564 29036
rect 1508 28982 1510 29034
rect 1510 28982 1562 29034
rect 1562 28982 1564 29034
rect 1508 28980 1564 28982
rect 1612 29034 1668 29036
rect 1612 28982 1614 29034
rect 1614 28982 1666 29034
rect 1666 28982 1668 29034
rect 1612 28980 1668 28982
rect 3780 29316 3836 29372
rect 3404 29034 3460 29036
rect 3404 28982 3406 29034
rect 3406 28982 3458 29034
rect 3458 28982 3460 29034
rect 3404 28980 3460 28982
rect 3508 29034 3564 29036
rect 3508 28982 3510 29034
rect 3510 28982 3562 29034
rect 3562 28982 3564 29034
rect 3508 28980 3564 28982
rect 3612 29034 3668 29036
rect 3612 28982 3614 29034
rect 3614 28982 3666 29034
rect 3666 28982 3668 29034
rect 3612 28980 3668 28982
rect 3668 28756 3724 28812
rect 1204 28420 1260 28476
rect 2404 28250 2460 28252
rect 2404 28198 2406 28250
rect 2406 28198 2458 28250
rect 2458 28198 2460 28250
rect 2404 28196 2460 28198
rect 2508 28250 2564 28252
rect 2508 28198 2510 28250
rect 2510 28198 2562 28250
rect 2562 28198 2564 28250
rect 2508 28196 2564 28198
rect 2612 28250 2668 28252
rect 2612 28198 2614 28250
rect 2614 28198 2666 28250
rect 2666 28198 2668 28250
rect 2612 28196 2668 28198
rect 756 26740 812 26796
rect 404 26682 460 26684
rect 404 26630 406 26682
rect 406 26630 458 26682
rect 458 26630 460 26682
rect 404 26628 460 26630
rect 508 26682 564 26684
rect 508 26630 510 26682
rect 510 26630 562 26682
rect 562 26630 564 26682
rect 508 26628 564 26630
rect 612 26682 668 26684
rect 612 26630 614 26682
rect 614 26630 666 26682
rect 666 26630 668 26682
rect 612 26628 668 26630
rect 404 25114 460 25116
rect 404 25062 406 25114
rect 406 25062 458 25114
rect 458 25062 460 25114
rect 404 25060 460 25062
rect 508 25114 564 25116
rect 508 25062 510 25114
rect 510 25062 562 25114
rect 562 25062 564 25114
rect 508 25060 564 25062
rect 612 25114 668 25116
rect 612 25062 614 25114
rect 614 25062 666 25114
rect 666 25062 668 25114
rect 612 25060 668 25062
rect 756 23950 812 23996
rect 756 23940 758 23950
rect 758 23940 810 23950
rect 810 23940 812 23950
rect 404 23546 460 23548
rect 404 23494 406 23546
rect 406 23494 458 23546
rect 458 23494 460 23546
rect 404 23492 460 23494
rect 508 23546 564 23548
rect 508 23494 510 23546
rect 510 23494 562 23546
rect 562 23494 564 23546
rect 508 23492 564 23494
rect 612 23546 668 23548
rect 612 23494 614 23546
rect 614 23494 666 23546
rect 666 23494 668 23546
rect 612 23492 668 23494
rect 404 21978 460 21980
rect 404 21926 406 21978
rect 406 21926 458 21978
rect 458 21926 460 21978
rect 404 21924 460 21926
rect 508 21978 564 21980
rect 508 21926 510 21978
rect 510 21926 562 21978
rect 562 21926 564 21978
rect 508 21924 564 21926
rect 612 21978 668 21980
rect 612 21926 614 21978
rect 614 21926 666 21978
rect 666 21926 668 21978
rect 612 21924 668 21926
rect 756 21588 812 21644
rect 404 20410 460 20412
rect 404 20358 406 20410
rect 406 20358 458 20410
rect 458 20358 460 20410
rect 404 20356 460 20358
rect 508 20410 564 20412
rect 508 20358 510 20410
rect 510 20358 562 20410
rect 562 20358 564 20410
rect 508 20356 564 20358
rect 612 20410 668 20412
rect 612 20358 614 20410
rect 614 20358 666 20410
rect 666 20358 668 20410
rect 612 20356 668 20358
rect 404 18842 460 18844
rect 404 18790 406 18842
rect 406 18790 458 18842
rect 458 18790 460 18842
rect 404 18788 460 18790
rect 508 18842 564 18844
rect 508 18790 510 18842
rect 510 18790 562 18842
rect 562 18790 564 18842
rect 508 18788 564 18790
rect 612 18842 668 18844
rect 612 18790 614 18842
rect 614 18790 666 18842
rect 666 18790 668 18842
rect 612 18788 668 18790
rect 404 17274 460 17276
rect 404 17222 406 17274
rect 406 17222 458 17274
rect 458 17222 460 17274
rect 404 17220 460 17222
rect 508 17274 564 17276
rect 508 17222 510 17274
rect 510 17222 562 17274
rect 562 17222 564 17274
rect 508 17220 564 17222
rect 612 17274 668 17276
rect 612 17222 614 17274
rect 614 17222 666 17274
rect 666 17222 668 17274
rect 612 17220 668 17222
rect 404 15706 460 15708
rect 404 15654 406 15706
rect 406 15654 458 15706
rect 458 15654 460 15706
rect 404 15652 460 15654
rect 508 15706 564 15708
rect 508 15654 510 15706
rect 510 15654 562 15706
rect 562 15654 564 15706
rect 508 15652 564 15654
rect 612 15706 668 15708
rect 612 15654 614 15706
rect 614 15654 666 15706
rect 666 15654 668 15706
rect 612 15652 668 15654
rect 404 14138 460 14140
rect 404 14086 406 14138
rect 406 14086 458 14138
rect 458 14086 460 14138
rect 404 14084 460 14086
rect 508 14138 564 14140
rect 508 14086 510 14138
rect 510 14086 562 14138
rect 562 14086 564 14138
rect 508 14084 564 14086
rect 612 14138 668 14140
rect 612 14086 614 14138
rect 614 14086 666 14138
rect 666 14086 668 14138
rect 612 14084 668 14086
rect 196 13972 252 14028
rect 196 13076 252 13132
rect 84 12404 140 12460
rect 404 12570 460 12572
rect 404 12518 406 12570
rect 406 12518 458 12570
rect 458 12518 460 12570
rect 404 12516 460 12518
rect 508 12570 564 12572
rect 508 12518 510 12570
rect 510 12518 562 12570
rect 562 12518 564 12570
rect 508 12516 564 12518
rect 612 12570 668 12572
rect 612 12518 614 12570
rect 614 12518 666 12570
rect 666 12518 668 12570
rect 612 12516 668 12518
rect 404 11002 460 11004
rect 404 10950 406 11002
rect 406 10950 458 11002
rect 458 10950 460 11002
rect 404 10948 460 10950
rect 508 11002 564 11004
rect 508 10950 510 11002
rect 510 10950 562 11002
rect 562 10950 564 11002
rect 508 10948 564 10950
rect 612 11002 668 11004
rect 612 10950 614 11002
rect 614 10950 666 11002
rect 666 10950 668 11002
rect 612 10948 668 10950
rect 196 9940 252 9996
rect 644 9994 700 9996
rect 644 9942 646 9994
rect 646 9942 698 9994
rect 698 9942 700 9994
rect 644 9940 700 9942
rect 196 9716 252 9772
rect 1764 27748 1820 27804
rect 1404 27466 1460 27468
rect 1404 27414 1406 27466
rect 1406 27414 1458 27466
rect 1458 27414 1460 27466
rect 1404 27412 1460 27414
rect 1508 27466 1564 27468
rect 1508 27414 1510 27466
rect 1510 27414 1562 27466
rect 1562 27414 1564 27466
rect 1508 27412 1564 27414
rect 1612 27466 1668 27468
rect 1612 27414 1614 27466
rect 1614 27414 1666 27466
rect 1666 27414 1668 27466
rect 1612 27412 1668 27414
rect 3444 27748 3500 27804
rect 3404 27466 3460 27468
rect 3404 27414 3406 27466
rect 3406 27414 3458 27466
rect 3458 27414 3460 27466
rect 3404 27412 3460 27414
rect 3508 27466 3564 27468
rect 3508 27414 3510 27466
rect 3510 27414 3562 27466
rect 3562 27414 3564 27466
rect 3508 27412 3564 27414
rect 3612 27466 3668 27468
rect 3612 27414 3614 27466
rect 3614 27414 3666 27466
rect 3666 27414 3668 27466
rect 3612 27412 3668 27414
rect 3668 27188 3724 27244
rect 4004 28756 4060 28812
rect 4340 31668 4396 31724
rect 4508 31722 4564 31724
rect 4508 31670 4510 31722
rect 4510 31670 4562 31722
rect 4562 31670 4564 31722
rect 4508 31668 4564 31670
rect 4788 31610 4844 31612
rect 4788 31558 4790 31610
rect 4790 31558 4842 31610
rect 4842 31558 4844 31610
rect 4788 31556 4844 31558
rect 4404 31386 4460 31388
rect 4404 31334 4406 31386
rect 4406 31334 4458 31386
rect 4458 31334 4460 31386
rect 4404 31332 4460 31334
rect 4508 31386 4564 31388
rect 4508 31334 4510 31386
rect 4510 31334 4562 31386
rect 4562 31334 4564 31386
rect 4508 31332 4564 31334
rect 4612 31386 4668 31388
rect 4612 31334 4614 31386
rect 4614 31334 4666 31386
rect 4666 31334 4668 31386
rect 4612 31332 4668 31334
rect 5124 31834 5180 31836
rect 5124 31782 5126 31834
rect 5126 31782 5178 31834
rect 5178 31782 5180 31834
rect 5124 31780 5180 31782
rect 5236 31668 5292 31724
rect 4116 30100 4172 30156
rect 3892 28420 3948 28476
rect 4004 27972 4060 28028
rect 4732 30938 4788 30940
rect 4732 30886 4734 30938
rect 4734 30886 4786 30938
rect 4786 30886 4788 30938
rect 4732 30884 4788 30886
rect 4900 30884 4956 30940
rect 4564 30324 4620 30380
rect 4340 29988 4396 30044
rect 4620 29988 4676 30044
rect 5460 30996 5516 31052
rect 5348 30884 5404 30940
rect 5404 30602 5460 30604
rect 5404 30550 5406 30602
rect 5406 30550 5458 30602
rect 5458 30550 5460 30602
rect 5404 30548 5460 30550
rect 5508 30602 5564 30604
rect 5508 30550 5510 30602
rect 5510 30550 5562 30602
rect 5562 30550 5564 30602
rect 5508 30548 5564 30550
rect 5612 30602 5668 30604
rect 5612 30550 5614 30602
rect 5614 30550 5666 30602
rect 5666 30550 5668 30602
rect 5612 30548 5668 30550
rect 4404 29818 4460 29820
rect 4404 29766 4406 29818
rect 4406 29766 4458 29818
rect 4458 29766 4460 29818
rect 4404 29764 4460 29766
rect 4508 29818 4564 29820
rect 4508 29766 4510 29818
rect 4510 29766 4562 29818
rect 4562 29766 4564 29818
rect 4508 29764 4564 29766
rect 4612 29818 4668 29820
rect 4612 29766 4614 29818
rect 4614 29766 4666 29818
rect 4666 29766 4668 29818
rect 4612 29764 4668 29766
rect 4900 29652 4956 29708
rect 4676 29204 4732 29260
rect 5012 29204 5068 29260
rect 5180 29258 5236 29260
rect 5180 29206 5182 29258
rect 5182 29206 5234 29258
rect 5234 29206 5236 29258
rect 5180 29204 5236 29206
rect 5796 29092 5852 29148
rect 5404 29034 5460 29036
rect 5404 28982 5406 29034
rect 5406 28982 5458 29034
rect 5458 28982 5460 29034
rect 5404 28980 5460 28982
rect 5508 29034 5564 29036
rect 5508 28982 5510 29034
rect 5510 28982 5562 29034
rect 5562 28982 5564 29034
rect 5508 28980 5564 28982
rect 5612 29034 5668 29036
rect 5612 28982 5614 29034
rect 5614 28982 5666 29034
rect 5666 28982 5668 29034
rect 5612 28980 5668 28982
rect 4404 28250 4460 28252
rect 4404 28198 4406 28250
rect 4406 28198 4458 28250
rect 4458 28198 4460 28250
rect 4404 28196 4460 28198
rect 4508 28250 4564 28252
rect 4508 28198 4510 28250
rect 4510 28198 4562 28250
rect 4562 28198 4564 28250
rect 4508 28196 4564 28198
rect 4612 28250 4668 28252
rect 4612 28198 4614 28250
rect 4614 28198 4666 28250
rect 4666 28198 4668 28250
rect 4612 28196 4668 28198
rect 4228 27188 4284 27244
rect 5236 27860 5292 27916
rect 1092 21476 1148 21532
rect 1204 26740 1260 26796
rect 2404 26682 2460 26684
rect 2404 26630 2406 26682
rect 2406 26630 2458 26682
rect 2458 26630 2460 26682
rect 2404 26628 2460 26630
rect 2508 26682 2564 26684
rect 2508 26630 2510 26682
rect 2510 26630 2562 26682
rect 2562 26630 2564 26682
rect 2508 26628 2564 26630
rect 2612 26682 2668 26684
rect 2612 26630 2614 26682
rect 2614 26630 2666 26682
rect 2666 26630 2668 26682
rect 2612 26628 2668 26630
rect 3332 26292 3388 26348
rect 3780 26628 3836 26684
rect 3780 26292 3836 26348
rect 3780 26122 3836 26124
rect 3780 26070 3782 26122
rect 3782 26070 3834 26122
rect 3834 26070 3836 26122
rect 3780 26068 3836 26070
rect 1404 25898 1460 25900
rect 1404 25846 1406 25898
rect 1406 25846 1458 25898
rect 1458 25846 1460 25898
rect 1404 25844 1460 25846
rect 1508 25898 1564 25900
rect 1508 25846 1510 25898
rect 1510 25846 1562 25898
rect 1562 25846 1564 25898
rect 1508 25844 1564 25846
rect 1612 25898 1668 25900
rect 1612 25846 1614 25898
rect 1614 25846 1666 25898
rect 1666 25846 1668 25898
rect 1612 25844 1668 25846
rect 3404 25898 3460 25900
rect 3404 25846 3406 25898
rect 3406 25846 3458 25898
rect 3458 25846 3460 25898
rect 3404 25844 3460 25846
rect 3508 25898 3564 25900
rect 3508 25846 3510 25898
rect 3510 25846 3562 25898
rect 3562 25846 3564 25898
rect 3508 25844 3564 25846
rect 3612 25898 3668 25900
rect 3612 25846 3614 25898
rect 3614 25846 3666 25898
rect 3666 25846 3668 25898
rect 3612 25844 3668 25846
rect 2404 25114 2460 25116
rect 2404 25062 2406 25114
rect 2406 25062 2458 25114
rect 2458 25062 2460 25114
rect 2404 25060 2460 25062
rect 2508 25114 2564 25116
rect 2508 25062 2510 25114
rect 2510 25062 2562 25114
rect 2562 25062 2564 25114
rect 2508 25060 2564 25062
rect 2612 25114 2668 25116
rect 2612 25062 2614 25114
rect 2614 25062 2666 25114
rect 2666 25062 2668 25114
rect 2612 25060 2668 25062
rect 3780 25060 3836 25116
rect 1404 24330 1460 24332
rect 1404 24278 1406 24330
rect 1406 24278 1458 24330
rect 1458 24278 1460 24330
rect 1404 24276 1460 24278
rect 1508 24330 1564 24332
rect 1508 24278 1510 24330
rect 1510 24278 1562 24330
rect 1562 24278 1564 24330
rect 1508 24276 1564 24278
rect 1612 24330 1668 24332
rect 1612 24278 1614 24330
rect 1614 24278 1666 24330
rect 1666 24278 1668 24330
rect 1612 24276 1668 24278
rect 3404 24330 3460 24332
rect 3404 24278 3406 24330
rect 3406 24278 3458 24330
rect 3458 24278 3460 24330
rect 3404 24276 3460 24278
rect 3508 24330 3564 24332
rect 3508 24278 3510 24330
rect 3510 24278 3562 24330
rect 3562 24278 3564 24330
rect 3508 24276 3564 24278
rect 3612 24330 3668 24332
rect 3612 24278 3614 24330
rect 3614 24278 3666 24330
rect 3666 24278 3668 24330
rect 3612 24276 3668 24278
rect 2404 23546 2460 23548
rect 2404 23494 2406 23546
rect 2406 23494 2458 23546
rect 2458 23494 2460 23546
rect 2404 23492 2460 23494
rect 2508 23546 2564 23548
rect 2508 23494 2510 23546
rect 2510 23494 2562 23546
rect 2562 23494 2564 23546
rect 2508 23492 2564 23494
rect 2612 23546 2668 23548
rect 2612 23494 2614 23546
rect 2614 23494 2666 23546
rect 2666 23494 2668 23546
rect 2612 23492 2668 23494
rect 2884 23268 2940 23324
rect 1404 22762 1460 22764
rect 1404 22710 1406 22762
rect 1406 22710 1458 22762
rect 1458 22710 1460 22762
rect 1404 22708 1460 22710
rect 1508 22762 1564 22764
rect 1508 22710 1510 22762
rect 1510 22710 1562 22762
rect 1562 22710 1564 22762
rect 1508 22708 1564 22710
rect 1612 22762 1668 22764
rect 1612 22710 1614 22762
rect 1614 22710 1666 22762
rect 1666 22710 1668 22762
rect 1612 22708 1668 22710
rect 1932 22148 1988 22204
rect 1428 21364 1484 21420
rect 1404 21194 1460 21196
rect 1404 21142 1406 21194
rect 1406 21142 1458 21194
rect 1458 21142 1460 21194
rect 1404 21140 1460 21142
rect 1508 21194 1564 21196
rect 1508 21142 1510 21194
rect 1510 21142 1562 21194
rect 1562 21142 1564 21194
rect 1508 21140 1564 21142
rect 1612 21194 1668 21196
rect 1612 21142 1614 21194
rect 1614 21142 1666 21194
rect 1666 21142 1668 21194
rect 1612 21140 1668 21142
rect 1404 19626 1460 19628
rect 1404 19574 1406 19626
rect 1406 19574 1458 19626
rect 1458 19574 1460 19626
rect 1404 19572 1460 19574
rect 1508 19626 1564 19628
rect 1508 19574 1510 19626
rect 1510 19574 1562 19626
rect 1562 19574 1564 19626
rect 1508 19572 1564 19574
rect 1612 19626 1668 19628
rect 1612 19574 1614 19626
rect 1614 19574 1666 19626
rect 1666 19574 1668 19626
rect 1612 19572 1668 19574
rect 2268 22314 2324 22316
rect 2268 22262 2270 22314
rect 2270 22262 2322 22314
rect 2322 22262 2324 22314
rect 2268 22260 2324 22262
rect 2716 22426 2772 22428
rect 2716 22374 2718 22426
rect 2718 22374 2770 22426
rect 2770 22374 2772 22426
rect 2716 22372 2772 22374
rect 2404 21978 2460 21980
rect 2404 21926 2406 21978
rect 2406 21926 2458 21978
rect 2458 21926 2460 21978
rect 2404 21924 2460 21926
rect 2508 21978 2564 21980
rect 2508 21926 2510 21978
rect 2510 21926 2562 21978
rect 2562 21926 2564 21978
rect 2508 21924 2564 21926
rect 2612 21978 2668 21980
rect 2612 21926 2614 21978
rect 2614 21926 2666 21978
rect 2666 21926 2668 21978
rect 2612 21924 2668 21926
rect 4116 26628 4172 26684
rect 5124 27748 5180 27804
rect 5796 27636 5852 27692
rect 5404 27466 5460 27468
rect 4788 27076 4844 27132
rect 4900 27188 4956 27244
rect 5124 27076 5180 27132
rect 5404 27414 5406 27466
rect 5406 27414 5458 27466
rect 5458 27414 5460 27466
rect 5404 27412 5460 27414
rect 5508 27466 5564 27468
rect 5508 27414 5510 27466
rect 5510 27414 5562 27466
rect 5562 27414 5564 27466
rect 5508 27412 5564 27414
rect 5612 27466 5668 27468
rect 5612 27414 5614 27466
rect 5614 27414 5666 27466
rect 5666 27414 5668 27466
rect 5612 27412 5668 27414
rect 4404 26682 4460 26684
rect 4404 26630 4406 26682
rect 4406 26630 4458 26682
rect 4458 26630 4460 26682
rect 4404 26628 4460 26630
rect 4508 26682 4564 26684
rect 4508 26630 4510 26682
rect 4510 26630 4562 26682
rect 4562 26630 4564 26682
rect 4508 26628 4564 26630
rect 4612 26682 4668 26684
rect 4612 26630 4614 26682
rect 4614 26630 4666 26682
rect 4666 26630 4668 26682
rect 4612 26628 4668 26630
rect 4900 26852 4956 26908
rect 4676 26404 4732 26460
rect 4396 26346 4452 26348
rect 4396 26294 4398 26346
rect 4398 26294 4450 26346
rect 4450 26294 4452 26346
rect 4396 26292 4452 26294
rect 4508 26180 4564 26236
rect 4340 26068 4396 26124
rect 4172 25956 4228 26012
rect 4340 25844 4396 25900
rect 4060 25562 4116 25564
rect 4060 25510 4062 25562
rect 4062 25510 4114 25562
rect 4114 25510 4116 25562
rect 4060 25508 4116 25510
rect 4508 25508 4564 25564
rect 4788 26346 4844 26348
rect 4788 26294 4790 26346
rect 4790 26294 4842 26346
rect 4842 26294 4844 26346
rect 4788 26292 4844 26294
rect 5012 26068 5068 26124
rect 4228 25060 4284 25116
rect 4404 25114 4460 25116
rect 4404 25062 4406 25114
rect 4406 25062 4458 25114
rect 4458 25062 4460 25114
rect 4404 25060 4460 25062
rect 4508 25114 4564 25116
rect 4508 25062 4510 25114
rect 4510 25062 4562 25114
rect 4562 25062 4564 25114
rect 4508 25060 4564 25062
rect 4612 25114 4668 25116
rect 4612 25062 4614 25114
rect 4614 25062 4666 25114
rect 4666 25062 4668 25114
rect 4612 25060 4668 25062
rect 3892 23940 3948 23996
rect 3404 22762 3460 22764
rect 3404 22710 3406 22762
rect 3406 22710 3458 22762
rect 3458 22710 3460 22762
rect 3404 22708 3460 22710
rect 3508 22762 3564 22764
rect 3508 22710 3510 22762
rect 3510 22710 3562 22762
rect 3562 22710 3564 22762
rect 3508 22708 3564 22710
rect 3612 22762 3668 22764
rect 3612 22710 3614 22762
rect 3614 22710 3666 22762
rect 3666 22710 3668 22762
rect 3612 22708 3668 22710
rect 3724 22484 3780 22540
rect 4004 23044 4060 23100
rect 4116 23828 4172 23884
rect 4620 23882 4676 23884
rect 4620 23830 4622 23882
rect 4622 23830 4674 23882
rect 4674 23830 4676 23882
rect 4620 23828 4676 23830
rect 3892 22372 3948 22428
rect 4004 22708 4060 22764
rect 3108 22148 3164 22204
rect 4404 23546 4460 23548
rect 4404 23494 4406 23546
rect 4406 23494 4458 23546
rect 4458 23494 4460 23546
rect 4404 23492 4460 23494
rect 4508 23546 4564 23548
rect 4508 23494 4510 23546
rect 4510 23494 4562 23546
rect 4562 23494 4564 23546
rect 4508 23492 4564 23494
rect 4612 23546 4668 23548
rect 4612 23494 4614 23546
rect 4614 23494 4666 23546
rect 4666 23494 4668 23546
rect 4612 23492 4668 23494
rect 5460 26740 5516 26796
rect 5348 26516 5404 26572
rect 5796 26068 5852 26124
rect 5404 25898 5460 25900
rect 5404 25846 5406 25898
rect 5406 25846 5458 25898
rect 5458 25846 5460 25898
rect 5404 25844 5460 25846
rect 5508 25898 5564 25900
rect 5508 25846 5510 25898
rect 5510 25846 5562 25898
rect 5562 25846 5564 25898
rect 5508 25844 5564 25846
rect 5612 25898 5668 25900
rect 5612 25846 5614 25898
rect 5614 25846 5666 25898
rect 5666 25846 5668 25898
rect 5612 25844 5668 25846
rect 5404 24330 5460 24332
rect 5404 24278 5406 24330
rect 5406 24278 5458 24330
rect 5458 24278 5460 24330
rect 5404 24276 5460 24278
rect 5508 24330 5564 24332
rect 5508 24278 5510 24330
rect 5510 24278 5562 24330
rect 5562 24278 5564 24330
rect 5508 24276 5564 24278
rect 5612 24330 5668 24332
rect 5612 24278 5614 24330
rect 5614 24278 5666 24330
rect 5666 24278 5668 24330
rect 5612 24276 5668 24278
rect 4676 23268 4732 23324
rect 4564 23098 4620 23100
rect 4564 23046 4566 23098
rect 4566 23046 4618 23098
rect 4618 23046 4620 23098
rect 4564 23044 4620 23046
rect 4956 23380 5012 23436
rect 5236 23828 5292 23884
rect 4228 22372 4284 22428
rect 1764 19348 1820 19404
rect 2100 20580 2156 20636
rect 1404 18058 1460 18060
rect 1404 18006 1406 18058
rect 1406 18006 1458 18058
rect 1458 18006 1460 18058
rect 1404 18004 1460 18006
rect 1508 18058 1564 18060
rect 1508 18006 1510 18058
rect 1510 18006 1562 18058
rect 1562 18006 1564 18058
rect 1508 18004 1564 18006
rect 1612 18058 1668 18060
rect 1612 18006 1614 18058
rect 1614 18006 1666 18058
rect 1666 18006 1668 18058
rect 1612 18004 1668 18006
rect 2404 20410 2460 20412
rect 2404 20358 2406 20410
rect 2406 20358 2458 20410
rect 2458 20358 2460 20410
rect 2404 20356 2460 20358
rect 2508 20410 2564 20412
rect 2508 20358 2510 20410
rect 2510 20358 2562 20410
rect 2562 20358 2564 20410
rect 2508 20356 2564 20358
rect 2612 20410 2668 20412
rect 2612 20358 2614 20410
rect 2614 20358 2666 20410
rect 2666 20358 2668 20410
rect 2612 20356 2668 20358
rect 3404 21194 3460 21196
rect 3404 21142 3406 21194
rect 3406 21142 3458 21194
rect 3458 21142 3460 21194
rect 3404 21140 3460 21142
rect 3508 21194 3564 21196
rect 3508 21142 3510 21194
rect 3510 21142 3562 21194
rect 3562 21142 3564 21194
rect 3508 21140 3564 21142
rect 3612 21194 3668 21196
rect 3612 21142 3614 21194
rect 3614 21142 3666 21194
rect 3666 21142 3668 21194
rect 3612 21140 3668 21142
rect 2268 19402 2324 19404
rect 2268 19350 2270 19402
rect 2270 19350 2322 19402
rect 2322 19350 2324 19402
rect 2268 19348 2324 19350
rect 2604 19402 2660 19404
rect 2604 19350 2606 19402
rect 2606 19350 2658 19402
rect 2658 19350 2660 19402
rect 2604 19348 2660 19350
rect 3404 19626 3460 19628
rect 3404 19574 3406 19626
rect 3406 19574 3458 19626
rect 3458 19574 3460 19626
rect 3404 19572 3460 19574
rect 3508 19626 3564 19628
rect 3508 19574 3510 19626
rect 3510 19574 3562 19626
rect 3562 19574 3564 19626
rect 3508 19572 3564 19574
rect 3612 19626 3668 19628
rect 3612 19574 3614 19626
rect 3614 19574 3666 19626
rect 3666 19574 3668 19626
rect 3612 19572 3668 19574
rect 2404 18842 2460 18844
rect 2404 18790 2406 18842
rect 2406 18790 2458 18842
rect 2458 18790 2460 18842
rect 2404 18788 2460 18790
rect 2508 18842 2564 18844
rect 2508 18790 2510 18842
rect 2510 18790 2562 18842
rect 2562 18790 2564 18842
rect 2508 18788 2564 18790
rect 2612 18842 2668 18844
rect 2612 18790 2614 18842
rect 2614 18790 2666 18842
rect 2666 18790 2668 18842
rect 2612 18788 2668 18790
rect 3404 18058 3460 18060
rect 3404 18006 3406 18058
rect 3406 18006 3458 18058
rect 3458 18006 3460 18058
rect 3404 18004 3460 18006
rect 3508 18058 3564 18060
rect 3508 18006 3510 18058
rect 3510 18006 3562 18058
rect 3562 18006 3564 18058
rect 3508 18004 3564 18006
rect 3612 18058 3668 18060
rect 3612 18006 3614 18058
rect 3614 18006 3666 18058
rect 3666 18006 3668 18058
rect 3612 18004 3668 18006
rect 4620 22820 4676 22876
rect 4620 22484 4676 22540
rect 4452 22148 4508 22204
rect 4404 21978 4460 21980
rect 4404 21926 4406 21978
rect 4406 21926 4458 21978
rect 4458 21926 4460 21978
rect 4404 21924 4460 21926
rect 4508 21978 4564 21980
rect 4508 21926 4510 21978
rect 4510 21926 4562 21978
rect 4562 21926 4564 21978
rect 4508 21924 4564 21926
rect 4612 21978 4668 21980
rect 4612 21926 4614 21978
rect 4614 21926 4666 21978
rect 4666 21926 4668 21978
rect 4612 21924 4668 21926
rect 5180 22932 5236 22988
rect 5796 23044 5852 23100
rect 5460 22866 5516 22922
rect 5404 22762 5460 22764
rect 5404 22710 5406 22762
rect 5406 22710 5458 22762
rect 5458 22710 5460 22762
rect 5404 22708 5460 22710
rect 5508 22762 5564 22764
rect 5508 22710 5510 22762
rect 5510 22710 5562 22762
rect 5562 22710 5564 22762
rect 5508 22708 5564 22710
rect 5612 22762 5668 22764
rect 5612 22710 5614 22762
rect 5614 22710 5666 22762
rect 5666 22710 5668 22762
rect 5612 22708 5668 22710
rect 5124 21812 5180 21868
rect 3892 21700 3948 21756
rect 4004 21364 4060 21420
rect 4452 21700 4508 21756
rect 4116 21252 4172 21308
rect 4676 21522 4678 21532
rect 4678 21522 4730 21532
rect 4730 21522 4732 21532
rect 4676 21476 4732 21522
rect 4452 21252 4508 21308
rect 4404 20410 4460 20412
rect 4404 20358 4406 20410
rect 4406 20358 4458 20410
rect 4458 20358 4460 20410
rect 4404 20356 4460 20358
rect 4508 20410 4564 20412
rect 4508 20358 4510 20410
rect 4510 20358 4562 20410
rect 4562 20358 4564 20410
rect 4508 20356 4564 20358
rect 4612 20410 4668 20412
rect 4612 20358 4614 20410
rect 4614 20358 4666 20410
rect 4666 20358 4668 20410
rect 4612 20356 4668 20358
rect 4404 18842 4460 18844
rect 4404 18790 4406 18842
rect 4406 18790 4458 18842
rect 4458 18790 4460 18842
rect 4404 18788 4460 18790
rect 4508 18842 4564 18844
rect 4508 18790 4510 18842
rect 4510 18790 4562 18842
rect 4562 18790 4564 18842
rect 4508 18788 4564 18790
rect 4612 18842 4668 18844
rect 4612 18790 4614 18842
rect 4614 18790 4666 18842
rect 4666 18790 4668 18842
rect 4612 18788 4668 18790
rect 3948 18394 4004 18396
rect 3948 18342 3950 18394
rect 3950 18342 4002 18394
rect 4002 18342 4004 18394
rect 3948 18340 4004 18342
rect 4172 18282 4228 18284
rect 4172 18230 4174 18282
rect 4174 18230 4226 18282
rect 4226 18230 4228 18282
rect 4172 18228 4228 18230
rect 3780 18004 3836 18060
rect 4284 17668 4340 17724
rect 4564 17780 4620 17836
rect 2772 17556 2828 17612
rect 2548 17498 2604 17500
rect 2548 17446 2550 17498
rect 2550 17446 2602 17498
rect 2602 17446 2604 17498
rect 2548 17444 2604 17446
rect 2404 17274 2460 17276
rect 2404 17222 2406 17274
rect 2406 17222 2458 17274
rect 2458 17222 2460 17274
rect 2404 17220 2460 17222
rect 2508 17274 2564 17276
rect 2508 17222 2510 17274
rect 2510 17222 2562 17274
rect 2562 17222 2564 17274
rect 2508 17220 2564 17222
rect 2612 17274 2668 17276
rect 2612 17222 2614 17274
rect 2614 17222 2666 17274
rect 2666 17222 2668 17274
rect 2612 17220 2668 17222
rect 3780 17556 3836 17612
rect 3500 16884 3556 16940
rect 4284 17498 4340 17500
rect 4284 17446 4286 17498
rect 4286 17446 4338 17498
rect 4338 17446 4340 17498
rect 4284 17444 4340 17446
rect 4404 17274 4460 17276
rect 4404 17222 4406 17274
rect 4406 17222 4458 17274
rect 4458 17222 4460 17274
rect 4404 17220 4460 17222
rect 4508 17274 4564 17276
rect 4508 17222 4510 17274
rect 4510 17222 4562 17274
rect 4562 17222 4564 17274
rect 4508 17220 4564 17222
rect 4612 17274 4668 17276
rect 4612 17222 4614 17274
rect 4614 17222 4666 17274
rect 4666 17222 4668 17274
rect 4612 17220 4668 17222
rect 4788 17108 4844 17164
rect 3948 16996 4004 17052
rect 4172 17050 4228 17052
rect 4172 16998 4174 17050
rect 4174 16998 4226 17050
rect 4226 16998 4228 17050
rect 4172 16996 4228 16998
rect 4732 16884 4788 16940
rect 2940 16826 2996 16828
rect 2940 16774 2942 16826
rect 2942 16774 2994 16826
rect 2994 16774 2996 16826
rect 2940 16772 2996 16774
rect 3780 16772 3836 16828
rect 4060 16772 4116 16828
rect 1932 16660 1988 16716
rect 1404 16490 1460 16492
rect 1404 16438 1406 16490
rect 1406 16438 1458 16490
rect 1458 16438 1460 16490
rect 1404 16436 1460 16438
rect 1508 16490 1564 16492
rect 1508 16438 1510 16490
rect 1510 16438 1562 16490
rect 1562 16438 1564 16490
rect 1508 16436 1564 16438
rect 1612 16490 1668 16492
rect 1612 16438 1614 16490
rect 1614 16438 1666 16490
rect 1666 16438 1668 16490
rect 1612 16436 1668 16438
rect 2548 16660 2604 16716
rect 3108 16660 3164 16716
rect 2380 16324 2436 16380
rect 2100 16212 2156 16268
rect 2100 16042 2156 16044
rect 2100 15990 2102 16042
rect 2102 15990 2154 16042
rect 2154 15990 2156 16042
rect 2100 15988 2156 15990
rect 1708 15876 1764 15932
rect 2548 16154 2604 16156
rect 2548 16102 2550 16154
rect 2550 16102 2602 16154
rect 2602 16102 2604 16154
rect 2548 16100 2604 16102
rect 2716 15876 2772 15932
rect 2404 15706 2460 15708
rect 2404 15654 2406 15706
rect 2406 15654 2458 15706
rect 2458 15654 2460 15706
rect 2404 15652 2460 15654
rect 2508 15706 2564 15708
rect 2508 15654 2510 15706
rect 2510 15654 2562 15706
rect 2562 15654 2564 15706
rect 2508 15652 2564 15654
rect 2612 15706 2668 15708
rect 2612 15654 2614 15706
rect 2614 15654 2666 15706
rect 2666 15654 2668 15706
rect 2612 15652 2668 15654
rect 1428 15326 1484 15372
rect 1428 15316 1430 15326
rect 1430 15316 1482 15326
rect 1482 15316 1484 15326
rect 3556 16714 3612 16716
rect 3556 16662 3558 16714
rect 3558 16662 3610 16714
rect 3610 16662 3612 16714
rect 3556 16660 3612 16662
rect 3404 16490 3460 16492
rect 3404 16438 3406 16490
rect 3406 16438 3458 16490
rect 3458 16438 3460 16490
rect 3404 16436 3460 16438
rect 3508 16490 3564 16492
rect 3508 16438 3510 16490
rect 3510 16438 3562 16490
rect 3562 16438 3564 16490
rect 3508 16436 3564 16438
rect 3612 16490 3668 16492
rect 3612 16438 3614 16490
rect 3614 16438 3666 16490
rect 3666 16438 3668 16490
rect 3612 16436 3668 16438
rect 3948 16266 4004 16268
rect 3948 16214 3950 16266
rect 3950 16214 4002 16266
rect 4002 16214 4004 16266
rect 3948 16212 4004 16214
rect 5180 21418 5236 21420
rect 5180 21366 5182 21418
rect 5182 21366 5234 21418
rect 5234 21366 5236 21418
rect 5180 21364 5236 21366
rect 5404 21194 5460 21196
rect 5404 21142 5406 21194
rect 5406 21142 5458 21194
rect 5458 21142 5460 21194
rect 5404 21140 5460 21142
rect 5508 21194 5564 21196
rect 5508 21142 5510 21194
rect 5510 21142 5562 21194
rect 5562 21142 5564 21194
rect 5508 21140 5564 21142
rect 5612 21194 5668 21196
rect 5612 21142 5614 21194
rect 5614 21142 5666 21194
rect 5666 21142 5668 21194
rect 5612 21140 5668 21142
rect 5236 20634 5292 20636
rect 5236 20582 5238 20634
rect 5238 20582 5290 20634
rect 5290 20582 5292 20634
rect 5236 20580 5292 20582
rect 5796 19684 5852 19740
rect 5404 19626 5460 19628
rect 5404 19574 5406 19626
rect 5406 19574 5458 19626
rect 5458 19574 5460 19626
rect 5404 19572 5460 19574
rect 5508 19626 5564 19628
rect 5508 19574 5510 19626
rect 5510 19574 5562 19626
rect 5562 19574 5564 19626
rect 5508 19572 5564 19574
rect 5612 19626 5668 19628
rect 5612 19574 5614 19626
rect 5614 19574 5666 19626
rect 5666 19574 5668 19626
rect 5612 19572 5668 19574
rect 5012 18900 5068 18956
rect 5012 18340 5068 18396
rect 5348 18452 5404 18508
rect 5180 18282 5236 18284
rect 5180 18230 5182 18282
rect 5182 18230 5234 18282
rect 5234 18230 5236 18282
rect 5180 18228 5236 18230
rect 5404 18058 5460 18060
rect 5404 18006 5406 18058
rect 5406 18006 5458 18058
rect 5458 18006 5460 18058
rect 5404 18004 5460 18006
rect 5508 18058 5564 18060
rect 5508 18006 5510 18058
rect 5510 18006 5562 18058
rect 5562 18006 5564 18058
rect 5508 18004 5564 18006
rect 5612 18058 5668 18060
rect 5612 18006 5614 18058
rect 5614 18006 5666 18058
rect 5666 18006 5668 18058
rect 5612 18004 5668 18006
rect 4900 16772 4956 16828
rect 5124 17668 5180 17724
rect 4732 16660 4788 16716
rect 3388 16100 3444 16156
rect 4452 16324 4508 16380
rect 5348 17444 5404 17500
rect 5684 16996 5740 17052
rect 5404 16490 5460 16492
rect 5404 16438 5406 16490
rect 5406 16438 5458 16490
rect 5458 16438 5460 16490
rect 5404 16436 5460 16438
rect 5508 16490 5564 16492
rect 5508 16438 5510 16490
rect 5510 16438 5562 16490
rect 5562 16438 5564 16490
rect 5508 16436 5564 16438
rect 5612 16490 5668 16492
rect 5612 16438 5614 16490
rect 5614 16438 5666 16490
rect 5666 16438 5668 16490
rect 5612 16436 5668 16438
rect 3388 15876 3444 15932
rect 3220 15316 3276 15372
rect 4676 16212 4732 16268
rect 4788 15988 4844 16044
rect 4956 16042 5012 16044
rect 4956 15990 4958 16042
rect 4958 15990 5010 16042
rect 5010 15990 5012 16042
rect 4956 15988 5012 15990
rect 4404 15706 4460 15708
rect 4404 15654 4406 15706
rect 4406 15654 4458 15706
rect 4458 15654 4460 15706
rect 4404 15652 4460 15654
rect 4508 15706 4564 15708
rect 4508 15654 4510 15706
rect 4510 15654 4562 15706
rect 4562 15654 4564 15706
rect 4508 15652 4564 15654
rect 4612 15706 4668 15708
rect 4612 15654 4614 15706
rect 4614 15654 4666 15706
rect 4666 15654 4668 15706
rect 4612 15652 4668 15654
rect 1404 14922 1460 14924
rect 1404 14870 1406 14922
rect 1406 14870 1458 14922
rect 1458 14870 1460 14922
rect 1404 14868 1460 14870
rect 1508 14922 1564 14924
rect 1508 14870 1510 14922
rect 1510 14870 1562 14922
rect 1562 14870 1564 14922
rect 1508 14868 1564 14870
rect 1612 14922 1668 14924
rect 1612 14870 1614 14922
rect 1614 14870 1666 14922
rect 1666 14870 1668 14922
rect 1612 14868 1668 14870
rect 3404 14922 3460 14924
rect 3404 14870 3406 14922
rect 3406 14870 3458 14922
rect 3458 14870 3460 14922
rect 3404 14868 3460 14870
rect 3508 14922 3564 14924
rect 3508 14870 3510 14922
rect 3510 14870 3562 14922
rect 3562 14870 3564 14922
rect 3508 14868 3564 14870
rect 3612 14922 3668 14924
rect 3612 14870 3614 14922
rect 3614 14870 3666 14922
rect 3666 14870 3668 14922
rect 3612 14868 3668 14870
rect 2156 14698 2212 14700
rect 2156 14646 2158 14698
rect 2158 14646 2210 14698
rect 2210 14646 2212 14698
rect 2156 14644 2212 14646
rect 2436 14644 2492 14700
rect 2404 14138 2460 14140
rect 2404 14086 2406 14138
rect 2406 14086 2458 14138
rect 2458 14086 2460 14138
rect 2404 14084 2460 14086
rect 2508 14138 2564 14140
rect 2508 14086 2510 14138
rect 2510 14086 2562 14138
rect 2562 14086 2564 14138
rect 2508 14084 2564 14086
rect 2612 14138 2668 14140
rect 2612 14086 2614 14138
rect 2614 14086 2666 14138
rect 2666 14086 2668 14138
rect 2612 14084 2668 14086
rect 2660 13860 2716 13916
rect 2324 13690 2380 13692
rect 2324 13638 2326 13690
rect 2326 13638 2378 13690
rect 2378 13638 2380 13690
rect 2324 13636 2380 13638
rect 2044 13578 2100 13580
rect 2044 13526 2046 13578
rect 2046 13526 2098 13578
rect 2098 13526 2100 13578
rect 2044 13524 2100 13526
rect 980 12404 1036 12460
rect 1092 13412 1148 13468
rect 868 9716 924 9772
rect 404 9434 460 9436
rect 404 9382 406 9434
rect 406 9382 458 9434
rect 458 9382 460 9434
rect 404 9380 460 9382
rect 508 9434 564 9436
rect 508 9382 510 9434
rect 510 9382 562 9434
rect 562 9382 564 9434
rect 508 9380 564 9382
rect 612 9434 668 9436
rect 612 9382 614 9434
rect 614 9382 666 9434
rect 666 9382 668 9434
rect 612 9380 668 9382
rect 756 9044 812 9100
rect 404 7866 460 7868
rect 404 7814 406 7866
rect 406 7814 458 7866
rect 458 7814 460 7866
rect 404 7812 460 7814
rect 508 7866 564 7868
rect 508 7814 510 7866
rect 510 7814 562 7866
rect 562 7814 564 7866
rect 508 7812 564 7814
rect 612 7866 668 7868
rect 612 7814 614 7866
rect 614 7814 666 7866
rect 666 7814 668 7866
rect 612 7812 668 7814
rect 404 6298 460 6300
rect 404 6246 406 6298
rect 406 6246 458 6298
rect 458 6246 460 6298
rect 404 6244 460 6246
rect 508 6298 564 6300
rect 508 6246 510 6298
rect 510 6246 562 6298
rect 562 6246 564 6298
rect 508 6244 564 6246
rect 612 6298 668 6300
rect 612 6246 614 6298
rect 614 6246 666 6298
rect 666 6246 668 6298
rect 612 6244 668 6246
rect 1404 13354 1460 13356
rect 1404 13302 1406 13354
rect 1406 13302 1458 13354
rect 1458 13302 1460 13354
rect 1404 13300 1460 13302
rect 1508 13354 1564 13356
rect 1508 13302 1510 13354
rect 1510 13302 1562 13354
rect 1562 13302 1564 13354
rect 1508 13300 1564 13302
rect 1612 13354 1668 13356
rect 1612 13302 1614 13354
rect 1614 13302 1666 13354
rect 1666 13302 1668 13354
rect 1612 13300 1668 13302
rect 1428 12964 1484 13020
rect 2492 13300 2548 13356
rect 1404 11786 1460 11788
rect 1404 11734 1406 11786
rect 1406 11734 1458 11786
rect 1458 11734 1460 11786
rect 1404 11732 1460 11734
rect 1508 11786 1564 11788
rect 1508 11734 1510 11786
rect 1510 11734 1562 11786
rect 1562 11734 1564 11786
rect 1508 11732 1564 11734
rect 1612 11786 1668 11788
rect 1612 11734 1614 11786
rect 1614 11734 1666 11786
rect 1666 11734 1668 11786
rect 1612 11732 1668 11734
rect 1404 10218 1460 10220
rect 1404 10166 1406 10218
rect 1406 10166 1458 10218
rect 1458 10166 1460 10218
rect 1404 10164 1460 10166
rect 1508 10218 1564 10220
rect 1508 10166 1510 10218
rect 1510 10166 1562 10218
rect 1562 10166 1564 10218
rect 1508 10164 1564 10166
rect 1612 10218 1668 10220
rect 1612 10166 1614 10218
rect 1614 10166 1666 10218
rect 1666 10166 1668 10218
rect 1612 10164 1668 10166
rect 1428 9835 1484 9884
rect 1428 9828 1430 9835
rect 1430 9828 1482 9835
rect 1482 9828 1484 9835
rect 1876 9156 1932 9212
rect 1204 9044 1260 9100
rect 1404 8650 1460 8652
rect 1404 8598 1406 8650
rect 1406 8598 1458 8650
rect 1458 8598 1460 8650
rect 1404 8596 1460 8598
rect 1508 8650 1564 8652
rect 1508 8598 1510 8650
rect 1510 8598 1562 8650
rect 1562 8598 1564 8650
rect 1508 8596 1564 8598
rect 1612 8650 1668 8652
rect 1612 8598 1614 8650
rect 1614 8598 1666 8650
rect 1666 8598 1668 8650
rect 1612 8596 1668 8598
rect 1092 8198 1094 8204
rect 1094 8198 1146 8204
rect 1146 8198 1148 8204
rect 1092 8148 1148 8198
rect 2828 13802 2884 13804
rect 2828 13750 2830 13802
rect 2830 13750 2882 13802
rect 2882 13750 2884 13802
rect 2828 13748 2884 13750
rect 3052 13300 3108 13356
rect 4228 15250 4230 15260
rect 4230 15250 4282 15260
rect 4282 15250 4284 15260
rect 4228 15204 4284 15250
rect 4676 15322 4732 15372
rect 4676 15316 4678 15322
rect 4678 15316 4730 15322
rect 4730 15316 4732 15322
rect 5348 16100 5404 16156
rect 4844 14586 4900 14588
rect 4844 14534 4846 14586
rect 4846 14534 4898 14586
rect 4898 14534 4900 14586
rect 4844 14532 4900 14534
rect 5796 15092 5852 15148
rect 5404 14922 5460 14924
rect 5404 14870 5406 14922
rect 5406 14870 5458 14922
rect 5458 14870 5460 14922
rect 5404 14868 5460 14870
rect 5508 14922 5564 14924
rect 5508 14870 5510 14922
rect 5510 14870 5562 14922
rect 5562 14870 5564 14922
rect 5508 14868 5564 14870
rect 5612 14922 5668 14924
rect 5612 14870 5614 14922
rect 5614 14870 5666 14922
rect 5666 14870 5668 14922
rect 5612 14868 5668 14870
rect 4676 14308 4732 14364
rect 5180 14308 5236 14364
rect 4404 14138 4460 14140
rect 4404 14086 4406 14138
rect 4406 14086 4458 14138
rect 4458 14086 4460 14138
rect 4404 14084 4460 14086
rect 4508 14138 4564 14140
rect 4508 14086 4510 14138
rect 4510 14086 4562 14138
rect 4562 14086 4564 14138
rect 4508 14084 4564 14086
rect 4612 14138 4668 14140
rect 4612 14086 4614 14138
rect 4614 14086 4666 14138
rect 4666 14086 4668 14138
rect 4612 14084 4668 14086
rect 4564 13860 4620 13916
rect 3780 13748 3836 13804
rect 3444 13578 3500 13580
rect 3444 13526 3446 13578
rect 3446 13526 3498 13578
rect 3498 13526 3500 13578
rect 3444 13524 3500 13526
rect 3404 13354 3460 13356
rect 3404 13302 3406 13354
rect 3406 13302 3458 13354
rect 3458 13302 3460 13354
rect 3404 13300 3460 13302
rect 3508 13354 3564 13356
rect 3508 13302 3510 13354
rect 3510 13302 3562 13354
rect 3562 13302 3564 13354
rect 3508 13300 3564 13302
rect 3612 13354 3668 13356
rect 3612 13302 3614 13354
rect 3614 13302 3666 13354
rect 3666 13302 3668 13354
rect 3612 13300 3668 13302
rect 4004 13578 4060 13580
rect 4004 13526 4006 13578
rect 4006 13526 4058 13578
rect 4058 13526 4060 13578
rect 4004 13524 4060 13526
rect 4452 13578 4508 13580
rect 4452 13526 4454 13578
rect 4454 13526 4506 13578
rect 4506 13526 4508 13578
rect 4452 13524 4508 13526
rect 4788 13914 4844 13916
rect 4788 13862 4790 13914
rect 4790 13862 4842 13914
rect 4842 13862 4844 13914
rect 4788 13860 4844 13862
rect 4900 13524 4956 13580
rect 4620 13188 4676 13244
rect 3780 12964 3836 13020
rect 2404 12570 2460 12572
rect 2404 12518 2406 12570
rect 2406 12518 2458 12570
rect 2458 12518 2460 12570
rect 2404 12516 2460 12518
rect 2508 12570 2564 12572
rect 2508 12518 2510 12570
rect 2510 12518 2562 12570
rect 2562 12518 2564 12570
rect 2508 12516 2564 12518
rect 2612 12570 2668 12572
rect 2612 12518 2614 12570
rect 2614 12518 2666 12570
rect 2666 12518 2668 12570
rect 2612 12516 2668 12518
rect 2404 11002 2460 11004
rect 2404 10950 2406 11002
rect 2406 10950 2458 11002
rect 2458 10950 2460 11002
rect 2404 10948 2460 10950
rect 2508 11002 2564 11004
rect 2508 10950 2510 11002
rect 2510 10950 2562 11002
rect 2562 10950 2564 11002
rect 2508 10948 2564 10950
rect 2612 11002 2668 11004
rect 2612 10950 2614 11002
rect 2614 10950 2666 11002
rect 2666 10950 2668 11002
rect 2612 10948 2668 10950
rect 2404 9434 2460 9436
rect 2404 9382 2406 9434
rect 2406 9382 2458 9434
rect 2458 9382 2460 9434
rect 2404 9380 2460 9382
rect 2508 9434 2564 9436
rect 2508 9382 2510 9434
rect 2510 9382 2562 9434
rect 2562 9382 2564 9434
rect 2508 9380 2564 9382
rect 2612 9434 2668 9436
rect 2612 9382 2614 9434
rect 2614 9382 2666 9434
rect 2666 9382 2668 9434
rect 2612 9380 2668 9382
rect 2660 9156 2716 9212
rect 2660 8986 2716 8988
rect 2660 8934 2662 8986
rect 2662 8934 2714 8986
rect 2714 8934 2716 8986
rect 2660 8932 2716 8934
rect 2380 8874 2436 8876
rect 2380 8822 2382 8874
rect 2382 8822 2434 8874
rect 2434 8822 2436 8874
rect 2380 8820 2436 8822
rect 2828 8874 2884 8876
rect 2828 8822 2830 8874
rect 2830 8822 2882 8874
rect 2882 8822 2884 8874
rect 2828 8820 2884 8822
rect 1404 7082 1460 7084
rect 1404 7030 1406 7082
rect 1406 7030 1458 7082
rect 1458 7030 1460 7082
rect 1404 7028 1460 7030
rect 1508 7082 1564 7084
rect 1508 7030 1510 7082
rect 1510 7030 1562 7082
rect 1562 7030 1564 7082
rect 1508 7028 1564 7030
rect 1612 7082 1668 7084
rect 1612 7030 1614 7082
rect 1614 7030 1666 7082
rect 1666 7030 1668 7082
rect 1612 7028 1668 7030
rect 980 6692 1036 6748
rect 644 4900 700 4956
rect 756 5012 812 5068
rect 404 4730 460 4732
rect 404 4678 406 4730
rect 406 4678 458 4730
rect 458 4678 460 4730
rect 404 4676 460 4678
rect 508 4730 564 4732
rect 508 4678 510 4730
rect 510 4678 562 4730
rect 562 4678 564 4730
rect 508 4676 564 4678
rect 612 4730 668 4732
rect 612 4678 614 4730
rect 614 4678 666 4730
rect 666 4678 668 4730
rect 612 4676 668 4678
rect 644 3556 700 3612
rect 1404 5514 1460 5516
rect 1404 5462 1406 5514
rect 1406 5462 1458 5514
rect 1458 5462 1460 5514
rect 1404 5460 1460 5462
rect 1508 5514 1564 5516
rect 1508 5462 1510 5514
rect 1510 5462 1562 5514
rect 1562 5462 1564 5514
rect 1508 5460 1564 5462
rect 1612 5514 1668 5516
rect 1612 5462 1614 5514
rect 1614 5462 1666 5514
rect 1666 5462 1668 5514
rect 1612 5460 1668 5462
rect 1204 4900 1260 4956
rect 980 3444 1036 3500
rect 1092 4788 1148 4844
rect 404 3162 460 3164
rect 404 3110 406 3162
rect 406 3110 458 3162
rect 458 3110 460 3162
rect 404 3108 460 3110
rect 508 3162 564 3164
rect 508 3110 510 3162
rect 510 3110 562 3162
rect 562 3110 564 3162
rect 508 3108 564 3110
rect 612 3162 668 3164
rect 612 3110 614 3162
rect 614 3110 666 3162
rect 666 3110 668 3162
rect 612 3108 668 3110
rect 404 1594 460 1596
rect 404 1542 406 1594
rect 406 1542 458 1594
rect 458 1542 460 1594
rect 404 1540 460 1542
rect 508 1594 564 1596
rect 508 1542 510 1594
rect 510 1542 562 1594
rect 562 1542 564 1594
rect 508 1540 564 1542
rect 612 1594 668 1596
rect 612 1542 614 1594
rect 614 1542 666 1594
rect 666 1542 668 1594
rect 612 1540 668 1542
rect 868 1764 924 1820
rect 1404 3946 1460 3948
rect 1404 3894 1406 3946
rect 1406 3894 1458 3946
rect 1458 3894 1460 3946
rect 1404 3892 1460 3894
rect 1508 3946 1564 3948
rect 1508 3894 1510 3946
rect 1510 3894 1562 3946
rect 1562 3894 1564 3946
rect 1508 3892 1564 3894
rect 1612 3946 1668 3948
rect 1612 3894 1614 3946
rect 1614 3894 1666 3946
rect 1666 3894 1668 3946
rect 1612 3892 1668 3894
rect 1316 3444 1372 3500
rect 2404 7866 2460 7868
rect 2404 7814 2406 7866
rect 2406 7814 2458 7866
rect 2458 7814 2460 7866
rect 2404 7812 2460 7814
rect 2508 7866 2564 7868
rect 2508 7814 2510 7866
rect 2510 7814 2562 7866
rect 2562 7814 2564 7866
rect 2508 7812 2564 7814
rect 2612 7866 2668 7868
rect 2612 7814 2614 7866
rect 2614 7814 2666 7866
rect 2666 7814 2668 7866
rect 2612 7812 2668 7814
rect 2404 6298 2460 6300
rect 2404 6246 2406 6298
rect 2406 6246 2458 6298
rect 2458 6246 2460 6298
rect 2404 6244 2460 6246
rect 2508 6298 2564 6300
rect 2508 6246 2510 6298
rect 2510 6246 2562 6298
rect 2562 6246 2564 6298
rect 2508 6244 2564 6246
rect 2612 6298 2668 6300
rect 2612 6246 2614 6298
rect 2614 6246 2666 6298
rect 2666 6246 2668 6298
rect 2612 6244 2668 6246
rect 3388 12906 3444 12908
rect 3388 12854 3390 12906
rect 3390 12854 3442 12906
rect 3442 12854 3444 12906
rect 3388 12852 3444 12854
rect 3404 11786 3460 11788
rect 3404 11734 3406 11786
rect 3406 11734 3458 11786
rect 3458 11734 3460 11786
rect 3404 11732 3460 11734
rect 3508 11786 3564 11788
rect 3508 11734 3510 11786
rect 3510 11734 3562 11786
rect 3562 11734 3564 11786
rect 3508 11732 3564 11734
rect 3612 11786 3668 11788
rect 3612 11734 3614 11786
rect 3614 11734 3666 11786
rect 3666 11734 3668 11786
rect 3612 11732 3668 11734
rect 3668 10724 3724 10780
rect 4284 12740 4340 12796
rect 4404 12570 4460 12572
rect 4404 12518 4406 12570
rect 4406 12518 4458 12570
rect 4458 12518 4460 12570
rect 4404 12516 4460 12518
rect 4508 12570 4564 12572
rect 4508 12518 4510 12570
rect 4510 12518 4562 12570
rect 4562 12518 4564 12570
rect 4508 12516 4564 12518
rect 4612 12570 4668 12572
rect 4612 12518 4614 12570
rect 4614 12518 4666 12570
rect 4666 12518 4668 12570
rect 4612 12516 4668 12518
rect 4060 12180 4116 12236
rect 4564 12180 4620 12236
rect 4676 12114 4678 12124
rect 4678 12114 4730 12124
rect 4730 12114 4732 12124
rect 4676 12068 4732 12114
rect 4900 12852 4956 12908
rect 5404 13354 5460 13356
rect 5404 13302 5406 13354
rect 5406 13302 5458 13354
rect 5458 13302 5460 13354
rect 5404 13300 5460 13302
rect 5508 13354 5564 13356
rect 5508 13302 5510 13354
rect 5510 13302 5562 13354
rect 5562 13302 5564 13354
rect 5508 13300 5564 13302
rect 5612 13354 5668 13356
rect 5612 13302 5614 13354
rect 5614 13302 5666 13354
rect 5666 13302 5668 13354
rect 5612 13300 5668 13302
rect 5236 13130 5292 13132
rect 5236 13078 5238 13130
rect 5238 13078 5290 13130
rect 5290 13078 5292 13130
rect 5236 13076 5292 13078
rect 5180 12234 5236 12236
rect 5180 12182 5182 12234
rect 5182 12182 5234 12234
rect 5234 12182 5236 12234
rect 5180 12180 5236 12182
rect 5796 12180 5852 12236
rect 5012 12068 5068 12124
rect 5404 11786 5460 11788
rect 5404 11734 5406 11786
rect 5406 11734 5458 11786
rect 5458 11734 5460 11786
rect 5404 11732 5460 11734
rect 5508 11786 5564 11788
rect 5508 11734 5510 11786
rect 5510 11734 5562 11786
rect 5562 11734 5564 11786
rect 5508 11732 5564 11734
rect 5612 11786 5668 11788
rect 5612 11734 5614 11786
rect 5614 11734 5666 11786
rect 5666 11734 5668 11786
rect 5612 11732 5668 11734
rect 4956 11338 5012 11340
rect 4956 11286 4958 11338
rect 4958 11286 5010 11338
rect 5010 11286 5012 11338
rect 4956 11284 5012 11286
rect 4228 10948 4284 11004
rect 4404 11002 4460 11004
rect 4404 10950 4406 11002
rect 4406 10950 4458 11002
rect 4458 10950 4460 11002
rect 4404 10948 4460 10950
rect 4508 11002 4564 11004
rect 4508 10950 4510 11002
rect 4510 10950 4562 11002
rect 4562 10950 4564 11002
rect 4508 10948 4564 10950
rect 4612 11002 4668 11004
rect 4612 10950 4614 11002
rect 4614 10950 4666 11002
rect 4666 10950 4668 11002
rect 4612 10948 4668 10950
rect 4564 10724 4620 10780
rect 4564 10554 4620 10556
rect 4564 10502 4566 10554
rect 4566 10502 4618 10554
rect 4618 10502 4620 10554
rect 4564 10500 4620 10502
rect 3444 10442 3500 10444
rect 3444 10390 3446 10442
rect 3446 10390 3498 10442
rect 3498 10390 3500 10442
rect 3444 10388 3500 10390
rect 4004 10388 4060 10444
rect 3404 10218 3460 10220
rect 3404 10166 3406 10218
rect 3406 10166 3458 10218
rect 3458 10166 3460 10218
rect 3404 10164 3460 10166
rect 3508 10218 3564 10220
rect 3508 10166 3510 10218
rect 3510 10166 3562 10218
rect 3562 10166 3564 10218
rect 3508 10164 3564 10166
rect 3612 10218 3668 10220
rect 3612 10166 3614 10218
rect 3614 10166 3666 10218
rect 3666 10166 3668 10218
rect 3612 10164 3668 10166
rect 3108 9828 3164 9884
rect 3388 9210 3444 9212
rect 3388 9158 3390 9210
rect 3390 9158 3442 9210
rect 3442 9158 3444 9210
rect 3388 9156 3444 9158
rect 3892 9156 3948 9212
rect 3164 9098 3220 9100
rect 3164 9046 3166 9098
rect 3166 9046 3218 9098
rect 3218 9046 3220 9098
rect 3164 9044 3220 9046
rect 3404 8650 3460 8652
rect 3404 8598 3406 8650
rect 3406 8598 3458 8650
rect 3458 8598 3460 8650
rect 3404 8596 3460 8598
rect 3508 8650 3564 8652
rect 3508 8598 3510 8650
rect 3510 8598 3562 8650
rect 3562 8598 3564 8650
rect 3508 8596 3564 8598
rect 3612 8650 3668 8652
rect 3612 8598 3614 8650
rect 3614 8598 3666 8650
rect 3666 8598 3668 8650
rect 3612 8596 3668 8598
rect 3780 7476 3836 7532
rect 5796 11284 5852 11340
rect 5404 10218 5460 10220
rect 5404 10166 5406 10218
rect 5406 10166 5458 10218
rect 5458 10166 5460 10218
rect 5404 10164 5460 10166
rect 5508 10218 5564 10220
rect 5508 10166 5510 10218
rect 5510 10166 5562 10218
rect 5562 10166 5564 10218
rect 5508 10164 5564 10166
rect 5612 10218 5668 10220
rect 5612 10166 5614 10218
rect 5614 10166 5666 10218
rect 5666 10166 5668 10218
rect 5612 10164 5668 10166
rect 4404 9434 4460 9436
rect 4404 9382 4406 9434
rect 4406 9382 4458 9434
rect 4458 9382 4460 9434
rect 4404 9380 4460 9382
rect 4508 9434 4564 9436
rect 4508 9382 4510 9434
rect 4510 9382 4562 9434
rect 4562 9382 4564 9434
rect 4508 9380 4564 9382
rect 4612 9434 4668 9436
rect 4612 9382 4614 9434
rect 4614 9382 4666 9434
rect 4666 9382 4668 9434
rect 4612 9380 4668 9382
rect 4620 9098 4676 9100
rect 4620 9046 4622 9098
rect 4622 9046 4674 9098
rect 4674 9046 4676 9098
rect 4620 9044 4676 9046
rect 4396 8932 4452 8988
rect 4228 8260 4284 8316
rect 4900 8260 4956 8316
rect 4452 8036 4508 8092
rect 4404 7866 4460 7868
rect 4404 7814 4406 7866
rect 4406 7814 4458 7866
rect 4458 7814 4460 7866
rect 4404 7812 4460 7814
rect 4508 7866 4564 7868
rect 4508 7814 4510 7866
rect 4510 7814 4562 7866
rect 4562 7814 4564 7866
rect 4508 7812 4564 7814
rect 4612 7866 4668 7868
rect 4612 7814 4614 7866
rect 4614 7814 4666 7866
rect 4666 7814 4668 7866
rect 4612 7812 4668 7814
rect 4452 7476 4508 7532
rect 4004 7252 4060 7308
rect 3404 7082 3460 7084
rect 3404 7030 3406 7082
rect 3406 7030 3458 7082
rect 3458 7030 3460 7082
rect 3404 7028 3460 7030
rect 3508 7082 3564 7084
rect 3508 7030 3510 7082
rect 3510 7030 3562 7082
rect 3562 7030 3564 7082
rect 3508 7028 3564 7030
rect 3612 7082 3668 7084
rect 3612 7030 3614 7082
rect 3614 7030 3666 7082
rect 3666 7030 3668 7082
rect 3612 7028 3668 7030
rect 4228 6692 4284 6748
rect 4404 6298 4460 6300
rect 4404 6246 4406 6298
rect 4406 6246 4458 6298
rect 4458 6246 4460 6298
rect 4404 6244 4460 6246
rect 4508 6298 4564 6300
rect 4508 6246 4510 6298
rect 4510 6246 4562 6298
rect 4562 6246 4564 6298
rect 4508 6244 4564 6246
rect 4612 6298 4668 6300
rect 4612 6246 4614 6298
rect 4614 6246 4666 6298
rect 4666 6246 4668 6298
rect 4612 6244 4668 6246
rect 2996 5796 3052 5852
rect 3556 5850 3612 5852
rect 3556 5798 3558 5850
rect 3558 5798 3610 5850
rect 3610 5798 3612 5850
rect 3556 5796 3612 5798
rect 3780 5796 3836 5852
rect 3404 5514 3460 5516
rect 3404 5462 3406 5514
rect 3406 5462 3458 5514
rect 3458 5462 3460 5514
rect 3404 5460 3460 5462
rect 3508 5514 3564 5516
rect 3508 5462 3510 5514
rect 3510 5462 3562 5514
rect 3562 5462 3564 5514
rect 3508 5460 3564 5462
rect 3612 5514 3668 5516
rect 3612 5462 3614 5514
rect 3614 5462 3666 5514
rect 3666 5462 3668 5514
rect 3612 5460 3668 5462
rect 4228 5796 4284 5852
rect 4396 5738 4452 5740
rect 4396 5686 4398 5738
rect 4398 5686 4450 5738
rect 4450 5686 4452 5738
rect 4396 5684 4452 5686
rect 5180 9098 5236 9100
rect 5180 9046 5182 9098
rect 5182 9046 5234 9098
rect 5234 9046 5236 9098
rect 5180 9044 5236 9046
rect 5404 8650 5460 8652
rect 5404 8598 5406 8650
rect 5406 8598 5458 8650
rect 5458 8598 5460 8650
rect 5404 8596 5460 8598
rect 5508 8650 5564 8652
rect 5508 8598 5510 8650
rect 5510 8598 5562 8650
rect 5562 8598 5564 8650
rect 5508 8596 5564 8598
rect 5612 8650 5668 8652
rect 5612 8598 5614 8650
rect 5614 8598 5666 8650
rect 5666 8598 5668 8650
rect 5612 8596 5668 8598
rect 5236 8426 5292 8428
rect 5236 8374 5238 8426
rect 5238 8374 5290 8426
rect 5290 8374 5292 8426
rect 5236 8372 5292 8374
rect 5012 8148 5068 8204
rect 5292 8036 5348 8092
rect 4900 5796 4956 5852
rect 5012 6692 5068 6748
rect 4228 5134 4284 5180
rect 4228 5124 4230 5134
rect 4230 5124 4282 5134
rect 4282 5124 4284 5134
rect 4620 5124 4676 5180
rect 2404 4730 2460 4732
rect 2404 4678 2406 4730
rect 2406 4678 2458 4730
rect 2458 4678 2460 4730
rect 2404 4676 2460 4678
rect 2508 4730 2564 4732
rect 2508 4678 2510 4730
rect 2510 4678 2562 4730
rect 2562 4678 2564 4730
rect 2508 4676 2564 4678
rect 2612 4730 2668 4732
rect 2612 4678 2614 4730
rect 2614 4678 2666 4730
rect 2666 4678 2668 4730
rect 2612 4676 2668 4678
rect 4404 4730 4460 4732
rect 4404 4678 4406 4730
rect 4406 4678 4458 4730
rect 4458 4678 4460 4730
rect 4404 4676 4460 4678
rect 4508 4730 4564 4732
rect 4508 4678 4510 4730
rect 4510 4678 4562 4730
rect 4562 4678 4564 4730
rect 4508 4676 4564 4678
rect 4612 4730 4668 4732
rect 4612 4678 4614 4730
rect 4614 4678 4666 4730
rect 4666 4678 4668 4730
rect 4612 4676 4668 4678
rect 3556 4340 3612 4396
rect 4396 4394 4452 4396
rect 4396 4342 4398 4394
rect 4398 4342 4450 4394
rect 4450 4342 4452 4394
rect 4396 4340 4452 4342
rect 4004 4228 4060 4284
rect 3780 4116 3836 4172
rect 3404 3946 3460 3948
rect 3404 3894 3406 3946
rect 3406 3894 3458 3946
rect 3458 3894 3460 3946
rect 3404 3892 3460 3894
rect 3508 3946 3564 3948
rect 3508 3894 3510 3946
rect 3510 3894 3562 3946
rect 3562 3894 3564 3946
rect 3508 3892 3564 3894
rect 3612 3946 3668 3948
rect 3612 3894 3614 3946
rect 3614 3894 3666 3946
rect 3666 3894 3668 3946
rect 3612 3892 3668 3894
rect 1764 3556 1820 3612
rect 3332 3444 3388 3500
rect 2404 3162 2460 3164
rect 2404 3110 2406 3162
rect 2406 3110 2458 3162
rect 2458 3110 2460 3162
rect 2404 3108 2460 3110
rect 2508 3162 2564 3164
rect 2508 3110 2510 3162
rect 2510 3110 2562 3162
rect 2562 3110 2564 3162
rect 2508 3108 2564 3110
rect 2612 3162 2668 3164
rect 2612 3110 2614 3162
rect 2614 3110 2666 3162
rect 2666 3110 2668 3162
rect 2612 3108 2668 3110
rect 2940 2884 2996 2940
rect 1428 2772 1484 2828
rect 1764 2772 1820 2828
rect 2324 2772 2380 2828
rect 1404 2378 1460 2380
rect 1404 2326 1406 2378
rect 1406 2326 1458 2378
rect 1458 2326 1460 2378
rect 1404 2324 1460 2326
rect 1508 2378 1564 2380
rect 1508 2326 1510 2378
rect 1510 2326 1562 2378
rect 1562 2326 1564 2378
rect 1508 2324 1564 2326
rect 1612 2378 1668 2380
rect 1612 2326 1614 2378
rect 1614 2326 1666 2378
rect 1666 2326 1668 2378
rect 1612 2324 1668 2326
rect 1764 2154 1820 2156
rect 1764 2102 1766 2154
rect 1766 2102 1818 2154
rect 1818 2102 1820 2154
rect 1764 2100 1820 2102
rect 1428 1818 1484 1820
rect 1428 1766 1430 1818
rect 1430 1766 1482 1818
rect 1482 1766 1484 1818
rect 1428 1764 1484 1766
rect 1404 810 1460 812
rect 1404 758 1406 810
rect 1406 758 1458 810
rect 1458 758 1460 810
rect 1404 756 1460 758
rect 1508 810 1564 812
rect 1508 758 1510 810
rect 1510 758 1562 810
rect 1562 758 1564 810
rect 1508 756 1564 758
rect 1612 810 1668 812
rect 1612 758 1614 810
rect 1614 758 1666 810
rect 1666 758 1668 810
rect 1612 756 1668 758
rect 2548 2548 2604 2604
rect 2772 2602 2828 2604
rect 2772 2550 2774 2602
rect 2774 2550 2826 2602
rect 2826 2550 2828 2602
rect 2772 2548 2828 2550
rect 2404 1594 2460 1596
rect 2404 1542 2406 1594
rect 2406 1542 2458 1594
rect 2458 1542 2460 1594
rect 2404 1540 2460 1542
rect 2508 1594 2564 1596
rect 2508 1542 2510 1594
rect 2510 1542 2562 1594
rect 2562 1542 2564 1594
rect 2508 1540 2564 1542
rect 2612 1594 2668 1596
rect 2612 1542 2614 1594
rect 2614 1542 2666 1594
rect 2666 1542 2668 1594
rect 2612 1540 2668 1542
rect 4228 4116 4284 4172
rect 5404 7082 5460 7084
rect 5404 7030 5406 7082
rect 5406 7030 5458 7082
rect 5458 7030 5460 7082
rect 5404 7028 5460 7030
rect 5508 7082 5564 7084
rect 5508 7030 5510 7082
rect 5510 7030 5562 7082
rect 5562 7030 5564 7082
rect 5508 7028 5564 7030
rect 5612 7082 5668 7084
rect 5612 7030 5614 7082
rect 5614 7030 5666 7082
rect 5666 7030 5668 7082
rect 5612 7028 5668 7030
rect 5404 5514 5460 5516
rect 5404 5462 5406 5514
rect 5406 5462 5458 5514
rect 5458 5462 5460 5514
rect 5404 5460 5460 5462
rect 5508 5514 5564 5516
rect 5508 5462 5510 5514
rect 5510 5462 5562 5514
rect 5562 5462 5564 5514
rect 5508 5460 5564 5462
rect 5612 5514 5668 5516
rect 5612 5462 5614 5514
rect 5614 5462 5666 5514
rect 5666 5462 5668 5514
rect 5612 5460 5668 5462
rect 5796 4788 5852 4844
rect 5124 4228 5180 4284
rect 4452 3498 4508 3500
rect 4452 3446 4454 3498
rect 4454 3446 4506 3498
rect 4506 3446 4508 3498
rect 4452 3444 4508 3446
rect 4404 3162 4460 3164
rect 4404 3110 4406 3162
rect 4406 3110 4458 3162
rect 4458 3110 4460 3162
rect 4404 3108 4460 3110
rect 4508 3162 4564 3164
rect 4508 3110 4510 3162
rect 4510 3110 4562 3162
rect 4562 3110 4564 3162
rect 4508 3108 4564 3110
rect 4612 3162 4668 3164
rect 4612 3110 4614 3162
rect 4614 3110 4666 3162
rect 4666 3110 4668 3162
rect 4612 3108 4668 3110
rect 4004 2884 4060 2940
rect 4396 2826 4452 2828
rect 4396 2774 4398 2826
rect 4398 2774 4450 2826
rect 4450 2774 4452 2826
rect 4396 2772 4452 2774
rect 3332 2714 3388 2716
rect 3332 2662 3334 2714
rect 3334 2662 3386 2714
rect 3386 2662 3388 2714
rect 3332 2660 3388 2662
rect 3668 2714 3724 2716
rect 3668 2662 3670 2714
rect 3670 2662 3722 2714
rect 3722 2662 3724 2714
rect 3668 2660 3724 2662
rect 3780 2548 3836 2604
rect 3404 2378 3460 2380
rect 3404 2326 3406 2378
rect 3406 2326 3458 2378
rect 3458 2326 3460 2378
rect 3404 2324 3460 2326
rect 3508 2378 3564 2380
rect 3508 2326 3510 2378
rect 3510 2326 3562 2378
rect 3562 2326 3564 2378
rect 3508 2324 3564 2326
rect 3612 2378 3668 2380
rect 3612 2326 3614 2378
rect 3614 2326 3666 2378
rect 3666 2326 3668 2378
rect 3612 2324 3668 2326
rect 3404 810 3460 812
rect 3404 758 3406 810
rect 3406 758 3458 810
rect 3458 758 3460 810
rect 3404 756 3460 758
rect 3508 810 3564 812
rect 3508 758 3510 810
rect 3510 758 3562 810
rect 3562 758 3564 810
rect 3508 756 3564 758
rect 3612 810 3668 812
rect 3612 758 3614 810
rect 3614 758 3666 810
rect 3666 758 3668 810
rect 3612 756 3668 758
rect 5404 3946 5460 3948
rect 5404 3894 5406 3946
rect 5406 3894 5458 3946
rect 5458 3894 5460 3946
rect 5404 3892 5460 3894
rect 5508 3946 5564 3948
rect 5508 3894 5510 3946
rect 5510 3894 5562 3946
rect 5562 3894 5564 3946
rect 5508 3892 5564 3894
rect 5612 3946 5668 3948
rect 5612 3894 5614 3946
rect 5614 3894 5666 3946
rect 5666 3894 5668 3946
rect 5612 3892 5668 3894
rect 5908 2660 5964 2716
rect 5404 2378 5460 2380
rect 5404 2326 5406 2378
rect 5406 2326 5458 2378
rect 5458 2326 5460 2378
rect 5404 2324 5460 2326
rect 5508 2378 5564 2380
rect 5508 2326 5510 2378
rect 5510 2326 5562 2378
rect 5562 2326 5564 2378
rect 5508 2324 5564 2326
rect 5612 2378 5668 2380
rect 5612 2326 5614 2378
rect 5614 2326 5666 2378
rect 5666 2326 5668 2378
rect 5612 2324 5668 2326
rect 5236 2100 5292 2156
rect 4404 1594 4460 1596
rect 4404 1542 4406 1594
rect 4406 1542 4458 1594
rect 4458 1542 4460 1594
rect 4404 1540 4460 1542
rect 4508 1594 4564 1596
rect 4508 1542 4510 1594
rect 4510 1542 4562 1594
rect 4562 1542 4564 1594
rect 4508 1540 4564 1542
rect 4612 1594 4668 1596
rect 4612 1542 4614 1594
rect 4614 1542 4666 1594
rect 4666 1542 4668 1594
rect 4612 1540 4668 1542
rect 5404 810 5460 812
rect 5404 758 5406 810
rect 5406 758 5458 810
rect 5458 758 5460 810
rect 5404 756 5460 758
rect 5508 810 5564 812
rect 5508 758 5510 810
rect 5510 758 5562 810
rect 5562 758 5564 810
rect 5508 756 5564 758
rect 5612 810 5668 812
rect 5612 758 5614 810
rect 5614 758 5666 810
rect 5666 758 5668 810
rect 5612 756 5668 758
<< metal3 >>
rect 1394 33684 1404 33740
rect 1460 33684 1508 33740
rect 1564 33684 1612 33740
rect 1668 33684 1678 33740
rect 3394 33684 3404 33740
rect 3460 33684 3508 33740
rect 3564 33684 3612 33740
rect 3668 33684 3678 33740
rect 5394 33684 5404 33740
rect 5460 33684 5508 33740
rect 5564 33684 5612 33740
rect 5668 33684 5678 33740
rect 3994 33236 4004 33292
rect 4060 33236 4620 33292
rect 4676 33236 4686 33292
rect 394 32900 404 32956
rect 460 32900 508 32956
rect 564 32900 612 32956
rect 668 32900 678 32956
rect 2394 32900 2404 32956
rect 2460 32900 2508 32956
rect 2564 32900 2612 32956
rect 2668 32900 2678 32956
rect 4394 32900 4404 32956
rect 4460 32900 4508 32956
rect 4564 32900 4612 32956
rect 4668 32900 4678 32956
rect 3378 32340 3388 32396
rect 3444 32340 4172 32396
rect 4116 32172 4172 32340
rect 1394 32116 1404 32172
rect 1460 32116 1508 32172
rect 1564 32116 1612 32172
rect 1668 32116 1678 32172
rect 3394 32116 3404 32172
rect 3460 32116 3508 32172
rect 3564 32116 3612 32172
rect 3668 32116 3678 32172
rect 4106 32116 4116 32172
rect 4172 32116 4732 32172
rect 4788 32116 4798 32172
rect 5394 32116 5404 32172
rect 5460 32116 5508 32172
rect 5564 32116 5612 32172
rect 5668 32116 5678 32172
rect 3210 32004 3220 32060
rect 3276 32004 3948 32060
rect 4004 32004 4014 32060
rect 2762 31892 2772 31948
rect 2828 31892 4564 31948
rect 3658 31780 3668 31836
rect 3724 31780 4228 31836
rect 4284 31780 4294 31836
rect 4508 31724 4564 31892
rect 5114 31780 5124 31836
rect 5180 31780 5796 31836
rect 5852 31780 5862 31836
rect 3994 31668 4004 31724
rect 4060 31668 4340 31724
rect 4396 31668 4406 31724
rect 4498 31668 4508 31724
rect 4564 31668 5236 31724
rect 5292 31668 5302 31724
rect 3882 31556 3892 31612
rect 3948 31556 4788 31612
rect 4844 31556 4854 31612
rect 394 31332 404 31388
rect 460 31332 508 31388
rect 564 31332 612 31388
rect 668 31332 678 31388
rect 2394 31332 2404 31388
rect 2460 31332 2508 31388
rect 2564 31332 2612 31388
rect 2668 31332 2678 31388
rect 4394 31332 4404 31388
rect 4460 31332 4508 31388
rect 4564 31332 4612 31388
rect 4668 31332 4678 31388
rect 746 31108 756 31164
rect 812 31108 3668 31164
rect 3724 31108 3734 31164
rect 4676 30996 4788 31052
rect 4844 30996 5460 31052
rect 5516 30996 5526 31052
rect 4676 30940 4732 30996
rect 3770 30884 3780 30940
rect 3836 30884 4732 30940
rect 4788 30884 4798 30940
rect 4890 30884 4900 30940
rect 4956 30884 5348 30940
rect 5404 30884 5414 30940
rect 1394 30548 1404 30604
rect 1460 30548 1508 30604
rect 1564 30548 1612 30604
rect 1668 30548 1678 30604
rect 3394 30548 3404 30604
rect 3460 30548 3508 30604
rect 3564 30548 3612 30604
rect 3668 30548 3678 30604
rect 5394 30548 5404 30604
rect 5460 30548 5508 30604
rect 5564 30548 5612 30604
rect 5668 30548 5678 30604
rect 4218 30324 4228 30380
rect 4284 30324 4564 30380
rect 4620 30324 4630 30380
rect 746 30100 756 30156
rect 812 30100 4116 30156
rect 4172 30100 4182 30156
rect 1866 29988 1876 30044
rect 1932 29988 4340 30044
rect 4396 29988 4406 30044
rect 4610 29988 4620 30044
rect 4676 29988 5012 30044
rect 5068 29988 5078 30044
rect 394 29764 404 29820
rect 460 29764 508 29820
rect 564 29764 612 29820
rect 668 29764 678 29820
rect 2394 29764 2404 29820
rect 2460 29764 2508 29820
rect 2564 29764 2612 29820
rect 2668 29764 2678 29820
rect 4394 29764 4404 29820
rect 4460 29764 4508 29820
rect 4564 29764 4612 29820
rect 4668 29764 4678 29820
rect 4862 29652 4900 29708
rect 4956 29652 4966 29708
rect 1418 29316 1428 29372
rect 1484 29316 3780 29372
rect 3836 29316 3846 29372
rect 1082 29204 1092 29260
rect 1148 29204 4676 29260
rect 4732 29204 5012 29260
rect 5068 29204 5180 29260
rect 5236 29204 5246 29260
rect 5114 29092 5124 29148
rect 5180 29092 5796 29148
rect 5852 29092 5862 29148
rect 1394 28980 1404 29036
rect 1460 28980 1508 29036
rect 1564 28980 1612 29036
rect 1668 28980 1678 29036
rect 3394 28980 3404 29036
rect 3460 28980 3508 29036
rect 3564 28980 3612 29036
rect 3668 28980 3678 29036
rect 5394 28980 5404 29036
rect 5460 28980 5508 29036
rect 5564 28980 5612 29036
rect 5668 28980 5678 29036
rect 3658 28756 3668 28812
rect 3724 28756 4004 28812
rect 4060 28756 4070 28812
rect 186 28420 196 28476
rect 252 28420 1204 28476
rect 1260 28420 1270 28476
rect 3882 28420 3892 28476
rect 3948 28420 3958 28476
rect 394 28196 404 28252
rect 460 28196 508 28252
rect 564 28196 612 28252
rect 668 28196 678 28252
rect 2394 28196 2404 28252
rect 2460 28196 2508 28252
rect 2564 28196 2612 28252
rect 2668 28196 2678 28252
rect 3892 28028 3948 28420
rect 4394 28196 4404 28252
rect 4460 28196 4508 28252
rect 4564 28196 4612 28252
rect 4668 28196 4678 28252
rect 3892 27972 4004 28028
rect 4060 27972 4070 28028
rect 3994 27860 4004 27916
rect 4060 27860 5236 27916
rect 5292 27860 5302 27916
rect 1754 27748 1764 27804
rect 1820 27748 3444 27804
rect 3500 27748 3892 27804
rect 3948 27748 5124 27804
rect 5180 27748 5190 27804
rect 5226 27636 5236 27692
rect 5292 27636 5796 27692
rect 5852 27636 5862 27692
rect 1394 27412 1404 27468
rect 1460 27412 1508 27468
rect 1564 27412 1612 27468
rect 1668 27412 1678 27468
rect 3394 27412 3404 27468
rect 3460 27412 3508 27468
rect 3564 27412 3612 27468
rect 3668 27412 3678 27468
rect 5394 27412 5404 27468
rect 5460 27412 5508 27468
rect 5564 27412 5612 27468
rect 5668 27412 5678 27468
rect 4778 27300 4788 27356
rect 4844 27300 4956 27356
rect 4900 27244 4956 27300
rect 3658 27188 3668 27244
rect 3724 27188 4228 27244
rect 4284 27188 4294 27244
rect 4890 27188 4900 27244
rect 4956 27188 4966 27244
rect 4750 27076 4788 27132
rect 4844 27076 4854 27132
rect 5002 27076 5012 27132
rect 5068 27076 5124 27132
rect 5180 27076 5190 27132
rect 4890 26852 4900 26908
rect 4956 26852 4966 26908
rect 4900 26796 4956 26852
rect 746 26740 756 26796
rect 812 26740 1204 26796
rect 1260 26740 1270 26796
rect 4900 26740 5460 26796
rect 5516 26740 5526 26796
rect 394 26628 404 26684
rect 460 26628 508 26684
rect 564 26628 612 26684
rect 668 26628 678 26684
rect 2394 26628 2404 26684
rect 2460 26628 2508 26684
rect 2564 26628 2612 26684
rect 2668 26628 2678 26684
rect 3770 26628 3780 26684
rect 3836 26628 4116 26684
rect 4172 26628 4182 26684
rect 4394 26628 4404 26684
rect 4460 26628 4508 26684
rect 4564 26628 4612 26684
rect 4668 26628 4678 26684
rect 4106 26516 4116 26572
rect 4172 26516 5348 26572
rect 5404 26516 5414 26572
rect 3994 26404 4004 26460
rect 4060 26404 4676 26460
rect 4732 26404 4742 26460
rect 3322 26292 3332 26348
rect 3388 26292 3780 26348
rect 3836 26292 3846 26348
rect 4106 26292 4116 26348
rect 4172 26292 4396 26348
rect 4452 26292 4462 26348
rect 4778 26292 4788 26348
rect 4844 26292 5796 26348
rect 5852 26292 5862 26348
rect 4498 26180 4508 26236
rect 4564 26180 4900 26236
rect 4956 26180 4966 26236
rect 3770 26068 3780 26124
rect 3836 26068 4340 26124
rect 4396 26068 4406 26124
rect 5002 26068 5012 26124
rect 5068 26068 5124 26124
rect 5180 26068 5190 26124
rect 5758 26068 5796 26124
rect 5852 26068 5862 26124
rect 4162 25956 4172 26012
rect 4228 25956 5012 26012
rect 5068 25956 5078 26012
rect 1394 25844 1404 25900
rect 1460 25844 1508 25900
rect 1564 25844 1612 25900
rect 1668 25844 1678 25900
rect 3394 25844 3404 25900
rect 3460 25844 3508 25900
rect 3564 25844 3612 25900
rect 3668 25844 3678 25900
rect 4218 25844 4228 25900
rect 4284 25844 4340 25900
rect 4396 25844 4406 25900
rect 5394 25844 5404 25900
rect 5460 25844 5508 25900
rect 5564 25844 5612 25900
rect 5668 25844 5678 25900
rect 4050 25508 4060 25564
rect 4116 25508 4508 25564
rect 4564 25508 4574 25564
rect 394 25060 404 25116
rect 460 25060 508 25116
rect 564 25060 612 25116
rect 668 25060 678 25116
rect 2394 25060 2404 25116
rect 2460 25060 2508 25116
rect 2564 25060 2612 25116
rect 2668 25060 2678 25116
rect 3770 25060 3780 25116
rect 3836 25060 3892 25116
rect 3948 25060 4228 25116
rect 4284 25060 4294 25116
rect 4394 25060 4404 25116
rect 4460 25060 4508 25116
rect 4564 25060 4612 25116
rect 4668 25060 4678 25116
rect 1394 24276 1404 24332
rect 1460 24276 1508 24332
rect 1564 24276 1612 24332
rect 1668 24276 1678 24332
rect 3394 24276 3404 24332
rect 3460 24276 3508 24332
rect 3564 24276 3612 24332
rect 3668 24276 3678 24332
rect 5394 24276 5404 24332
rect 5460 24276 5508 24332
rect 5564 24276 5612 24332
rect 5668 24276 5678 24332
rect 746 23940 756 23996
rect 812 23940 3892 23996
rect 3948 23940 4172 23996
rect 4116 23884 4172 23940
rect 4106 23828 4116 23884
rect 4172 23828 4620 23884
rect 4676 23828 4686 23884
rect 5226 23828 5236 23884
rect 5292 23828 5796 23884
rect 5852 23828 5862 23884
rect 394 23492 404 23548
rect 460 23492 508 23548
rect 564 23492 612 23548
rect 668 23492 678 23548
rect 2394 23492 2404 23548
rect 2460 23492 2508 23548
rect 2564 23492 2612 23548
rect 2668 23492 2678 23548
rect 4394 23492 4404 23548
rect 4460 23492 4508 23548
rect 4564 23492 4612 23548
rect 4668 23492 4678 23548
rect 4676 23380 4956 23436
rect 5012 23380 5022 23436
rect 4676 23324 4732 23380
rect 2874 23268 2884 23324
rect 2940 23268 3388 23324
rect 4666 23268 4676 23324
rect 4732 23268 4742 23324
rect 3332 23100 3388 23268
rect 3332 23044 4004 23100
rect 4060 23044 4564 23100
rect 4620 23044 4630 23100
rect 5786 23044 5796 23100
rect 5852 23044 5908 23100
rect 5964 23044 5974 23100
rect 4004 22932 5180 22988
rect 5236 22932 5246 22988
rect 4004 22764 4060 22932
rect 5450 22876 5460 22922
rect 4610 22820 4620 22876
rect 4676 22820 5012 22876
rect 5068 22820 5078 22876
rect 5226 22820 5236 22876
rect 5292 22866 5460 22876
rect 5516 22866 5526 22922
rect 5292 22820 5516 22866
rect 1394 22708 1404 22764
rect 1460 22708 1508 22764
rect 1564 22708 1612 22764
rect 1668 22708 1678 22764
rect 3394 22708 3404 22764
rect 3460 22708 3508 22764
rect 3564 22708 3612 22764
rect 3668 22708 3678 22764
rect 3994 22708 4004 22764
rect 4060 22708 4070 22764
rect 5394 22708 5404 22764
rect 5460 22708 5508 22764
rect 5564 22708 5612 22764
rect 5668 22708 5678 22764
rect 4004 22652 4060 22708
rect 3332 22596 4060 22652
rect 3332 22428 3388 22596
rect 3714 22484 3724 22540
rect 3780 22484 4620 22540
rect 4676 22484 4686 22540
rect 2436 22372 2716 22428
rect 2772 22372 3388 22428
rect 3882 22372 3892 22428
rect 3948 22372 4228 22428
rect 4284 22372 4294 22428
rect 2436 22316 2492 22372
rect 2258 22260 2268 22316
rect 2324 22260 2492 22316
rect 1922 22148 1932 22204
rect 1988 22148 3108 22204
rect 3164 22148 3174 22204
rect 4228 22148 4452 22204
rect 4508 22148 4518 22204
rect 394 21924 404 21980
rect 460 21924 508 21980
rect 564 21924 612 21980
rect 668 21924 678 21980
rect 2394 21924 2404 21980
rect 2460 21924 2508 21980
rect 2564 21924 2612 21980
rect 2668 21924 2678 21980
rect 4228 21756 4284 22148
rect 4394 21924 4404 21980
rect 4460 21924 4508 21980
rect 4564 21924 4612 21980
rect 4668 21924 4678 21980
rect 5114 21812 5124 21868
rect 5180 21812 5190 21868
rect 1092 21700 3892 21756
rect 3948 21700 3958 21756
rect 4228 21700 4452 21756
rect 4508 21700 4518 21756
rect 1092 21644 1148 21700
rect 5124 21644 5180 21812
rect 746 21588 756 21644
rect 812 21588 1092 21644
rect 1148 21588 1158 21644
rect 3882 21588 3892 21644
rect 3948 21588 5180 21644
rect 1082 21476 1092 21532
rect 1148 21476 4004 21532
rect 4060 21476 4676 21532
rect 4732 21476 4742 21532
rect 4676 21420 4732 21476
rect 1418 21364 1428 21420
rect 1484 21364 4004 21420
rect 4060 21364 4070 21420
rect 4676 21364 5180 21420
rect 5236 21364 5246 21420
rect 4106 21252 4116 21308
rect 4172 21252 4452 21308
rect 4508 21252 4518 21308
rect 1394 21140 1404 21196
rect 1460 21140 1508 21196
rect 1564 21140 1612 21196
rect 1668 21140 1678 21196
rect 3394 21140 3404 21196
rect 3460 21140 3508 21196
rect 3564 21140 3612 21196
rect 3668 21140 3678 21196
rect 5394 21140 5404 21196
rect 5460 21140 5508 21196
rect 5564 21140 5612 21196
rect 5668 21140 5678 21196
rect 2090 20580 2100 20636
rect 2156 20580 5236 20636
rect 5292 20580 5302 20636
rect 394 20356 404 20412
rect 460 20356 508 20412
rect 564 20356 612 20412
rect 668 20356 678 20412
rect 2394 20356 2404 20412
rect 2460 20356 2508 20412
rect 2564 20356 2612 20412
rect 2668 20356 2678 20412
rect 4394 20356 4404 20412
rect 4460 20356 4508 20412
rect 4564 20356 4612 20412
rect 4668 20356 4678 20412
rect 5758 19684 5796 19740
rect 5852 19684 5862 19740
rect 1394 19572 1404 19628
rect 1460 19572 1508 19628
rect 1564 19572 1612 19628
rect 1668 19572 1678 19628
rect 3394 19572 3404 19628
rect 3460 19572 3508 19628
rect 3564 19572 3612 19628
rect 3668 19572 3678 19628
rect 5394 19572 5404 19628
rect 5460 19572 5508 19628
rect 5564 19572 5612 19628
rect 5668 19572 5678 19628
rect 1754 19348 1764 19404
rect 1820 19348 2100 19404
rect 2156 19348 2268 19404
rect 2324 19348 2604 19404
rect 2660 19348 2670 19404
rect 5002 18900 5012 18956
rect 5068 18900 6000 18956
rect 394 18788 404 18844
rect 460 18788 508 18844
rect 564 18788 612 18844
rect 668 18788 678 18844
rect 2394 18788 2404 18844
rect 2460 18788 2508 18844
rect 2564 18788 2612 18844
rect 2668 18788 2678 18844
rect 4394 18788 4404 18844
rect 4460 18788 4508 18844
rect 4564 18788 4612 18844
rect 4668 18788 4678 18844
rect 5338 18452 5348 18508
rect 5404 18452 6000 18508
rect 3938 18340 3948 18396
rect 4004 18340 5012 18396
rect 5068 18340 5078 18396
rect 4162 18228 4172 18284
rect 4228 18228 5180 18284
rect 5236 18228 5852 18284
rect 5796 18060 5852 18228
rect 1394 18004 1404 18060
rect 1460 18004 1508 18060
rect 1564 18004 1612 18060
rect 1668 18004 1678 18060
rect 3394 18004 3404 18060
rect 3460 18004 3508 18060
rect 3564 18004 3612 18060
rect 3668 18004 3678 18060
rect 3770 18004 3780 18060
rect 3836 18004 4228 18060
rect 4284 18004 4294 18060
rect 5394 18004 5404 18060
rect 5460 18004 5508 18060
rect 5564 18004 5612 18060
rect 5668 18004 5678 18060
rect 5796 18032 6000 18060
rect 5800 18004 6000 18032
rect 2772 17780 4564 17836
rect 4620 17780 4788 17836
rect 4844 17780 4854 17836
rect 2772 17612 2828 17780
rect 4274 17668 4284 17724
rect 4340 17668 5124 17724
rect 5180 17668 5190 17724
rect 2762 17556 2772 17612
rect 2828 17556 2838 17612
rect 3770 17556 3780 17612
rect 3836 17556 6000 17612
rect 2538 17444 2548 17500
rect 2604 17444 2772 17500
rect 2828 17444 2838 17500
rect 4274 17444 4284 17500
rect 4340 17444 5348 17500
rect 5404 17444 5414 17500
rect 394 17220 404 17276
rect 460 17220 508 17276
rect 564 17220 612 17276
rect 668 17220 678 17276
rect 2394 17220 2404 17276
rect 2460 17220 2508 17276
rect 2564 17220 2612 17276
rect 2668 17220 2678 17276
rect 4394 17220 4404 17276
rect 4460 17220 4508 17276
rect 4564 17220 4612 17276
rect 4668 17220 4678 17276
rect 4778 17108 4788 17164
rect 4844 17108 6000 17164
rect 970 16996 980 17052
rect 1036 16996 3948 17052
rect 4004 16996 4014 17052
rect 4162 16996 4172 17052
rect 4228 16996 5684 17052
rect 5740 16996 5750 17052
rect 3490 16884 3500 16940
rect 3556 16884 4732 16940
rect 4788 16884 4798 16940
rect 2930 16772 2940 16828
rect 2996 16772 3780 16828
rect 3836 16772 3846 16828
rect 4050 16772 4060 16828
rect 4116 16772 4900 16828
rect 4956 16772 4966 16828
rect 1922 16660 1932 16716
rect 1988 16660 2548 16716
rect 2604 16660 2614 16716
rect 3098 16660 3108 16716
rect 3164 16660 3556 16716
rect 3612 16660 3622 16716
rect 4722 16660 4732 16716
rect 4788 16660 6000 16716
rect 1394 16436 1404 16492
rect 1460 16436 1508 16492
rect 1564 16436 1612 16492
rect 1668 16436 1678 16492
rect 3394 16436 3404 16492
rect 3460 16436 3508 16492
rect 3564 16436 3612 16492
rect 3668 16436 3678 16492
rect 5394 16436 5404 16492
rect 5460 16436 5508 16492
rect 5564 16436 5612 16492
rect 5668 16436 5678 16492
rect 2370 16324 2380 16380
rect 2436 16324 4452 16380
rect 4508 16324 4518 16380
rect 2090 16212 2100 16268
rect 2156 16212 3948 16268
rect 4004 16212 4676 16268
rect 4732 16212 4742 16268
rect 5002 16212 5012 16268
rect 5068 16212 5078 16268
rect 5226 16212 5236 16268
rect 5292 16212 6000 16268
rect 5012 16156 5068 16212
rect 2538 16100 2548 16156
rect 2604 16100 2772 16156
rect 2828 16100 2838 16156
rect 3378 16100 3388 16156
rect 3444 16100 5348 16156
rect 5404 16100 5414 16156
rect 2090 15988 2100 16044
rect 2156 15988 4788 16044
rect 4844 15988 4854 16044
rect 4946 15988 4956 16044
rect 5068 15988 5078 16044
rect 1698 15876 1708 15932
rect 1764 15876 2716 15932
rect 2772 15876 3388 15932
rect 3444 15876 3454 15932
rect 4778 15764 4788 15820
rect 4844 15764 6000 15820
rect 394 15652 404 15708
rect 460 15652 508 15708
rect 564 15652 612 15708
rect 668 15652 678 15708
rect 2394 15652 2404 15708
rect 2460 15652 2508 15708
rect 2564 15652 2612 15708
rect 2668 15652 2678 15708
rect 4394 15652 4404 15708
rect 4460 15652 4508 15708
rect 4564 15652 4612 15708
rect 4668 15652 4678 15708
rect 1418 15316 1428 15372
rect 1484 15316 3220 15372
rect 3276 15316 3286 15372
rect 3994 15316 4004 15372
rect 4060 15316 4676 15372
rect 4732 15316 4742 15372
rect 4106 15204 4116 15260
rect 4172 15204 4228 15260
rect 4284 15204 4294 15260
rect 5786 15092 5796 15148
rect 5852 15092 5908 15148
rect 5964 15092 5974 15148
rect 1394 14868 1404 14924
rect 1460 14868 1508 14924
rect 1564 14868 1612 14924
rect 1668 14868 1678 14924
rect 3394 14868 3404 14924
rect 3460 14868 3508 14924
rect 3564 14868 3612 14924
rect 3668 14868 3678 14924
rect 5394 14868 5404 14924
rect 5460 14868 5508 14924
rect 5564 14868 5612 14924
rect 5668 14868 5678 14924
rect 2090 14644 2100 14700
rect 2212 14644 2436 14700
rect 2492 14644 2502 14700
rect 4834 14532 4844 14588
rect 4956 14532 4966 14588
rect 4666 14308 4676 14364
rect 4732 14308 5180 14364
rect 5236 14308 5246 14364
rect 394 14084 404 14140
rect 460 14084 508 14140
rect 564 14084 612 14140
rect 668 14084 678 14140
rect 2394 14084 2404 14140
rect 2460 14084 2508 14140
rect 2564 14084 2612 14140
rect 2668 14084 2678 14140
rect 4394 14084 4404 14140
rect 4460 14084 4508 14140
rect 4564 14084 4612 14140
rect 4668 14084 4678 14140
rect 186 13972 196 14028
rect 252 13972 4620 14028
rect 4564 13916 4620 13972
rect 2090 13860 2100 13916
rect 2156 13860 2660 13916
rect 2716 13860 2726 13916
rect 4554 13860 4564 13916
rect 4620 13860 4630 13916
rect 4750 13860 4788 13916
rect 4844 13860 4854 13916
rect 2818 13748 2828 13804
rect 2884 13748 3780 13804
rect 3836 13748 4116 13804
rect 4172 13748 4182 13804
rect 2314 13636 2324 13692
rect 2380 13636 2772 13692
rect 2828 13636 2838 13692
rect 2034 13524 2044 13580
rect 1054 13412 1092 13468
rect 1148 13412 1158 13468
rect 2100 13356 2156 13580
rect 3434 13524 3444 13580
rect 3500 13524 4004 13580
rect 4060 13524 4070 13580
rect 4442 13524 4452 13580
rect 4508 13524 4900 13580
rect 4956 13524 4966 13580
rect 1394 13300 1404 13356
rect 1460 13300 1508 13356
rect 1564 13300 1612 13356
rect 1668 13300 1678 13356
rect 2100 13300 2492 13356
rect 2548 13300 3052 13356
rect 3108 13244 3164 13356
rect 3394 13300 3404 13356
rect 3460 13300 3508 13356
rect 3564 13300 3612 13356
rect 3668 13300 3678 13356
rect 5394 13300 5404 13356
rect 5460 13300 5508 13356
rect 5564 13300 5612 13356
rect 5668 13300 5678 13356
rect 3108 13188 4620 13244
rect 4676 13188 5124 13244
rect 5180 13188 5190 13244
rect 158 13076 196 13132
rect 252 13076 262 13132
rect 5198 13076 5236 13132
rect 5292 13076 5302 13132
rect 1418 12964 1428 13020
rect 1484 12964 3780 13020
rect 3836 12964 3846 13020
rect 3378 12852 3388 12908
rect 3444 12852 4900 12908
rect 4956 12852 4966 12908
rect 4106 12740 4116 12796
rect 4172 12740 4284 12796
rect 4340 12740 4350 12796
rect 394 12516 404 12572
rect 460 12516 508 12572
rect 564 12516 612 12572
rect 668 12516 678 12572
rect 2394 12516 2404 12572
rect 2460 12516 2508 12572
rect 2564 12516 2612 12572
rect 2668 12516 2678 12572
rect 4394 12516 4404 12572
rect 4460 12516 4508 12572
rect 4564 12516 4612 12572
rect 4668 12516 4678 12572
rect 74 12404 84 12460
rect 140 12404 980 12460
rect 1036 12404 1046 12460
rect 4050 12180 4060 12236
rect 4116 12180 4564 12236
rect 4620 12180 5180 12236
rect 5236 12180 5796 12236
rect 5852 12180 5862 12236
rect 4666 12068 4676 12124
rect 4732 12068 5012 12124
rect 5068 12068 5078 12124
rect 1394 11732 1404 11788
rect 1460 11732 1508 11788
rect 1564 11732 1612 11788
rect 1668 11732 1678 11788
rect 3394 11732 3404 11788
rect 3460 11732 3508 11788
rect 3564 11732 3612 11788
rect 3668 11732 3678 11788
rect 5394 11732 5404 11788
rect 5460 11732 5508 11788
rect 5564 11732 5612 11788
rect 5668 11732 5678 11788
rect 4946 11284 4956 11340
rect 5012 11284 5796 11340
rect 5852 11284 5862 11340
rect 394 10948 404 11004
rect 460 10948 508 11004
rect 564 10948 612 11004
rect 668 10948 678 11004
rect 2394 10948 2404 11004
rect 2460 10948 2508 11004
rect 2564 10948 2612 11004
rect 2668 10948 2678 11004
rect 3994 10948 4004 11004
rect 4060 10948 4228 11004
rect 4284 10948 4294 11004
rect 4394 10948 4404 11004
rect 4460 10948 4508 11004
rect 4564 10948 4612 11004
rect 4668 10948 4678 11004
rect 3658 10724 3668 10780
rect 3724 10724 4564 10780
rect 4620 10724 4630 10780
rect 2762 10500 2772 10556
rect 2828 10500 4564 10556
rect 4620 10500 4630 10556
rect 3434 10388 3444 10444
rect 3500 10388 4004 10444
rect 4060 10388 4070 10444
rect 1394 10164 1404 10220
rect 1460 10164 1508 10220
rect 1564 10164 1612 10220
rect 1668 10164 1678 10220
rect 3394 10164 3404 10220
rect 3460 10164 3508 10220
rect 3564 10164 3612 10220
rect 3668 10164 3678 10220
rect 5394 10164 5404 10220
rect 5460 10164 5508 10220
rect 5564 10164 5612 10220
rect 5668 10164 5678 10220
rect 186 9940 196 9996
rect 252 9940 644 9996
rect 700 9940 710 9996
rect 1418 9828 1428 9884
rect 1484 9828 3108 9884
rect 3164 9828 3174 9884
rect 186 9716 196 9772
rect 252 9716 868 9772
rect 924 9716 934 9772
rect 394 9380 404 9436
rect 460 9380 508 9436
rect 564 9380 612 9436
rect 668 9380 678 9436
rect 2394 9380 2404 9436
rect 2460 9380 2508 9436
rect 2564 9380 2612 9436
rect 2668 9380 2678 9436
rect 4394 9380 4404 9436
rect 4460 9380 4508 9436
rect 4564 9380 4612 9436
rect 4668 9380 4678 9436
rect 1866 9156 1876 9212
rect 1932 9156 2660 9212
rect 2716 9156 2726 9212
rect 3378 9156 3388 9212
rect 3444 9156 3892 9212
rect 3948 9156 4844 9212
rect 4788 9100 4844 9156
rect 746 9044 756 9100
rect 812 9044 1204 9100
rect 1260 9044 1270 9100
rect 3154 9044 3164 9100
rect 3220 9044 4116 9100
rect 4172 9044 4620 9100
rect 4676 9044 4686 9100
rect 4788 9044 5180 9100
rect 5236 9044 5796 9100
rect 5852 9044 5862 9100
rect 2650 8932 2660 8988
rect 2716 8932 2772 8988
rect 2828 8932 2838 8988
rect 3882 8932 3892 8988
rect 3948 8932 4396 8988
rect 4452 8932 4462 8988
rect 3892 8876 3948 8932
rect 2370 8820 2380 8876
rect 2436 8820 2828 8876
rect 2884 8820 3948 8876
rect 1394 8596 1404 8652
rect 1460 8596 1508 8652
rect 1564 8596 1612 8652
rect 1668 8596 1678 8652
rect 3394 8596 3404 8652
rect 3460 8596 3508 8652
rect 3564 8596 3612 8652
rect 3668 8596 3678 8652
rect 5394 8596 5404 8652
rect 5460 8596 5508 8652
rect 5564 8596 5612 8652
rect 5668 8596 5678 8652
rect 186 8372 196 8428
rect 252 8372 5236 8428
rect 5292 8372 5302 8428
rect 4218 8260 4228 8316
rect 4284 8260 4900 8316
rect 4956 8260 4966 8316
rect 1082 8148 1092 8204
rect 1148 8148 5012 8204
rect 5068 8148 5078 8204
rect 4442 8036 4452 8092
rect 4508 8036 5292 8092
rect 5348 8036 5358 8092
rect 394 7812 404 7868
rect 460 7812 508 7868
rect 564 7812 612 7868
rect 668 7812 678 7868
rect 2394 7812 2404 7868
rect 2460 7812 2508 7868
rect 2564 7812 2612 7868
rect 2668 7812 2678 7868
rect 4394 7812 4404 7868
rect 4460 7812 4508 7868
rect 4564 7812 4612 7868
rect 4668 7812 4678 7868
rect 3770 7476 3780 7532
rect 3836 7476 4452 7532
rect 4508 7476 4518 7532
rect 2762 7252 2772 7308
rect 2828 7252 4004 7308
rect 4060 7252 4070 7308
rect 1394 7028 1404 7084
rect 1460 7028 1508 7084
rect 1564 7028 1612 7084
rect 1668 7028 1678 7084
rect 3394 7028 3404 7084
rect 3460 7028 3508 7084
rect 3564 7028 3612 7084
rect 3668 7028 3678 7084
rect 5394 7028 5404 7084
rect 5460 7028 5508 7084
rect 5564 7028 5612 7084
rect 5668 7028 5678 7084
rect 942 6692 980 6748
rect 1036 6692 1046 6748
rect 4190 6692 4228 6748
rect 4284 6692 4294 6748
rect 4974 6692 5012 6748
rect 5068 6692 5078 6748
rect 394 6244 404 6300
rect 460 6244 508 6300
rect 564 6244 612 6300
rect 668 6244 678 6300
rect 2394 6244 2404 6300
rect 2460 6244 2508 6300
rect 2564 6244 2612 6300
rect 2668 6244 2678 6300
rect 4394 6244 4404 6300
rect 4460 6244 4508 6300
rect 4564 6244 4612 6300
rect 4668 6244 4678 6300
rect 2986 5796 2996 5852
rect 3052 5796 3556 5852
rect 3612 5796 3622 5852
rect 3770 5796 3780 5852
rect 3836 5796 4228 5852
rect 4284 5796 4900 5852
rect 4956 5796 4966 5852
rect 3556 5740 3612 5796
rect 3556 5684 4396 5740
rect 4452 5684 4462 5740
rect 1394 5460 1404 5516
rect 1460 5460 1508 5516
rect 1564 5460 1612 5516
rect 1668 5460 1678 5516
rect 3394 5460 3404 5516
rect 3460 5460 3508 5516
rect 3564 5460 3612 5516
rect 3668 5460 3678 5516
rect 5394 5460 5404 5516
rect 5460 5460 5508 5516
rect 5564 5460 5612 5516
rect 5668 5460 5678 5516
rect 4218 5124 4228 5180
rect 4284 5124 4620 5180
rect 4676 5124 4686 5180
rect 4228 5068 4284 5124
rect 746 5012 756 5068
rect 812 5012 4284 5068
rect 634 4900 644 4956
rect 700 4900 1204 4956
rect 1260 4900 1270 4956
rect 1082 4788 1092 4844
rect 1148 4788 5796 4844
rect 5852 4788 5862 4844
rect 394 4676 404 4732
rect 460 4676 508 4732
rect 564 4676 612 4732
rect 668 4676 678 4732
rect 2394 4676 2404 4732
rect 2460 4676 2508 4732
rect 2564 4676 2612 4732
rect 2668 4676 2678 4732
rect 4394 4676 4404 4732
rect 4460 4676 4508 4732
rect 4564 4676 4612 4732
rect 4668 4676 4678 4732
rect 3546 4340 3556 4396
rect 3612 4340 4228 4396
rect 4284 4340 4396 4396
rect 4452 4340 4462 4396
rect 3994 4228 4004 4284
rect 4060 4228 5124 4284
rect 5180 4228 5190 4284
rect 3770 4116 3780 4172
rect 3836 4116 4004 4172
rect 4060 4116 4228 4172
rect 4284 4116 4294 4172
rect 1394 3892 1404 3948
rect 1460 3892 1508 3948
rect 1564 3892 1612 3948
rect 1668 3892 1678 3948
rect 3394 3892 3404 3948
rect 3460 3892 3508 3948
rect 3564 3892 3612 3948
rect 3668 3892 3678 3948
rect 5394 3892 5404 3948
rect 5460 3892 5508 3948
rect 5564 3892 5612 3948
rect 5668 3892 5678 3948
rect 634 3556 644 3612
rect 700 3556 1764 3612
rect 1820 3556 1830 3612
rect 970 3444 980 3500
rect 1036 3444 1316 3500
rect 1372 3444 1382 3500
rect 3322 3444 3332 3500
rect 3388 3444 4452 3500
rect 4508 3444 4518 3500
rect 394 3108 404 3164
rect 460 3108 508 3164
rect 564 3108 612 3164
rect 668 3108 678 3164
rect 2394 3108 2404 3164
rect 2460 3108 2508 3164
rect 2564 3108 2612 3164
rect 2668 3108 2678 3164
rect 4394 3108 4404 3164
rect 4460 3108 4508 3164
rect 4564 3108 4612 3164
rect 4668 3108 4678 3164
rect 2930 2884 2940 2940
rect 2996 2884 4004 2940
rect 4060 2884 4070 2940
rect 1418 2772 1428 2828
rect 1484 2772 1764 2828
rect 1820 2772 2324 2828
rect 2380 2772 4228 2828
rect 4284 2772 4396 2828
rect 4452 2772 4462 2828
rect 2548 2660 3332 2716
rect 3388 2660 3398 2716
rect 3658 2660 3668 2716
rect 3724 2660 5908 2716
rect 5964 2660 5974 2716
rect 2548 2604 2604 2660
rect 2538 2548 2548 2604
rect 2604 2548 2614 2604
rect 2762 2548 2772 2604
rect 2828 2548 3780 2604
rect 3836 2548 3846 2604
rect 1394 2324 1404 2380
rect 1460 2324 1508 2380
rect 1564 2324 1612 2380
rect 1668 2324 1678 2380
rect 3394 2324 3404 2380
rect 3460 2324 3508 2380
rect 3564 2324 3612 2380
rect 3668 2324 3678 2380
rect 5394 2324 5404 2380
rect 5460 2324 5508 2380
rect 5564 2324 5612 2380
rect 5668 2324 5678 2380
rect 1754 2100 1764 2156
rect 1820 2100 5236 2156
rect 5292 2100 5302 2156
rect 858 1764 868 1820
rect 924 1764 1428 1820
rect 1484 1764 1494 1820
rect 394 1540 404 1596
rect 460 1540 508 1596
rect 564 1540 612 1596
rect 668 1540 678 1596
rect 2394 1540 2404 1596
rect 2460 1540 2508 1596
rect 2564 1540 2612 1596
rect 2668 1540 2678 1596
rect 4394 1540 4404 1596
rect 4460 1540 4508 1596
rect 4564 1540 4612 1596
rect 4668 1540 4678 1596
rect 1394 756 1404 812
rect 1460 756 1508 812
rect 1564 756 1612 812
rect 1668 756 1678 812
rect 3394 756 3404 812
rect 3460 756 3508 812
rect 3564 756 3612 812
rect 3668 756 3678 812
rect 5394 756 5404 812
rect 5460 756 5508 812
rect 5564 756 5612 812
rect 5668 756 5678 812
<< via3 >>
rect 1404 33684 1460 33740
rect 1508 33684 1564 33740
rect 1612 33684 1668 33740
rect 3404 33684 3460 33740
rect 3508 33684 3564 33740
rect 3612 33684 3668 33740
rect 5404 33684 5460 33740
rect 5508 33684 5564 33740
rect 5612 33684 5668 33740
rect 404 32900 460 32956
rect 508 32900 564 32956
rect 612 32900 668 32956
rect 2404 32900 2460 32956
rect 2508 32900 2564 32956
rect 2612 32900 2668 32956
rect 4404 32900 4460 32956
rect 4508 32900 4564 32956
rect 4612 32900 4668 32956
rect 1404 32116 1460 32172
rect 1508 32116 1564 32172
rect 1612 32116 1668 32172
rect 3404 32116 3460 32172
rect 3508 32116 3564 32172
rect 3612 32116 3668 32172
rect 4116 32116 4172 32172
rect 5404 32116 5460 32172
rect 5508 32116 5564 32172
rect 5612 32116 5668 32172
rect 5796 31780 5852 31836
rect 404 31332 460 31388
rect 508 31332 564 31388
rect 612 31332 668 31388
rect 2404 31332 2460 31388
rect 2508 31332 2564 31388
rect 2612 31332 2668 31388
rect 4404 31332 4460 31388
rect 4508 31332 4564 31388
rect 4612 31332 4668 31388
rect 4788 30996 4844 31052
rect 1404 30548 1460 30604
rect 1508 30548 1564 30604
rect 1612 30548 1668 30604
rect 3404 30548 3460 30604
rect 3508 30548 3564 30604
rect 3612 30548 3668 30604
rect 5404 30548 5460 30604
rect 5508 30548 5564 30604
rect 5612 30548 5668 30604
rect 4228 30324 4284 30380
rect 5012 29988 5068 30044
rect 404 29764 460 29820
rect 508 29764 564 29820
rect 612 29764 668 29820
rect 2404 29764 2460 29820
rect 2508 29764 2564 29820
rect 2612 29764 2668 29820
rect 4404 29764 4460 29820
rect 4508 29764 4564 29820
rect 4612 29764 4668 29820
rect 4900 29652 4956 29708
rect 5124 29092 5180 29148
rect 1404 28980 1460 29036
rect 1508 28980 1564 29036
rect 1612 28980 1668 29036
rect 3404 28980 3460 29036
rect 3508 28980 3564 29036
rect 3612 28980 3668 29036
rect 5404 28980 5460 29036
rect 5508 28980 5564 29036
rect 5612 28980 5668 29036
rect 404 28196 460 28252
rect 508 28196 564 28252
rect 612 28196 668 28252
rect 2404 28196 2460 28252
rect 2508 28196 2564 28252
rect 2612 28196 2668 28252
rect 4404 28196 4460 28252
rect 4508 28196 4564 28252
rect 4612 28196 4668 28252
rect 4004 27860 4060 27916
rect 3892 27748 3948 27804
rect 5236 27636 5292 27692
rect 1404 27412 1460 27468
rect 1508 27412 1564 27468
rect 1612 27412 1668 27468
rect 3404 27412 3460 27468
rect 3508 27412 3564 27468
rect 3612 27412 3668 27468
rect 5404 27412 5460 27468
rect 5508 27412 5564 27468
rect 5612 27412 5668 27468
rect 4788 27300 4844 27356
rect 4788 27076 4844 27132
rect 5012 27076 5068 27132
rect 404 26628 460 26684
rect 508 26628 564 26684
rect 612 26628 668 26684
rect 2404 26628 2460 26684
rect 2508 26628 2564 26684
rect 2612 26628 2668 26684
rect 4404 26628 4460 26684
rect 4508 26628 4564 26684
rect 4612 26628 4668 26684
rect 4116 26516 4172 26572
rect 4004 26404 4060 26460
rect 4116 26292 4172 26348
rect 5796 26292 5852 26348
rect 4900 26180 4956 26236
rect 5124 26068 5180 26124
rect 5796 26068 5852 26124
rect 5012 25956 5068 26012
rect 1404 25844 1460 25900
rect 1508 25844 1564 25900
rect 1612 25844 1668 25900
rect 3404 25844 3460 25900
rect 3508 25844 3564 25900
rect 3612 25844 3668 25900
rect 4228 25844 4284 25900
rect 5404 25844 5460 25900
rect 5508 25844 5564 25900
rect 5612 25844 5668 25900
rect 404 25060 460 25116
rect 508 25060 564 25116
rect 612 25060 668 25116
rect 2404 25060 2460 25116
rect 2508 25060 2564 25116
rect 2612 25060 2668 25116
rect 3892 25060 3948 25116
rect 4404 25060 4460 25116
rect 4508 25060 4564 25116
rect 4612 25060 4668 25116
rect 1404 24276 1460 24332
rect 1508 24276 1564 24332
rect 1612 24276 1668 24332
rect 3404 24276 3460 24332
rect 3508 24276 3564 24332
rect 3612 24276 3668 24332
rect 5404 24276 5460 24332
rect 5508 24276 5564 24332
rect 5612 24276 5668 24332
rect 5796 23828 5852 23884
rect 404 23492 460 23548
rect 508 23492 564 23548
rect 612 23492 668 23548
rect 2404 23492 2460 23548
rect 2508 23492 2564 23548
rect 2612 23492 2668 23548
rect 4404 23492 4460 23548
rect 4508 23492 4564 23548
rect 4612 23492 4668 23548
rect 5908 23044 5964 23100
rect 5012 22820 5068 22876
rect 5236 22820 5292 22876
rect 1404 22708 1460 22764
rect 1508 22708 1564 22764
rect 1612 22708 1668 22764
rect 3404 22708 3460 22764
rect 3508 22708 3564 22764
rect 3612 22708 3668 22764
rect 5404 22708 5460 22764
rect 5508 22708 5564 22764
rect 5612 22708 5668 22764
rect 4228 22372 4284 22428
rect 404 21924 460 21980
rect 508 21924 564 21980
rect 612 21924 668 21980
rect 2404 21924 2460 21980
rect 2508 21924 2564 21980
rect 2612 21924 2668 21980
rect 4404 21924 4460 21980
rect 4508 21924 4564 21980
rect 4612 21924 4668 21980
rect 1092 21588 1148 21644
rect 3892 21588 3948 21644
rect 4004 21476 4060 21532
rect 1404 21140 1460 21196
rect 1508 21140 1564 21196
rect 1612 21140 1668 21196
rect 3404 21140 3460 21196
rect 3508 21140 3564 21196
rect 3612 21140 3668 21196
rect 5404 21140 5460 21196
rect 5508 21140 5564 21196
rect 5612 21140 5668 21196
rect 404 20356 460 20412
rect 508 20356 564 20412
rect 612 20356 668 20412
rect 2404 20356 2460 20412
rect 2508 20356 2564 20412
rect 2612 20356 2668 20412
rect 4404 20356 4460 20412
rect 4508 20356 4564 20412
rect 4612 20356 4668 20412
rect 5796 19684 5852 19740
rect 1404 19572 1460 19628
rect 1508 19572 1564 19628
rect 1612 19572 1668 19628
rect 3404 19572 3460 19628
rect 3508 19572 3564 19628
rect 3612 19572 3668 19628
rect 5404 19572 5460 19628
rect 5508 19572 5564 19628
rect 5612 19572 5668 19628
rect 2100 19348 2156 19404
rect 404 18788 460 18844
rect 508 18788 564 18844
rect 612 18788 668 18844
rect 2404 18788 2460 18844
rect 2508 18788 2564 18844
rect 2612 18788 2668 18844
rect 4404 18788 4460 18844
rect 4508 18788 4564 18844
rect 4612 18788 4668 18844
rect 1404 18004 1460 18060
rect 1508 18004 1564 18060
rect 1612 18004 1668 18060
rect 3404 18004 3460 18060
rect 3508 18004 3564 18060
rect 3612 18004 3668 18060
rect 4228 18004 4284 18060
rect 5404 18004 5460 18060
rect 5508 18004 5564 18060
rect 5612 18004 5668 18060
rect 4788 17780 4844 17836
rect 2772 17444 2828 17500
rect 404 17220 460 17276
rect 508 17220 564 17276
rect 612 17220 668 17276
rect 2404 17220 2460 17276
rect 2508 17220 2564 17276
rect 2612 17220 2668 17276
rect 4404 17220 4460 17276
rect 4508 17220 4564 17276
rect 4612 17220 4668 17276
rect 980 16996 1036 17052
rect 1404 16436 1460 16492
rect 1508 16436 1564 16492
rect 1612 16436 1668 16492
rect 3404 16436 3460 16492
rect 3508 16436 3564 16492
rect 3612 16436 3668 16492
rect 5404 16436 5460 16492
rect 5508 16436 5564 16492
rect 5612 16436 5668 16492
rect 5012 16212 5068 16268
rect 5236 16212 5292 16268
rect 2772 16100 2828 16156
rect 5012 15988 5068 16044
rect 4788 15764 4844 15820
rect 404 15652 460 15708
rect 508 15652 564 15708
rect 612 15652 668 15708
rect 2404 15652 2460 15708
rect 2508 15652 2564 15708
rect 2612 15652 2668 15708
rect 4404 15652 4460 15708
rect 4508 15652 4564 15708
rect 4612 15652 4668 15708
rect 4004 15316 4060 15372
rect 4116 15204 4172 15260
rect 5908 15092 5964 15148
rect 1404 14868 1460 14924
rect 1508 14868 1564 14924
rect 1612 14868 1668 14924
rect 3404 14868 3460 14924
rect 3508 14868 3564 14924
rect 3612 14868 3668 14924
rect 5404 14868 5460 14924
rect 5508 14868 5564 14924
rect 5612 14868 5668 14924
rect 2100 14644 2156 14700
rect 4900 14532 4956 14588
rect 404 14084 460 14140
rect 508 14084 564 14140
rect 612 14084 668 14140
rect 2404 14084 2460 14140
rect 2508 14084 2564 14140
rect 2612 14084 2668 14140
rect 4404 14084 4460 14140
rect 4508 14084 4564 14140
rect 4612 14084 4668 14140
rect 2100 13860 2156 13916
rect 4788 13860 4844 13916
rect 4116 13748 4172 13804
rect 2772 13636 2828 13692
rect 1092 13412 1148 13468
rect 1404 13300 1460 13356
rect 1508 13300 1564 13356
rect 1612 13300 1668 13356
rect 3404 13300 3460 13356
rect 3508 13300 3564 13356
rect 3612 13300 3668 13356
rect 5404 13300 5460 13356
rect 5508 13300 5564 13356
rect 5612 13300 5668 13356
rect 5124 13188 5180 13244
rect 196 13076 252 13132
rect 5236 13076 5292 13132
rect 4116 12740 4172 12796
rect 404 12516 460 12572
rect 508 12516 564 12572
rect 612 12516 668 12572
rect 2404 12516 2460 12572
rect 2508 12516 2564 12572
rect 2612 12516 2668 12572
rect 4404 12516 4460 12572
rect 4508 12516 4564 12572
rect 4612 12516 4668 12572
rect 1404 11732 1460 11788
rect 1508 11732 1564 11788
rect 1612 11732 1668 11788
rect 3404 11732 3460 11788
rect 3508 11732 3564 11788
rect 3612 11732 3668 11788
rect 5404 11732 5460 11788
rect 5508 11732 5564 11788
rect 5612 11732 5668 11788
rect 404 10948 460 11004
rect 508 10948 564 11004
rect 612 10948 668 11004
rect 2404 10948 2460 11004
rect 2508 10948 2564 11004
rect 2612 10948 2668 11004
rect 4004 10948 4060 11004
rect 4404 10948 4460 11004
rect 4508 10948 4564 11004
rect 4612 10948 4668 11004
rect 2772 10500 2828 10556
rect 1404 10164 1460 10220
rect 1508 10164 1564 10220
rect 1612 10164 1668 10220
rect 3404 10164 3460 10220
rect 3508 10164 3564 10220
rect 3612 10164 3668 10220
rect 5404 10164 5460 10220
rect 5508 10164 5564 10220
rect 5612 10164 5668 10220
rect 404 9380 460 9436
rect 508 9380 564 9436
rect 612 9380 668 9436
rect 2404 9380 2460 9436
rect 2508 9380 2564 9436
rect 2612 9380 2668 9436
rect 4404 9380 4460 9436
rect 4508 9380 4564 9436
rect 4612 9380 4668 9436
rect 4116 9044 4172 9100
rect 5796 9044 5852 9100
rect 2772 8932 2828 8988
rect 3892 8932 3948 8988
rect 1404 8596 1460 8652
rect 1508 8596 1564 8652
rect 1612 8596 1668 8652
rect 3404 8596 3460 8652
rect 3508 8596 3564 8652
rect 3612 8596 3668 8652
rect 5404 8596 5460 8652
rect 5508 8596 5564 8652
rect 5612 8596 5668 8652
rect 196 8372 252 8428
rect 404 7812 460 7868
rect 508 7812 564 7868
rect 612 7812 668 7868
rect 2404 7812 2460 7868
rect 2508 7812 2564 7868
rect 2612 7812 2668 7868
rect 4404 7812 4460 7868
rect 4508 7812 4564 7868
rect 4612 7812 4668 7868
rect 2772 7252 2828 7308
rect 1404 7028 1460 7084
rect 1508 7028 1564 7084
rect 1612 7028 1668 7084
rect 3404 7028 3460 7084
rect 3508 7028 3564 7084
rect 3612 7028 3668 7084
rect 5404 7028 5460 7084
rect 5508 7028 5564 7084
rect 5612 7028 5668 7084
rect 980 6692 1036 6748
rect 4228 6692 4284 6748
rect 5012 6692 5068 6748
rect 404 6244 460 6300
rect 508 6244 564 6300
rect 612 6244 668 6300
rect 2404 6244 2460 6300
rect 2508 6244 2564 6300
rect 2612 6244 2668 6300
rect 4404 6244 4460 6300
rect 4508 6244 4564 6300
rect 4612 6244 4668 6300
rect 1404 5460 1460 5516
rect 1508 5460 1564 5516
rect 1612 5460 1668 5516
rect 3404 5460 3460 5516
rect 3508 5460 3564 5516
rect 3612 5460 3668 5516
rect 5404 5460 5460 5516
rect 5508 5460 5564 5516
rect 5612 5460 5668 5516
rect 404 4676 460 4732
rect 508 4676 564 4732
rect 612 4676 668 4732
rect 2404 4676 2460 4732
rect 2508 4676 2564 4732
rect 2612 4676 2668 4732
rect 4404 4676 4460 4732
rect 4508 4676 4564 4732
rect 4612 4676 4668 4732
rect 4228 4340 4284 4396
rect 4004 4116 4060 4172
rect 1404 3892 1460 3948
rect 1508 3892 1564 3948
rect 1612 3892 1668 3948
rect 3404 3892 3460 3948
rect 3508 3892 3564 3948
rect 3612 3892 3668 3948
rect 5404 3892 5460 3948
rect 5508 3892 5564 3948
rect 5612 3892 5668 3948
rect 404 3108 460 3164
rect 508 3108 564 3164
rect 612 3108 668 3164
rect 2404 3108 2460 3164
rect 2508 3108 2564 3164
rect 2612 3108 2668 3164
rect 4404 3108 4460 3164
rect 4508 3108 4564 3164
rect 4612 3108 4668 3164
rect 4228 2772 4284 2828
rect 1404 2324 1460 2380
rect 1508 2324 1564 2380
rect 1612 2324 1668 2380
rect 3404 2324 3460 2380
rect 3508 2324 3564 2380
rect 3612 2324 3668 2380
rect 5404 2324 5460 2380
rect 5508 2324 5564 2380
rect 5612 2324 5668 2380
rect 404 1540 460 1596
rect 508 1540 564 1596
rect 612 1540 668 1596
rect 2404 1540 2460 1596
rect 2508 1540 2564 1596
rect 2612 1540 2668 1596
rect 4404 1540 4460 1596
rect 4508 1540 4564 1596
rect 4612 1540 4668 1596
rect 1404 756 1460 812
rect 1508 756 1564 812
rect 1612 756 1668 812
rect 3404 756 3460 812
rect 3508 756 3564 812
rect 3612 756 3668 812
rect 5404 756 5460 812
rect 5508 756 5564 812
rect 5612 756 5668 812
<< metal4 >>
rect 376 32956 696 33772
rect 376 32900 404 32956
rect 460 32900 508 32956
rect 564 32900 612 32956
rect 668 32900 696 32956
rect 376 31388 696 32900
rect 376 31332 404 31388
rect 460 31332 508 31388
rect 564 31332 612 31388
rect 668 31332 696 31388
rect 376 29820 696 31332
rect 376 29764 404 29820
rect 460 29764 508 29820
rect 564 29764 612 29820
rect 668 29764 696 29820
rect 376 29216 696 29764
rect 376 29160 404 29216
rect 460 29160 508 29216
rect 564 29160 612 29216
rect 668 29160 696 29216
rect 376 29112 696 29160
rect 376 29056 404 29112
rect 460 29056 508 29112
rect 564 29056 612 29112
rect 668 29056 696 29112
rect 376 29008 696 29056
rect 376 28952 404 29008
rect 460 28952 508 29008
rect 564 28952 612 29008
rect 668 28952 696 29008
rect 376 28252 696 28952
rect 376 28196 404 28252
rect 460 28196 508 28252
rect 564 28196 612 28252
rect 668 28196 696 28252
rect 376 26684 696 28196
rect 376 26628 404 26684
rect 460 26628 508 26684
rect 564 26628 612 26684
rect 668 26628 696 26684
rect 376 25116 696 26628
rect 376 25060 404 25116
rect 460 25060 508 25116
rect 564 25060 612 25116
rect 668 25060 696 25116
rect 376 23548 696 25060
rect 376 23492 404 23548
rect 460 23492 508 23548
rect 564 23492 612 23548
rect 668 23492 696 23548
rect 376 22216 696 23492
rect 376 22160 404 22216
rect 460 22160 508 22216
rect 564 22160 612 22216
rect 668 22160 696 22216
rect 376 22112 696 22160
rect 376 22056 404 22112
rect 460 22056 508 22112
rect 564 22056 612 22112
rect 668 22056 696 22112
rect 376 22008 696 22056
rect 376 21924 404 22008
rect 460 21924 508 22008
rect 564 21924 612 22008
rect 668 21924 696 22008
rect 376 20412 696 21924
rect 1376 33740 1696 33772
rect 1376 33684 1404 33740
rect 1460 33684 1508 33740
rect 1564 33684 1612 33740
rect 1668 33684 1696 33740
rect 1376 32716 1696 33684
rect 1376 32660 1404 32716
rect 1460 32660 1508 32716
rect 1564 32660 1612 32716
rect 1668 32660 1696 32716
rect 1376 32612 1696 32660
rect 1376 32556 1404 32612
rect 1460 32556 1508 32612
rect 1564 32556 1612 32612
rect 1668 32556 1696 32612
rect 1376 32508 1696 32556
rect 1376 32452 1404 32508
rect 1460 32452 1508 32508
rect 1564 32452 1612 32508
rect 1668 32452 1696 32508
rect 1376 32172 1696 32452
rect 1376 32116 1404 32172
rect 1460 32116 1508 32172
rect 1564 32116 1612 32172
rect 1668 32116 1696 32172
rect 1376 30604 1696 32116
rect 1376 30548 1404 30604
rect 1460 30548 1508 30604
rect 1564 30548 1612 30604
rect 1668 30548 1696 30604
rect 1376 29036 1696 30548
rect 1376 28980 1404 29036
rect 1460 28980 1508 29036
rect 1564 28980 1612 29036
rect 1668 28980 1696 29036
rect 1376 27468 1696 28980
rect 1376 27412 1404 27468
rect 1460 27412 1508 27468
rect 1564 27412 1612 27468
rect 1668 27412 1696 27468
rect 1376 25900 1696 27412
rect 1376 25844 1404 25900
rect 1460 25844 1508 25900
rect 1564 25844 1612 25900
rect 1668 25844 1696 25900
rect 1376 25716 1696 25844
rect 1376 25660 1404 25716
rect 1460 25660 1508 25716
rect 1564 25660 1612 25716
rect 1668 25660 1696 25716
rect 1376 25612 1696 25660
rect 1376 25556 1404 25612
rect 1460 25556 1508 25612
rect 1564 25556 1612 25612
rect 1668 25556 1696 25612
rect 1376 25508 1696 25556
rect 1376 25452 1404 25508
rect 1460 25452 1508 25508
rect 1564 25452 1612 25508
rect 1668 25452 1696 25508
rect 1376 24332 1696 25452
rect 1376 24276 1404 24332
rect 1460 24276 1508 24332
rect 1564 24276 1612 24332
rect 1668 24276 1696 24332
rect 1376 22764 1696 24276
rect 1376 22708 1404 22764
rect 1460 22708 1508 22764
rect 1564 22708 1612 22764
rect 1668 22708 1696 22764
rect 376 20356 404 20412
rect 460 20356 508 20412
rect 564 20356 612 20412
rect 668 20356 696 20412
rect 376 18844 696 20356
rect 376 18788 404 18844
rect 460 18788 508 18844
rect 564 18788 612 18844
rect 668 18788 696 18844
rect 376 17276 696 18788
rect 376 17220 404 17276
rect 460 17220 508 17276
rect 564 17220 612 17276
rect 668 17220 696 17276
rect 376 15708 696 17220
rect 1092 21644 1148 21654
rect 376 15652 404 15708
rect 460 15652 508 15708
rect 564 15652 612 15708
rect 668 15652 696 15708
rect 376 15216 696 15652
rect 376 15160 404 15216
rect 460 15160 508 15216
rect 564 15160 612 15216
rect 668 15160 696 15216
rect 376 15112 696 15160
rect 376 15056 404 15112
rect 460 15056 508 15112
rect 564 15056 612 15112
rect 668 15056 696 15112
rect 376 15008 696 15056
rect 376 14952 404 15008
rect 460 14952 508 15008
rect 564 14952 612 15008
rect 668 14952 696 15008
rect 376 14140 696 14952
rect 376 14084 404 14140
rect 460 14084 508 14140
rect 564 14084 612 14140
rect 668 14084 696 14140
rect 196 13132 252 13142
rect 196 8428 252 13076
rect 196 8362 252 8372
rect 376 12572 696 14084
rect 376 12516 404 12572
rect 460 12516 508 12572
rect 564 12516 612 12572
rect 668 12516 696 12572
rect 376 11004 696 12516
rect 376 10948 404 11004
rect 460 10948 508 11004
rect 564 10948 612 11004
rect 668 10948 696 11004
rect 376 9436 696 10948
rect 376 9380 404 9436
rect 460 9380 508 9436
rect 564 9380 612 9436
rect 668 9380 696 9436
rect 376 8216 696 9380
rect 376 8160 404 8216
rect 460 8160 508 8216
rect 564 8160 612 8216
rect 668 8160 696 8216
rect 376 8112 696 8160
rect 376 8056 404 8112
rect 460 8056 508 8112
rect 564 8056 612 8112
rect 668 8056 696 8112
rect 376 8008 696 8056
rect 376 7952 404 8008
rect 460 7952 508 8008
rect 564 7952 612 8008
rect 668 7952 696 8008
rect 376 7868 696 7952
rect 376 7812 404 7868
rect 460 7812 508 7868
rect 564 7812 612 7868
rect 668 7812 696 7868
rect 376 6300 696 7812
rect 980 17052 1036 17062
rect 980 6748 1036 16996
rect 1092 13468 1148 21588
rect 1092 13402 1148 13412
rect 1376 21196 1696 22708
rect 1376 21140 1404 21196
rect 1460 21140 1508 21196
rect 1564 21140 1612 21196
rect 1668 21140 1696 21196
rect 1376 19628 1696 21140
rect 1376 19572 1404 19628
rect 1460 19572 1508 19628
rect 1564 19572 1612 19628
rect 1668 19572 1696 19628
rect 1376 18716 1696 19572
rect 2376 32956 2696 33772
rect 2376 32900 2404 32956
rect 2460 32900 2508 32956
rect 2564 32900 2612 32956
rect 2668 32900 2696 32956
rect 2376 31388 2696 32900
rect 2376 31332 2404 31388
rect 2460 31332 2508 31388
rect 2564 31332 2612 31388
rect 2668 31332 2696 31388
rect 2376 29820 2696 31332
rect 2376 29764 2404 29820
rect 2460 29764 2508 29820
rect 2564 29764 2612 29820
rect 2668 29764 2696 29820
rect 2376 29216 2696 29764
rect 2376 29160 2404 29216
rect 2460 29160 2508 29216
rect 2564 29160 2612 29216
rect 2668 29160 2696 29216
rect 2376 29112 2696 29160
rect 2376 29056 2404 29112
rect 2460 29056 2508 29112
rect 2564 29056 2612 29112
rect 2668 29056 2696 29112
rect 2376 29008 2696 29056
rect 2376 28952 2404 29008
rect 2460 28952 2508 29008
rect 2564 28952 2612 29008
rect 2668 28952 2696 29008
rect 2376 28252 2696 28952
rect 2376 28196 2404 28252
rect 2460 28196 2508 28252
rect 2564 28196 2612 28252
rect 2668 28196 2696 28252
rect 2376 26684 2696 28196
rect 2376 26628 2404 26684
rect 2460 26628 2508 26684
rect 2564 26628 2612 26684
rect 2668 26628 2696 26684
rect 2376 25116 2696 26628
rect 2376 25060 2404 25116
rect 2460 25060 2508 25116
rect 2564 25060 2612 25116
rect 2668 25060 2696 25116
rect 2376 23548 2696 25060
rect 2376 23492 2404 23548
rect 2460 23492 2508 23548
rect 2564 23492 2612 23548
rect 2668 23492 2696 23548
rect 2376 22216 2696 23492
rect 2376 22160 2404 22216
rect 2460 22160 2508 22216
rect 2564 22160 2612 22216
rect 2668 22160 2696 22216
rect 2376 22112 2696 22160
rect 2376 22056 2404 22112
rect 2460 22056 2508 22112
rect 2564 22056 2612 22112
rect 2668 22056 2696 22112
rect 2376 22008 2696 22056
rect 2376 21924 2404 22008
rect 2460 21924 2508 22008
rect 2564 21924 2612 22008
rect 2668 21924 2696 22008
rect 2376 20412 2696 21924
rect 2376 20356 2404 20412
rect 2460 20356 2508 20412
rect 2564 20356 2612 20412
rect 2668 20356 2696 20412
rect 1376 18660 1404 18716
rect 1460 18660 1508 18716
rect 1564 18660 1612 18716
rect 1668 18660 1696 18716
rect 1376 18612 1696 18660
rect 1376 18556 1404 18612
rect 1460 18556 1508 18612
rect 1564 18556 1612 18612
rect 1668 18556 1696 18612
rect 1376 18508 1696 18556
rect 1376 18452 1404 18508
rect 1460 18452 1508 18508
rect 1564 18452 1612 18508
rect 1668 18452 1696 18508
rect 1376 18060 1696 18452
rect 1376 18004 1404 18060
rect 1460 18004 1508 18060
rect 1564 18004 1612 18060
rect 1668 18004 1696 18060
rect 1376 16492 1696 18004
rect 1376 16436 1404 16492
rect 1460 16436 1508 16492
rect 1564 16436 1612 16492
rect 1668 16436 1696 16492
rect 1376 14924 1696 16436
rect 1376 14868 1404 14924
rect 1460 14868 1508 14924
rect 1564 14868 1612 14924
rect 1668 14868 1696 14924
rect 980 6682 1036 6692
rect 1376 13356 1696 14868
rect 2100 19404 2156 19414
rect 2100 14700 2156 19348
rect 2100 13916 2156 14644
rect 2100 13850 2156 13860
rect 2376 18844 2696 20356
rect 2376 18788 2404 18844
rect 2460 18788 2508 18844
rect 2564 18788 2612 18844
rect 2668 18788 2696 18844
rect 2376 17276 2696 18788
rect 3376 33740 3696 33772
rect 3376 33684 3404 33740
rect 3460 33684 3508 33740
rect 3564 33684 3612 33740
rect 3668 33684 3696 33740
rect 3376 32716 3696 33684
rect 3376 32660 3404 32716
rect 3460 32660 3508 32716
rect 3564 32660 3612 32716
rect 3668 32660 3696 32716
rect 3376 32612 3696 32660
rect 3376 32556 3404 32612
rect 3460 32556 3508 32612
rect 3564 32556 3612 32612
rect 3668 32556 3696 32612
rect 3376 32508 3696 32556
rect 3376 32452 3404 32508
rect 3460 32452 3508 32508
rect 3564 32452 3612 32508
rect 3668 32452 3696 32508
rect 3376 32172 3696 32452
rect 4376 32956 4696 33772
rect 4376 32900 4404 32956
rect 4460 32900 4508 32956
rect 4564 32900 4612 32956
rect 4668 32900 4696 32956
rect 3376 32116 3404 32172
rect 3460 32116 3508 32172
rect 3564 32116 3612 32172
rect 3668 32116 3696 32172
rect 3376 30604 3696 32116
rect 3376 30548 3404 30604
rect 3460 30548 3508 30604
rect 3564 30548 3612 30604
rect 3668 30548 3696 30604
rect 3376 29036 3696 30548
rect 3376 28980 3404 29036
rect 3460 28980 3508 29036
rect 3564 28980 3612 29036
rect 3668 28980 3696 29036
rect 3376 27468 3696 28980
rect 4116 32172 4172 32182
rect 4004 27916 4060 27926
rect 3376 27412 3404 27468
rect 3460 27412 3508 27468
rect 3564 27412 3612 27468
rect 3668 27412 3696 27468
rect 3376 25900 3696 27412
rect 3376 25844 3404 25900
rect 3460 25844 3508 25900
rect 3564 25844 3612 25900
rect 3668 25844 3696 25900
rect 3376 25716 3696 25844
rect 3376 25660 3404 25716
rect 3460 25660 3508 25716
rect 3564 25660 3612 25716
rect 3668 25660 3696 25716
rect 3376 25612 3696 25660
rect 3376 25556 3404 25612
rect 3460 25556 3508 25612
rect 3564 25556 3612 25612
rect 3668 25556 3696 25612
rect 3376 25508 3696 25556
rect 3376 25452 3404 25508
rect 3460 25452 3508 25508
rect 3564 25452 3612 25508
rect 3668 25452 3696 25508
rect 3376 24332 3696 25452
rect 3892 27804 3948 27814
rect 3892 25116 3948 27748
rect 4004 26460 4060 27860
rect 4004 26394 4060 26404
rect 4116 26572 4172 32116
rect 4376 31388 4696 32900
rect 4376 31332 4404 31388
rect 4460 31332 4508 31388
rect 4564 31332 4612 31388
rect 4668 31332 4696 31388
rect 4116 26348 4172 26516
rect 4116 26282 4172 26292
rect 4228 30380 4284 30390
rect 4228 25900 4284 30324
rect 4228 25834 4284 25844
rect 4376 29820 4696 31332
rect 5376 33740 5696 33772
rect 5376 33684 5404 33740
rect 5460 33684 5508 33740
rect 5564 33684 5612 33740
rect 5668 33684 5696 33740
rect 5376 32716 5696 33684
rect 5376 32660 5404 32716
rect 5460 32660 5508 32716
rect 5564 32660 5612 32716
rect 5668 32660 5696 32716
rect 5376 32612 5696 32660
rect 5376 32556 5404 32612
rect 5460 32556 5508 32612
rect 5564 32556 5612 32612
rect 5668 32556 5696 32612
rect 5376 32508 5696 32556
rect 5376 32452 5404 32508
rect 5460 32452 5508 32508
rect 5564 32452 5612 32508
rect 5668 32452 5696 32508
rect 5376 32172 5696 32452
rect 5376 32116 5404 32172
rect 5460 32116 5508 32172
rect 5564 32116 5612 32172
rect 5668 32116 5696 32172
rect 4376 29764 4404 29820
rect 4460 29764 4508 29820
rect 4564 29764 4612 29820
rect 4668 29764 4696 29820
rect 4376 29216 4696 29764
rect 4376 29160 4404 29216
rect 4460 29160 4508 29216
rect 4564 29160 4612 29216
rect 4668 29160 4696 29216
rect 4376 29112 4696 29160
rect 4376 29056 4404 29112
rect 4460 29056 4508 29112
rect 4564 29056 4612 29112
rect 4668 29056 4696 29112
rect 4376 29008 4696 29056
rect 4376 28952 4404 29008
rect 4460 28952 4508 29008
rect 4564 28952 4612 29008
rect 4668 28952 4696 29008
rect 4376 28252 4696 28952
rect 4376 28196 4404 28252
rect 4460 28196 4508 28252
rect 4564 28196 4612 28252
rect 4668 28196 4696 28252
rect 4376 26684 4696 28196
rect 4788 31052 4844 31062
rect 4788 27356 4844 30996
rect 5376 30604 5696 32116
rect 5376 30548 5404 30604
rect 5460 30548 5508 30604
rect 5564 30548 5612 30604
rect 5668 30548 5696 30604
rect 5012 30044 5068 30054
rect 4788 27290 4844 27300
rect 4900 29708 4956 29718
rect 4376 26628 4404 26684
rect 4460 26628 4508 26684
rect 4564 26628 4612 26684
rect 4668 26628 4696 26684
rect 3892 25050 3948 25060
rect 4376 25116 4696 26628
rect 4376 25060 4404 25116
rect 4460 25060 4508 25116
rect 4564 25060 4612 25116
rect 4668 25060 4696 25116
rect 3376 24276 3404 24332
rect 3460 24276 3508 24332
rect 3564 24276 3612 24332
rect 3668 24276 3696 24332
rect 3376 22764 3696 24276
rect 3376 22708 3404 22764
rect 3460 22708 3508 22764
rect 3564 22708 3612 22764
rect 3668 22708 3696 22764
rect 3376 21196 3696 22708
rect 4376 23548 4696 25060
rect 4376 23492 4404 23548
rect 4460 23492 4508 23548
rect 4564 23492 4612 23548
rect 4668 23492 4696 23548
rect 4228 22428 4284 22438
rect 4228 21868 4284 22372
rect 4116 21812 4284 21868
rect 4376 22216 4696 23492
rect 4376 22160 4404 22216
rect 4460 22160 4508 22216
rect 4564 22160 4612 22216
rect 4668 22160 4696 22216
rect 4376 22112 4696 22160
rect 4376 22056 4404 22112
rect 4460 22056 4508 22112
rect 4564 22056 4612 22112
rect 4668 22056 4696 22112
rect 4376 22008 4696 22056
rect 4376 21924 4404 22008
rect 4460 21924 4508 22008
rect 4564 21924 4612 22008
rect 4668 21924 4696 22008
rect 3376 21140 3404 21196
rect 3460 21140 3508 21196
rect 3564 21140 3612 21196
rect 3668 21140 3696 21196
rect 3376 19628 3696 21140
rect 3376 19572 3404 19628
rect 3460 19572 3508 19628
rect 3564 19572 3612 19628
rect 3668 19572 3696 19628
rect 3376 18716 3696 19572
rect 3376 18660 3404 18716
rect 3460 18660 3508 18716
rect 3564 18660 3612 18716
rect 3668 18660 3696 18716
rect 3376 18612 3696 18660
rect 3376 18556 3404 18612
rect 3460 18556 3508 18612
rect 3564 18556 3612 18612
rect 3668 18556 3696 18612
rect 3376 18508 3696 18556
rect 3376 18452 3404 18508
rect 3460 18452 3508 18508
rect 3564 18452 3612 18508
rect 3668 18452 3696 18508
rect 3376 18060 3696 18452
rect 3376 18004 3404 18060
rect 3460 18004 3508 18060
rect 3564 18004 3612 18060
rect 3668 18004 3696 18060
rect 2376 17220 2404 17276
rect 2460 17220 2508 17276
rect 2564 17220 2612 17276
rect 2668 17220 2696 17276
rect 2376 15708 2696 17220
rect 2376 15652 2404 15708
rect 2460 15652 2508 15708
rect 2564 15652 2612 15708
rect 2668 15652 2696 15708
rect 2376 15216 2696 15652
rect 2376 15160 2404 15216
rect 2460 15160 2508 15216
rect 2564 15160 2612 15216
rect 2668 15160 2696 15216
rect 2376 15112 2696 15160
rect 2376 15056 2404 15112
rect 2460 15056 2508 15112
rect 2564 15056 2612 15112
rect 2668 15056 2696 15112
rect 2376 15008 2696 15056
rect 2376 14952 2404 15008
rect 2460 14952 2508 15008
rect 2564 14952 2612 15008
rect 2668 14952 2696 15008
rect 2376 14140 2696 14952
rect 2376 14084 2404 14140
rect 2460 14084 2508 14140
rect 2564 14084 2612 14140
rect 2668 14084 2696 14140
rect 1376 13300 1404 13356
rect 1460 13300 1508 13356
rect 1564 13300 1612 13356
rect 1668 13300 1696 13356
rect 1376 11788 1696 13300
rect 1376 11732 1404 11788
rect 1460 11732 1508 11788
rect 1564 11732 1612 11788
rect 1668 11732 1696 11788
rect 1376 11716 1696 11732
rect 1376 11660 1404 11716
rect 1460 11660 1508 11716
rect 1564 11660 1612 11716
rect 1668 11660 1696 11716
rect 1376 11612 1696 11660
rect 1376 11556 1404 11612
rect 1460 11556 1508 11612
rect 1564 11556 1612 11612
rect 1668 11556 1696 11612
rect 1376 11508 1696 11556
rect 1376 11452 1404 11508
rect 1460 11452 1508 11508
rect 1564 11452 1612 11508
rect 1668 11452 1696 11508
rect 1376 10220 1696 11452
rect 1376 10164 1404 10220
rect 1460 10164 1508 10220
rect 1564 10164 1612 10220
rect 1668 10164 1696 10220
rect 1376 8652 1696 10164
rect 1376 8596 1404 8652
rect 1460 8596 1508 8652
rect 1564 8596 1612 8652
rect 1668 8596 1696 8652
rect 1376 7084 1696 8596
rect 1376 7028 1404 7084
rect 1460 7028 1508 7084
rect 1564 7028 1612 7084
rect 1668 7028 1696 7084
rect 376 6244 404 6300
rect 460 6244 508 6300
rect 564 6244 612 6300
rect 668 6244 696 6300
rect 376 4732 696 6244
rect 376 4676 404 4732
rect 460 4676 508 4732
rect 564 4676 612 4732
rect 668 4676 696 4732
rect 376 3164 696 4676
rect 376 3108 404 3164
rect 460 3108 508 3164
rect 564 3108 612 3164
rect 668 3108 696 3164
rect 376 1596 696 3108
rect 376 1540 404 1596
rect 460 1540 508 1596
rect 564 1540 612 1596
rect 668 1540 696 1596
rect 376 1216 696 1540
rect 376 1160 404 1216
rect 460 1160 508 1216
rect 564 1160 612 1216
rect 668 1160 696 1216
rect 376 1112 696 1160
rect 376 1056 404 1112
rect 460 1056 508 1112
rect 564 1056 612 1112
rect 668 1056 696 1112
rect 376 1008 696 1056
rect 376 952 404 1008
rect 460 952 508 1008
rect 564 952 612 1008
rect 668 952 696 1008
rect 376 724 696 952
rect 1376 5516 1696 7028
rect 1376 5460 1404 5516
rect 1460 5460 1508 5516
rect 1564 5460 1612 5516
rect 1668 5460 1696 5516
rect 1376 4716 1696 5460
rect 1376 4660 1404 4716
rect 1460 4660 1508 4716
rect 1564 4660 1612 4716
rect 1668 4660 1696 4716
rect 1376 4612 1696 4660
rect 1376 4556 1404 4612
rect 1460 4556 1508 4612
rect 1564 4556 1612 4612
rect 1668 4556 1696 4612
rect 1376 4508 1696 4556
rect 1376 4452 1404 4508
rect 1460 4452 1508 4508
rect 1564 4452 1612 4508
rect 1668 4452 1696 4508
rect 1376 3948 1696 4452
rect 1376 3892 1404 3948
rect 1460 3892 1508 3948
rect 1564 3892 1612 3948
rect 1668 3892 1696 3948
rect 1376 2380 1696 3892
rect 1376 2324 1404 2380
rect 1460 2324 1508 2380
rect 1564 2324 1612 2380
rect 1668 2324 1696 2380
rect 1376 812 1696 2324
rect 1376 756 1404 812
rect 1460 756 1508 812
rect 1564 756 1612 812
rect 1668 756 1696 812
rect 1376 724 1696 756
rect 2376 12572 2696 14084
rect 2376 12516 2404 12572
rect 2460 12516 2508 12572
rect 2564 12516 2612 12572
rect 2668 12516 2696 12572
rect 2376 11004 2696 12516
rect 2376 10948 2404 11004
rect 2460 10948 2508 11004
rect 2564 10948 2612 11004
rect 2668 10948 2696 11004
rect 2376 9436 2696 10948
rect 2376 9380 2404 9436
rect 2460 9380 2508 9436
rect 2564 9380 2612 9436
rect 2668 9380 2696 9436
rect 2376 8216 2696 9380
rect 2376 8160 2404 8216
rect 2460 8160 2508 8216
rect 2564 8160 2612 8216
rect 2668 8160 2696 8216
rect 2376 8112 2696 8160
rect 2376 8056 2404 8112
rect 2460 8056 2508 8112
rect 2564 8056 2612 8112
rect 2668 8056 2696 8112
rect 2376 8008 2696 8056
rect 2376 7952 2404 8008
rect 2460 7952 2508 8008
rect 2564 7952 2612 8008
rect 2668 7952 2696 8008
rect 2376 7868 2696 7952
rect 2376 7812 2404 7868
rect 2460 7812 2508 7868
rect 2564 7812 2612 7868
rect 2668 7812 2696 7868
rect 2376 6300 2696 7812
rect 2772 17500 2828 17510
rect 2772 16156 2828 17444
rect 2772 13692 2828 16100
rect 2772 10556 2828 13636
rect 2772 8988 2828 10500
rect 2772 7308 2828 8932
rect 2772 7242 2828 7252
rect 3376 16492 3696 18004
rect 3376 16436 3404 16492
rect 3460 16436 3508 16492
rect 3564 16436 3612 16492
rect 3668 16436 3696 16492
rect 3376 14924 3696 16436
rect 3376 14868 3404 14924
rect 3460 14868 3508 14924
rect 3564 14868 3612 14924
rect 3668 14868 3696 14924
rect 3376 13356 3696 14868
rect 3376 13300 3404 13356
rect 3460 13300 3508 13356
rect 3564 13300 3612 13356
rect 3668 13300 3696 13356
rect 3376 11788 3696 13300
rect 3376 11732 3404 11788
rect 3460 11732 3508 11788
rect 3564 11732 3612 11788
rect 3668 11732 3696 11788
rect 3376 11716 3696 11732
rect 3376 11660 3404 11716
rect 3460 11660 3508 11716
rect 3564 11660 3612 11716
rect 3668 11660 3696 11716
rect 3376 11612 3696 11660
rect 3376 11556 3404 11612
rect 3460 11556 3508 11612
rect 3564 11556 3612 11612
rect 3668 11556 3696 11612
rect 3376 11508 3696 11556
rect 3376 11452 3404 11508
rect 3460 11452 3508 11508
rect 3564 11452 3612 11508
rect 3668 11452 3696 11508
rect 3376 10220 3696 11452
rect 3376 10164 3404 10220
rect 3460 10164 3508 10220
rect 3564 10164 3612 10220
rect 3668 10164 3696 10220
rect 3376 8652 3696 10164
rect 3892 21644 3948 21654
rect 3892 8988 3948 21588
rect 4004 21532 4060 21542
rect 4004 15372 4060 21476
rect 4004 15306 4060 15316
rect 4116 15260 4172 21812
rect 4376 20412 4696 21924
rect 4376 20356 4404 20412
rect 4460 20356 4508 20412
rect 4564 20356 4612 20412
rect 4668 20356 4696 20412
rect 4376 18844 4696 20356
rect 4376 18788 4404 18844
rect 4460 18788 4508 18844
rect 4564 18788 4612 18844
rect 4668 18788 4696 18844
rect 4116 15194 4172 15204
rect 4228 18060 4284 18070
rect 4116 13804 4172 13814
rect 4116 12796 4172 13748
rect 3892 8922 3948 8932
rect 4004 11004 4060 11014
rect 3376 8596 3404 8652
rect 3460 8596 3508 8652
rect 3564 8596 3612 8652
rect 3668 8596 3696 8652
rect 2376 6244 2404 6300
rect 2460 6244 2508 6300
rect 2564 6244 2612 6300
rect 2668 6244 2696 6300
rect 2376 4732 2696 6244
rect 2376 4676 2404 4732
rect 2460 4676 2508 4732
rect 2564 4676 2612 4732
rect 2668 4676 2696 4732
rect 2376 3164 2696 4676
rect 2376 3108 2404 3164
rect 2460 3108 2508 3164
rect 2564 3108 2612 3164
rect 2668 3108 2696 3164
rect 2376 1596 2696 3108
rect 2376 1540 2404 1596
rect 2460 1540 2508 1596
rect 2564 1540 2612 1596
rect 2668 1540 2696 1596
rect 2376 1216 2696 1540
rect 2376 1160 2404 1216
rect 2460 1160 2508 1216
rect 2564 1160 2612 1216
rect 2668 1160 2696 1216
rect 2376 1112 2696 1160
rect 2376 1056 2404 1112
rect 2460 1056 2508 1112
rect 2564 1056 2612 1112
rect 2668 1056 2696 1112
rect 2376 1008 2696 1056
rect 2376 952 2404 1008
rect 2460 952 2508 1008
rect 2564 952 2612 1008
rect 2668 952 2696 1008
rect 2376 724 2696 952
rect 3376 7084 3696 8596
rect 3376 7028 3404 7084
rect 3460 7028 3508 7084
rect 3564 7028 3612 7084
rect 3668 7028 3696 7084
rect 3376 5516 3696 7028
rect 3376 5460 3404 5516
rect 3460 5460 3508 5516
rect 3564 5460 3612 5516
rect 3668 5460 3696 5516
rect 3376 4716 3696 5460
rect 3376 4660 3404 4716
rect 3460 4660 3508 4716
rect 3564 4660 3612 4716
rect 3668 4660 3696 4716
rect 3376 4612 3696 4660
rect 3376 4556 3404 4612
rect 3460 4556 3508 4612
rect 3564 4556 3612 4612
rect 3668 4556 3696 4612
rect 3376 4508 3696 4556
rect 3376 4452 3404 4508
rect 3460 4452 3508 4508
rect 3564 4452 3612 4508
rect 3668 4452 3696 4508
rect 3376 3948 3696 4452
rect 4004 4172 4060 10948
rect 4116 9100 4172 12740
rect 4116 9034 4172 9044
rect 4228 6748 4284 18004
rect 4228 6682 4284 6692
rect 4376 17276 4696 18788
rect 4376 17220 4404 17276
rect 4460 17220 4508 17276
rect 4564 17220 4612 17276
rect 4668 17220 4696 17276
rect 4376 15708 4696 17220
rect 4788 27132 4844 27142
rect 4788 17836 4844 27076
rect 4900 26236 4956 29652
rect 4900 26170 4956 26180
rect 5012 27132 5068 29988
rect 5012 26012 5068 27076
rect 5124 29148 5180 29158
rect 5124 26124 5180 29092
rect 5376 29036 5696 30548
rect 5376 28980 5404 29036
rect 5460 28980 5508 29036
rect 5564 28980 5612 29036
rect 5668 28980 5696 29036
rect 5124 26058 5180 26068
rect 5236 27692 5292 27702
rect 5012 22876 5068 25956
rect 5236 23740 5292 27636
rect 5012 22810 5068 22820
rect 5124 23684 5292 23740
rect 5376 27468 5696 28980
rect 5376 27412 5404 27468
rect 5460 27412 5508 27468
rect 5564 27412 5612 27468
rect 5668 27412 5696 27468
rect 5376 25900 5696 27412
rect 5796 31836 5852 31846
rect 5796 26348 5852 31780
rect 5796 26282 5852 26292
rect 5376 25844 5404 25900
rect 5460 25844 5508 25900
rect 5564 25844 5612 25900
rect 5668 25844 5696 25900
rect 5376 25716 5696 25844
rect 5376 25660 5404 25716
rect 5460 25660 5508 25716
rect 5564 25660 5612 25716
rect 5668 25660 5696 25716
rect 5376 25612 5696 25660
rect 5376 25556 5404 25612
rect 5460 25556 5508 25612
rect 5564 25556 5612 25612
rect 5668 25556 5696 25612
rect 5376 25508 5696 25556
rect 5376 25452 5404 25508
rect 5460 25452 5508 25508
rect 5564 25452 5612 25508
rect 5668 25452 5696 25508
rect 5376 24332 5696 25452
rect 5376 24276 5404 24332
rect 5460 24276 5508 24332
rect 5564 24276 5612 24332
rect 5668 24276 5696 24332
rect 5124 21868 5180 23684
rect 4788 16044 4844 17780
rect 5012 21812 5180 21868
rect 5236 22876 5292 22886
rect 5012 16268 5068 21812
rect 5236 17708 5292 22820
rect 5012 16202 5068 16212
rect 5124 17652 5292 17708
rect 5376 22764 5696 24276
rect 5796 26124 5852 26134
rect 5796 23884 5852 26068
rect 5796 23818 5852 23828
rect 5376 22708 5404 22764
rect 5460 22708 5508 22764
rect 5564 22708 5612 22764
rect 5668 22708 5696 22764
rect 5376 21196 5696 22708
rect 5376 21140 5404 21196
rect 5460 21140 5508 21196
rect 5564 21140 5612 21196
rect 5668 21140 5696 21196
rect 5376 19628 5696 21140
rect 5908 23100 5964 23110
rect 5376 19572 5404 19628
rect 5460 19572 5508 19628
rect 5564 19572 5612 19628
rect 5668 19572 5696 19628
rect 5376 18716 5696 19572
rect 5376 18660 5404 18716
rect 5460 18660 5508 18716
rect 5564 18660 5612 18716
rect 5668 18660 5696 18716
rect 5376 18612 5696 18660
rect 5376 18556 5404 18612
rect 5460 18556 5508 18612
rect 5564 18556 5612 18612
rect 5668 18556 5696 18612
rect 5376 18508 5696 18556
rect 5376 18452 5404 18508
rect 5460 18452 5508 18508
rect 5564 18452 5612 18508
rect 5668 18452 5696 18508
rect 5376 18060 5696 18452
rect 5376 18004 5404 18060
rect 5460 18004 5508 18060
rect 5564 18004 5612 18060
rect 5668 18004 5696 18060
rect 5012 16044 5068 16054
rect 4788 15988 4956 16044
rect 4376 15652 4404 15708
rect 4460 15652 4508 15708
rect 4564 15652 4612 15708
rect 4668 15652 4696 15708
rect 4376 15216 4696 15652
rect 4376 15160 4404 15216
rect 4460 15160 4508 15216
rect 4564 15160 4612 15216
rect 4668 15160 4696 15216
rect 4376 15112 4696 15160
rect 4376 15056 4404 15112
rect 4460 15056 4508 15112
rect 4564 15056 4612 15112
rect 4668 15056 4696 15112
rect 4376 15008 4696 15056
rect 4376 14952 4404 15008
rect 4460 14952 4508 15008
rect 4564 14952 4612 15008
rect 4668 14952 4696 15008
rect 4376 14140 4696 14952
rect 4376 14084 4404 14140
rect 4460 14084 4508 14140
rect 4564 14084 4612 14140
rect 4668 14084 4696 14140
rect 4376 12572 4696 14084
rect 4788 15820 4844 15830
rect 4788 13916 4844 15764
rect 4900 14588 4956 15988
rect 4900 14522 4956 14532
rect 4788 13850 4844 13860
rect 4376 12516 4404 12572
rect 4460 12516 4508 12572
rect 4564 12516 4612 12572
rect 4668 12516 4696 12572
rect 4376 11004 4696 12516
rect 4376 10948 4404 11004
rect 4460 10948 4508 11004
rect 4564 10948 4612 11004
rect 4668 10948 4696 11004
rect 4376 9436 4696 10948
rect 4376 9380 4404 9436
rect 4460 9380 4508 9436
rect 4564 9380 4612 9436
rect 4668 9380 4696 9436
rect 4376 8216 4696 9380
rect 4376 8160 4404 8216
rect 4460 8160 4508 8216
rect 4564 8160 4612 8216
rect 4668 8160 4696 8216
rect 4376 8112 4696 8160
rect 4376 8056 4404 8112
rect 4460 8056 4508 8112
rect 4564 8056 4612 8112
rect 4668 8056 4696 8112
rect 4376 8008 4696 8056
rect 4376 7952 4404 8008
rect 4460 7952 4508 8008
rect 4564 7952 4612 8008
rect 4668 7952 4696 8008
rect 4376 7868 4696 7952
rect 4376 7812 4404 7868
rect 4460 7812 4508 7868
rect 4564 7812 4612 7868
rect 4668 7812 4696 7868
rect 4376 6300 4696 7812
rect 5012 6748 5068 15988
rect 5124 13244 5180 17652
rect 5376 16492 5696 18004
rect 5376 16436 5404 16492
rect 5460 16436 5508 16492
rect 5564 16436 5612 16492
rect 5668 16436 5696 16492
rect 5124 13178 5180 13188
rect 5236 16268 5292 16278
rect 5236 13132 5292 16212
rect 5236 13066 5292 13076
rect 5376 14924 5696 16436
rect 5376 14868 5404 14924
rect 5460 14868 5508 14924
rect 5564 14868 5612 14924
rect 5668 14868 5696 14924
rect 5376 13356 5696 14868
rect 5376 13300 5404 13356
rect 5460 13300 5508 13356
rect 5564 13300 5612 13356
rect 5668 13300 5696 13356
rect 5012 6682 5068 6692
rect 5376 11788 5696 13300
rect 5376 11732 5404 11788
rect 5460 11732 5508 11788
rect 5564 11732 5612 11788
rect 5668 11732 5696 11788
rect 5376 11716 5696 11732
rect 5376 11660 5404 11716
rect 5460 11660 5508 11716
rect 5564 11660 5612 11716
rect 5668 11660 5696 11716
rect 5376 11612 5696 11660
rect 5376 11556 5404 11612
rect 5460 11556 5508 11612
rect 5564 11556 5612 11612
rect 5668 11556 5696 11612
rect 5376 11508 5696 11556
rect 5376 11452 5404 11508
rect 5460 11452 5508 11508
rect 5564 11452 5612 11508
rect 5668 11452 5696 11508
rect 5376 10220 5696 11452
rect 5376 10164 5404 10220
rect 5460 10164 5508 10220
rect 5564 10164 5612 10220
rect 5668 10164 5696 10220
rect 5376 8652 5696 10164
rect 5796 19740 5852 19750
rect 5796 9100 5852 19684
rect 5908 15148 5964 23044
rect 5908 15082 5964 15092
rect 5796 9034 5852 9044
rect 5376 8596 5404 8652
rect 5460 8596 5508 8652
rect 5564 8596 5612 8652
rect 5668 8596 5696 8652
rect 5376 7084 5696 8596
rect 5376 7028 5404 7084
rect 5460 7028 5508 7084
rect 5564 7028 5612 7084
rect 5668 7028 5696 7084
rect 4376 6244 4404 6300
rect 4460 6244 4508 6300
rect 4564 6244 4612 6300
rect 4668 6244 4696 6300
rect 4376 4732 4696 6244
rect 4376 4676 4404 4732
rect 4460 4676 4508 4732
rect 4564 4676 4612 4732
rect 4668 4676 4696 4732
rect 4004 4106 4060 4116
rect 4228 4396 4284 4406
rect 3376 3892 3404 3948
rect 3460 3892 3508 3948
rect 3564 3892 3612 3948
rect 3668 3892 3696 3948
rect 3376 2380 3696 3892
rect 4228 2828 4284 4340
rect 4228 2762 4284 2772
rect 4376 3164 4696 4676
rect 4376 3108 4404 3164
rect 4460 3108 4508 3164
rect 4564 3108 4612 3164
rect 4668 3108 4696 3164
rect 3376 2324 3404 2380
rect 3460 2324 3508 2380
rect 3564 2324 3612 2380
rect 3668 2324 3696 2380
rect 3376 812 3696 2324
rect 3376 756 3404 812
rect 3460 756 3508 812
rect 3564 756 3612 812
rect 3668 756 3696 812
rect 3376 724 3696 756
rect 4376 1596 4696 3108
rect 4376 1540 4404 1596
rect 4460 1540 4508 1596
rect 4564 1540 4612 1596
rect 4668 1540 4696 1596
rect 4376 1216 4696 1540
rect 4376 1160 4404 1216
rect 4460 1160 4508 1216
rect 4564 1160 4612 1216
rect 4668 1160 4696 1216
rect 4376 1112 4696 1160
rect 4376 1056 4404 1112
rect 4460 1056 4508 1112
rect 4564 1056 4612 1112
rect 4668 1056 4696 1112
rect 4376 1008 4696 1056
rect 4376 952 4404 1008
rect 4460 952 4508 1008
rect 4564 952 4612 1008
rect 4668 952 4696 1008
rect 4376 724 4696 952
rect 5376 5516 5696 7028
rect 5376 5460 5404 5516
rect 5460 5460 5508 5516
rect 5564 5460 5612 5516
rect 5668 5460 5696 5516
rect 5376 4716 5696 5460
rect 5376 4660 5404 4716
rect 5460 4660 5508 4716
rect 5564 4660 5612 4716
rect 5668 4660 5696 4716
rect 5376 4612 5696 4660
rect 5376 4556 5404 4612
rect 5460 4556 5508 4612
rect 5564 4556 5612 4612
rect 5668 4556 5696 4612
rect 5376 4508 5696 4556
rect 5376 4452 5404 4508
rect 5460 4452 5508 4508
rect 5564 4452 5612 4508
rect 5668 4452 5696 4508
rect 5376 3948 5696 4452
rect 5376 3892 5404 3948
rect 5460 3892 5508 3948
rect 5564 3892 5612 3948
rect 5668 3892 5696 3948
rect 5376 2380 5696 3892
rect 5376 2324 5404 2380
rect 5460 2324 5508 2380
rect 5564 2324 5612 2380
rect 5668 2324 5696 2380
rect 5376 812 5696 2324
rect 5376 756 5404 812
rect 5460 756 5508 812
rect 5564 756 5612 812
rect 5668 756 5696 812
rect 5376 724 5696 756
<< via4 >>
rect 404 29160 460 29216
rect 508 29160 564 29216
rect 612 29160 668 29216
rect 404 29056 460 29112
rect 508 29056 564 29112
rect 612 29056 668 29112
rect 404 28952 460 29008
rect 508 28952 564 29008
rect 612 28952 668 29008
rect 404 22160 460 22216
rect 508 22160 564 22216
rect 612 22160 668 22216
rect 404 22056 460 22112
rect 508 22056 564 22112
rect 612 22056 668 22112
rect 404 21980 460 22008
rect 404 21952 460 21980
rect 508 21980 564 22008
rect 508 21952 564 21980
rect 612 21980 668 22008
rect 612 21952 668 21980
rect 1404 32660 1460 32716
rect 1508 32660 1564 32716
rect 1612 32660 1668 32716
rect 1404 32556 1460 32612
rect 1508 32556 1564 32612
rect 1612 32556 1668 32612
rect 1404 32452 1460 32508
rect 1508 32452 1564 32508
rect 1612 32452 1668 32508
rect 1404 25660 1460 25716
rect 1508 25660 1564 25716
rect 1612 25660 1668 25716
rect 1404 25556 1460 25612
rect 1508 25556 1564 25612
rect 1612 25556 1668 25612
rect 1404 25452 1460 25508
rect 1508 25452 1564 25508
rect 1612 25452 1668 25508
rect 404 15160 460 15216
rect 508 15160 564 15216
rect 612 15160 668 15216
rect 404 15056 460 15112
rect 508 15056 564 15112
rect 612 15056 668 15112
rect 404 14952 460 15008
rect 508 14952 564 15008
rect 612 14952 668 15008
rect 404 8160 460 8216
rect 508 8160 564 8216
rect 612 8160 668 8216
rect 404 8056 460 8112
rect 508 8056 564 8112
rect 612 8056 668 8112
rect 404 7952 460 8008
rect 508 7952 564 8008
rect 612 7952 668 8008
rect 2404 29160 2460 29216
rect 2508 29160 2564 29216
rect 2612 29160 2668 29216
rect 2404 29056 2460 29112
rect 2508 29056 2564 29112
rect 2612 29056 2668 29112
rect 2404 28952 2460 29008
rect 2508 28952 2564 29008
rect 2612 28952 2668 29008
rect 2404 22160 2460 22216
rect 2508 22160 2564 22216
rect 2612 22160 2668 22216
rect 2404 22056 2460 22112
rect 2508 22056 2564 22112
rect 2612 22056 2668 22112
rect 2404 21980 2460 22008
rect 2404 21952 2460 21980
rect 2508 21980 2564 22008
rect 2508 21952 2564 21980
rect 2612 21980 2668 22008
rect 2612 21952 2668 21980
rect 1404 18660 1460 18716
rect 1508 18660 1564 18716
rect 1612 18660 1668 18716
rect 1404 18556 1460 18612
rect 1508 18556 1564 18612
rect 1612 18556 1668 18612
rect 1404 18452 1460 18508
rect 1508 18452 1564 18508
rect 1612 18452 1668 18508
rect 3404 32660 3460 32716
rect 3508 32660 3564 32716
rect 3612 32660 3668 32716
rect 3404 32556 3460 32612
rect 3508 32556 3564 32612
rect 3612 32556 3668 32612
rect 3404 32452 3460 32508
rect 3508 32452 3564 32508
rect 3612 32452 3668 32508
rect 3404 25660 3460 25716
rect 3508 25660 3564 25716
rect 3612 25660 3668 25716
rect 3404 25556 3460 25612
rect 3508 25556 3564 25612
rect 3612 25556 3668 25612
rect 3404 25452 3460 25508
rect 3508 25452 3564 25508
rect 3612 25452 3668 25508
rect 5404 32660 5460 32716
rect 5508 32660 5564 32716
rect 5612 32660 5668 32716
rect 5404 32556 5460 32612
rect 5508 32556 5564 32612
rect 5612 32556 5668 32612
rect 5404 32452 5460 32508
rect 5508 32452 5564 32508
rect 5612 32452 5668 32508
rect 4404 29160 4460 29216
rect 4508 29160 4564 29216
rect 4612 29160 4668 29216
rect 4404 29056 4460 29112
rect 4508 29056 4564 29112
rect 4612 29056 4668 29112
rect 4404 28952 4460 29008
rect 4508 28952 4564 29008
rect 4612 28952 4668 29008
rect 4404 22160 4460 22216
rect 4508 22160 4564 22216
rect 4612 22160 4668 22216
rect 4404 22056 4460 22112
rect 4508 22056 4564 22112
rect 4612 22056 4668 22112
rect 4404 21980 4460 22008
rect 4404 21952 4460 21980
rect 4508 21980 4564 22008
rect 4508 21952 4564 21980
rect 4612 21980 4668 22008
rect 4612 21952 4668 21980
rect 3404 18660 3460 18716
rect 3508 18660 3564 18716
rect 3612 18660 3668 18716
rect 3404 18556 3460 18612
rect 3508 18556 3564 18612
rect 3612 18556 3668 18612
rect 3404 18452 3460 18508
rect 3508 18452 3564 18508
rect 3612 18452 3668 18508
rect 2404 15160 2460 15216
rect 2508 15160 2564 15216
rect 2612 15160 2668 15216
rect 2404 15056 2460 15112
rect 2508 15056 2564 15112
rect 2612 15056 2668 15112
rect 2404 14952 2460 15008
rect 2508 14952 2564 15008
rect 2612 14952 2668 15008
rect 1404 11660 1460 11716
rect 1508 11660 1564 11716
rect 1612 11660 1668 11716
rect 1404 11556 1460 11612
rect 1508 11556 1564 11612
rect 1612 11556 1668 11612
rect 1404 11452 1460 11508
rect 1508 11452 1564 11508
rect 1612 11452 1668 11508
rect 404 1160 460 1216
rect 508 1160 564 1216
rect 612 1160 668 1216
rect 404 1056 460 1112
rect 508 1056 564 1112
rect 612 1056 668 1112
rect 404 952 460 1008
rect 508 952 564 1008
rect 612 952 668 1008
rect 1404 4660 1460 4716
rect 1508 4660 1564 4716
rect 1612 4660 1668 4716
rect 1404 4556 1460 4612
rect 1508 4556 1564 4612
rect 1612 4556 1668 4612
rect 1404 4452 1460 4508
rect 1508 4452 1564 4508
rect 1612 4452 1668 4508
rect 2404 8160 2460 8216
rect 2508 8160 2564 8216
rect 2612 8160 2668 8216
rect 2404 8056 2460 8112
rect 2508 8056 2564 8112
rect 2612 8056 2668 8112
rect 2404 7952 2460 8008
rect 2508 7952 2564 8008
rect 2612 7952 2668 8008
rect 3404 11660 3460 11716
rect 3508 11660 3564 11716
rect 3612 11660 3668 11716
rect 3404 11556 3460 11612
rect 3508 11556 3564 11612
rect 3612 11556 3668 11612
rect 3404 11452 3460 11508
rect 3508 11452 3564 11508
rect 3612 11452 3668 11508
rect 2404 1160 2460 1216
rect 2508 1160 2564 1216
rect 2612 1160 2668 1216
rect 2404 1056 2460 1112
rect 2508 1056 2564 1112
rect 2612 1056 2668 1112
rect 2404 952 2460 1008
rect 2508 952 2564 1008
rect 2612 952 2668 1008
rect 3404 4660 3460 4716
rect 3508 4660 3564 4716
rect 3612 4660 3668 4716
rect 3404 4556 3460 4612
rect 3508 4556 3564 4612
rect 3612 4556 3668 4612
rect 3404 4452 3460 4508
rect 3508 4452 3564 4508
rect 3612 4452 3668 4508
rect 5404 25660 5460 25716
rect 5508 25660 5564 25716
rect 5612 25660 5668 25716
rect 5404 25556 5460 25612
rect 5508 25556 5564 25612
rect 5612 25556 5668 25612
rect 5404 25452 5460 25508
rect 5508 25452 5564 25508
rect 5612 25452 5668 25508
rect 5404 18660 5460 18716
rect 5508 18660 5564 18716
rect 5612 18660 5668 18716
rect 5404 18556 5460 18612
rect 5508 18556 5564 18612
rect 5612 18556 5668 18612
rect 5404 18452 5460 18508
rect 5508 18452 5564 18508
rect 5612 18452 5668 18508
rect 4404 15160 4460 15216
rect 4508 15160 4564 15216
rect 4612 15160 4668 15216
rect 4404 15056 4460 15112
rect 4508 15056 4564 15112
rect 4612 15056 4668 15112
rect 4404 14952 4460 15008
rect 4508 14952 4564 15008
rect 4612 14952 4668 15008
rect 4404 8160 4460 8216
rect 4508 8160 4564 8216
rect 4612 8160 4668 8216
rect 4404 8056 4460 8112
rect 4508 8056 4564 8112
rect 4612 8056 4668 8112
rect 4404 7952 4460 8008
rect 4508 7952 4564 8008
rect 4612 7952 4668 8008
rect 5404 11660 5460 11716
rect 5508 11660 5564 11716
rect 5612 11660 5668 11716
rect 5404 11556 5460 11612
rect 5508 11556 5564 11612
rect 5612 11556 5668 11612
rect 5404 11452 5460 11508
rect 5508 11452 5564 11508
rect 5612 11452 5668 11508
rect 4404 1160 4460 1216
rect 4508 1160 4564 1216
rect 4612 1160 4668 1216
rect 4404 1056 4460 1112
rect 4508 1056 4564 1112
rect 4612 1056 4668 1112
rect 4404 952 4460 1008
rect 4508 952 4564 1008
rect 4612 952 4668 1008
rect 5404 4660 5460 4716
rect 5508 4660 5564 4716
rect 5612 4660 5668 4716
rect 5404 4556 5460 4612
rect 5508 4556 5564 4612
rect 5612 4556 5668 4612
rect 5404 4452 5460 4508
rect 5508 4452 5564 4508
rect 5612 4452 5668 4508
<< metal5 >>
rect 276 32716 5696 32744
rect 276 32660 1404 32716
rect 1460 32660 1508 32716
rect 1564 32660 1612 32716
rect 1668 32660 3404 32716
rect 3460 32660 3508 32716
rect 3564 32660 3612 32716
rect 3668 32660 5404 32716
rect 5460 32660 5508 32716
rect 5564 32660 5612 32716
rect 5668 32660 5696 32716
rect 276 32612 5696 32660
rect 276 32556 1404 32612
rect 1460 32556 1508 32612
rect 1564 32556 1612 32612
rect 1668 32556 3404 32612
rect 3460 32556 3508 32612
rect 3564 32556 3612 32612
rect 3668 32556 5404 32612
rect 5460 32556 5508 32612
rect 5564 32556 5612 32612
rect 5668 32556 5696 32612
rect 276 32508 5696 32556
rect 276 32452 1404 32508
rect 1460 32452 1508 32508
rect 1564 32452 1612 32508
rect 1668 32452 3404 32508
rect 3460 32452 3508 32508
rect 3564 32452 3612 32508
rect 3668 32452 5404 32508
rect 5460 32452 5508 32508
rect 5564 32452 5612 32508
rect 5668 32452 5696 32508
rect 276 32424 5696 32452
rect 276 29216 5660 29244
rect 276 29160 404 29216
rect 460 29160 508 29216
rect 564 29160 612 29216
rect 668 29160 2404 29216
rect 2460 29160 2508 29216
rect 2564 29160 2612 29216
rect 2668 29160 4404 29216
rect 4460 29160 4508 29216
rect 4564 29160 4612 29216
rect 4668 29160 5660 29216
rect 276 29112 5660 29160
rect 276 29056 404 29112
rect 460 29056 508 29112
rect 564 29056 612 29112
rect 668 29056 2404 29112
rect 2460 29056 2508 29112
rect 2564 29056 2612 29112
rect 2668 29056 4404 29112
rect 4460 29056 4508 29112
rect 4564 29056 4612 29112
rect 4668 29056 5660 29112
rect 276 29008 5660 29056
rect 276 28952 404 29008
rect 460 28952 508 29008
rect 564 28952 612 29008
rect 668 28952 2404 29008
rect 2460 28952 2508 29008
rect 2564 28952 2612 29008
rect 2668 28952 4404 29008
rect 4460 28952 4508 29008
rect 4564 28952 4612 29008
rect 4668 28952 5660 29008
rect 276 28924 5660 28952
rect 276 25716 5696 25744
rect 276 25660 1404 25716
rect 1460 25660 1508 25716
rect 1564 25660 1612 25716
rect 1668 25660 3404 25716
rect 3460 25660 3508 25716
rect 3564 25660 3612 25716
rect 3668 25660 5404 25716
rect 5460 25660 5508 25716
rect 5564 25660 5612 25716
rect 5668 25660 5696 25716
rect 276 25612 5696 25660
rect 276 25556 1404 25612
rect 1460 25556 1508 25612
rect 1564 25556 1612 25612
rect 1668 25556 3404 25612
rect 3460 25556 3508 25612
rect 3564 25556 3612 25612
rect 3668 25556 5404 25612
rect 5460 25556 5508 25612
rect 5564 25556 5612 25612
rect 5668 25556 5696 25612
rect 276 25508 5696 25556
rect 276 25452 1404 25508
rect 1460 25452 1508 25508
rect 1564 25452 1612 25508
rect 1668 25452 3404 25508
rect 3460 25452 3508 25508
rect 3564 25452 3612 25508
rect 3668 25452 5404 25508
rect 5460 25452 5508 25508
rect 5564 25452 5612 25508
rect 5668 25452 5696 25508
rect 276 25424 5696 25452
rect 276 22216 5660 22244
rect 276 22160 404 22216
rect 460 22160 508 22216
rect 564 22160 612 22216
rect 668 22160 2404 22216
rect 2460 22160 2508 22216
rect 2564 22160 2612 22216
rect 2668 22160 4404 22216
rect 4460 22160 4508 22216
rect 4564 22160 4612 22216
rect 4668 22160 5660 22216
rect 276 22112 5660 22160
rect 276 22056 404 22112
rect 460 22056 508 22112
rect 564 22056 612 22112
rect 668 22056 2404 22112
rect 2460 22056 2508 22112
rect 2564 22056 2612 22112
rect 2668 22056 4404 22112
rect 4460 22056 4508 22112
rect 4564 22056 4612 22112
rect 4668 22056 5660 22112
rect 276 22008 5660 22056
rect 276 21952 404 22008
rect 460 21952 508 22008
rect 564 21952 612 22008
rect 668 21952 2404 22008
rect 2460 21952 2508 22008
rect 2564 21952 2612 22008
rect 2668 21952 4404 22008
rect 4460 21952 4508 22008
rect 4564 21952 4612 22008
rect 4668 21952 5660 22008
rect 276 21924 5660 21952
rect 276 18716 5696 18744
rect 276 18660 1404 18716
rect 1460 18660 1508 18716
rect 1564 18660 1612 18716
rect 1668 18660 3404 18716
rect 3460 18660 3508 18716
rect 3564 18660 3612 18716
rect 3668 18660 5404 18716
rect 5460 18660 5508 18716
rect 5564 18660 5612 18716
rect 5668 18660 5696 18716
rect 276 18612 5696 18660
rect 276 18556 1404 18612
rect 1460 18556 1508 18612
rect 1564 18556 1612 18612
rect 1668 18556 3404 18612
rect 3460 18556 3508 18612
rect 3564 18556 3612 18612
rect 3668 18556 5404 18612
rect 5460 18556 5508 18612
rect 5564 18556 5612 18612
rect 5668 18556 5696 18612
rect 276 18508 5696 18556
rect 276 18452 1404 18508
rect 1460 18452 1508 18508
rect 1564 18452 1612 18508
rect 1668 18452 3404 18508
rect 3460 18452 3508 18508
rect 3564 18452 3612 18508
rect 3668 18452 5404 18508
rect 5460 18452 5508 18508
rect 5564 18452 5612 18508
rect 5668 18452 5696 18508
rect 276 18424 5696 18452
rect 276 15216 5660 15244
rect 276 15160 404 15216
rect 460 15160 508 15216
rect 564 15160 612 15216
rect 668 15160 2404 15216
rect 2460 15160 2508 15216
rect 2564 15160 2612 15216
rect 2668 15160 4404 15216
rect 4460 15160 4508 15216
rect 4564 15160 4612 15216
rect 4668 15160 5660 15216
rect 276 15112 5660 15160
rect 276 15056 404 15112
rect 460 15056 508 15112
rect 564 15056 612 15112
rect 668 15056 2404 15112
rect 2460 15056 2508 15112
rect 2564 15056 2612 15112
rect 2668 15056 4404 15112
rect 4460 15056 4508 15112
rect 4564 15056 4612 15112
rect 4668 15056 5660 15112
rect 276 15008 5660 15056
rect 276 14952 404 15008
rect 460 14952 508 15008
rect 564 14952 612 15008
rect 668 14952 2404 15008
rect 2460 14952 2508 15008
rect 2564 14952 2612 15008
rect 2668 14952 4404 15008
rect 4460 14952 4508 15008
rect 4564 14952 4612 15008
rect 4668 14952 5660 15008
rect 276 14924 5660 14952
rect 276 11716 5696 11744
rect 276 11660 1404 11716
rect 1460 11660 1508 11716
rect 1564 11660 1612 11716
rect 1668 11660 3404 11716
rect 3460 11660 3508 11716
rect 3564 11660 3612 11716
rect 3668 11660 5404 11716
rect 5460 11660 5508 11716
rect 5564 11660 5612 11716
rect 5668 11660 5696 11716
rect 276 11612 5696 11660
rect 276 11556 1404 11612
rect 1460 11556 1508 11612
rect 1564 11556 1612 11612
rect 1668 11556 3404 11612
rect 3460 11556 3508 11612
rect 3564 11556 3612 11612
rect 3668 11556 5404 11612
rect 5460 11556 5508 11612
rect 5564 11556 5612 11612
rect 5668 11556 5696 11612
rect 276 11508 5696 11556
rect 276 11452 1404 11508
rect 1460 11452 1508 11508
rect 1564 11452 1612 11508
rect 1668 11452 3404 11508
rect 3460 11452 3508 11508
rect 3564 11452 3612 11508
rect 3668 11452 5404 11508
rect 5460 11452 5508 11508
rect 5564 11452 5612 11508
rect 5668 11452 5696 11508
rect 276 11424 5696 11452
rect 276 8216 5660 8244
rect 276 8160 404 8216
rect 460 8160 508 8216
rect 564 8160 612 8216
rect 668 8160 2404 8216
rect 2460 8160 2508 8216
rect 2564 8160 2612 8216
rect 2668 8160 4404 8216
rect 4460 8160 4508 8216
rect 4564 8160 4612 8216
rect 4668 8160 5660 8216
rect 276 8112 5660 8160
rect 276 8056 404 8112
rect 460 8056 508 8112
rect 564 8056 612 8112
rect 668 8056 2404 8112
rect 2460 8056 2508 8112
rect 2564 8056 2612 8112
rect 2668 8056 4404 8112
rect 4460 8056 4508 8112
rect 4564 8056 4612 8112
rect 4668 8056 5660 8112
rect 276 8008 5660 8056
rect 276 7952 404 8008
rect 460 7952 508 8008
rect 564 7952 612 8008
rect 668 7952 2404 8008
rect 2460 7952 2508 8008
rect 2564 7952 2612 8008
rect 2668 7952 4404 8008
rect 4460 7952 4508 8008
rect 4564 7952 4612 8008
rect 4668 7952 5660 8008
rect 276 7924 5660 7952
rect 276 4716 5696 4744
rect 276 4660 1404 4716
rect 1460 4660 1508 4716
rect 1564 4660 1612 4716
rect 1668 4660 3404 4716
rect 3460 4660 3508 4716
rect 3564 4660 3612 4716
rect 3668 4660 5404 4716
rect 5460 4660 5508 4716
rect 5564 4660 5612 4716
rect 5668 4660 5696 4716
rect 276 4612 5696 4660
rect 276 4556 1404 4612
rect 1460 4556 1508 4612
rect 1564 4556 1612 4612
rect 1668 4556 3404 4612
rect 3460 4556 3508 4612
rect 3564 4556 3612 4612
rect 3668 4556 5404 4612
rect 5460 4556 5508 4612
rect 5564 4556 5612 4612
rect 5668 4556 5696 4612
rect 276 4508 5696 4556
rect 276 4452 1404 4508
rect 1460 4452 1508 4508
rect 1564 4452 1612 4508
rect 1668 4452 3404 4508
rect 3460 4452 3508 4508
rect 3564 4452 3612 4508
rect 3668 4452 5404 4508
rect 5460 4452 5508 4508
rect 5564 4452 5612 4508
rect 5668 4452 5696 4508
rect 276 4424 5696 4452
rect 276 1216 5660 1244
rect 276 1160 404 1216
rect 460 1160 508 1216
rect 564 1160 612 1216
rect 668 1160 2404 1216
rect 2460 1160 2508 1216
rect 2564 1160 2612 1216
rect 2668 1160 4404 1216
rect 4460 1160 4508 1216
rect 4564 1160 4612 1216
rect 4668 1160 5660 1216
rect 276 1112 5660 1160
rect 276 1056 404 1112
rect 460 1056 508 1112
rect 564 1056 612 1112
rect 668 1056 2404 1112
rect 2460 1056 2508 1112
rect 2564 1056 2612 1112
rect 2668 1056 4404 1112
rect 4460 1056 4508 1112
rect 4564 1056 4612 1112
rect 4668 1056 5660 1112
rect 276 1008 5660 1056
rect 276 952 404 1008
rect 460 952 508 1008
rect 564 952 612 1008
rect 668 952 2404 1008
rect 2460 952 2508 1008
rect 2564 952 2612 1008
rect 2668 952 4404 1008
rect 4460 952 4508 1008
rect 4564 952 4612 1008
rect 4668 952 5660 1008
rect 276 924 5660 952
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__A2 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 3808 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__047__I
timestamp 1654395037
transform 1 0 5152 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I0
timestamp 1654395037
transform -1 0 4032 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I1
timestamp 1654395037
transform -1 0 5376 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1654395037
transform 1 0 1904 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__A2
timestamp 1654395037
transform -1 0 5376 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1654395037
transform 1 0 2240 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__A2
timestamp 1654395037
transform -1 0 3472 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__A2
timestamp 1654395037
transform 1 0 5152 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__A2
timestamp 1654395037
transform -1 0 4144 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__A2
timestamp 1654395037
transform -1 0 5376 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__A2
timestamp 1654395037
transform -1 0 3920 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__A2
timestamp 1654395037
transform 1 0 5152 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__A2
timestamp 1654395037
transform 1 0 4928 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__A2
timestamp 1654395037
transform 1 0 5152 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__A2
timestamp 1654395037
transform -1 0 2352 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1654395037
transform 1 0 2128 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__A2
timestamp 1654395037
transform -1 0 5376 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__A2
timestamp 1654395037
transform -1 0 1792 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__A2
timestamp 1654395037
transform -1 0 4704 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__A2
timestamp 1654395037
transform -1 0 2128 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__A2
timestamp 1654395037
transform 1 0 5152 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__A2
timestamp 1654395037
transform 1 0 3472 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__A2
timestamp 1654395037
transform 1 0 5152 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__A2
timestamp 1654395037
transform -1 0 5152 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__A2
timestamp 1654395037
transform -1 0 5376 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__A2
timestamp 1654395037
transform -1 0 2464 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__CLK
timestamp 1654395037
transform 1 0 5152 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__CLK
timestamp 1654395037
transform 1 0 5152 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__CLK
timestamp 1654395037
transform 1 0 4480 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__CLK
timestamp 1654395037
transform 1 0 5152 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__CLK
timestamp 1654395037
transform 1 0 5152 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__CLK
timestamp 1654395037
transform 1 0 5152 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__CLK
timestamp 1654395037
transform 1 0 5152 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__CLK
timestamp 1654395037
transform 1 0 5152 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__CLK
timestamp 1654395037
transform 1 0 5152 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__CLK
timestamp 1654395037
transform 1 0 5152 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__CLK
timestamp 1654395037
transform 1 0 3472 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__D
timestamp 1654395037
transform 1 0 4144 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__RN
timestamp 1654395037
transform 1 0 4368 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__CLK
timestamp 1654395037
transform 1 0 4592 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__RN
timestamp 1654395037
transform 1 0 3920 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__CLK
timestamp 1654395037
transform 1 0 4144 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__RN
timestamp 1654395037
transform 1 0 5152 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__CLK
timestamp 1654395037
transform 1 0 3136 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__RN
timestamp 1654395037
transform 1 0 5152 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__CLK
timestamp 1654395037
transform 1 0 4592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__RN
timestamp 1654395037
transform 1 0 4368 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__CLK
timestamp 1654395037
transform 1 0 4592 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__RN
timestamp 1654395037
transform 1 0 4368 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__CLK
timestamp 1654395037
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__RN
timestamp 1654395037
transform 1 0 4368 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__CLK
timestamp 1654395037
transform 1 0 4592 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__RN
timestamp 1654395037
transform 1 0 4368 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__CLK
timestamp 1654395037
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__RN
timestamp 1654395037
transform 1 0 4368 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__CLK
timestamp 1654395037
transform -1 0 4816 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__RN
timestamp 1654395037
transform 1 0 4368 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__I
timestamp 1654395037
transform 1 0 3360 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__I
timestamp 1654395037
transform -1 0 2464 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__I
timestamp 1654395037
transform 1 0 5040 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__I
timestamp 1654395037
transform 1 0 2912 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__I
timestamp 1654395037
transform 1 0 4928 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 560 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4144 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_38 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4592 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4816 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_43
timestamp 1654395037
transform 1 0 5152 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1654395037
transform 1 0 560 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_6
timestamp 1654395037
transform 1 0 1008 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_8
timestamp 1654395037
transform 1 0 1232 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_15
timestamp 1654395037
transform 1 0 2016 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_19 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 2464 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_35 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4256 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_43
timestamp 1654395037
transform 1 0 5152 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_2
timestamp 1654395037
transform 1 0 560 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_4
timestamp 1654395037
transform 1 0 784 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_25
timestamp 1654395037
transform 1 0 3136 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_32
timestamp 1654395037
transform 1 0 3920 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_40
timestamp 1654395037
transform 1 0 4816 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_43
timestamp 1654395037
transform 1 0 5152 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_44
timestamp 1654395037
transform 1 0 5264 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_40
timestamp 1654395037
transform 1 0 4816 0 1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_43
timestamp 1654395037
transform 1 0 5152 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_40
timestamp 1654395037
transform 1 0 4816 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_44
timestamp 1654395037
transform 1 0 5264 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_40
timestamp 1654395037
transform 1 0 4816 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_43
timestamp 1654395037
transform 1 0 5152 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1654395037
transform 1 0 560 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_34
timestamp 1654395037
transform 1 0 4144 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_42
timestamp 1654395037
transform 1 0 5040 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_2
timestamp 1654395037
transform 1 0 560 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_18
timestamp 1654395037
transform 1 0 2352 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_26
timestamp 1654395037
transform 1 0 3248 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_2
timestamp 1654395037
transform 1 0 560 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1654395037
transform 1 0 560 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_10
timestamp 1654395037
transform 1 0 1456 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_14
timestamp 1654395037
transform 1 0 1904 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_16
timestamp 1654395037
transform 1 0 2128 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_40
timestamp 1654395037
transform 1 0 4816 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_2
timestamp 1654395037
transform 1 0 560 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_18
timestamp 1654395037
transform 1 0 2352 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_12_22
timestamp 1654395037
transform 1 0 2800 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_2
timestamp 1654395037
transform 1 0 560 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_10
timestamp 1654395037
transform 1 0 1456 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_2
timestamp 1654395037
transform 1 0 560 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_10
timestamp 1654395037
transform 1 0 1456 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_2
timestamp 1654395037
transform 1 0 560 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_10
timestamp 1654395037
transform 1 0 1456 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_17_14
timestamp 1654395037
transform 1 0 1904 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_17_24
timestamp 1654395037
transform 1 0 3024 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_2
timestamp 1654395037
transform 1 0 560 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_10
timestamp 1654395037
transform 1 0 1456 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_2
timestamp 1654395037
transform 1 0 560 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_10
timestamp 1654395037
transform 1 0 1456 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_20_14
timestamp 1654395037
transform 1 0 1904 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_2
timestamp 1654395037
transform 1 0 560 0 -1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_18
timestamp 1654395037
transform 1 0 2352 0 -1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_25
timestamp 1654395037
transform 1 0 3136 0 -1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_2
timestamp 1654395037
transform 1 0 560 0 1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_18
timestamp 1654395037
transform 1 0 2352 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_26
timestamp 1654395037
transform 1 0 3248 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_30
timestamp 1654395037
transform 1 0 3696 0 1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_2
timestamp 1654395037
transform 1 0 560 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_10
timestamp 1654395037
transform 1 0 1456 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_23_14
timestamp 1654395037
transform 1 0 1904 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_16
timestamp 1654395037
transform 1 0 2128 0 -1 19600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_23
timestamp 1654395037
transform 1 0 2912 0 -1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_2
timestamp 1654395037
transform 1 0 560 0 1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_24_18
timestamp 1654395037
transform 1 0 2352 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_20
timestamp 1654395037
transform 1 0 2576 0 1 19600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_27
timestamp 1654395037
transform 1 0 3360 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_24_31
timestamp 1654395037
transform 1 0 3808 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_33
timestamp 1654395037
transform 1 0 4032 0 1 19600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_40
timestamp 1654395037
transform 1 0 4816 0 1 19600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_2
timestamp 1654395037
transform 1 0 560 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_2
timestamp 1654395037
transform 1 0 560 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_10
timestamp 1654395037
transform 1 0 1456 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_40
timestamp 1654395037
transform 1 0 4816 0 -1 24304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1654395037
transform 1 0 560 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_30_34
timestamp 1654395037
transform 1 0 4144 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_40
timestamp 1654395037
transform 1 0 4816 0 1 24304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_2
timestamp 1654395037
transform 1 0 560 0 -1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_18
timestamp 1654395037
transform 1 0 2352 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_26
timestamp 1654395037
transform 1 0 3248 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_31_30
timestamp 1654395037
transform 1 0 3696 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_2
timestamp 1654395037
transform 1 0 560 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_18
timestamp 1654395037
transform 1 0 2352 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_32_22
timestamp 1654395037
transform 1 0 2800 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_24
timestamp 1654395037
transform 1 0 3024 0 1 25872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_44
timestamp 1654395037
transform 1 0 5264 0 -1 27440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_2
timestamp 1654395037
transform 1 0 560 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_36
timestamp 1654395037
transform 1 0 4368 0 -1 30576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_36
timestamp 1654395037
transform 1 0 4368 0 -1 32144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_2
timestamp 1654395037
transform 1 0 560 0 1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_18
timestamp 1654395037
transform 1 0 2352 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_2
timestamp 1654395037
transform 1 0 560 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_40
timestamp 1654395037
transform 1 0 4816 0 -1 33712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 336 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1654395037
transform -1 0 5600 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1654395037
transform 1 0 336 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1654395037
transform -1 0 5600 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1654395037
transform 1 0 336 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1654395037
transform -1 0 5600 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1654395037
transform 1 0 336 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1654395037
transform -1 0 5600 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1654395037
transform 1 0 336 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1654395037
transform -1 0 5600 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1654395037
transform 1 0 336 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1654395037
transform -1 0 5600 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1654395037
transform 1 0 336 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1654395037
transform -1 0 5600 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1654395037
transform 1 0 336 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1654395037
transform -1 0 5600 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1654395037
transform 1 0 336 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1654395037
transform -1 0 5600 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1654395037
transform 1 0 336 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1654395037
transform -1 0 5600 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1654395037
transform 1 0 336 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1654395037
transform -1 0 5600 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1654395037
transform 1 0 336 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1654395037
transform -1 0 5600 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1654395037
transform 1 0 336 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1654395037
transform -1 0 5600 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1654395037
transform 1 0 336 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1654395037
transform -1 0 5600 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1654395037
transform 1 0 336 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1654395037
transform -1 0 5600 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1654395037
transform 1 0 336 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1654395037
transform -1 0 5600 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1654395037
transform 1 0 336 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1654395037
transform -1 0 5600 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1654395037
transform 1 0 336 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1654395037
transform -1 0 5600 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1654395037
transform 1 0 336 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1654395037
transform -1 0 5600 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1654395037
transform 1 0 336 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1654395037
transform -1 0 5600 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1654395037
transform 1 0 336 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1654395037
transform -1 0 5600 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1654395037
transform 1 0 336 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1654395037
transform -1 0 5600 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1654395037
transform 1 0 336 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1654395037
transform -1 0 5600 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1654395037
transform 1 0 336 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1654395037
transform -1 0 5600 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1654395037
transform 1 0 336 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1654395037
transform -1 0 5600 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1654395037
transform 1 0 336 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1654395037
transform -1 0 5600 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1654395037
transform 1 0 336 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1654395037
transform -1 0 5600 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1654395037
transform 1 0 336 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1654395037
transform -1 0 5600 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1654395037
transform 1 0 336 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1654395037
transform -1 0 5600 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1654395037
transform 1 0 336 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1654395037
transform -1 0 5600 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1654395037
transform 1 0 336 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1654395037
transform -1 0 5600 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1654395037
transform 1 0 336 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1654395037
transform -1 0 5600 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1654395037
transform 1 0 336 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1654395037
transform -1 0 5600 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1654395037
transform 1 0 336 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1654395037
transform -1 0 5600 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1654395037
transform 1 0 336 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1654395037
transform -1 0 5600 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1654395037
transform 1 0 336 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1654395037
transform -1 0 5600 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1654395037
transform 1 0 336 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1654395037
transform -1 0 5600 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1654395037
transform 1 0 336 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1654395037
transform -1 0 5600 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1654395037
transform 1 0 336 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1654395037
transform -1 0 5600 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1654395037
transform 1 0 336 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1654395037
transform -1 0 5600 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1654395037
transform 1 0 336 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1654395037
transform -1 0 5600 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1654395037
transform 1 0 336 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1654395037
transform -1 0 5600 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_84
timestamp 1654395037
transform 1 0 4928 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_85
timestamp 1654395037
transform 1 0 4928 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86
timestamp 1654395037
transform 1 0 4928 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1654395037
transform 1 0 4928 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1654395037
transform 1 0 4928 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1654395037
transform 1 0 4928 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1654395037
transform 1 0 4928 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1654395037
transform 1 0 4928 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1654395037
transform 1 0 4928 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1654395037
transform 1 0 4928 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1654395037
transform 1 0 4928 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1654395037
transform 1 0 4928 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1654395037
transform 1 0 4928 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1654395037
transform 1 0 4928 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1654395037
transform 1 0 4928 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1654395037
transform 1 0 4928 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1654395037
transform 1 0 4928 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1654395037
transform 1 0 4928 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1654395037
transform 1 0 4928 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1654395037
transform 1 0 4928 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1654395037
transform 1 0 4928 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1654395037
transform 1 0 4928 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _044_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 4256 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _045_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 3136 0 1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _046_
timestamp 1654395037
transform 1 0 1792 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _047_
timestamp 1654395037
transform 1 0 4032 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _048_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4704 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _049_
timestamp 1654395037
transform 1 0 2128 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _050_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4256 0 -1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _051_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 2016 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _052_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 3696 0 -1 18032
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _053_
timestamp 1654395037
transform -1 0 1568 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _054_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 4928 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _055_
timestamp 1654395037
transform -1 0 3920 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _056_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 2912 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _057_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4032 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _058_
timestamp 1654395037
transform -1 0 5376 0 -1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _059_
timestamp 1654395037
transform 1 0 2464 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _060_
timestamp 1654395037
transform 1 0 2688 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _061_
timestamp 1654395037
transform -1 0 4928 0 1 32144
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _062_
timestamp 1654395037
transform 1 0 4480 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _063_
timestamp 1654395037
transform -1 0 5376 0 -1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _064_
timestamp 1654395037
transform -1 0 4704 0 -1 25872
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _065_
timestamp 1654395037
transform -1 0 5264 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _066_
timestamp 1654395037
transform -1 0 4032 0 1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _067_
timestamp 1654395037
transform -1 0 4928 0 1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _068_
timestamp 1654395037
transform 1 0 4480 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _069_
timestamp 1654395037
transform -1 0 5376 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _070_
timestamp 1654395037
transform -1 0 4928 0 1 22736
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _071_
timestamp 1654395037
transform 1 0 3584 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _072_
timestamp 1654395037
transform -1 0 4816 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _073_
timestamp 1654395037
transform -1 0 2912 0 -1 22736
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _074_
timestamp 1654395037
transform 1 0 2352 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _075_
timestamp 1654395037
transform -1 0 3808 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _076_
timestamp 1654395037
transform -1 0 3808 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _077_
timestamp 1654395037
transform -1 0 3136 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _078_
timestamp 1654395037
transform -1 0 2912 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _079_
timestamp 1654395037
transform 1 0 2688 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _080_
timestamp 1654395037
transform -1 0 4256 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _081_
timestamp 1654395037
transform -1 0 2688 0 1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _082_
timestamp 1654395037
transform 1 0 3024 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _083_
timestamp 1654395037
transform 1 0 4256 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _084_
timestamp 1654395037
transform 1 0 3696 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _085_
timestamp 1654395037
transform -1 0 4480 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _086_
timestamp 1654395037
transform 1 0 3696 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _087_
timestamp 1654395037
transform -1 0 4928 0 1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _088_
timestamp 1654395037
transform -1 0 4816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _089_
timestamp 1654395037
transform -1 0 3696 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _090_
timestamp 1654395037
transform -1 0 3024 0 1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _091_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 560 0 1 27440
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _092_
timestamp 1654395037
transform 1 0 1008 0 -1 29008
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _093_
timestamp 1654395037
transform -1 0 4928 0 1 29008
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _094_
timestamp 1654395037
transform 1 0 1008 0 -1 21168
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _095_
timestamp 1654395037
transform -1 0 4928 0 1 21168
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _096_
timestamp 1654395037
transform -1 0 4928 0 1 14896
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _097_
timestamp 1654395037
transform -1 0 4928 0 1 11760
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _098_
timestamp 1654395037
transform 1 0 1008 0 -1 8624
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _099_
timestamp 1654395037
transform 1 0 560 0 -1 11760
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _100_
timestamp 1654395037
transform -1 0 4928 0 -1 10192
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _101_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 4368 0 -1 32144
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _102_
timestamp 1654395037
transform -1 0 4368 0 1 30576
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _103_
timestamp 1654395037
transform 1 0 560 0 -1 30576
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _104_
timestamp 1654395037
transform -1 0 4368 0 -1 27440
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _105_
timestamp 1654395037
transform 1 0 560 0 -1 24304
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _106_
timestamp 1654395037
transform -1 0 4368 0 1 22736
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _107_
timestamp 1654395037
transform 1 0 560 0 1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _108_
timestamp 1654395037
transform -1 0 4368 0 -1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _109_
timestamp 1654395037
transform 1 0 560 0 1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _110_
timestamp 1654395037
transform -1 0 4368 0 -1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1654395037
transform 1 0 4256 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1654395037
transform 1 0 1568 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1654395037
transform -1 0 5040 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1654395037
transform 1 0 2240 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1654395037
transform 1 0 4704 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  const_source_one pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 3248 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  const_source_zero pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4480 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  data_delay_1 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1904 0 -1 13328
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  data_delay_2
timestamp 1654395037
transform 1 0 3248 0 -1 14896
box -86 -86 1542 870
<< labels >>
flabel metal4 s 376 724 696 33772 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 2376 724 2696 33772 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 4376 724 4696 33772 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 276 924 5660 1244 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 276 7924 5660 8244 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 276 14924 5660 15244 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 276 21924 5660 22244 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 276 28924 5660 29244 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 1376 724 1696 33772 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 3376 724 3696 33772 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 5376 724 5696 33772 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 276 4424 5696 4744 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 276 11424 5696 11744 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 276 18424 5696 18744 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 276 25424 5696 25744 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 276 32424 5696 32744 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal2 s 5900 34944 6100 35000 0 FreeSans 448 0 0 0 gpio_defaults[0]
port 2 nsew signal input
flabel metal2 s 5900 33488 6100 33544 0 FreeSans 448 0 0 0 gpio_defaults[1]
port 3 nsew signal input
flabel metal2 s 5900 31926 6100 31982 0 FreeSans 448 0 0 0 gpio_defaults[2]
port 4 nsew signal input
flabel metal2 s 5900 30470 6100 30526 0 FreeSans 448 0 0 0 gpio_defaults[3]
port 5 nsew signal input
flabel metal2 s 5900 28906 6100 28962 0 FreeSans 448 0 0 0 gpio_defaults[4]
port 6 nsew signal input
flabel metal2 s 5900 27450 6100 27506 0 FreeSans 448 0 0 0 gpio_defaults[5]
port 7 nsew signal input
flabel metal2 s 5900 25886 6100 25942 0 FreeSans 448 0 0 0 gpio_defaults[6]
port 8 nsew signal input
flabel metal2 s 5900 24430 6100 24486 0 FreeSans 448 0 0 0 gpio_defaults[7]
port 9 nsew signal input
flabel metal2 s 5900 22866 6100 22922 0 FreeSans 448 0 0 0 gpio_defaults[8]
port 10 nsew signal input
flabel metal2 s 5900 21410 6100 21466 0 FreeSans 448 0 0 0 gpio_defaults[9]
port 11 nsew signal input
flabel metal3 s 5800 15764 6000 15820 0 FreeSans 448 0 0 0 mgmt_gpio_in
port 12 nsew signal tristate
flabel metal3 s 5800 17556 6000 17612 0 FreeSans 448 0 0 0 mgmt_gpio_oeb
port 13 nsew signal input
flabel metal3 s 5800 18452 6000 18508 0 FreeSans 448 0 0 0 mgmt_gpio_out
port 14 nsew signal input
flabel metal3 s 5800 16660 6000 16716 0 FreeSans 448 0 0 0 one
port 15 nsew signal tristate
flabel metal2 s -100 13502 100 13578 0 FreeSans 448 0 0 0 pad_gpio_drive_sel[0]
port 16 nsew signal tristate
flabel metal2 s -100 13360 100 13436 0 FreeSans 448 0 0 0 pad_gpio_drive_sel[1]
port 17 nsew signal tristate
flabel metal2 s -100 752 100 828 0 FreeSans 448 0 0 0 pad_gpio_in
port 18 nsew signal input
flabel metal2 s -100 12647 100 12723 0 FreeSans 448 0 0 0 pad_gpio_inen
port 19 nsew signal tristate
flabel metal2 s -100 1044 100 1120 0 FreeSans 448 0 0 0 pad_gpio_out
port 20 nsew signal tristate
flabel metal2 s -100 898 100 974 0 FreeSans 448 0 0 0 pad_gpio_outen
port 21 nsew signal tristate
flabel metal2 s -100 12858 100 12934 0 FreeSans 448 0 0 0 pad_gpio_pulldown_sel
port 22 nsew signal tristate
flabel metal2 s -100 13731 100 13807 0 FreeSans 448 0 0 0 pad_gpio_pullup_sel
port 23 nsew signal tristate
flabel metal2 s -100 14252 100 14328 0 FreeSans 448 0 0 0 pad_gpio_schmitt_sel
port 24 nsew signal tristate
flabel metal2 s -100 1190 100 1266 0 FreeSans 448 0 0 0 pad_gpio_slew_sel
port 25 nsew signal tristate
flabel metal2 s 2212 34600 2268 35200 0 FreeSans 448 90 0 0 resetn
port 26 nsew signal input
flabel metal2 s 2212 -200 2268 400 0 FreeSans 448 90 0 0 resetn_out
port 27 nsew signal tristate
flabel metal2 s 3108 34600 3164 35200 0 FreeSans 448 90 0 0 serial_clock
port 28 nsew signal input
flabel metal2 s 3108 -200 3164 400 0 FreeSans 448 90 0 0 serial_clock_out
port 29 nsew signal tristate
flabel metal2 s 3556 34600 3612 35200 0 FreeSans 448 90 0 0 serial_data_in
port 30 nsew signal input
flabel metal2 s 2660 -200 2716 400 0 FreeSans 448 90 0 0 serial_data_out
port 31 nsew signal tristate
flabel metal2 s 2660 34600 2716 35200 0 FreeSans 448 90 0 0 serial_load
port 32 nsew signal input
flabel metal2 s 3556 -200 3612 400 0 FreeSans 448 90 0 0 serial_load_out
port 33 nsew signal tristate
flabel metal3 s 5800 16212 6000 16268 0 FreeSans 448 0 0 0 user_gpio_in
port 34 nsew signal tristate
flabel metal3 s 5800 18004 6000 18060 0 FreeSans 448 0 0 0 user_gpio_oeb
port 35 nsew signal input
flabel metal3 s 5800 18900 6000 18956 0 FreeSans 448 0 0 0 user_gpio_out
port 36 nsew signal input
flabel metal3 s 5800 17108 6000 17164 0 FreeSans 448 0 0 0 zero
port 37 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 6000 35000
<< end >>
