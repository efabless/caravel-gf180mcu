* NGSPICE file created from caravel_clocking.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

.subckt caravel_clocking VDD VSS core_clk ext_clk ext_clk_sel ext_reset pll_clk pll_clk90
+ resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
X_501_ _501_/D _350_/S _242_/Z _501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_294_ _312_/B _431_/B _338_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_363_ _501_/Q _407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_432_ _432_/A1 _432_/A2 _432_/B _433_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_415_ _489_/Q _415_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_346_ _340_/B _468_/Q _346_/A3 _346_/B _468_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_277_ _456_/Q _313_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_329_ _324_/B _465_/Q _336_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__365__A2 _360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__492__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__445__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_500_ _500_/D _350_/S _242_/Z _500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_362_ _361_/Z _478_/Q _362_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_431_ _432_/A1 _432_/A2 _431_/B _432_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__445__CLKN _233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_293_ _301_/A1 _291_/Z _331_/C _459_/Q _298_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_414_ _414_/I _488_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_276_ _458_/Q _459_/Q _299_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_345_ _340_/B _467_/Q _468_/Q _346_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ _271_/I _226_/I _260_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_328_ _430_/A1 _335_/B _323_/Z _331_/C _330_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_output12_I _233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__312__B _312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__491__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I pll_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_292_ _311_/B _331_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_430_ _430_/A1 _335_/B _466_/Q _226_/Z _432_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_361_ _500_/Q _361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__265__A2 _312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__496__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_413_ _422_/C _413_/A2 _413_/B _414_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__238__A2 _500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_275_ _311_/B _301_/A1 _289_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_344_ _344_/A1 _312_/B _344_/B _346_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__410__A2 _358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__469__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__459__CLKN input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__448__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_327_ _464_/Q _430_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_258_ _456_/Q _271_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_360_ _360_/I _360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_291_ _270_/I _458_/Q _291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_489_ _489_/D _350_/S input4/Z _489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__481__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_412_ _370_/Z _486_/Q _360_/Z _488_/Q _413_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_343_ _469_/Q _344_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_274_ _280_/I _220_/Z _279_/C _301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__490__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__238__A3 input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__458__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_257_ _257_/I _455_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_326_ _283_/C _326_/A2 _326_/A3 _464_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_309_ _462_/Q _461_/Q _318_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__458__CLKN input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput12 _233_/Z core_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__295__I _312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__440__A1 _435_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_488_ _488_/D _350_/S input4/Z _488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_290_ _290_/I _458_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_411_ _358_/I _411_/A2 _411_/A3 _411_/B _487_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__239__B _499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_273_ _462_/Q _463_/Q _279_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_342_ _342_/I _467_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__471__CLK _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_325_ _337_/C _325_/A2 _326_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_256_ _455_/Q _256_/A2 _257_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__494__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_239_ _501_/Q _500_/Q _499_/Q _360_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_308_ _260_/I _316_/A2 _308_/A3 _308_/B _461_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_1_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput13 _247_/Z resetb_sync VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__457__CLKN input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__499__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__422__A2 _360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_487_ _487_/D _350_/S input4/Z _487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XANTENNA_input1_I ext_clk_sel VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_410_ _370_/Z _358_/Z _411_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_272_ _473_/Q _280_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_341_ _340_/B _344_/B _341_/B _342_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__340__A1 _285_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__398__A1 _500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_324_ _335_/B _323_/Z _324_/B _325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_255_ _224_/B _467_/Q _340_/A2 _256_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_238_ _501_/Q _500_/Q input4/Z _241_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_307_ _260_/I _316_/A2 _461_/Q _308_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput14 _244_/Z user_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_486_ _486_/D _350_/S input4/Z _486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XANTENNA__435__C _435_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_340_ _285_/I _340_/A2 _340_/B _344_/B _341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_271_ _271_/I _311_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__398__A2 _499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_469_ _469_/D _350_/S input3/Z _469_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_254_ _469_/Q _468_/Q _340_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_323_ _466_/Q _323_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_237_ _426_/A1 _384_/A1 _480_/Q _241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_306_ _311_/B _304_/Z _306_/B _308_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__451__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__407__A1 _361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_485_ _485_/D _350_/S input4/Z _485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XANTENNA__474__CLK _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__455__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_270_ _270_/I _283_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_399_ _382_/B _399_/A2 _400_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_468_ _468_/D _350_/S input3/Z _468_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_3_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_322_ _465_/Q _335_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_253_ _253_/I _450_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_236_ _500_/Q _384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_305_ _461_/Q _311_/B _306_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__425__A2 _358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__416__A2 _358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__407__A2 _499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_484_ _484_/D _350_/S input4/Z _484_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_398_ _500_/Q _499_/Q _399_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__500__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_467_ _467_/D _350_/S input3/Z _467_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_4_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__464__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_252_ _450_/Q _249_/Z _252_/B _253_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_321_ _324_/B _260_/Z _326_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_235_ _501_/Q _426_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_304_ _224_/B _474_/Q _304_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_483_ _483_/D _350_/S input4/Z _483_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
X_397_ _422_/C _395_/Z _397_/A3 _485_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_466_ _466_/D _350_/S input3/Z _466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_251_ _450_/Q _249_/Z _251_/B _252_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_320_ _464_/Q _324_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_449_ _449_/D _350_/S input3/Z _449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_234_ _499_/Q _378_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_303_ _462_/Q _463_/Q _313_/C _316_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__454__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__477__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_482_ _482_/D _350_/S input4/Z _482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_396_ _371_/Z _396_/A2 _485_/Q _397_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_465_ _465_/D _350_/S input3/Z _465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_2_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_250_ _481_/Q _251_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_448_ _448_/D _350_/S input3/Z _449_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_379_ _435_/C _251_/B _380_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__236__I _500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ _233_/I _233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__456__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_302_ _331_/C _300_/Z _302_/A3 _460_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__364__A1 _407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__346__A1 _340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__467__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_481_ _481_/D _350_/S input4/Z _481_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__467__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_464_ _464_/D _350_/S input3/Z _464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_395_ _485_/Q _371_/Z _396_/A2 _395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_447_ _447_/D _350_/S _233_/Z _447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
X_378_ _378_/I _435_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_232_ _231_/Z _230_/Z _449_/Q _233_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_301_ _301_/A1 _301_/A2 _460_/Q _302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input8_I sel2[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__282__A1 _340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_480_ _480_/D _350_/S input4/Z _480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__501__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_394_ _369_/I _394_/A2 _396_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_463_ _463_/D _350_/S input3/Z _463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_446_ _447_/Q _350_/S _233_/Z _446_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XFILLER_13_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_377_ _380_/A1 _394_/A2 _377_/B _428_/C _380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_231_ ext_clk _451_/Q _449_/D _231_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_300_ _460_/Q _301_/A1 _301_/A2 _300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_429_ _429_/A1 _429_/A2 _429_/A3 _491_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput1 ext_clk_sel _245_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__490__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__361__I _500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__495__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__486__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_393_ _393_/A1 _429_/A1 _393_/A3 _484_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_462_ _462_/D _350_/S input3/Z _462_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XANTENNA__468__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__459__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_445_ _446_/Q _350_/S _233_/Z _445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
X_376_ _382_/B _360_/Z _428_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_230_ _230_/I _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_359_ _477_/Q _365_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_428_ _491_/Q _428_/A2 _428_/B _428_/C _429_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__450__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__465__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 ext_reset input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__480__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_392_ _428_/C _377_/B _394_/A2 _392_/A4 _393_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_461_ _461_/D _350_/S input3/Z _461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_375_ _481_/Q _382_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_444_ _444_/I _495_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_358_ _358_/I _358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_427_ _491_/Q _427_/A2 _428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__376__A2 _360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 pll_clk input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_289_ _458_/Q _289_/I1 _289_/S _290_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__294__A1 _312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__421__A1 _361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__285__I _285_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I sel2[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_391_ _426_/A1 _369_/I _392_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_460_ _460_/D _350_/S input3/Z _460_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
X_374_ _488_/Q _370_/Z _377_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_443_ _495_/Q _443_/A2 _444_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__470__CLK _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__493__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_426_ _426_/A1 _415_/Z _490_/Q _428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput4 pll_clk90 input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_357_ _419_/B _360_/I _358_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__378__I _378_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_288_ _288_/A1 _288_/A2 _287_/Z _313_/C _289_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_409_ _419_/B _409_/A2 _406_/Z _413_/B _411_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_2_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__340__B _340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__498__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__489__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_390_ _407_/B _251_/B _429_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__330__A1 _285_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__463__CLKN input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_442_ _378_/I _494_/Q _493_/Q _443_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_373_ _483_/Q _484_/Q _394_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__379__A1 _435_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 resetb _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_425_ _491_/Q _358_/Z _429_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_356_ _481_/Q _419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_287_ _457_/Q _458_/Q _287_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_408_ _382_/B _408_/A2 _413_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_339_ _467_/Q _344_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__412__A3 _360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_372_ _419_/B _371_/Z _385_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_441_ _435_/C _494_/Q _441_/A3 _441_/B _494_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__462__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__312__A2 _285_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_424_ _424_/I _490_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_355_ _355_/I _480_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_286_ _270_/I _299_/A2 _313_/C _288_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput6 sel2[0] _496_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__221__A1 input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__462__CLKN input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_407_ _361_/Z _499_/Q _407_/B _408_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__442__A1 _378_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_269_ _457_/Q _270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_338_ _338_/A1 _338_/A2 _338_/A3 _466_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__450__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__406__A1 _407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__473__CLK _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I pll_clk90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_440_ _435_/C _493_/Q _494_/Q _441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_371_ _488_/Q _370_/Z _360_/I _371_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_1_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_423_ _358_/Z _423_/A2 _423_/B _424_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_354_ _480_/Q _354_/A2 _355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__470__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_285_ _285_/I _288_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 sel2[1] _497_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__461__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_406_ _407_/B _361_/Z _378_/I _406_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_268_ _268_/I _456_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_337_ _323_/Z _337_/A2 _337_/B _337_/C _338_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__461__CLKN input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 sel[1] _471_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__406__A2 _361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_370_ _487_/Q _370_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_499_ _499_/D _350_/S _242_/Z _499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_422_ _415_/Z _360_/Z _490_/Q _422_/C _423_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_284_ _284_/I _457_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_353_ _378_/I _495_/Q _494_/Q _439_/B _354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput8 sel2[2] _498_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_405_ _487_/Q _486_/Q _409_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_336_ _323_/Z _336_/A2 _337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_267_ _260_/Z _267_/A2 _268_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput11 sel[2] _472_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_319_ _319_/I _463_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__460__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__406__A3 _378_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__460__CLKN input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_498_ _498_/D _350_/S _242_/Z _501_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_421_ _361_/Z _421_/A2 _427_/A2 _422_/C _423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_352_ _493_/Q _439_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 sel[0] _470_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_283_ _283_/A1 _289_/S _283_/B _283_/C _284_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__453__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_404_ _404_/I _486_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__436__A1 _435_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_335_ _335_/A1 _324_/B _335_/B _337_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_266_ _266_/A1 _226_/Z _263_/Z _265_/Z _267_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__476__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_249_ _419_/A1 _490_/Q _491_/Q _360_/I _249_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_318_ _337_/C _318_/A2 _313_/B _431_/B _318_/C _319_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__491__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__474__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input10_I sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__482__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_497_ _497_/D _350_/S _242_/Z _500_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__473__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I ext_reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__464__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_351_ _351_/I _476_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_420_ _415_/Z _490_/Q _427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_282_ _340_/B _431_/B _283_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__390__A1 _407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_403_ _486_/Q _403_/I1 _403_/S _404_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_334_ _323_/Z _260_/Z _338_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_265_ _454_/Q _312_/B _265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_248_ _489_/Q _419_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__350__S _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__345__A1 _340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_317_ _463_/Q _431_/B _318_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__234__I _499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__350__I1 ext_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__466__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__489__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_496_ _496_/D _350_/S _242_/Z _499_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_350_ _476_/Q ext_clk _350_/S _351_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_281_ _456_/Q _431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_479_ _501_/Q input4/Z _479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_402_ _358_/I _411_/A2 _403_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_264_ _475_/Q _312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_333_ _333_/I _465_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__488__CLKN input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_316_ _260_/I _316_/A2 _314_/Z _316_/B _462_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_247_ _247_/I _247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__477__D _499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__456__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_495_ _495_/D _350_/S input4/Z _495_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__479__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__232__I1 _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_280_ _280_/I _340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_478_ _500_/Q input4/Z _478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__439__A1 _407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_401_ _488_/Q _370_/Z _382_/B _411_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_263_ _453_/Q _285_/I _263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_332_ _260_/Z _332_/A2 _332_/B _333_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__487__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_246_ input2/Z _445_/Q _247_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_315_ _462_/Q _260_/Z _316_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__487__CLKN input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__263__A2 _285_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_229_ _229_/A1 _229_/A2 _226_/Z _228_/Z _230_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__494__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__449__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_494_ _494_/D _350_/S input4/Z _494_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_5_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_477_ _499_/Q input4/Z _477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__366__A1 _358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_400_ _486_/Q _251_/B _400_/B _403_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__469__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_331_ _324_/B _226_/Z _335_/B _331_/C _332_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_262_ _474_/Q _285_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_245_ _245_/I _448_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_314_ _314_/A1 _314_/A2 _314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__471__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_228_ _460_/Q _432_/A1 _228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__486__CLKN input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_493_ _493_/D _350_/S input4/Z _493_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_476_ _476_/D input3/Z _476_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_330_ _285_/I _330_/A2 _336_/A2 _331_/C _332_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_261_ _452_/Q _266_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_459_ _459_/D _350_/S input3/Z _459_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_244_ _244_/I _244_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_313_ _280_/I _220_/Z _313_/B _313_/C _314_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_227_ _492_/Q _432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_492_ _492_/D _350_/S input3/Z _492_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__485__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__407__B _407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_475_ _475_/D _350_/S _230_/Z _475_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__492__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__485__CLKN input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_260_ _260_/I _260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_389_ _371_/Z _387_/Z _422_/C _484_/Q _393_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_458_ _458_/D _350_/S input3/Z _458_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
X_243_ _231_/Z _242_/Z _449_/Q _244_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_312_ _280_/I _285_/I _312_/B _313_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__488__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__239__A2 _500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_226_ _226_/I _226_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__449__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_491_ _491_/D _350_/S input4/Z _491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_474_ _474_/D _350_/S _230_/Z _474_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_388_ _419_/B _422_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_457_ _457_/D _350_/S input3/Z _457_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_242_ _242_/I _242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_311_ _318_/A2 _310_/Z _311_/B _314_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__484__CLKN input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_225_ _474_/Q _475_/Q _473_/Q _226_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input9_I sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_490_ _490_/D _350_/S input4/Z _490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_473_ _473_/D _350_/S _230_/Z _473_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_456_ _456_/D _350_/S input3/Z _456_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__441__A1 _435_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_387_ _483_/Q _369_/I _387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_310_ _462_/Q _461_/Q _310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_241_ _378_/I _241_/A2 _241_/A3 _360_/I _241_/B2 _242_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__423__A1 _358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_439_ _407_/B _439_/A2 _439_/B _441_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__483__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_224_ _455_/Q _224_/A2 _224_/B _229_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__472__CLK _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__483__CLKN input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__495__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_472_ _472_/D _350_/S _230_/Z _475_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__451__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_386_ _386_/I _483_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_455_ _455_/D _350_/S input3/Z _455_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_240_ _485_/Q _450_/Q _241_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_438_ _495_/Q _439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_369_ _369_/I _380_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_223_ _473_/Q _224_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__341__A1 _340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__497__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_447__15 _447_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__482__CLKN input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_471_ _471_/D _350_/S _230_/Z _474_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_454_ _475_/Q input3/Z _454_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_385_ _483_/Q _385_/I1 _385_/S _386_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_437_ _437_/I _493_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_299_ _270_/I _299_/A2 _301_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_368_ _482_/Q _369_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_222_ _474_/Q _475_/Q _224_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__241__A1 _378_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input7_I sel2[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_470_ _470_/D _350_/S _230_/Z _473_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_384_ _384_/A1 _384_/A2 _383_/Z _251_/B _385_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__435__A1 _361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__452__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_453_ _474_/Q input3/Z _453_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__475__CLK _230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_367_ _367_/I _481_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_436_ _435_/C _439_/B _436_/B _437_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_298_ _298_/A1 _338_/A1 _298_/A3 _459_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_221_ input3/Z _220_/Z _229_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_419_ _419_/A1 _490_/Q _491_/Q _419_/B _421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_3_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__481__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__472__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__463__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_452_ _473_/Q input3/Z _452_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_383_ _483_/Q _482_/Q _383_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__480__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__353__A1 _378_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__362__A1 _361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__417__A2 _360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_366_ _358_/Z _366_/A2 _367_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_435_ _361_/Z _435_/A2 _439_/B _435_/C _436_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_297_ _279_/C _299_/A2 _337_/C _297_/A4 _298_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_3_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_220_ _474_/Q _475_/Q _220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_418_ _249_/Z _380_/C _418_/A3 _417_/Z _489_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_349_ _349_/I _469_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__465__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__231__I0 ext_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_451_ _476_/Q _350_/S input3/Z _451_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_382_ _369_/I _394_/A2 _382_/B _384_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_434_ _495_/Q _494_/Q _435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_365_ _365_/A1 _360_/Z _362_/Z _364_/Z _366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_296_ _335_/A1 _270_/I _297_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__344__A2 _312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_417_ _415_/Z _360_/Z _417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__447__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ _469_/Q _348_/A2 _349_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_279_ _283_/A1 _299_/A2 _337_/C _279_/C _283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__455__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__447__CLKN _233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__478__CLK input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I resetb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_450_ _450_/D _350_/S input4/Z _450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_381_ _381_/I _482_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_433_ _433_/I _492_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_364_ _407_/B _479_/Q _364_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_295_ _312_/B _335_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_416_ _415_/Z _358_/Z _418_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_347_ _280_/I _468_/Q _467_/Q _348_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_278_ _313_/C _226_/Z _337_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__484__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__475__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__446__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__493__SETN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__466__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__457__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__448__RN _350_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__478__D _500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__446__CLKN _233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_380_ _380_/A1 _385_/S _380_/B _380_/C _381_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__468__CLK input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

