magic
tech gf180mcuC
magscale 1 10
timestamp 1655473345
<< checkpaint >>
rect -1976 -1926 27112 10716
<< obsm1 >>
rect 90 99 25112 8716
<< metal2 >>
rect 24889 6817 25108 7017
rect 24890 6342 25109 6542
<< obsm2 >>
rect 343 7077 24890 8714
rect 343 6757 24829 7077
rect 343 6602 24890 6757
rect 343 6282 24830 6602
rect 343 5473 24890 6282
<< obsm3 >>
rect 3923 5808 17907 8714
<< obsm4 >>
rect 3923 427 17907 8714
<< metal5 >>
rect 24 7914 3963 8714
rect 24 5884 4003 6684
<< obsm5 >>
rect 4063 7814 17907 8714
rect 3963 6784 17907 7814
rect 4103 5784 17907 6784
rect 3963 74 17907 5784
<< labels >>
rlabel metal5 s 24 7914 3963 8714 6 VDD
port 1 nsew
rlabel metal5 s 24 5884 4003 6684 6 VSS
port 2 nsew
rlabel metal2 s 24890 6342 25109 6542 6 porb
port 3 nsew
rlabel metal2 s 24889 6817 25108 7017 6 por
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 25156 8716
string GDS_END 304670
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 218002
string LEFclass BLOCK
string LEFview TRUE
<< end >>
