VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO housekeeping
  CLASS BLOCK ;
  FOREIGN housekeeping ;
  ORIGIN 0.000 0.000 ;
  SIZE 520.000 BY 780.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -0.880 8.080 0.720 768.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 8.080 520.560 9.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 766.480 520.560 768.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 518.960 8.080 520.560 768.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.240 4.780 23.840 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.040 4.780 100.640 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 4.780 177.440 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 4.780 254.240 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 4.780 331.040 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 4.780 407.840 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 4.780 484.640 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 21.290 523.860 22.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 81.290 523.860 82.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 141.290 523.860 142.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 201.290 523.860 202.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 261.290 523.860 262.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 321.290 523.860 322.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 381.290 523.860 382.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 441.290 523.860 442.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 501.290 523.860 502.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 561.290 523.860 562.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 621.290 523.860 622.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 681.290 523.860 682.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 741.290 523.860 742.890 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -4.180 4.780 -2.580 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 4.780 523.860 6.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 769.780 523.860 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 522.260 4.780 523.860 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 25.540 4.780 27.140 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.340 4.780 103.940 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 4.780 180.740 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.940 4.780 257.540 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 4.780 334.340 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.540 4.780 411.140 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 4.780 487.940 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 51.290 523.860 52.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 111.290 523.860 112.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 171.290 523.860 172.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 231.290 523.860 232.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 291.290 523.860 292.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 351.290 523.860 352.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 411.290 523.860 412.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 471.290 523.860 472.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 531.290 523.860 532.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 591.290 523.860 592.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 651.290 523.860 652.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 711.290 523.860 712.890 ;
    END
  END VSS
  PIN debug_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.960 4.000 23.520 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.280 4.000 35.840 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 4.000 42.000 ;
    END
  END debug_out
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.920 4.000 60.480 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END irq[2]
  PIN mask_rev_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END mask_rev_in[0]
  PIN mask_rev_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.280 0.000 385.840 4.000 ;
    END
  END mask_rev_in[10]
  PIN mask_rev_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END mask_rev_in[11]
  PIN mask_rev_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 0.000 397.040 4.000 ;
    END
  END mask_rev_in[12]
  PIN mask_rev_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END mask_rev_in[13]
  PIN mask_rev_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 0.000 408.240 4.000 ;
    END
  END mask_rev_in[14]
  PIN mask_rev_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END mask_rev_in[15]
  PIN mask_rev_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END mask_rev_in[16]
  PIN mask_rev_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END mask_rev_in[17]
  PIN mask_rev_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 0.000 430.640 4.000 ;
    END
  END mask_rev_in[18]
  PIN mask_rev_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 0.000 436.240 4.000 ;
    END
  END mask_rev_in[19]
  PIN mask_rev_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 0.000 335.440 4.000 ;
    END
  END mask_rev_in[1]
  PIN mask_rev_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 0.000 441.840 4.000 ;
    END
  END mask_rev_in[20]
  PIN mask_rev_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 0.000 447.440 4.000 ;
    END
  END mask_rev_in[21]
  PIN mask_rev_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 452.480 0.000 453.040 4.000 ;
    END
  END mask_rev_in[22]
  PIN mask_rev_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END mask_rev_in[23]
  PIN mask_rev_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 0.000 464.240 4.000 ;
    END
  END mask_rev_in[24]
  PIN mask_rev_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END mask_rev_in[25]
  PIN mask_rev_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.880 0.000 475.440 4.000 ;
    END
  END mask_rev_in[26]
  PIN mask_rev_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 0.000 481.040 4.000 ;
    END
  END mask_rev_in[27]
  PIN mask_rev_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 0.000 486.640 4.000 ;
    END
  END mask_rev_in[28]
  PIN mask_rev_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 0.000 492.240 4.000 ;
    END
  END mask_rev_in[29]
  PIN mask_rev_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END mask_rev_in[2]
  PIN mask_rev_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 0.000 497.840 4.000 ;
    END
  END mask_rev_in[30]
  PIN mask_rev_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 0.000 503.440 4.000 ;
    END
  END mask_rev_in[31]
  PIN mask_rev_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END mask_rev_in[3]
  PIN mask_rev_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 4.000 ;
    END
  END mask_rev_in[4]
  PIN mask_rev_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END mask_rev_in[5]
  PIN mask_rev_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 0.000 363.440 4.000 ;
    END
  END mask_rev_in[6]
  PIN mask_rev_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END mask_rev_in[7]
  PIN mask_rev_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 0.000 374.640 4.000 ;
    END
  END mask_rev_in[8]
  PIN mask_rev_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END mask_rev_in[9]
  PIN mgmt_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 72.240 520.000 72.800 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 425.040 520.000 425.600 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 460.320 520.000 460.880 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 495.600 520.000 496.160 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 530.880 520.000 531.440 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 566.160 520.000 566.720 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 601.440 520.000 602.000 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 636.720 520.000 637.280 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 672.000 520.000 672.560 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 707.280 520.000 707.840 ;
    END
  END mgmt_gpio_in[18]
  PIN mgmt_gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 742.560 520.000 743.120 ;
    END
  END mgmt_gpio_in[19]
  PIN mgmt_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 107.520 520.000 108.080 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 429.520 4.000 430.080 ;
    END
  END mgmt_gpio_in[20]
  PIN mgmt_gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END mgmt_gpio_in[21]
  PIN mgmt_gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 466.480 4.000 467.040 ;
    END
  END mgmt_gpio_in[22]
  PIN mgmt_gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 484.960 4.000 485.520 ;
    END
  END mgmt_gpio_in[23]
  PIN mgmt_gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 503.440 4.000 504.000 ;
    END
  END mgmt_gpio_in[24]
  PIN mgmt_gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END mgmt_gpio_in[25]
  PIN mgmt_gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.400 4.000 540.960 ;
    END
  END mgmt_gpio_in[26]
  PIN mgmt_gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 558.880 4.000 559.440 ;
    END
  END mgmt_gpio_in[27]
  PIN mgmt_gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.360 4.000 577.920 ;
    END
  END mgmt_gpio_in[28]
  PIN mgmt_gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 595.840 4.000 596.400 ;
    END
  END mgmt_gpio_in[29]
  PIN mgmt_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 142.800 520.000 143.360 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.320 4.000 614.880 ;
    END
  END mgmt_gpio_in[30]
  PIN mgmt_gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.800 4.000 633.360 ;
    END
  END mgmt_gpio_in[31]
  PIN mgmt_gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.280 4.000 651.840 ;
    END
  END mgmt_gpio_in[32]
  PIN mgmt_gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 669.760 4.000 670.320 ;
    END
  END mgmt_gpio_in[33]
  PIN mgmt_gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.240 4.000 688.800 ;
    END
  END mgmt_gpio_in[34]
  PIN mgmt_gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 706.720 4.000 707.280 ;
    END
  END mgmt_gpio_in[35]
  PIN mgmt_gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.200 4.000 725.760 ;
    END
  END mgmt_gpio_in[36]
  PIN mgmt_gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 743.680 4.000 744.240 ;
    END
  END mgmt_gpio_in[37]
  PIN mgmt_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 178.080 520.000 178.640 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 213.360 520.000 213.920 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 248.640 520.000 249.200 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 283.920 520.000 284.480 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 319.200 520.000 319.760 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 354.480 520.000 355.040 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 389.760 520.000 390.320 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 84.000 520.000 84.560 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 436.800 520.000 437.360 ;
    END
  END mgmt_gpio_oeb[10]
  PIN mgmt_gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 472.080 520.000 472.640 ;
    END
  END mgmt_gpio_oeb[11]
  PIN mgmt_gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 507.360 520.000 507.920 ;
    END
  END mgmt_gpio_oeb[12]
  PIN mgmt_gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 542.640 520.000 543.200 ;
    END
  END mgmt_gpio_oeb[13]
  PIN mgmt_gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 577.920 520.000 578.480 ;
    END
  END mgmt_gpio_oeb[14]
  PIN mgmt_gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 613.200 520.000 613.760 ;
    END
  END mgmt_gpio_oeb[15]
  PIN mgmt_gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 648.480 520.000 649.040 ;
    END
  END mgmt_gpio_oeb[16]
  PIN mgmt_gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 683.760 520.000 684.320 ;
    END
  END mgmt_gpio_oeb[17]
  PIN mgmt_gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 719.040 520.000 719.600 ;
    END
  END mgmt_gpio_oeb[18]
  PIN mgmt_gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 754.320 520.000 754.880 ;
    END
  END mgmt_gpio_oeb[19]
  PIN mgmt_gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 119.280 520.000 119.840 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.680 4.000 436.240 ;
    END
  END mgmt_gpio_oeb[20]
  PIN mgmt_gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.160 4.000 454.720 ;
    END
  END mgmt_gpio_oeb[21]
  PIN mgmt_gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 472.640 4.000 473.200 ;
    END
  END mgmt_gpio_oeb[22]
  PIN mgmt_gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.120 4.000 491.680 ;
    END
  END mgmt_gpio_oeb[23]
  PIN mgmt_gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END mgmt_gpio_oeb[24]
  PIN mgmt_gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 528.080 4.000 528.640 ;
    END
  END mgmt_gpio_oeb[25]
  PIN mgmt_gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 546.560 4.000 547.120 ;
    END
  END mgmt_gpio_oeb[26]
  PIN mgmt_gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 565.040 4.000 565.600 ;
    END
  END mgmt_gpio_oeb[27]
  PIN mgmt_gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 583.520 4.000 584.080 ;
    END
  END mgmt_gpio_oeb[28]
  PIN mgmt_gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.000 4.000 602.560 ;
    END
  END mgmt_gpio_oeb[29]
  PIN mgmt_gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 154.560 520.000 155.120 ;
    END
  END mgmt_gpio_oeb[2]
  PIN mgmt_gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 620.480 4.000 621.040 ;
    END
  END mgmt_gpio_oeb[30]
  PIN mgmt_gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.960 4.000 639.520 ;
    END
  END mgmt_gpio_oeb[31]
  PIN mgmt_gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 657.440 4.000 658.000 ;
    END
  END mgmt_gpio_oeb[32]
  PIN mgmt_gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.920 4.000 676.480 ;
    END
  END mgmt_gpio_oeb[33]
  PIN mgmt_gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.400 4.000 694.960 ;
    END
  END mgmt_gpio_oeb[34]
  PIN mgmt_gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 712.880 4.000 713.440 ;
    END
  END mgmt_gpio_oeb[35]
  PIN mgmt_gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 731.360 4.000 731.920 ;
    END
  END mgmt_gpio_oeb[36]
  PIN mgmt_gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 749.840 4.000 750.400 ;
    END
  END mgmt_gpio_oeb[37]
  PIN mgmt_gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 189.840 520.000 190.400 ;
    END
  END mgmt_gpio_oeb[3]
  PIN mgmt_gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 225.120 520.000 225.680 ;
    END
  END mgmt_gpio_oeb[4]
  PIN mgmt_gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 260.400 520.000 260.960 ;
    END
  END mgmt_gpio_oeb[5]
  PIN mgmt_gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 295.680 520.000 296.240 ;
    END
  END mgmt_gpio_oeb[6]
  PIN mgmt_gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 330.960 520.000 331.520 ;
    END
  END mgmt_gpio_oeb[7]
  PIN mgmt_gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 366.240 520.000 366.800 ;
    END
  END mgmt_gpio_oeb[8]
  PIN mgmt_gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 401.520 520.000 402.080 ;
    END
  END mgmt_gpio_oeb[9]
  PIN mgmt_gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 95.760 520.000 96.320 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 448.560 520.000 449.120 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 483.840 520.000 484.400 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 519.120 520.000 519.680 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 554.400 520.000 554.960 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 589.680 520.000 590.240 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 624.960 520.000 625.520 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 660.240 520.000 660.800 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 695.520 520.000 696.080 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 730.800 520.000 731.360 ;
    END
  END mgmt_gpio_out[18]
  PIN mgmt_gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 766.080 520.000 766.640 ;
    END
  END mgmt_gpio_out[19]
  PIN mgmt_gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 131.040 520.000 131.600 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 441.840 4.000 442.400 ;
    END
  END mgmt_gpio_out[20]
  PIN mgmt_gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 4.000 460.880 ;
    END
  END mgmt_gpio_out[21]
  PIN mgmt_gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 478.800 4.000 479.360 ;
    END
  END mgmt_gpio_out[22]
  PIN mgmt_gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 497.280 4.000 497.840 ;
    END
  END mgmt_gpio_out[23]
  PIN mgmt_gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.760 4.000 516.320 ;
    END
  END mgmt_gpio_out[24]
  PIN mgmt_gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END mgmt_gpio_out[25]
  PIN mgmt_gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.720 4.000 553.280 ;
    END
  END mgmt_gpio_out[26]
  PIN mgmt_gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END mgmt_gpio_out[27]
  PIN mgmt_gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.680 4.000 590.240 ;
    END
  END mgmt_gpio_out[28]
  PIN mgmt_gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 4.000 608.720 ;
    END
  END mgmt_gpio_out[29]
  PIN mgmt_gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 166.320 520.000 166.880 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 626.640 4.000 627.200 ;
    END
  END mgmt_gpio_out[30]
  PIN mgmt_gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END mgmt_gpio_out[31]
  PIN mgmt_gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 663.600 4.000 664.160 ;
    END
  END mgmt_gpio_out[32]
  PIN mgmt_gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END mgmt_gpio_out[33]
  PIN mgmt_gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 700.560 4.000 701.120 ;
    END
  END mgmt_gpio_out[34]
  PIN mgmt_gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 719.040 4.000 719.600 ;
    END
  END mgmt_gpio_out[35]
  PIN mgmt_gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 737.520 4.000 738.080 ;
    END
  END mgmt_gpio_out[36]
  PIN mgmt_gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.000 4.000 756.560 ;
    END
  END mgmt_gpio_out[37]
  PIN mgmt_gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 201.600 520.000 202.160 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 236.880 520.000 237.440 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 272.160 520.000 272.720 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 307.440 520.000 308.000 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 342.720 520.000 343.280 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 378.000 520.000 378.560 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 413.280 520.000 413.840 ;
    END
  END mgmt_gpio_out[9]
  PIN pad_flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 0.000 16.240 4.000 ;
    END
  END pad_flash_clk
  PIN pad_flash_clk_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 0.000 21.840 4.000 ;
    END
  END pad_flash_clk_oe
  PIN pad_flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END pad_flash_csb
  PIN pad_flash_csb_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 4.000 ;
    END
  END pad_flash_csb_oe
  PIN pad_flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END pad_flash_io0_di
  PIN pad_flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END pad_flash_io0_do
  PIN pad_flash_io0_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END pad_flash_io0_ie
  PIN pad_flash_io0_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 4.000 ;
    END
  END pad_flash_io0_oe
  PIN pad_flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END pad_flash_io1_di
  PIN pad_flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END pad_flash_io1_do
  PIN pad_flash_io1_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 4.000 ;
    END
  END pad_flash_io1_ie
  PIN pad_flash_io1_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END pad_flash_io1_oe
  PIN pll90_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 4.000 ;
    END
  END pll90_sel[0]
  PIN pll90_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END pll90_sel[1]
  PIN pll90_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END pll90_sel[2]
  PIN pll_bypass
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END pll_bypass
  PIN pll_dco_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 4.000 ;
    END
  END pll_dco_ena
  PIN pll_div[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END pll_div[0]
  PIN pll_div[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END pll_div[1]
  PIN pll_div[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END pll_div[2]
  PIN pll_div[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 4.000 ;
    END
  END pll_div[3]
  PIN pll_div[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END pll_div[4]
  PIN pll_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END pll_ena
  PIN pll_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 4.000 ;
    END
  END pll_sel[0]
  PIN pll_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END pll_sel[1]
  PIN pll_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END pll_sel[2]
  PIN pll_trim[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END pll_trim[0]
  PIN pll_trim[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END pll_trim[10]
  PIN pll_trim[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 0.000 229.040 4.000 ;
    END
  END pll_trim[11]
  PIN pll_trim[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END pll_trim[12]
  PIN pll_trim[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END pll_trim[13]
  PIN pll_trim[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END pll_trim[14]
  PIN pll_trim[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 0.000 251.440 4.000 ;
    END
  END pll_trim[15]
  PIN pll_trim[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END pll_trim[16]
  PIN pll_trim[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END pll_trim[17]
  PIN pll_trim[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END pll_trim[18]
  PIN pll_trim[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 0.000 273.840 4.000 ;
    END
  END pll_trim[19]
  PIN pll_trim[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 4.000 ;
    END
  END pll_trim[1]
  PIN pll_trim[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END pll_trim[20]
  PIN pll_trim[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END pll_trim[21]
  PIN pll_trim[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END pll_trim[22]
  PIN pll_trim[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 0.000 296.240 4.000 ;
    END
  END pll_trim[23]
  PIN pll_trim[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 0.000 301.840 4.000 ;
    END
  END pll_trim[24]
  PIN pll_trim[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END pll_trim[25]
  PIN pll_trim[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END pll_trim[2]
  PIN pll_trim[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 0.000 184.240 4.000 ;
    END
  END pll_trim[3]
  PIN pll_trim[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 4.000 ;
    END
  END pll_trim[4]
  PIN pll_trim[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END pll_trim[5]
  PIN pll_trim[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 4.000 ;
    END
  END pll_trim[6]
  PIN pll_trim[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 0.000 206.640 4.000 ;
    END
  END pll_trim[7]
  PIN pll_trim[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END pll_trim[8]
  PIN pll_trim[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END pll_trim[9]
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END porb
  PIN pwr_ctrl_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END pwr_ctrl_out
  PIN qspi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END qspi_enabled
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 4.000 ;
    END
  END reset
  PIN ser_rx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.200 4.000 109.760 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.040 4.000 103.600 ;
    END
  END ser_tx
  PIN serial_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 13.440 520.000 14.000 ;
    END
  END serial_clock
  PIN serial_data_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 48.720 520.000 49.280 ;
    END
  END serial_data_1
  PIN serial_data_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 60.480 520.000 61.040 ;
    END
  END serial_data_2
  PIN serial_load
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 36.960 520.000 37.520 ;
    END
  END serial_load
  PIN serial_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 516.000 25.200 520.000 25.760 ;
    END
  END serial_resetn
  PIN spi_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.560 4.000 85.120 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.880 4.000 97.440 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.240 4.000 72.800 ;
    END
  END spi_sdoenb
  PIN spimemio_flash_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 343.280 4.000 343.840 ;
    END
  END spimemio_flash_clk
  PIN spimemio_flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.440 4.000 350.000 ;
    END
  END spimemio_flash_csb
  PIN spimemio_flash_io0_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.600 4.000 356.160 ;
    END
  END spimemio_flash_io0_di
  PIN spimemio_flash_io0_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 361.760 4.000 362.320 ;
    END
  END spimemio_flash_io0_do
  PIN spimemio_flash_io0_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 367.920 4.000 368.480 ;
    END
  END spimemio_flash_io0_oeb
  PIN spimemio_flash_io1_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END spimemio_flash_io1_di
  PIN spimemio_flash_io1_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.240 4.000 380.800 ;
    END
  END spimemio_flash_io1_do
  PIN spimemio_flash_io1_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END spimemio_flash_io1_oeb
  PIN spimemio_flash_io2_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.560 4.000 393.120 ;
    END
  END spimemio_flash_io2_di
  PIN spimemio_flash_io2_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.720 4.000 399.280 ;
    END
  END spimemio_flash_io2_do
  PIN spimemio_flash_io2_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 404.880 4.000 405.440 ;
    END
  END spimemio_flash_io2_oeb
  PIN spimemio_flash_io3_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 411.040 4.000 411.600 ;
    END
  END spimemio_flash_io3_di
  PIN spimemio_flash_io3_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.200 4.000 417.760 ;
    END
  END spimemio_flash_io3_do
  PIN spimemio_flash_io3_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END spimemio_flash_io3_oeb
  PIN trap
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.600 4.000 48.160 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 121.520 4.000 122.080 ;
    END
  END uart_enabled
  PIN user_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END user_clock
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.840 4.000 134.400 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.400 776.000 8.960 780.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.200 776.000 81.760 780.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 776.000 89.040 780.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.760 776.000 96.320 780.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 776.000 103.600 780.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.320 776.000 110.880 780.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 776.000 118.160 780.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.880 776.000 125.440 780.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 776.000 132.720 780.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 139.440 776.000 140.000 780.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 776.000 147.280 780.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 776.000 16.240 780.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.000 776.000 154.560 780.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 776.000 161.840 780.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.560 776.000 169.120 780.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 776.000 176.400 780.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.120 776.000 183.680 780.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 776.000 190.960 780.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.680 776.000 198.240 780.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 776.000 205.520 780.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.240 776.000 212.800 780.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 776.000 220.080 780.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.960 776.000 23.520 780.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.800 776.000 227.360 780.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 776.000 234.640 780.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 776.000 30.800 780.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.520 776.000 38.080 780.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 776.000 45.360 780.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.080 776.000 52.640 780.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 776.000 59.920 780.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.640 776.000 67.200 780.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 776.000 74.480 780.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 0.000 318.640 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 776.000 511.280 780.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.360 776.000 241.920 780.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 314.160 776.000 314.720 780.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 776.000 322.000 780.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 776.000 329.280 780.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 776.000 336.560 780.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.280 776.000 343.840 780.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.560 776.000 351.120 780.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.840 776.000 358.400 780.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 776.000 365.680 780.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.400 776.000 372.960 780.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 776.000 380.240 780.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 776.000 249.200 780.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.960 776.000 387.520 780.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 776.000 394.800 780.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 401.520 776.000 402.080 780.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 776.000 409.360 780.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.080 776.000 416.640 780.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 776.000 423.920 780.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.640 776.000 431.200 780.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 776.000 438.480 780.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.200 776.000 445.760 780.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 452.480 776.000 453.040 780.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.920 776.000 256.480 780.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 459.760 776.000 460.320 780.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 776.000 467.600 780.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 776.000 263.760 780.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 270.480 776.000 271.040 780.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 776.000 278.320 780.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.040 776.000 285.600 780.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 776.000 292.880 780.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.600 776.000 300.160 780.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 776.000 307.440 780.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.160 4.000 146.720 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.760 4.000 208.320 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 4.000 214.480 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.080 4.000 220.640 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.240 4.000 226.800 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.400 4.000 232.960 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.720 4.000 245.280 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.880 4.000 251.440 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.040 4.000 257.600 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.360 4.000 269.920 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.680 4.000 282.240 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 287.840 4.000 288.400 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 4.000 294.560 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 300.160 4.000 300.720 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.320 4.000 306.880 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.640 4.000 319.200 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.480 4.000 159.040 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.960 4.000 331.520 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.120 4.000 337.680 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.800 4.000 171.360 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.120 4.000 183.680 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.440 4.000 196.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END wb_dat_o[9]
  PIN wb_rstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 0.000 324.240 4.000 ;
    END
  END wb_rstn_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.320 776.000 474.880 780.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 776.000 482.160 780.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 488.880 776.000 489.440 780.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 776.000 496.720 780.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.440 776.000 504.000 780.000 ;
    END
  END wb_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 512.960 762.010 ;
      LAYER Metal2 ;
        RECT 3.500 775.700 8.100 776.580 ;
        RECT 9.260 775.700 15.380 776.580 ;
        RECT 16.540 775.700 22.660 776.580 ;
        RECT 23.820 775.700 29.940 776.580 ;
        RECT 31.100 775.700 37.220 776.580 ;
        RECT 38.380 775.700 44.500 776.580 ;
        RECT 45.660 775.700 51.780 776.580 ;
        RECT 52.940 775.700 59.060 776.580 ;
        RECT 60.220 775.700 66.340 776.580 ;
        RECT 67.500 775.700 73.620 776.580 ;
        RECT 74.780 775.700 80.900 776.580 ;
        RECT 82.060 775.700 88.180 776.580 ;
        RECT 89.340 775.700 95.460 776.580 ;
        RECT 96.620 775.700 102.740 776.580 ;
        RECT 103.900 775.700 110.020 776.580 ;
        RECT 111.180 775.700 117.300 776.580 ;
        RECT 118.460 775.700 124.580 776.580 ;
        RECT 125.740 775.700 131.860 776.580 ;
        RECT 133.020 775.700 139.140 776.580 ;
        RECT 140.300 775.700 146.420 776.580 ;
        RECT 147.580 775.700 153.700 776.580 ;
        RECT 154.860 775.700 160.980 776.580 ;
        RECT 162.140 775.700 168.260 776.580 ;
        RECT 169.420 775.700 175.540 776.580 ;
        RECT 176.700 775.700 182.820 776.580 ;
        RECT 183.980 775.700 190.100 776.580 ;
        RECT 191.260 775.700 197.380 776.580 ;
        RECT 198.540 775.700 204.660 776.580 ;
        RECT 205.820 775.700 211.940 776.580 ;
        RECT 213.100 775.700 219.220 776.580 ;
        RECT 220.380 775.700 226.500 776.580 ;
        RECT 227.660 775.700 233.780 776.580 ;
        RECT 234.940 775.700 241.060 776.580 ;
        RECT 242.220 775.700 248.340 776.580 ;
        RECT 249.500 775.700 255.620 776.580 ;
        RECT 256.780 775.700 262.900 776.580 ;
        RECT 264.060 775.700 270.180 776.580 ;
        RECT 271.340 775.700 277.460 776.580 ;
        RECT 278.620 775.700 284.740 776.580 ;
        RECT 285.900 775.700 292.020 776.580 ;
        RECT 293.180 775.700 299.300 776.580 ;
        RECT 300.460 775.700 306.580 776.580 ;
        RECT 307.740 775.700 313.860 776.580 ;
        RECT 315.020 775.700 321.140 776.580 ;
        RECT 322.300 775.700 328.420 776.580 ;
        RECT 329.580 775.700 335.700 776.580 ;
        RECT 336.860 775.700 342.980 776.580 ;
        RECT 344.140 775.700 350.260 776.580 ;
        RECT 351.420 775.700 357.540 776.580 ;
        RECT 358.700 775.700 364.820 776.580 ;
        RECT 365.980 775.700 372.100 776.580 ;
        RECT 373.260 775.700 379.380 776.580 ;
        RECT 380.540 775.700 386.660 776.580 ;
        RECT 387.820 775.700 393.940 776.580 ;
        RECT 395.100 775.700 401.220 776.580 ;
        RECT 402.380 775.700 408.500 776.580 ;
        RECT 409.660 775.700 415.780 776.580 ;
        RECT 416.940 775.700 423.060 776.580 ;
        RECT 424.220 775.700 430.340 776.580 ;
        RECT 431.500 775.700 437.620 776.580 ;
        RECT 438.780 775.700 444.900 776.580 ;
        RECT 446.060 775.700 452.180 776.580 ;
        RECT 453.340 775.700 459.460 776.580 ;
        RECT 460.620 775.700 466.740 776.580 ;
        RECT 467.900 775.700 474.020 776.580 ;
        RECT 475.180 775.700 481.300 776.580 ;
        RECT 482.460 775.700 488.580 776.580 ;
        RECT 489.740 775.700 495.860 776.580 ;
        RECT 497.020 775.700 503.140 776.580 ;
        RECT 504.300 775.700 510.420 776.580 ;
        RECT 511.580 775.700 516.180 776.580 ;
        RECT 3.500 4.300 516.180 775.700 ;
        RECT 3.500 3.500 9.780 4.300 ;
        RECT 10.940 3.500 15.380 4.300 ;
        RECT 16.540 3.500 20.980 4.300 ;
        RECT 22.140 3.500 26.580 4.300 ;
        RECT 27.740 3.500 32.180 4.300 ;
        RECT 33.340 3.500 37.780 4.300 ;
        RECT 38.940 3.500 43.380 4.300 ;
        RECT 44.540 3.500 48.980 4.300 ;
        RECT 50.140 3.500 54.580 4.300 ;
        RECT 55.740 3.500 60.180 4.300 ;
        RECT 61.340 3.500 65.780 4.300 ;
        RECT 66.940 3.500 71.380 4.300 ;
        RECT 72.540 3.500 76.980 4.300 ;
        RECT 78.140 3.500 82.580 4.300 ;
        RECT 83.740 3.500 88.180 4.300 ;
        RECT 89.340 3.500 93.780 4.300 ;
        RECT 94.940 3.500 99.380 4.300 ;
        RECT 100.540 3.500 104.980 4.300 ;
        RECT 106.140 3.500 110.580 4.300 ;
        RECT 111.740 3.500 116.180 4.300 ;
        RECT 117.340 3.500 121.780 4.300 ;
        RECT 122.940 3.500 127.380 4.300 ;
        RECT 128.540 3.500 132.980 4.300 ;
        RECT 134.140 3.500 138.580 4.300 ;
        RECT 139.740 3.500 144.180 4.300 ;
        RECT 145.340 3.500 149.780 4.300 ;
        RECT 150.940 3.500 155.380 4.300 ;
        RECT 156.540 3.500 160.980 4.300 ;
        RECT 162.140 3.500 166.580 4.300 ;
        RECT 167.740 3.500 172.180 4.300 ;
        RECT 173.340 3.500 177.780 4.300 ;
        RECT 178.940 3.500 183.380 4.300 ;
        RECT 184.540 3.500 188.980 4.300 ;
        RECT 190.140 3.500 194.580 4.300 ;
        RECT 195.740 3.500 200.180 4.300 ;
        RECT 201.340 3.500 205.780 4.300 ;
        RECT 206.940 3.500 211.380 4.300 ;
        RECT 212.540 3.500 216.980 4.300 ;
        RECT 218.140 3.500 222.580 4.300 ;
        RECT 223.740 3.500 228.180 4.300 ;
        RECT 229.340 3.500 233.780 4.300 ;
        RECT 234.940 3.500 239.380 4.300 ;
        RECT 240.540 3.500 244.980 4.300 ;
        RECT 246.140 3.500 250.580 4.300 ;
        RECT 251.740 3.500 256.180 4.300 ;
        RECT 257.340 3.500 261.780 4.300 ;
        RECT 262.940 3.500 267.380 4.300 ;
        RECT 268.540 3.500 272.980 4.300 ;
        RECT 274.140 3.500 278.580 4.300 ;
        RECT 279.740 3.500 284.180 4.300 ;
        RECT 285.340 3.500 289.780 4.300 ;
        RECT 290.940 3.500 295.380 4.300 ;
        RECT 296.540 3.500 300.980 4.300 ;
        RECT 302.140 3.500 306.580 4.300 ;
        RECT 307.740 3.500 312.180 4.300 ;
        RECT 313.340 3.500 317.780 4.300 ;
        RECT 318.940 3.500 323.380 4.300 ;
        RECT 324.540 3.500 328.980 4.300 ;
        RECT 330.140 3.500 334.580 4.300 ;
        RECT 335.740 3.500 340.180 4.300 ;
        RECT 341.340 3.500 345.780 4.300 ;
        RECT 346.940 3.500 351.380 4.300 ;
        RECT 352.540 3.500 356.980 4.300 ;
        RECT 358.140 3.500 362.580 4.300 ;
        RECT 363.740 3.500 368.180 4.300 ;
        RECT 369.340 3.500 373.780 4.300 ;
        RECT 374.940 3.500 379.380 4.300 ;
        RECT 380.540 3.500 384.980 4.300 ;
        RECT 386.140 3.500 390.580 4.300 ;
        RECT 391.740 3.500 396.180 4.300 ;
        RECT 397.340 3.500 401.780 4.300 ;
        RECT 402.940 3.500 407.380 4.300 ;
        RECT 408.540 3.500 412.980 4.300 ;
        RECT 414.140 3.500 418.580 4.300 ;
        RECT 419.740 3.500 424.180 4.300 ;
        RECT 425.340 3.500 429.780 4.300 ;
        RECT 430.940 3.500 435.380 4.300 ;
        RECT 436.540 3.500 440.980 4.300 ;
        RECT 442.140 3.500 446.580 4.300 ;
        RECT 447.740 3.500 452.180 4.300 ;
        RECT 453.340 3.500 457.780 4.300 ;
        RECT 458.940 3.500 463.380 4.300 ;
        RECT 464.540 3.500 468.980 4.300 ;
        RECT 470.140 3.500 474.580 4.300 ;
        RECT 475.740 3.500 480.180 4.300 ;
        RECT 481.340 3.500 485.780 4.300 ;
        RECT 486.940 3.500 491.380 4.300 ;
        RECT 492.540 3.500 496.980 4.300 ;
        RECT 498.140 3.500 502.580 4.300 ;
        RECT 503.740 3.500 508.180 4.300 ;
        RECT 509.340 3.500 516.180 4.300 ;
      LAYER Metal3 ;
        RECT 3.450 766.940 516.740 767.620 ;
        RECT 3.450 765.780 515.700 766.940 ;
        RECT 3.450 756.860 516.740 765.780 ;
        RECT 4.300 755.700 516.740 756.860 ;
        RECT 3.450 755.180 516.740 755.700 ;
        RECT 3.450 754.020 515.700 755.180 ;
        RECT 3.450 750.700 516.740 754.020 ;
        RECT 4.300 749.540 516.740 750.700 ;
        RECT 3.450 744.540 516.740 749.540 ;
        RECT 4.300 743.420 516.740 744.540 ;
        RECT 4.300 743.380 515.700 743.420 ;
        RECT 3.450 742.260 515.700 743.380 ;
        RECT 3.450 738.380 516.740 742.260 ;
        RECT 4.300 737.220 516.740 738.380 ;
        RECT 3.450 732.220 516.740 737.220 ;
        RECT 4.300 731.660 516.740 732.220 ;
        RECT 4.300 731.060 515.700 731.660 ;
        RECT 3.450 730.500 515.700 731.060 ;
        RECT 3.450 726.060 516.740 730.500 ;
        RECT 4.300 724.900 516.740 726.060 ;
        RECT 3.450 719.900 516.740 724.900 ;
        RECT 4.300 718.740 515.700 719.900 ;
        RECT 3.450 713.740 516.740 718.740 ;
        RECT 4.300 712.580 516.740 713.740 ;
        RECT 3.450 708.140 516.740 712.580 ;
        RECT 3.450 707.580 515.700 708.140 ;
        RECT 4.300 706.980 515.700 707.580 ;
        RECT 4.300 706.420 516.740 706.980 ;
        RECT 3.450 701.420 516.740 706.420 ;
        RECT 4.300 700.260 516.740 701.420 ;
        RECT 3.450 696.380 516.740 700.260 ;
        RECT 3.450 695.260 515.700 696.380 ;
        RECT 4.300 695.220 515.700 695.260 ;
        RECT 4.300 694.100 516.740 695.220 ;
        RECT 3.450 689.100 516.740 694.100 ;
        RECT 4.300 687.940 516.740 689.100 ;
        RECT 3.450 684.620 516.740 687.940 ;
        RECT 3.450 683.460 515.700 684.620 ;
        RECT 3.450 682.940 516.740 683.460 ;
        RECT 4.300 681.780 516.740 682.940 ;
        RECT 3.450 676.780 516.740 681.780 ;
        RECT 4.300 675.620 516.740 676.780 ;
        RECT 3.450 672.860 516.740 675.620 ;
        RECT 3.450 671.700 515.700 672.860 ;
        RECT 3.450 670.620 516.740 671.700 ;
        RECT 4.300 669.460 516.740 670.620 ;
        RECT 3.450 664.460 516.740 669.460 ;
        RECT 4.300 663.300 516.740 664.460 ;
        RECT 3.450 661.100 516.740 663.300 ;
        RECT 3.450 659.940 515.700 661.100 ;
        RECT 3.450 658.300 516.740 659.940 ;
        RECT 4.300 657.140 516.740 658.300 ;
        RECT 3.450 652.140 516.740 657.140 ;
        RECT 4.300 650.980 516.740 652.140 ;
        RECT 3.450 649.340 516.740 650.980 ;
        RECT 3.450 648.180 515.700 649.340 ;
        RECT 3.450 645.980 516.740 648.180 ;
        RECT 4.300 644.820 516.740 645.980 ;
        RECT 3.450 639.820 516.740 644.820 ;
        RECT 4.300 638.660 516.740 639.820 ;
        RECT 3.450 637.580 516.740 638.660 ;
        RECT 3.450 636.420 515.700 637.580 ;
        RECT 3.450 633.660 516.740 636.420 ;
        RECT 4.300 632.500 516.740 633.660 ;
        RECT 3.450 627.500 516.740 632.500 ;
        RECT 4.300 626.340 516.740 627.500 ;
        RECT 3.450 625.820 516.740 626.340 ;
        RECT 3.450 624.660 515.700 625.820 ;
        RECT 3.450 621.340 516.740 624.660 ;
        RECT 4.300 620.180 516.740 621.340 ;
        RECT 3.450 615.180 516.740 620.180 ;
        RECT 4.300 614.060 516.740 615.180 ;
        RECT 4.300 614.020 515.700 614.060 ;
        RECT 3.450 612.900 515.700 614.020 ;
        RECT 3.450 609.020 516.740 612.900 ;
        RECT 4.300 607.860 516.740 609.020 ;
        RECT 3.450 602.860 516.740 607.860 ;
        RECT 4.300 602.300 516.740 602.860 ;
        RECT 4.300 601.700 515.700 602.300 ;
        RECT 3.450 601.140 515.700 601.700 ;
        RECT 3.450 596.700 516.740 601.140 ;
        RECT 4.300 595.540 516.740 596.700 ;
        RECT 3.450 590.540 516.740 595.540 ;
        RECT 4.300 589.380 515.700 590.540 ;
        RECT 3.450 584.380 516.740 589.380 ;
        RECT 4.300 583.220 516.740 584.380 ;
        RECT 3.450 578.780 516.740 583.220 ;
        RECT 3.450 578.220 515.700 578.780 ;
        RECT 4.300 577.620 515.700 578.220 ;
        RECT 4.300 577.060 516.740 577.620 ;
        RECT 3.450 572.060 516.740 577.060 ;
        RECT 4.300 570.900 516.740 572.060 ;
        RECT 3.450 567.020 516.740 570.900 ;
        RECT 3.450 565.900 515.700 567.020 ;
        RECT 4.300 565.860 515.700 565.900 ;
        RECT 4.300 564.740 516.740 565.860 ;
        RECT 3.450 559.740 516.740 564.740 ;
        RECT 4.300 558.580 516.740 559.740 ;
        RECT 3.450 555.260 516.740 558.580 ;
        RECT 3.450 554.100 515.700 555.260 ;
        RECT 3.450 553.580 516.740 554.100 ;
        RECT 4.300 552.420 516.740 553.580 ;
        RECT 3.450 547.420 516.740 552.420 ;
        RECT 4.300 546.260 516.740 547.420 ;
        RECT 3.450 543.500 516.740 546.260 ;
        RECT 3.450 542.340 515.700 543.500 ;
        RECT 3.450 541.260 516.740 542.340 ;
        RECT 4.300 540.100 516.740 541.260 ;
        RECT 3.450 535.100 516.740 540.100 ;
        RECT 4.300 533.940 516.740 535.100 ;
        RECT 3.450 531.740 516.740 533.940 ;
        RECT 3.450 530.580 515.700 531.740 ;
        RECT 3.450 528.940 516.740 530.580 ;
        RECT 4.300 527.780 516.740 528.940 ;
        RECT 3.450 522.780 516.740 527.780 ;
        RECT 4.300 521.620 516.740 522.780 ;
        RECT 3.450 519.980 516.740 521.620 ;
        RECT 3.450 518.820 515.700 519.980 ;
        RECT 3.450 516.620 516.740 518.820 ;
        RECT 4.300 515.460 516.740 516.620 ;
        RECT 3.450 510.460 516.740 515.460 ;
        RECT 4.300 509.300 516.740 510.460 ;
        RECT 3.450 508.220 516.740 509.300 ;
        RECT 3.450 507.060 515.700 508.220 ;
        RECT 3.450 504.300 516.740 507.060 ;
        RECT 4.300 503.140 516.740 504.300 ;
        RECT 3.450 498.140 516.740 503.140 ;
        RECT 4.300 496.980 516.740 498.140 ;
        RECT 3.450 496.460 516.740 496.980 ;
        RECT 3.450 495.300 515.700 496.460 ;
        RECT 3.450 491.980 516.740 495.300 ;
        RECT 4.300 490.820 516.740 491.980 ;
        RECT 3.450 485.820 516.740 490.820 ;
        RECT 4.300 484.700 516.740 485.820 ;
        RECT 4.300 484.660 515.700 484.700 ;
        RECT 3.450 483.540 515.700 484.660 ;
        RECT 3.450 479.660 516.740 483.540 ;
        RECT 4.300 478.500 516.740 479.660 ;
        RECT 3.450 473.500 516.740 478.500 ;
        RECT 4.300 472.940 516.740 473.500 ;
        RECT 4.300 472.340 515.700 472.940 ;
        RECT 3.450 471.780 515.700 472.340 ;
        RECT 3.450 467.340 516.740 471.780 ;
        RECT 4.300 466.180 516.740 467.340 ;
        RECT 3.450 461.180 516.740 466.180 ;
        RECT 4.300 460.020 515.700 461.180 ;
        RECT 3.450 455.020 516.740 460.020 ;
        RECT 4.300 453.860 516.740 455.020 ;
        RECT 3.450 449.420 516.740 453.860 ;
        RECT 3.450 448.860 515.700 449.420 ;
        RECT 4.300 448.260 515.700 448.860 ;
        RECT 4.300 447.700 516.740 448.260 ;
        RECT 3.450 442.700 516.740 447.700 ;
        RECT 4.300 441.540 516.740 442.700 ;
        RECT 3.450 437.660 516.740 441.540 ;
        RECT 3.450 436.540 515.700 437.660 ;
        RECT 4.300 436.500 515.700 436.540 ;
        RECT 4.300 435.380 516.740 436.500 ;
        RECT 3.450 430.380 516.740 435.380 ;
        RECT 4.300 429.220 516.740 430.380 ;
        RECT 3.450 425.900 516.740 429.220 ;
        RECT 3.450 424.740 515.700 425.900 ;
        RECT 3.450 424.220 516.740 424.740 ;
        RECT 4.300 423.060 516.740 424.220 ;
        RECT 3.450 418.060 516.740 423.060 ;
        RECT 4.300 416.900 516.740 418.060 ;
        RECT 3.450 414.140 516.740 416.900 ;
        RECT 3.450 412.980 515.700 414.140 ;
        RECT 3.450 411.900 516.740 412.980 ;
        RECT 4.300 410.740 516.740 411.900 ;
        RECT 3.450 405.740 516.740 410.740 ;
        RECT 4.300 404.580 516.740 405.740 ;
        RECT 3.450 402.380 516.740 404.580 ;
        RECT 3.450 401.220 515.700 402.380 ;
        RECT 3.450 399.580 516.740 401.220 ;
        RECT 4.300 398.420 516.740 399.580 ;
        RECT 3.450 393.420 516.740 398.420 ;
        RECT 4.300 392.260 516.740 393.420 ;
        RECT 3.450 390.620 516.740 392.260 ;
        RECT 3.450 389.460 515.700 390.620 ;
        RECT 3.450 387.260 516.740 389.460 ;
        RECT 4.300 386.100 516.740 387.260 ;
        RECT 3.450 381.100 516.740 386.100 ;
        RECT 4.300 379.940 516.740 381.100 ;
        RECT 3.450 378.860 516.740 379.940 ;
        RECT 3.450 377.700 515.700 378.860 ;
        RECT 3.450 374.940 516.740 377.700 ;
        RECT 4.300 373.780 516.740 374.940 ;
        RECT 3.450 368.780 516.740 373.780 ;
        RECT 4.300 367.620 516.740 368.780 ;
        RECT 3.450 367.100 516.740 367.620 ;
        RECT 3.450 365.940 515.700 367.100 ;
        RECT 3.450 362.620 516.740 365.940 ;
        RECT 4.300 361.460 516.740 362.620 ;
        RECT 3.450 356.460 516.740 361.460 ;
        RECT 4.300 355.340 516.740 356.460 ;
        RECT 4.300 355.300 515.700 355.340 ;
        RECT 3.450 354.180 515.700 355.300 ;
        RECT 3.450 350.300 516.740 354.180 ;
        RECT 4.300 349.140 516.740 350.300 ;
        RECT 3.450 344.140 516.740 349.140 ;
        RECT 4.300 343.580 516.740 344.140 ;
        RECT 4.300 342.980 515.700 343.580 ;
        RECT 3.450 342.420 515.700 342.980 ;
        RECT 3.450 337.980 516.740 342.420 ;
        RECT 4.300 336.820 516.740 337.980 ;
        RECT 3.450 331.820 516.740 336.820 ;
        RECT 4.300 330.660 515.700 331.820 ;
        RECT 3.450 325.660 516.740 330.660 ;
        RECT 4.300 324.500 516.740 325.660 ;
        RECT 3.450 320.060 516.740 324.500 ;
        RECT 3.450 319.500 515.700 320.060 ;
        RECT 4.300 318.900 515.700 319.500 ;
        RECT 4.300 318.340 516.740 318.900 ;
        RECT 3.450 313.340 516.740 318.340 ;
        RECT 4.300 312.180 516.740 313.340 ;
        RECT 3.450 308.300 516.740 312.180 ;
        RECT 3.450 307.180 515.700 308.300 ;
        RECT 4.300 307.140 515.700 307.180 ;
        RECT 4.300 306.020 516.740 307.140 ;
        RECT 3.450 301.020 516.740 306.020 ;
        RECT 4.300 299.860 516.740 301.020 ;
        RECT 3.450 296.540 516.740 299.860 ;
        RECT 3.450 295.380 515.700 296.540 ;
        RECT 3.450 294.860 516.740 295.380 ;
        RECT 4.300 293.700 516.740 294.860 ;
        RECT 3.450 288.700 516.740 293.700 ;
        RECT 4.300 287.540 516.740 288.700 ;
        RECT 3.450 284.780 516.740 287.540 ;
        RECT 3.450 283.620 515.700 284.780 ;
        RECT 3.450 282.540 516.740 283.620 ;
        RECT 4.300 281.380 516.740 282.540 ;
        RECT 3.450 276.380 516.740 281.380 ;
        RECT 4.300 275.220 516.740 276.380 ;
        RECT 3.450 273.020 516.740 275.220 ;
        RECT 3.450 271.860 515.700 273.020 ;
        RECT 3.450 270.220 516.740 271.860 ;
        RECT 4.300 269.060 516.740 270.220 ;
        RECT 3.450 264.060 516.740 269.060 ;
        RECT 4.300 262.900 516.740 264.060 ;
        RECT 3.450 261.260 516.740 262.900 ;
        RECT 3.450 260.100 515.700 261.260 ;
        RECT 3.450 257.900 516.740 260.100 ;
        RECT 4.300 256.740 516.740 257.900 ;
        RECT 3.450 251.740 516.740 256.740 ;
        RECT 4.300 250.580 516.740 251.740 ;
        RECT 3.450 249.500 516.740 250.580 ;
        RECT 3.450 248.340 515.700 249.500 ;
        RECT 3.450 245.580 516.740 248.340 ;
        RECT 4.300 244.420 516.740 245.580 ;
        RECT 3.450 239.420 516.740 244.420 ;
        RECT 4.300 238.260 516.740 239.420 ;
        RECT 3.450 237.740 516.740 238.260 ;
        RECT 3.450 236.580 515.700 237.740 ;
        RECT 3.450 233.260 516.740 236.580 ;
        RECT 4.300 232.100 516.740 233.260 ;
        RECT 3.450 227.100 516.740 232.100 ;
        RECT 4.300 225.980 516.740 227.100 ;
        RECT 4.300 225.940 515.700 225.980 ;
        RECT 3.450 224.820 515.700 225.940 ;
        RECT 3.450 220.940 516.740 224.820 ;
        RECT 4.300 219.780 516.740 220.940 ;
        RECT 3.450 214.780 516.740 219.780 ;
        RECT 4.300 214.220 516.740 214.780 ;
        RECT 4.300 213.620 515.700 214.220 ;
        RECT 3.450 213.060 515.700 213.620 ;
        RECT 3.450 208.620 516.740 213.060 ;
        RECT 4.300 207.460 516.740 208.620 ;
        RECT 3.450 202.460 516.740 207.460 ;
        RECT 4.300 201.300 515.700 202.460 ;
        RECT 3.450 196.300 516.740 201.300 ;
        RECT 4.300 195.140 516.740 196.300 ;
        RECT 3.450 190.700 516.740 195.140 ;
        RECT 3.450 190.140 515.700 190.700 ;
        RECT 4.300 189.540 515.700 190.140 ;
        RECT 4.300 188.980 516.740 189.540 ;
        RECT 3.450 183.980 516.740 188.980 ;
        RECT 4.300 182.820 516.740 183.980 ;
        RECT 3.450 178.940 516.740 182.820 ;
        RECT 3.450 177.820 515.700 178.940 ;
        RECT 4.300 177.780 515.700 177.820 ;
        RECT 4.300 176.660 516.740 177.780 ;
        RECT 3.450 171.660 516.740 176.660 ;
        RECT 4.300 170.500 516.740 171.660 ;
        RECT 3.450 167.180 516.740 170.500 ;
        RECT 3.450 166.020 515.700 167.180 ;
        RECT 3.450 165.500 516.740 166.020 ;
        RECT 4.300 164.340 516.740 165.500 ;
        RECT 3.450 159.340 516.740 164.340 ;
        RECT 4.300 158.180 516.740 159.340 ;
        RECT 3.450 155.420 516.740 158.180 ;
        RECT 3.450 154.260 515.700 155.420 ;
        RECT 3.450 153.180 516.740 154.260 ;
        RECT 4.300 152.020 516.740 153.180 ;
        RECT 3.450 147.020 516.740 152.020 ;
        RECT 4.300 145.860 516.740 147.020 ;
        RECT 3.450 143.660 516.740 145.860 ;
        RECT 3.450 142.500 515.700 143.660 ;
        RECT 3.450 140.860 516.740 142.500 ;
        RECT 4.300 139.700 516.740 140.860 ;
        RECT 3.450 134.700 516.740 139.700 ;
        RECT 4.300 133.540 516.740 134.700 ;
        RECT 3.450 131.900 516.740 133.540 ;
        RECT 3.450 130.740 515.700 131.900 ;
        RECT 3.450 128.540 516.740 130.740 ;
        RECT 4.300 127.380 516.740 128.540 ;
        RECT 3.450 122.380 516.740 127.380 ;
        RECT 4.300 121.220 516.740 122.380 ;
        RECT 3.450 120.140 516.740 121.220 ;
        RECT 3.450 118.980 515.700 120.140 ;
        RECT 3.450 116.220 516.740 118.980 ;
        RECT 4.300 115.060 516.740 116.220 ;
        RECT 3.450 110.060 516.740 115.060 ;
        RECT 4.300 108.900 516.740 110.060 ;
        RECT 3.450 108.380 516.740 108.900 ;
        RECT 3.450 107.220 515.700 108.380 ;
        RECT 3.450 103.900 516.740 107.220 ;
        RECT 4.300 102.740 516.740 103.900 ;
        RECT 3.450 97.740 516.740 102.740 ;
        RECT 4.300 96.620 516.740 97.740 ;
        RECT 4.300 96.580 515.700 96.620 ;
        RECT 3.450 95.460 515.700 96.580 ;
        RECT 3.450 91.580 516.740 95.460 ;
        RECT 4.300 90.420 516.740 91.580 ;
        RECT 3.450 85.420 516.740 90.420 ;
        RECT 4.300 84.860 516.740 85.420 ;
        RECT 4.300 84.260 515.700 84.860 ;
        RECT 3.450 83.700 515.700 84.260 ;
        RECT 3.450 79.260 516.740 83.700 ;
        RECT 4.300 78.100 516.740 79.260 ;
        RECT 3.450 73.100 516.740 78.100 ;
        RECT 4.300 71.940 515.700 73.100 ;
        RECT 3.450 66.940 516.740 71.940 ;
        RECT 4.300 65.780 516.740 66.940 ;
        RECT 3.450 61.340 516.740 65.780 ;
        RECT 3.450 60.780 515.700 61.340 ;
        RECT 4.300 60.180 515.700 60.780 ;
        RECT 4.300 59.620 516.740 60.180 ;
        RECT 3.450 54.620 516.740 59.620 ;
        RECT 4.300 53.460 516.740 54.620 ;
        RECT 3.450 49.580 516.740 53.460 ;
        RECT 3.450 48.460 515.700 49.580 ;
        RECT 4.300 48.420 515.700 48.460 ;
        RECT 4.300 47.300 516.740 48.420 ;
        RECT 3.450 42.300 516.740 47.300 ;
        RECT 4.300 41.140 516.740 42.300 ;
        RECT 3.450 37.820 516.740 41.140 ;
        RECT 3.450 36.660 515.700 37.820 ;
        RECT 3.450 36.140 516.740 36.660 ;
        RECT 4.300 34.980 516.740 36.140 ;
        RECT 3.450 29.980 516.740 34.980 ;
        RECT 4.300 28.820 516.740 29.980 ;
        RECT 3.450 26.060 516.740 28.820 ;
        RECT 3.450 24.900 515.700 26.060 ;
        RECT 3.450 23.820 516.740 24.900 ;
        RECT 4.300 22.660 516.740 23.820 ;
        RECT 3.450 14.300 516.740 22.660 ;
        RECT 3.450 13.140 515.700 14.300 ;
        RECT 3.450 8.540 516.740 13.140 ;
      LAYER Metal4 ;
        RECT 5.180 16.330 21.940 765.430 ;
        RECT 24.140 16.330 25.240 765.430 ;
        RECT 27.440 16.330 98.740 765.430 ;
        RECT 100.940 16.330 102.040 765.430 ;
        RECT 104.240 16.330 175.540 765.430 ;
        RECT 177.740 16.330 178.840 765.430 ;
        RECT 181.040 16.330 252.340 765.430 ;
        RECT 254.540 16.330 255.640 765.430 ;
        RECT 257.840 16.330 329.140 765.430 ;
        RECT 331.340 16.330 332.440 765.430 ;
        RECT 334.640 16.330 405.940 765.430 ;
        RECT 408.140 16.330 409.240 765.430 ;
        RECT 411.440 16.330 482.740 765.430 ;
        RECT 484.940 16.330 486.040 765.430 ;
        RECT 488.240 16.330 511.140 765.430 ;
      LAYER Metal5 ;
        RECT 6.220 743.390 510.100 758.740 ;
        RECT 6.220 713.390 510.100 740.790 ;
        RECT 6.220 683.390 510.100 710.790 ;
        RECT 6.220 653.390 510.100 680.790 ;
        RECT 6.220 623.390 510.100 650.790 ;
        RECT 6.220 593.390 510.100 620.790 ;
        RECT 6.220 563.390 510.100 590.790 ;
        RECT 6.220 533.390 510.100 560.790 ;
        RECT 6.220 503.390 510.100 530.790 ;
        RECT 6.220 473.390 510.100 500.790 ;
        RECT 6.220 443.390 510.100 470.790 ;
        RECT 6.220 413.390 510.100 440.790 ;
        RECT 6.220 383.390 510.100 410.790 ;
        RECT 6.220 353.390 510.100 380.790 ;
        RECT 6.220 323.390 510.100 350.790 ;
        RECT 6.220 293.390 510.100 320.790 ;
        RECT 6.220 263.390 510.100 290.790 ;
        RECT 6.220 233.390 510.100 260.790 ;
        RECT 6.220 203.390 510.100 230.790 ;
        RECT 6.220 173.390 510.100 200.790 ;
        RECT 6.220 143.390 510.100 170.790 ;
        RECT 6.220 113.390 510.100 140.790 ;
        RECT 6.220 83.390 510.100 110.790 ;
        RECT 6.220 53.390 510.100 80.790 ;
        RECT 6.220 28.060 510.100 50.790 ;
  END
END housekeeping
END LIBRARY

