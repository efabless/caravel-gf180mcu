* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_100_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6914_ _6914_/D _7218_/RN _6914_/CLK _7329_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ _6845_/D _7170_/RN _6845_/CLK _6845_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3988_ _3988_/I0 _6658_/Q _3988_/S _6658_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6776_ _6776_/D _7218_/RN _6776_/CLK _6776_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5727_ hold2/Z hold117/Z _5727_/S _5727_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5658_ hold655/Z hold291/Z hold56/Z _7013_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4609_ _4601_/Z _5285_/B _4607_/Z _5021_/B _4612_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5589_ hold151/Z hold48/Z _5592_/S _5589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold362 _7271_/Q hold362/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7328_ _7328_/I _7328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold351 _5624_/Z _6983_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold340 _5633_/Z _6991_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold384 _7210_/Q hold384/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold395 _5594_/Z _6956_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7259_ _7259_/D _7260_/RN _7260_/CLK _7259_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold373 _7091_/Q hold373/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_461 net813_461/I _6704_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_472 net413_59/I _6693_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_494 net413_88/I _6671_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_483 net813_483/I _6682_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f__1062_ clkbuf_0__1062_/Z _4309_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _5420_/A3 _5420_/A2 _5270_/A1 _4761_/I _4960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_91_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _5315_/A2 _4524_/Z _4675_/Z _4700_/Z _4891_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3911_ _3485_/Z _3525_/Z _3913_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _7170_/RN _6652_/A2 _6630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3842_ _3519_/Z _3537_/Z _3950_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6561_ _6561_/A1 _7261_/Q _6833_/D _6561_/B2 _6562_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3773_ _3773_/A1 _3773_/A2 _3773_/A3 _3773_/A4 _3773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5512_ hold291/Z hold839/Z _5512_/S _5512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6492_ _6492_/A1 _6492_/A2 _6492_/A3 _6492_/A4 _6492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _5443_/A1 _5245_/Z _5444_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_161_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5374_ _5374_/A1 _5374_/A2 _5374_/A3 _5374_/A4 _5374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7113_ _7113_/D _7237_/RN _7113_/CLK _7113_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4325_ hold291/Z hold897/Z _4325_/S _4325_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4256_ hold91/Z hold452/Z _4261_/S _4256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7044_ _7044_/D _7258_/RN _7044_/CLK _7044_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_95_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4187_ hold291/Z hold745/Z _4187_/S _4187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6828_ _6828_/D _7279_/RN _7279_/CLK _6828_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _6759_/D _7258_/RN _6759_/CLK _7314_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold170 _7066_/Q hold170/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold181 _4156_/Z _6704_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold192 _7073_/Q hold192/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_59_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5090_ _5090_/A1 _5090_/A2 _5400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4110_ hold65/Z hold282/Z _4118_/S _4110_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4041_ _3425_/S _7283_/Q _4041_/A3 _4041_/B1 _3409_/Z _6733_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_151_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_3_0__1359_ clkbuf_0__1359_/Z _4073__7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_49_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _5992_/A1 _5991_/Z _5995_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4943_ _4759_/Z _4903_/Z _5330_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_91_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4874_ _4641_/Z _4833_/Z _4874_/B _4874_/C _4876_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_32_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6613_ hold909/Z hold291/Z _6613_/S _6613_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3825_ _3519_/Z _3527_/Z _3933_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3756_ _6685_/Q _3945_/C2 _3941_/A2 _7161_/Q _3757_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6544_ _6711_/Q _5948_/Z _6261_/Z _6810_/Q _6546_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _6475_/I _6476_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _3401_/I _4369_/Z _5172_/B _5172_/C _5426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_118_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3687_ _3687_/A1 _3687_/A2 _3687_/A3 _3686_/Z _3687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_133_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput253 _4079_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput242 _7311_/Z mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput220 _4062_/Z mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput231 _7308_/Z mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5357_ _5357_/A1 _5357_/A2 _5357_/A3 _5357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_58_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput264 _6880_/Q pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput286 _6673_/Q pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput275 _6679_/Q pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _5288_/A1 _5468_/A2 _5288_/B _5288_/C _5292_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_114_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput297 _6892_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _6567_/I0 _6814_/Q _4312_/S _6814_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4239_ _4238_/Z hold795/Z _4245_/S _4239_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7027_ _7027_/D _7258_/RN _7027_/CLK _7027_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_28_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4590_ _4454_/Z _4878_/A2 _5364_/B _4586_/Z _4590_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3610_ _6571_/I0 _6874_/Q _3898_/S _3610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _3485_/Z _3540_/Z _4210_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_171_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold928 _5684_/Z _7036_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold917 _7094_/Q hold917/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold906 _4352_/Z _6852_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_31_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3472_ _3472_/I0 hold14/Z hold54/I hold15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_127_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold939 _7150_/Q hold939/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6260_ _6260_/A1 _6260_/A2 _6260_/A3 _6259_/Z _6260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_170_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _4892_/B _4683_/Z _5211_/B _5211_/C _5396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_130_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6191_ _7076_/Q _5965_/Z _5980_/Z _6694_/Q _5967_/Z _6720_/Q _6193_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5142_ _5281_/C _4539_/I _4817_/Z _5287_/B _4547_/Z _5470_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_9_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5073_ _4699_/Z _5255_/B _5073_/B _5335_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_111_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ _4024_/I _6731_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5975_ _7044_/Q _7228_/Q _7227_/Q _6211_/A2 _5975_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _5324_/A1 _4926_/A2 _4926_/B _4929_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _4614_/Z _4833_/Z _5289_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet563_219 net763_423/I _7006_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _3537_/Z _3617_/Z _5728_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet563_208 net563_225/I _7017_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4788_ _5414_/A2 _5218_/B _5125_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6527_ _6554_/A1 _6521_/Z _6526_/Z _6527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_174_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3739_ _3739_/A1 _3739_/A2 _3739_/A3 _3739_/A4 _3739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6458_ _7116_/Q _6240_/Z _6297_/Z _6704_/Q _6459_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5409_ _5334_/Z _5409_/A2 _5448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6389_ _7031_/Q _6269_/Z _6273_/Z hold69/I _6390_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_102_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5760_ hold955/Z hold291/Z _5766_/S _5760_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5691_ hold334/Z hold2/Z _5691_/S _5691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4711_ _5302_/B _5099_/A1 _5099_/A2 _4703_/Z _4711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4642_ _5315_/A1 _5315_/A2 _4551_/Z _5364_/B _5038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_30_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4573_ _4551_/Z _5364_/B _5471_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_129_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold703 _6893_/Q hold703/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7292_ _7292_/D _6646_/Z _7305_/CLK _7292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_171_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3524_ _3509_/Z _3523_/Z _3957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6312_ _6989_/Q _6533_/A2 _6533_/A3 _6533_/A4 _6318_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold725 _6711_/Q hold725/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold714 _4336_/Z _6841_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold736 _4355_/Z _6854_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3455_ hold11/Z hold19/Z _3460_/S _7289_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold769 _6762_/Q hold769/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6243_ _6484_/A2 _6533_/A4 _6285_/A2 _6302_/A4 _6243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold747 _6838_/Q hold747/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold758 _4181_/Z _6721_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_118_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3386_ _7228_/Q _6021_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_6174_ _7067_/Q _5985_/Z _6000_/Z _7133_/Q _6174_/C _6180_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5125_ _5317_/A1 _5123_/Z _5125_/A3 _5126_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_69_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _4699_/Z _5051_/Z _5056_/B _5056_/C _5057_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_85_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4007_ _3990_/I _4006_/Z _4008_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54__1359_ net663_324/I net413_95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_134__1359_ net513_165/I net713_385/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_179_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5958_ _7228_/Q _7227_/Q _6210_/C _6210_/A2 _5958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_25_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _4500_/Z _5072_/A4 _4436_/B _4494_/Z _4909_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_179_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5889_ hold48/Z hold749/Z _5892_/S _5889_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold41 hold41/I hold41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_88_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold30 hold30/I hold30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold52 hold52/I hold52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold63 hold63/I hold63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold74 hold74/I hold74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_57_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold96 hold96/I hold96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold85 hold85/I hold85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_35_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _4067_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_5 _6811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6930_ _6930_/D _7256_/RN _6930_/CLK _6930_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_94_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _6861_/D _7279_/RN _7269_/CLK _6861_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5812_ _3515_/Z _3552_/Z _5520_/C _5820_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_63_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6792_ _6792_/D _7265_/CLK _6792_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ hold91/Z hold590/Z _5748_/S _5743_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5674_ _5674_/A1 hold32/Z hold33/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_31_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4625_ _4887_/A1 _4868_/A1 _4551_/Z _5364_/B _4625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4556_ _4528_/Z _4536_/Z _4556_/A3 _4547_/Z _4556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold500 _7219_/Q hold500/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold511 _6688_/Q hold511/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold522 _5789_/Z _7129_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold533 _7145_/Q hold533/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3507_ hold320/Z _3497_/I _3501_/Z _3489_/I _3507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold544 _6686_/Q hold544/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7275_ _7275_/D _7279_/RN _7279_/CLK _7275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4487_ _4687_/A2 _4687_/A3 _5220_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold555 _5744_/Z _7089_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold588 _7038_/Q hold588/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold577 _5704_/Z _7054_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold566 _7006_/Q hold566/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3438_ input58/Z _3438_/I1 _3438_/S _7295_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold599 _5869_/Z _7200_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6226_ _6727_/Q _5994_/I _6226_/B _6227_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_140_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6157_ _7116_/Q _5984_/Z _5997_/Z _7100_/Q _7074_/Q _5980_/Z _6158_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3369_ _7007_/Q _3369_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5108_ _5400_/A1 _5108_/A2 _5310_/C _5107_/I _5108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_57_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ _6088_/I _6089_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5039_ _5035_/Z _5036_/Z _5205_/C _5039_/A4 _5040_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput120 wb_adr_i[3] _4456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_163_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput142 wb_dat_i[22] _6597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput131 wb_dat_i[12] _6591_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput153 wb_dat_i[3] _3396_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_103_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput164 wb_sel_i[3] _6575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_60_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4410_ _4412_/B _4412_/C _5003_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_172_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _5390_/A1 _5390_/A2 _5350_/Z _5390_/A4 _5390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_172_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _3529_/Z hold674/Z _5520_/C _4341_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_28_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7060_ _7060_/D _7258_/RN _7060_/CLK _7060_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4272_ _4103_/I hold681/Z _4273_/S _4272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6011_ _6011_/A1 _6558_/S _6011_/B1 _6310_/A3 _7241_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_113_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6913_ _6913_/D _7218_/RN _6913_/CLK _7328_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _6844_/D _7170_/RN _6844_/CLK _6844_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3987_ _6733_/Q _3972_/Z _3987_/A3 _3987_/B _3988_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_6775_ _6775_/D _7218_/RN _6775_/CLK _6775_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ hold12/Z hold172/Z _5727_/S _5726_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5657_ hold262/Z hold227/Z hold56/Z _7012_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4608_ _4551_/Z _4501_/B _4853_/A1 _5364_/B _5021_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_151_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5588_ hold101/Z hold65/Z _5592_/S _5588_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7327_ _7327_/I _7327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4539_ _4539_/I _5281_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_117_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold341 _7047_/Q hold341/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold330 _5862_/Z _7194_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold352 _7169_/Q hold352/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold363 _4105_/Z hold363/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_120_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _7258_/D _7258_/RN _7258_/CLK _7258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold385 _5880_/Z _7210_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold396 _6988_/Q hold396/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold374 _5746_/Z _7091_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6209_ _7297_/Q _5969_/Z _6227_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7189_ _7189_/D _7237_/RN _7189_/CLK _7189_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_131_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet813_462 net813_464/I _6703_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_473 net813_473/I _6692_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_484 net813_488/I _6681_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_495 net413_88/I _6670_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _4890_/I _5259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3910_ _6932_/Q _3910_/A2 _3953_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3841_ _6695_/Q _4143_/A1 _3868_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6560_ _6561_/B2 _6559_/Z _6561_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3772_ _7216_/Q _3912_/A2 _3930_/A2 _7128_/Q _3773_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_186_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5511_ hold227/Z hold380/Z _5512_/S _5511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6491_ _7173_/Q _5948_/Z _6261_/Z _6963_/Q _6266_/Z _7019_/Q _6492_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5442_ _5056_/C _5442_/A2 _5442_/A3 _5442_/A4 _5442_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_121_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5373_ _5287_/C _4551_/Z _5287_/B _5373_/B _5374_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_160_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7112_ _7112_/D _7256_/RN _7112_/CLK _7112_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4324_ _4103_/I hold853/Z _4325_/S _4324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7043_ _7043_/D _7256_/RN _7043_/CLK _7043_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4255_ hold291/Z hold817/Z _4261_/S _4255_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4186_ _4103_/I hold705/Z _4187_/S _4186_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _6827_/D _7279_/RN _7278_/CLK _6833_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_11_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6758_ _6758_/D _7258_/RN _6758_/CLK _7313_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5709_ hold127/Z hold2/Z _5709_/S _5709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6689_ _6689_/D _7008_/RN _6689_/CLK _6689_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_164_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold171 _5717_/Z _7066_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold160 _5625_/Z _6984_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold193 _5725_/Z _7073_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold182 _7331_/I hold182/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_78_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4040_ _4040_/I _6734_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _7231_/Q _7228_/Q _7227_/Q _5991_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_52_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4942_ _4939_/Z _4942_/A2 _5062_/B _4948_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_52_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_90 net413_91/I _7135_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4873_ _4641_/Z _5051_/S _5287_/B _4681_/Z _4874_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6612_ hold877/Z _4103_/I _6613_/S _6612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3824_ _3529_/Z _3653_/Z _3935_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_159_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3755_ _6951_/Q _5584_/A1 _3956_/A2 _7121_/Q _7145_/Q _3951_/C1 _3757_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6543_ _6852_/Q _6274_/Z _6285_/Z _6693_/Q _6707_/Q _6254_/Z _6546_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6474_ _6744_/Q _7256_/Q _6474_/B _6475_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3686_ _3686_/A1 _3686_/A2 _3686_/A3 _3686_/A4 _3686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _5425_/A1 _5425_/A2 _5425_/A3 _5425_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xoutput210 _4056_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput232 _7329_/Z mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput221 _7319_/Z mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput243 _4059_/Z mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5356_ _5356_/A1 _5387_/A2 _5356_/B _5356_/C _5357_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput254 _7332_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput276 _6680_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput265 _6881_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5287_ _4554_/Z _4683_/Z _5287_/B _5287_/C _5487_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_101_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput298 _3907_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4307_ _6566_/I0 _6813_/Q _4312_/S _6813_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput287 _6889_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4238_ hold411/Z hold48/Z _4244_/S _4238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7026_ _7026_/D _7258_/RN _7026_/CLK _7026_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4169_ hold291/Z hold915/Z _4169_/S _4169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3540_ _3653_/A1 _3617_/A1 hold673/Z _3492_/Z _3540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_182_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold918 _5750_/Z _7094_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold907 _7077_/Q hold907/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_31_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5210_ _5209_/Z _5208_/Z _5417_/A1 _5210_/A4 _5210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3471_ _3471_/I _3472_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold929 _7158_/Q hold929/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6190_ _6716_/Q _5997_/Z _6014_/Z _6809_/Q _6193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5141_ _5293_/A1 _4614_/Z _5289_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _4500_/Z _4906_/Z _5078_/A2 _5072_/A4 _5072_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_96_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4023_ _4023_/A1 _4022_/Z _4024_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5974_ _5974_/A1 _5974_/A2 _5974_/A3 _5974_/A4 _5983_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4925_ _5083_/B _5080_/C _5370_/B _4926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_100_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4856_ _4614_/Z _4817_/Z _4858_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet563_209 net613_256/I _7016_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3807_ _3509_/Z _3519_/Z _3923_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4787_ _5220_/B2 _5092_/A1 _4787_/A3 _4491_/B _4787_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6526_ _6526_/A1 _6526_/A2 _6526_/A3 _6526_/A4 _6526_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_180_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3738_ input67/Z _4227_/S _4244_/S input38/Z _5701_/A1 _7055_/Q _3739_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _7188_/Q _6282_/Z _6293_/Z _7156_/Q _6296_/Z _7164_/Q _6465_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3669_ hold71/I _5584_/A1 _3959_/B1 _6671_/Q _3673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5408_ _4761_/I _5245_/Z _5481_/B1 _4908_/Z _5408_/C _5409_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_162_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6388_ _6943_/Q _6245_/Z _6288_/Z _7121_/Q _6390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_14__1359_ _4073__7/I _4073__11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5339_ _5261_/I _5338_/Z _5262_/Z _5339_/A4 _5340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7009_ _7009_/D _7260_/RN _7009_/CLK _7009_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7279_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_188_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ hold440/Z hold12/Z _5691_/S _5690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ _4694_/Z _4703_/Z _5308_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4641_ _5281_/C _4467_/B _4472_/B _4501_/B _4641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_128_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4572_ _4572_/I _5472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_129_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7291_ _7291_/D _6645_/Z _7304_/CLK _7291_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_157_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3523_ hold320/Z _3617_/A1 _3501_/Z _3489_/I _3523_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6311_ _6973_/Q _6484_/A2 _6311_/A3 _6533_/A2 _6327_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold726 _4166_/Z _6711_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold704 _5518_/Z _6893_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold715 _6720_/Q hold715/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold737 _6846_/Q hold737/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3454_ hold1/Z hold11/Z _3460_/S _7290_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold748 _4331_/Z _6838_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6242_ _7110_/Q _6240_/Z _6241_/Z _7044_/Q _6260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold759 _6850_/Q hold759/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_157_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6173_ _6173_/I _6174_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3385_ _7231_/Q _6210_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
XFILLER_112_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _5414_/A2 _4784_/Z _5124_/B _5317_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_85_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5055_ _5130_/B2 _5420_/A2 _4367_/Z _5291_/C _5055_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_84_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4006_ _5900_/A1 _5911_/A1 _7225_/Q _7224_/Q _4006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_84_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5957_ _3990_/I _6745_/Q _5957_/S _6558_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_80_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_1__1359_ net763_436/I net763_445/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4908_ _5324_/A1 _4759_/Z _4494_/Z _4496_/Z _4908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_80_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5888_ hold65/Z hold629/Z _5892_/S _5888_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4839_ _4887_/A1 _5414_/A2 _5399_/A2 _5287_/B _5369_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6509_ _6692_/Q _6285_/Z _6299_/Z _6857_/Q _6511_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold31 hold31/I hold31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold20 hold20/I hold20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold64 hold64/I hold64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold42 hold42/I hold42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_76_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold53 hold53/I hold53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_91_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold86 hold86/I hold86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold97 hold97/I hold97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold75 hold75/I hold75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_56_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_6 _4336_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60__1359_ net513_170/I net763_435/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6860_ _6860_/D _7279_/RN _7278_/CLK _6860_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ hold2/Z hold308/Z _5811_/S _5811_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _6791_/D _7265_/CLK _6791_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_290 _4073__5/I _6935_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5742_ hold291/Z hold984/Z _5748_/S _5742_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ hold209/Z hold2/Z _5673_/S _5673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4441_/B _5281_/C _4436_/B _4501_/B _4624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_117_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4555_ _5129_/A3 _4835_/A2 _4555_/B _4555_/C _4556_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold501 _5890_/Z _7219_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold523 _7185_/Q hold523/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold534 _5807_/Z _7145_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3506_ _3485_/Z _3505_/Z _3909_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold545 _4133_/Z _6686_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold512 _4135_/Z _6688_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4486_ _4486_/A1 _4483_/B _4486_/B1 _4484_/Z _5312_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7274_ _7274_/D _7279_/RN _7279_/CLK _7274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold556 _6974_/Q hold556/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold578 _6684_/Q hold578/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold567 _5650_/Z _7006_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3437_ _3442_/B _6663_/Q _6664_/Q _6665_/Q _3438_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_89_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold589 _5686_/Z _7038_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6225_ _6800_/Q _5958_/Z _5967_/Z _6721_/Q _6227_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_170_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3368_ hold75/I _3368_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6156_ _7156_/Q _5960_/Z _5965_/Z _6704_/Q _6006_/Z _7172_/Q _6158_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_98_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _5107_/I _5309_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3299_ _6665_/Q _3465_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6087_ _6555_/C _7243_/Q _6087_/B _6088_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _5038_/A1 _4606_/Z _5003_/Z _5038_/B _5205_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_2728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6989_ _6989_/D _7008_/RN _6989_/CLK _6989_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_167_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput110 wb_adr_i[23] _4026_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_150_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput143 wb_dat_i[23] _6600_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput132 wb_dat_i[13] _6594_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput154 wb_dat_i[4] _3397_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput121 wb_adr_i[4] _4460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_0_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput165 wb_stb_i _4032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4340_ hold291/Z hold763/Z _4340_/S _4340_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4271_ _5520_/C _3527_/Z _5513_/A3 _5839_/A3 _4273_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_98_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6010_ _6010_/A1 _6010_/A2 _6924_/Q _6201_/A3 _6011_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_100_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6912_ _6912_/D _7218_/RN _6912_/CLK _7327_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6843_ _6843_/D _7170_/RN _6843_/CLK _6843_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3986_ _7305_/Q _3415_/Z _6658_/Q _3987_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6774_ _6774_/D _7218_/RN _6774_/CLK _6774_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5725_ hold20/Z hold192/Z _5727_/S _5725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5656_ _5656_/A1 hold32/Z hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4607_ _4607_/A1 _4570_/Z _4606_/Z _4501_/B _4607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_11_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold320 _3493_/Z hold320/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5587_ hold196/Z hold91/Z _5592_/S _5587_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7326_ _7326_/I _7326_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4538_ _5288_/B _4467_/B _4472_/B _4539_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_105_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold331 _7031_/Q hold331/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold353 _5834_/Z _7169_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold342 _7211_/Q hold342/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold386 _7062_/Q hold386/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ _7257_/D _7258_/RN _7258_/CLK _7257_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ _4459_/Z _4469_/A2 _4690_/B _4690_/C _4786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_77_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold364 _5527_/Z _6900_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold375 _6929_/Q hold375/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold397 _5630_/Z _6988_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6208_ _7249_/Q _6208_/I1 _6558_/S _7249_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7188_ _7188_/D _7237_/RN _7188_/CLK _7188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_3204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6139_ _7058_/Q _6210_/A2 _6210_/B _6210_/C _6155_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_485 net813_488/I _6680_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_463 net813_463/I _6702_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_452 net813_453/I _6713_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_474 net813_475/I _6691_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_496 net413_88/I _6669_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ _3537_/Z _3680_/Z _4143_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3771_ _7070_/Q _3943_/A2 _3945_/B1 _7088_/Q _3773_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5510_ _3521_/Z _3527_/Z _5520_/C _5512_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_145_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6490_ _7085_/Q _6290_/Z _6302_/Z _7093_/Q _6490_/C _6492_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_173_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5441_ _5437_/Z _5440_/Z _5441_/B _5463_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_145_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5372_ _5372_/A1 _5139_/Z _5055_/Z _5372_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7111_ _7111_/D _7237_/RN _7111_/CLK _7111_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4323_ _3509_/Z _5821_/A3 _5513_/A3 _5520_/C _4325_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7042_ _7042_/D _7256_/RN _7042_/CLK _7042_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4254_ hold227/Z hold482/Z _4261_/S _4254_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4185_ _5520_/C _3537_/Z _5513_/A3 _5839_/A3 _4187_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_94_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6826_ _6826_/D _7279_/RN _7279_/CLK _6826_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_149_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6757_ _6757_/D _7258_/RN _6757_/CLK _6757_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3969_ _3427_/Z _6663_/Q _6664_/Q _3970_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5708_ hold670/Z hold12/Z _5709_/S _5708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6688_ _6688_/D _7008_/RN _6688_/CLK _6688_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_12_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_3_0__1359_ clkbuf_4_10_0__1359_/Z clkbuf_opt_3_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5639_ _6996_/Q hold227/Z _5646_/S _5639_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold161 _6942_/Q hold161/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7309_ _7309_/I _7309_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold150 _4250_/Z _6766_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold172 _7074_/Q hold172/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold183 _4249_/Z _6765_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold194 _7080_/Q hold194/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _7020_/Q _6211_/A2 _6002_/A2 _6956_/Q _6211_/B1 _6988_/Q _5992_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4941_ _5464_/A1 _5410_/A1 _5062_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet413_80 net413_80/I _7145_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4872_ _4872_/A1 _5215_/C _5117_/A2 _5215_/B _4874_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4073__50 _4073__50/I _7175_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_91 net413_91/I _7134_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3823_ _6981_/Q _3901_/A2 _3889_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_21_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ _6611_/A1 hold32/Z _6613_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ _6542_/A1 _6542_/A2 _6542_/A3 _6542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_3754_ _7137_/Q _3951_/A2 _3954_/B1 input23/Z _3754_/C _3757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6473_ _6466_/Z _6472_/Z _6473_/B1 _6286_/Z _6555_/C _6474_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3685_ hold86/I _3957_/A2 _3941_/B1 _7171_/Q _3686_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xoutput200 _4050_/Z mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_146_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5424_ _5489_/A1 _5423_/Z _5427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput233 _7330_/Z mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput211 _7313_/Z mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput222 _7320_/Z mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput244 _7312_/Z mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5355_ _5437_/A2 _5350_/Z _5352_/Z _5354_/Z _5355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput255 _4077_/ZN pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput266 _6882_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput277 _6681_/Q pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5286_ _5286_/A1 _5374_/A3 _5374_/A2 _5292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_102_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput299 _4085_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput288 _6890_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4306_ _6565_/I0 _6812_/Q _4312_/S _6812_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4237_ _4236_/Z hold787/Z _4245_/S _4237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7025_ hold81/Z _7260_/RN _7025_/CLK hold80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_74_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7260_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4168_ _4103_/I hold865/Z _4169_/S _4168_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4099_ hold23/Z _6608_/I0 hold54/I hold24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_56_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_117__1359_ net613_261/I net413_83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_169_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _6809_/D _7008_/RN _6809_/CLK _6809_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold919 _7102_/Q hold919/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold908 _5730_/Z _7077_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3470_ _6660_/Q _6733_/Q _6661_/Q _3471_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_155_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5140_ _5293_/A1 _4549_/Z _5147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _4376_/Z _5071_/A2 _5257_/A1 _4699_/Z _5408_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4022_ _7282_/Q _3409_/Z _4022_/A3 _6730_/Q _4022_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5973_ _7012_/Q _5971_/Z _5972_/Z _6940_/Q _5974_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4924_ _5259_/A1 _5337_/A2 _5258_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_166_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4855_ _5287_/C _4844_/Z _4855_/B _4855_/C _4858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_159_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ _4786_/A1 _4786_/A2 _4786_/A3 _5137_/B1 _4787_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3806_ _3509_/Z _3535_/Z _3924_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_158_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3737_ _6927_/Q _3935_/A2 _3916_/A2 _7153_/Q _3912_/B1 _6886_/Q _3739_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6525_ _6694_/Q _6248_/Z _6300_/Z _6720_/Q _6526_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ hold52/I _6253_/Z _6272_/Z _7204_/Q _6456_/C _6465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_109_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3668_ hold78/I _3923_/C1 _3956_/A2 hold76/I _3668_/C _3674_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_115_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _5406_/Z _5454_/A2 _5419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3599_ _7011_/Q _3934_/A2 _5683_/A1 _7043_/Q _7051_/Q _3952_/A2 _3601_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6387_ _7047_/Q _6241_/Z _6251_/Z _6983_/Q _6268_/Z _6951_/Q _6390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5338_ _5332_/Z _5334_/Z _5447_/A1 _5338_/A4 _5338_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_161_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5269_ _4454_/Z _5269_/A2 _4651_/Z _4675_/Z _5464_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7008_ _7008_/D _7008_/RN _7008_/CLK _7008_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_100__1359_ clkbuf_4_5_0__1359_/Z net413_78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4640_ _5315_/A1 _5315_/A2 _5468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_83__1359_ net413_62/I net413_73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ _4549_/Z _4570_/Z _4572_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6310_ _6308_/Z _6310_/A2 _6310_/A3 _6558_/S _6310_/B2 _7251_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_171_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7290_ _7290_/D _6644_/Z _4072_/B2 hold1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold727 _6933_/Q hold727/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3522_ _3509_/Z _3521_/Z _3910_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold716 _4180_/Z _6720_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold705 _6724_/Q hold705/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3453_ _4041_/B1 _3442_/B _6732_/Q _3460_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_170_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6241_ _7235_/Q _7234_/Q _6300_/A2 _6533_/A2 _6241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold749 _7218_/Q hold749/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold738 _6840_/Q hold738/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6172_ _6979_/Q _5964_/Z _6014_/Z _6963_/Q _5999_/Z _7035_/Q _6173_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5123_ _5456_/A1 _5220_/B2 _5312_/A2 _5137_/B1 _5123_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_69_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3384_ _6786_/Q _6555_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_111_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _5370_/B _5258_/A2 _4977_/Z _5323_/B _5324_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_57_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4005_ _4005_/A1 _4003_/Z _5945_/A1 _6901_/Q _6743_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xnet663_350 net413_66/I _6867_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5956_ _5957_/S _6745_/Q _6310_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_80_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _4759_/Z _4906_/Z _5257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_179_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5887_ hold91/Z hold240/Z _5892_/S _5887_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4838_ _4555_/C _4876_/A2 _4838_/B1 _5291_/C _4841_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_154_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4769_ _4703_/Z _4764_/Z _5117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_5_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _6724_/Q _6240_/Z _6247_/Z _6728_/Q _6511_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_136_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _6434_/Z _6439_/A2 _6439_/A3 _6439_/A4 _6439_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_150_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold32 hold55/Z hold32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_88_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold10 hold10/I hold10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold21 hold21/I hold21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold54 hold54/I hold54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_152_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold65 hold65/I hold65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold43 hold43/I hold43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold98 hold98/I hold98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold87 hold87/I hold87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold76 hold76/I hold76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_17_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_7 _5495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5810_ hold12/Z hold488/Z _5811_/S _5810_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6790_ _6790_/D _7008_/RN _6790_/CLK _6790_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_291 net413_81/I _6934_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5741_ hold227/Z hold639/Z _5748_/S _5741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet613_280 net713_394/I _6945_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_188_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5672_ hold265/Z hold12/Z _5673_/S _5672_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4623_ _4887_/A1 _4868_/A1 _5376_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_135_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4554_ _3401_/I _3402_/I _4456_/B _5051_/S _4554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold502 _7195_/Q hold502/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7273_ _7273_/D _7279_/RN _7279_/CLK _7273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold524 _5852_/Z _7185_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold535 _7201_/Q hold535/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3505_ _3617_/A1 _3501_/Z _3489_/I _3492_/Z _3505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold513 _7030_/Q hold513/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4485_ _4381_/Z _4485_/A2 _4486_/B1 _4424_/B _4687_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold546 _7104_/Q hold546/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold557 _5614_/Z _6974_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold579 _4131_/Z _6684_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6224_ _6719_/Q _5960_/Z _5965_/Z _7077_/Q _6006_/Z _6711_/Q _6227_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold568 _6998_/Q hold568/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3436_ _6665_/Q _6664_/Q _6663_/Q _3898_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_131_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3367_ _7023_/Q _3367_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6155_ _6155_/A1 _6155_/A2 _6155_/A3 _6155_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_58_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6086_ _6073_/Z _6085_/Z _6392_/B1 _6168_/C _6555_/C _6087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5106_ _5106_/A1 _5106_/A2 _5107_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3298_ hold22/Z hold23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5037_ _5039_/A4 _5036_/Z _5357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6988_ _6988_/D _7258_/RN _6988_/CLK _6988_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_167_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ _6745_/Q _5939_/A2 _5913_/I _6282_/A2 _7233_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_40_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput111 wb_adr_i[24] _4029_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput100 wb_adr_i[14] _4386_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput144 wb_dat_i[24] _6579_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput133 wb_dat_i[14] _6597_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput122 wb_adr_i[5] _4436_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_89_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput166 wb_we_i _6575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xinput155 wb_dat_i[5] _3398_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ hold256/Z hold2/Z _4270_/S _4270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ _6911_/D _7218_/RN _6911_/CLK _7326_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6842_ _6842_/D _7170_/RN _6842_/CLK _6842_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_90_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3985_ _3984_/Z _6659_/Q _3988_/S _6659_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6773_ _6773_/D _7218_/RN _6773_/CLK _6773_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ hold48/Z hold414/Z _5727_/S _5724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ hold327/Z hold2/Z _5655_/S _5655_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4606_ _4648_/A2 _4467_/B _4648_/A1 _4606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_175_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7325_ _7325_/I _7325_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold310 _7085_/Q hold310/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5586_ hold697/Z hold291/Z _5592_/S _5586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4537_ _4441_/B _4501_/B _5399_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_144_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold332 _6979_/Q hold332/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold343 _5881_/Z _7211_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_11_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold321 _3904_/Z hold321/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold387 _5713_/Z _7062_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7256_ _7256_/D _7256_/RN _7258_/CLK _7256_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4468_ _4467_/B _4736_/A1 _4468_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xhold365 _7041_/Q hold365/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold354 _7134_/Q hold354/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold376 _5563_/Z _6929_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3419_ _4041_/B1 _6730_/Q _7304_/Q _3421_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_120_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7187_ _7187_/D _7256_/RN _7187_/CLK _7187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold398 _6698_/Q hold398/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6207_ _6207_/I _6208_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4399_ _4402_/B _4483_/B _4026_/B _4026_/C _4399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_98_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6138_ _7108_/Q _5967_/Z _6147_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_58_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1010 _7294_/Q _3440_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_97_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _7063_/Q _5985_/Z _6084_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_3249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_464 net813_464/I _6701_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_453 net813_453/I _6712_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_475 net813_475/I _6690_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_497 net413_88/I _6668_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_486 net813_489/I _6679_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3770_ _7160_/Q _3941_/A2 _5503_/A2 _3904_/A2 _3770_/C _3773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_73_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _5440_/A1 _5357_/Z _5388_/Z _5440_/A4 _5440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_157_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _5371_/A1 _5287_/B _5470_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_126_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ _7110_/D _7218_/RN _7110_/CLK _7110_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4322_ hold291/Z hold775/Z _4322_/S _4322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4253_ _3485_/Z _3540_/Z _6652_/A2 hold24/Z _4261_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7041_ _7041_/D _7258_/RN _7041_/CLK _7041_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_141_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4184_ hold899/Z hold291/Z _4184_/S _4184_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7258_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6825_ _6825_/D _7008_/RN _6825_/CLK _6825_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3968_ _6665_/Q _3967_/Z _6665_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6756_ _6756_/D _7258_/RN _6756_/CLK _6756_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ hold378/Z hold20/Z _5709_/S _5707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _6687_/D _7008_/RN _6687_/CLK _6687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3899_ _3898_/Z _3899_/I1 _3899_/S _6869_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5638_ _5638_/A1 hold32/Z _5646_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_152_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5569_ hold91/Z hold506/Z _5574_/S _5569_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold151 _6952_/Q hold151/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7308_ _7308_/I _7308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold140 _5835_/Z _7170_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold162 _5578_/Z _6942_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold184 _6703_/Q hold184/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold173 _5726_/Z _7074_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold195 _5734_/Z _7080_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7239_ _7239_/D _7256_/RN _4067_/I1 _7239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4940_ _4421_/Z _5410_/A1 _4942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet413_70 net413_79/I _7155_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_92 net413_95/I _7133_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__40 net413_96/I _7185_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4871_ _4641_/Z _4817_/Z _5117_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet413_81 net413_81/I _7144_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__51 _4073__51/I _7174_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _6610_/A1 _6610_/A2 _6610_/A3 _6610_/A4 _7279_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3822_ _6788_/Q _4274_/A1 _3947_/B1 _6717_/Q _3873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ _6725_/Q _6240_/Z _6248_/Z _6695_/Q _6542_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3753_ _3753_/I _3754_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6472_ _6554_/A1 _6472_/A2 _6472_/A3 _6472_/A4 _6472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3684_ hold82/I _3916_/A2 _5528_/S _3683_/Z _3686_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xoutput201 _4049_/Z mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _5423_/A1 _5423_/A2 _5377_/Z _5422_/Z _5423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_134_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput234 _4053_/Z mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5354_ _5354_/A1 _5354_/A2 _5354_/A3 _5354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput212 _7314_/Z mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput223 _7321_/Z mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput245 _4058_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput256 _4077_/I pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4305_ _6564_/I0 _6811_/Q _4312_/S _6811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput267 _6876_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5285_ _4598_/Z _4683_/Z _5285_/B _5374_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_114_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput278 _6666_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput289 _6684_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4236_ hold458/Z hold65/Z _4244_/S _4236_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7024_ hold94/Z _7260_/RN _7024_/CLK hold93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4167_ _3535_/Z _3537_/Z _5520_/C _4169_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_4098_ _7235_/RN _6657_/A2 _4098_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_167_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6808_ _6808_/D _6818_/CLK _6808_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6739_ _6739_/D _7218_/RN _6739_/CLK _7319_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold909 _7297_/Q hold909/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5070_ _5070_/A1 _5070_/A2 _5334_/A1 _5070_/A4 _5074_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4021_ _4021_/I _6746_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_123__1359_ net613_261/I _4073__39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ _7228_/Q _6210_/C _6015_/A3 _6210_/A2 _5972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4923_ _4423_/Z _4923_/A2 _4923_/B _5080_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_52_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4854_ _4422_/Z _5414_/A2 _4614_/Z _4483_/B _4855_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4785_ _4808_/A2 _5220_/B2 _5092_/A1 _4491_/B _5124_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3805_ _3519_/Z _3552_/Z _3912_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3736_ _7217_/Q _3912_/A2 _4194_/A1 input55/Z _3948_/C1 input64/Z _3739_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6524_ _6690_/Q _6257_/Z _6275_/Z _6849_/Q _6526_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _7084_/Q _6290_/Z _6299_/Z _7058_/Q _6466_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3667_ _3667_/I _3668_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5406_ _5406_/A1 _5404_/Z _5406_/A3 _4799_/Z _5406_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3598_ _7165_/Q _3941_/A2 _3947_/A2 _7101_/Q _7059_/Q _5701_/A1 _3601_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6386_ _7023_/Q _6235_/Z _6243_/Z _7007_/Q _6265_/Z _6999_/Q _6391_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_47_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5337_ _5337_/A1 _5337_/A2 _5337_/B _5337_/C _5449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_87_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ _5368_/A1 _4650_/Z _5172_/C _5268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_130_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7007_ _7007_/D _7258_/RN _7007_/CLK _7007_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4219_ hold67/Z hold65/Z _4227_/S _4219_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5199_ _5191_/Z _5196_/Z _5390_/A2 _5476_/A2 _5199_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_69_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4570_ _5270_/A1 _4454_/Z _5364_/B _4570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3521_ _3489_/I _3492_/Z _3497_/I _3501_/Z _3521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_183_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold717 _7132_/Q hold717/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold728 _5568_/Z _6933_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold706 _4186_/Z _6724_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3452_ _3451_/Z _7291_/Q _3452_/S _7291_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6240_ _7236_/Q _6533_/A4 _6302_/A4 _6533_/A3 _6240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold739 _6825_/Q hold739/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6171_ _7149_/Q _5987_/Z _6002_/Z _7093_/Q _6003_/Z _7165_/Q _6181_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3383_ _7077_/Q _3866_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _5456_/A1 _5231_/A2 _5122_/B _5213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5053_ _5325_/B _5078_/A2 _5060_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ _4005_/A1 _4003_/Z _5894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_351 net413_64/I _6866_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_340 net413_75/I _6885_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5955_ _5954_/Z _7240_/Q _5955_/S _7240_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _4494_/Z _5259_/A1 _4496_/Z _4407_/Z _4906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_179_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5886_ hold291/Z hold937/Z _5892_/S _5886_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4837_ _5278_/C _4784_/Z _4838_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4768_ _4510_/Z _4764_/Z _4770_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_5_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4699_ _5420_/A3 _4835_/A2 _4456_/B _3402_/I _4699_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6507_ _6726_/Q _6253_/Z _6296_/Z _6714_/Q _6511_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3719_ _3719_/A1 _3719_/A2 _3719_/A3 _3719_/A4 _3719_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ hold78/I _6290_/Z _6302_/Z _7091_/Q _6438_/C _6439_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_162_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6369_ _6967_/Q _6262_/Z _6391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold22 hold22/I hold22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold11 hold11/I hold11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold55 hold55/I hold55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_102_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold33 hold33/I hold33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold44 hold44/I hold44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_91_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold99 hold99/I hold99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold77 hold77/I hold77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold88 hold88/I hold88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold66 hold66/I hold66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_57_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_8 _5500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5740_ _3515_/Z _3537_/Z hold24/Z _5748_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_50_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_270 net613_284/I _6955_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_281 net813_492/I _6944_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_292 net413_91/I _6933_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5671_ hold80/Z hold20/Z _5673_/S hold81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4622_ _4622_/A1 _5029_/B _5353_/B _4627_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_4553_ _4836_/A4 _4454_/Z _5370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_129_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4484_ _4381_/Z _4385_/Z _4387_/Z _4424_/B _4484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7272_ _7272_/D _7279_/RN _7279_/CLK _7272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold525 _7113_/Q hold525/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold536 _5870_/Z _7201_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold514 _7203_/Q hold514/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold503 _5863_/Z _7195_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3504_ _5857_/A2 _5857_/A3 _5647_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3435_ _3435_/A1 _3435_/A2 _7298_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold558 _7177_/Q hold558/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold547 _5761_/Z _7104_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold569 _5641_/Z _6998_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6223_ _6691_/Q _5985_/Z _6014_/Z _6810_/Q _6228_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_143_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3366_ _7031_/Q _3366_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6154_ _7018_/Q _5971_/Z _6005_/Z _7042_/Q _7050_/Q _6019_/Z _6155_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3297_ _7291_/Q _3451_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6085_ _6078_/Z _6085_/A2 _6085_/A3 _6084_/Z _6085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5105_ _5105_/A1 _5104_/Z _5310_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_57_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5036_ _5356_/C _5389_/C _5328_/A1 _5356_/B _5036_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6987_ _6987_/D _7258_/RN _6987_/CLK _6987_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _6484_/A2 _6302_/A3 _5939_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5869_ hold91/Z hold598/Z _5874_/S _5869_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 wb_adr_i[15] _4386_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput145 wb_dat_i[25] _6582_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput134 wb_dat_i[15] _6600_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput123 wb_adr_i[6] _4472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput112 wb_adr_i[25] _3334_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput156 wb_dat_i[6] _3399_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_57_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7278_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_6_0__1359_ clkbuf_0__1359_/Z net613_261/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_43_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6910_ _6910_/D _7218_/RN _6910_/CLK _7325_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _6841_/D _7170_/RN _6841_/CLK _6841_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_51_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ _3983_/Z _6658_/Q _6733_/Q _3984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6772_ _6772_/D _7256_/RN _6772_/CLK _6772_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ hold65/Z hold254/Z _5727_/S _5723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5654_ hold267/Z hold12/Z _5655_/S _5654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4605_ _4638_/A2 _4648_/B _5356_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_163_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold311 _5739_/Z _7085_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7324_ _7324_/I _7324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5585_ hold360/Z hold227/Z _5592_/S _5585_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold300 _6677_/Q hold300/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4536_ _5414_/A2 _4501_/B _4472_/B _4524_/Z _4536_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold333 _5619_/Z _6979_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold344 _6999_/Q hold344/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_11_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold322 hold322/I _6894_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7255_ _7255_/D _7256_/RN _7258_/CLK _7255_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4467_ _4467_/A1 _4555_/B _4467_/B _4690_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_89_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold366 _5689_/Z _7041_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold355 _5795_/Z _7134_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold377 _7017_/Q hold377/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4398_ _5002_/A3 _5002_/A4 _5165_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3418_ _3417_/Z _7305_/Q _3988_/S _7305_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold388 _7181_/Q hold388/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7186_ _7186_/D _7256_/RN _7186_/CLK _7186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold399 _4150_/Z _6698_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6206_ _6555_/C _7248_/Q _6206_/B _6207_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3349_ _7161_/Q _3349_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6137_ _7246_/Q _6136_/Z _6558_/S _7246_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1000 _6869_/Q _3899_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold1011 _7282_/Q _4041_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_100_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ _7145_/Q _7231_/Q _6210_/B _6068_/A4 _6076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_85_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _5191_/A3 _5019_/A2 _5390_/A1 _5019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_2527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_465 _4073__15/I _6700_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_476 net813_483/I _6689_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_454 net813_455/I _6711_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_487 net813_487/I _6678_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_498 net813_499/I _6667_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5370_ _5370_/A1 _5172_/B _5370_/B _5370_/C _5371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_113_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4321_ hold227/Z hold574/Z _4322_/S _4321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4252_ hold20/Z hold600/Z _4252_/S _4252_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7040_ _7040_/D _7218_/RN _7040_/CLK _7040_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4183_ hold863/Z _4103_/I _4184_/S _4183_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6824_ _6824_/D _7008_/RN _6824_/CLK _6824_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_177_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3967_ _3427_/Z _6663_/Q _6664_/Q _3967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6755_ _6755_/D _7258_/RN _6755_/CLK _6755_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5706_ hold490/Z hold48/Z _5709_/S _5706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6686_ _6686_/D _7008_/RN _6686_/CLK _6686_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3898_ _6565_/I0 _6868_/Q _3898_/S _3898_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ hold2/Z hold302/Z _5637_/S _5637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5568_ hold291/Z hold727/Z _5574_/S _5568_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4519_ _5170_/A2 _5269_/A2 _5328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold130 _5883_/Z _7213_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold141 _7157_/Q hold141/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7307_ _7307_/I _7307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold152 _5589_/Z _6952_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold185 _4155_/Z _6703_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold174 _7204_/Q hold174/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7238_ _7238_/D _7238_/RN _7260_/CLK _7238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold163 _6673_/Q hold163/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5499_ hold470/Z hold291/Z _5502_/S _5499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold196 _6950_/Q hold196/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_101_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7169_ _7169_/D _7218_/RN _7169_/CLK _7169_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7__1359_ clkbuf_4_2_0__1359_/Z net413_63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_60 net413_60/I _7165_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_93 net413_93/I _7132_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4870_ _5293_/B _4844_/Z _5215_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4073__30 _4073__6/I _7195_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__41 _4073__41/I _7184_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_71 _4073__3/I _7154_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_82 net413_83/I _7143_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3821_ _3537_/Z _3653_/Z _3947_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6540_ _6867_/Q _6272_/Z _6293_/Z _6719_/Q _6540_/C _6547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_60_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_66__1359_ net513_170/I net613_294/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_146__1359_ net763_436/I net813_491/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3752_ hold69/I _3923_/A2 _3959_/B1 _6669_/Q _5656_/A1 hold75/I _3753_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_118_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ hold45/I _6245_/Z _6273_/Z _6978_/Q _7124_/Q _6288_/Z _6472_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3683_ _7250_/Q hold39/I _6900_/Q _3683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5422_ _5034_/B _4866_/Z _5422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xoutput235 _4054_/Z mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ _5353_/A1 _5387_/A2 _5353_/B _5354_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput213 _4068_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput224 _7322_/Z mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput202 _3376_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput246 _4057_/Z mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4304_ _6829_/Q _7279_/RN _4312_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xoutput257 _6886_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput268 _6883_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5284_ _5284_/A1 _5369_/B _5284_/A3 _5277_/I _5286_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_99_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput279 _6667_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4235_ _4234_/Z hold807/Z _4245_/S _4235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7023_ _7023_/D _7260_/RN _7023_/CLK _7023_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_96_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4166_ hold291/Z hold725/Z _4166_/S _4166_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4097_ _4097_/A1 _4415_/B _6828_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _6807_/D _6818_/CLK _6807_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4999_ _4999_/A1 _4999_/A2 _4998_/Z _5341_/B _5000_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_6738_ _6738_/D _7256_/RN _6738_/CLK _7318_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6669_ _6669_/D _7238_/RN _6669_/CLK _6669_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_165_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4020_ _4014_/Z _4020_/A2 _6746_/Q _4003_/Z _4021_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_84_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _7228_/Q _7227_/Q _6211_/B1 _6210_/A2 _5971_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_64_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4922_ _4373_/Z _4385_/Z _4922_/A3 _4922_/A4 _4923_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_45_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _4853_/A1 _5287_/B _4784_/Z _4501_/B _4853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4784_ _5420_/A3 _3402_/I _4456_/B _5051_/S _4784_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3804_ _6842_/Q _3930_/B1 _3884_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_119_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3735_ _7113_/Q _3917_/A2 _5674_/A1 _7031_/Q _3735_/C _3760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6523_ _6866_/Q _6272_/Z _6290_/Z _6708_/Q _6526_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_147_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6454_ _7100_/Q _6250_/Z _6302_/Z _7092_/Q _6292_/Z _7148_/Q _6466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5405_ _5454_/A1 _4791_/Z _5126_/I _5406_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_106_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3666_ _6929_/Q _3935_/A2 _5656_/A1 _7017_/Q _3667_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _6385_/A1 _6385_/A2 _6385_/A3 _6384_/Z _6385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3597_ _6681_/Q _3546_/Z _3945_/C2 _6689_/Q _3913_/A2 input19/Z _3601_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5336_ _5412_/A1 _5412_/A3 _5338_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_142_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _4898_/C _5428_/A4 _4893_/Z _5267_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_125_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7006_ _7006_/D _7260_/RN _7006_/CLK _7006_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4218_ _4217_/Z hold582/Z _4228_/S _4218_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5198_ _5309_/B2 _5205_/A1 _5351_/C _5205_/B1 _5198_/C _5476_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_83_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4149_ _3507_/Z _3537_/Z _5520_/C _4157_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_28_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3520_ _3485_/Z _3519_/Z _4225_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_7_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold718 _5792_/Z _7132_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_128_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold707 _6690_/Q hold707/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3451_ _3451_/I0 input58/Z _6730_/Q _3451_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold729 _6788_/Q hold729/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6170_ _6971_/Q _5979_/Z _5981_/Z _6939_/Q _5996_/Z _7085_/Q _6181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3382_ _6785_/Q _6528_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_111_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5121_ _5121_/A1 _4876_/C _5457_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _4936_/I _5051_/Z _5064_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_78_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4003_ _5954_/A3 _7225_/Q _7226_/Q _7223_/Q _4003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet663_341 net813_487/I _6884_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_330 net663_330/I _6895_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5954_ _7223_/Q _5954_/A2 _5954_/A3 _6746_/Q _5954_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_81_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _4467_/B _4495_/Z _5263_/A2 _5324_/A1 _4905_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5885_ _4103_/I hold967/Z _5892_/S _5885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _5420_/A3 _4549_/Z _3402_/I _4836_/A4 _4836_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_166_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _4716_/Z _4764_/Z _5118_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6506_ _6820_/Q _6262_/Z _6269_/Z _6847_/Q _6512_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4698_ _5097_/A1 _4704_/A2 _4698_/B _5094_/B _4714_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3718_ input16/Z _3913_/A2 _3945_/B1 _7090_/Q _3719_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3649_ _3648_/Z hold999/Z _3899_/S _6874_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6437_ _6437_/I _6438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6368_ _7145_/Q _6292_/Z _6383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_103_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ _5392_/B _4801_/Z _5319_/A3 _5319_/A4 _5319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_102_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold23 hold23/I hold23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6299_ _7236_/Q _6533_/A3 _6452_/A4 _6302_/A4 _6299_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold12 hold12/I hold12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_49_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold56 hold56/I hold56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold34 hold34/I hold34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold45 hold45/I hold45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold67 hold67/I hold67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold78 hold78/I hold78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold89 hold89/I hold89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_90_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_9 _5502_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7269_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_260 _4073__27/I _6965_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_282 net713_394/I _6943_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_271 net613_275/I _6954_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5670_ hold93/Z hold48/Z _5673_/S hold94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet613_293 net413_83/I _6932_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _4367_/Z _4555_/B _5291_/C _5353_/A1 _5353_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_148_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _4549_/Z _4551_/Z _5011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7271_ _7271_/D _7279_/RN _7279_/CLK _7271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold526 _5771_/Z _7113_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4483_ _4489_/A1 _4692_/B _4483_/B _4687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold515 _5872_/Z _7203_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3503_ _3497_/I hold673/Z _5857_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold504 _7007_/Q hold504/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3434_ _3442_/B _3409_/Z _3434_/B _3435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_132_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold559 _5843_/Z _7177_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold548 _6903_/Q hold548/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold537 _6700_/Q hold537/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6222_ _6823_/Q _5964_/Z _5999_/Z _6848_/Q _6729_/Q _6000_/Z _6228_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_143_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3365_ _7039_/Q _3365_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6153_ hold45/I _5972_/Z _6021_/Z _7002_/Q _6155_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3296_ _7294_/Q _4084_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5104_ _5104_/A1 _5139_/A3 _5094_/B _5104_/A4 _5104_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6084_ _6084_/A1 _6084_/A2 _6084_/A3 _6084_/A4 _6084_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ _5035_/A1 _5032_/Z _5204_/C _5035_/A4 _5035_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_73_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6986_ _6986_/D _7258_/RN _6986_/CLK _6986_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_25_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5937_ _6279_/A3 _7233_/Q _6302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_53_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5868_ hold291/Z hold986/Z _5874_/S _5868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ _4422_/Z _4624_/Z _4673_/Z _4483_/B _4819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5799_ hold48/Z hold99/Z _5802_/S _5799_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput102 wb_adr_i[16] _4391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput135 wb_dat_i[16] _6579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput113 wb_adr_i[26] _4031_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput124 wb_adr_i[7] _4501_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_163_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput146 wb_dat_i[26] _6585_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput157 wb_dat_i[7] _3400_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _6840_/D _7008_/RN _6840_/CLK _6840_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6771_ _6771_/D _7256_/RN _6771_/CLK _6771_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3983_ _6659_/Q _3972_/Z _3983_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5722_ hold91/Z hold402/Z _5727_/S _5722_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5653_ hold371/Z hold20/Z _5655_/S _5653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4604_ _4501_/B _4604_/A2 _4604_/A3 _4604_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5584_ _5584_/A1 hold32/Z _5592_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4535_ _5414_/A2 _4534_/Z _5323_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7323_ _7323_/I _7323_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold301 _4123_/Z _6677_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold334 _7043_/Q hold334/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold312 _7125_/Q hold312/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold323 _7161_/Q hold323/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7254_ _7254_/D _7256_/RN _7258_/CLK _7254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold356 _6916_/Q hold356/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4466_ _4454_/Z _4367_/Z _4363_/Z _4690_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_116_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold345 _5642_/Z _6999_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold367 _7187_/Q hold367/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold378 _7057_/Q hold378/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4397_ _5002_/A3 _5002_/A4 _4397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3417_ _3416_/Z _7304_/Q _6733_/Q _3417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7185_ _7185_/D _7237_/RN _7185_/CLK _7185_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold389 _5847_/Z _7181_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6205_ _6193_/Z _6204_/Z _6528_/B1 _6168_/C _6555_/C _6206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3348_ _7169_/Q _3348_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6136_ _6136_/I0 _7245_/Q _6555_/C _6136_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1012 _7282_/Q _3425_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1001 _6870_/Q _3799_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XTAP_3229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6067_ _6067_/A1 _5991_/Z _6072_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5018_ _5389_/B _5439_/B2 _5018_/B _5390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet813_466 net813_466/I _6699_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_455 net813_455/I _6710_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_499 net813_499/I _6666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_488 net813_488/I _6677_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_477 net813_481/I _6688_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6969_ hold44/Z _7260_/RN _6969_/CLK _6969_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_167_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold890 _4290_/Z _6799_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_67_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ hold24/Z _3535_/Z hold42/Z hold6/Z _4322_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_141_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4251_ hold48/Z hold616/Z _4252_/S _4251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4182_ _4182_/A1 hold32/Z _4184_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_68_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_106__1359_ net413_62/I net413_54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_89__1359_ net513_175/I net763_420/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_169_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6823_ _6823_/D _7008_/RN _6823_/CLK _6823_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _6754_/D _7260_/RN _6754_/CLK _7312_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3966_ _3966_/I _6868_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ hold723/Z hold65/Z _5709_/S _5705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6685_ _6685_/D _7008_/RN _6685_/CLK _6685_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_176_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5636_ hold12/Z hold279/Z _5637_/S _5636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3897_ _3897_/A1 _3897_/A2 _3855_/Z _3896_/Z _6565_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_164_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ hold227/Z hold627/Z _5574_/S _5567_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold131 _7117_/Q hold131/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold120 _5892_/Z _7221_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4518_ _4835_/A2 _4456_/B _5269_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_117_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold142 _5820_/Z _7157_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold153 _6944_/Q hold153/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ hold472/Z _4103_/I _5502_/S _5498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4449_ _4853_/A1 _5464_/A1 _4501_/B _4451_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_160_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7237_ _7237_/D _7237_/RN _7258_/CLK _7237_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold175 _5873_/Z _7204_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold186 _7212_/Q hold186/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold164 _4118_/Z _6673_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_137_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold197 _5587_/Z _6950_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_113_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7168_ _7168_/D _7256_/RN _7168_/CLK _7168_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_3004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7099_ _7099_/D _7237_/RN _7099_/CLK _7099_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_74_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ hold82/I _5960_/Z _6133_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_3037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet413_61 net413_77/I _7164_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_94 net413_95/I _7131_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__20 _4073__9/I _7205_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_72 net413_72/I _7153_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__31 net413_64/I _7194_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__42 net413_57/I _7183_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_83 net413_83/I _7142_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ _3527_/Z _3578_/Z _4274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3751_ _3751_/A1 _3751_/A2 _3732_/Z _3751_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_158_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _7050_/Q _6241_/Z _6251_/Z _6986_/Q _6268_/Z hold50/I _6472_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_9_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3682_ hold62/I _5638_/A1 _3912_/B1 _6888_/Q _3686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_127_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _5420_/Z _5421_/A2 _5421_/A3 _5421_/A4 _5489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_64_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _5191_/Z _5352_/A2 _5285_/B _5020_/Z _5352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput214 _4067_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xoutput225 _7323_/Z mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput203 _3375_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput236 _7331_/Z mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput258 _6887_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput247 _4075_/Z pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4303_ hold895/Z hold291/Z _4303_/S _4303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5283_ _5278_/C _4554_/Z _5283_/B _5471_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_87_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7022_ _7022_/D _7260_/RN _7022_/CLK _7022_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xoutput269 _6884_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4234_ hold448/Z hold91/Z _4244_/S _4234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _4103_/I hold662/Z _4166_/S _4165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4096_ _4097_/A1 _4096_/A2 _6829_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _6806_/D _6818_/CLK _6806_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4998_ _5340_/A1 _4998_/A2 _5262_/A2 _5343_/A2 _4998_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_56_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6737_ _6737_/D _7256_/RN _6737_/CLK _7317_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3949_ _3949_/A1 _3949_/A2 _3949_/A3 _3949_/A4 _3949_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_164_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6668_ _6668_/D _7238_/RN _6668_/CLK _6668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6599_ _6599_/I0 _7276_/Q _6602_/S _7276_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5619_ hold2/Z hold332/Z _5619_/S _5619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_72__1359_ net513_167/I net563_246/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5970_ _7102_/Q _5967_/Z _5969_/Z _7118_/Q _5974_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4921_ _4920_/Z _4890_/I _4926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_79_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _4852_/A1 _5106_/A2 _4852_/A3 _4855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_127_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3803_ _3529_/Z _3680_/Z _3930_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4783_ _4836_/A4 _4530_/I _5137_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3734_ _3734_/I _3735_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6522_ _6696_/Q _6282_/Z _6302_/Z _6712_/Q _6526_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _7066_/Q _6257_/Z _6275_/Z _7042_/Q _6300_/Z _7108_/Q _6466_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3665_ _7009_/Q _3934_/A2 _3954_/A2 hold27/I _3674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ _5404_/A1 _5314_/Z _5404_/A3 _5404_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6384_ _6384_/A1 _6384_/A2 _6380_/Z _6383_/Z _6384_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3596_ _3592_/Z _3596_/A2 _3596_/A3 _3596_/A4 _3596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5335_ _4908_/Z _5245_/Z _5481_/B1 _4905_/Z _5335_/C _5447_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_130_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _5265_/Z _5341_/B _4994_/Z _5266_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_142_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4217_ hold97/Z hold91/Z _4227_/S _4217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7005_ _7005_/D _7008_/RN _7005_/CLK _7005_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5197_ _5346_/A2 _5349_/A1 _5276_/C _5205_/A1 _5197_/C _5390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_84_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ hold869/Z hold291/Z _4148_/S _4148_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ _4079_/I _4079_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7265_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_182_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold719 _6777_/Q hold719/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold708 _4138_/Z _6690_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3450_ _3450_/A1 _3450_/A2 _7292_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_171_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3381_ _6931_/Q _6500_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5120_ _5118_/Z _5238_/A1 _5127_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5051_ _4698_/B _5343_/A1 _5051_/S _5051_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_123_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4002_ _7225_/Q _7226_/Q _5954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_320 _4073__49/I _6905_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_342 net413_75/I _6883_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_331 net763_427/I _6894_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5953_ _5953_/I0 _7239_/Q _5955_/S _7239_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _5263_/A2 _4903_/Z _5255_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5884_ _3485_/Z _3515_/Z _5520_/C _5892_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_178_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4835_ _4555_/C _4835_/A2 _5129_/A3 _5420_/A2 _5368_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4766_ _4766_/A1 _4766_/A2 _4762_/Z _4765_/Z _4770_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3717_ _6928_/Q _3935_/A2 _3943_/A2 _7072_/Q _6895_/Q _5528_/S _3719_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6505_ _6853_/Q _6241_/Z _6297_/Z _7076_/Q _6512_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_147_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4697_ _4467_/B _4463_/Z _5302_/B _5099_/A2 _4697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_14_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ hold58/I _6292_/Z _6300_/Z _7107_/Q _6437_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3648_ _6570_/I0 _6873_/Q _3898_/S _3648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6367_ _7253_/Q _6367_/I1 _6558_/S _7253_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3579_ _3533_/Z _3578_/Z _3959_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_121_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5318_ _5318_/A1 _5314_/Z _5316_/Z _5318_/A4 _5320_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_96_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6298_ _7158_/Q _6296_/Z _6297_/Z _6698_/Q _6298_/C _6307_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold13 hold13/I hold13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5249_ _5410_/A1 _5245_/Z _5250_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_152_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold24 hold24/I hold24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold46 hold46/I hold46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold35 hold35/I hold35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_188_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold68 hold68/I hold68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold57 hold57/I hold57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold79 hold79/I hold79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_283 net713_394/I _6942_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_272 net613_275/I _6953_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_261 net613_261/I _6964_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_188_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_294 net613_294/I _6931_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4620_ _4557_/Z _4604_/Z _5353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4551_ _5129_/A3 _5051_/S _3401_/I _3402_/I _4551_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4482_ _4381_/Z _4485_/A2 _4390_/Z _5170_/A3 _4486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_171_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7270_ _7270_/D _7279_/RN _7279_/CLK _7270_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold516 _6921_/Q hold516/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3502_ _3617_/A1 _3501_/Z _3904_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold527 _7178_/Q hold527/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold505 _5651_/Z _7007_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3433_ _3427_/Z _3433_/A2 _3433_/B _3435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_171_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold549 _5533_/Z _6903_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold538 _4152_/Z _6700_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6221_ _6725_/Q _5984_/Z _5997_/Z _6717_/Q _6695_/Q _5980_/Z _6228_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_131_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6152_ _6152_/A1 _6152_/A2 _6152_/A3 _6152_/A4 _6152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3364_ _7047_/Q _3364_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5103_ _5103_/A1 _5101_/Z _5103_/A3 _5308_/A2 _5108_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ _7283_/Q _4022_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6083_ hold69/I _5964_/Z _5999_/Z _7031_/Q _6084_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _5190_/A2 _4604_/Z _5003_/Z _5034_/B _5204_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ hold21/Z _7260_/RN _6985_/CLK _6985_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5936_ _6745_/Q _7233_/Q _7232_/Q _5936_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_15_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ hold227/Z hold660/Z _5874_/S _5867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4818_ _4624_/Z _4817_/Z _5313_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5798_ hold65/Z hold155/Z _5802_/S _5798_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4749_ _4703_/Z _5230_/B _5313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_162_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6419_ _6744_/Q _7254_/Q _6419_/B _6420_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_89_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput136 wb_dat_i[17] _6582_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput103 wb_adr_i[17] _4391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput114 wb_adr_i[27] _4027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput125 wb_adr_i[8] _4388_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput147 wb_dat_i[27] _6588_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput158 wb_dat_i[8] _6579_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3982_ _3981_/Z _6660_/Q _3988_/S _6660_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6770_ _6770_/D _7256_/RN _6770_/CLK _6770_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5721_ hold291/Z hold982/Z _5727_/S _5721_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ hold495/Z hold48/Z _5655_/S _5652_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4603_ _4580_/B _4604_/A3 _5351_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_49__1359_ net413_93/I net413_80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5583_ _6947_/Q hold2/Z _5583_/S hold3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4534_ _4782_/A1 _4736_/A3 _4736_/A1 _4436_/B _4534_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7322_ _7322_/I _7322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold302 _6995_/Q hold302/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold335 _5691_/Z _7043_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold313 _5784_/Z _7125_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold324 _5825_/Z _7161_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7253_ _7253_/D _7256_/RN _7258_/CLK _7253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold357 _5549_/Z _6916_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4465_ _5315_/A1 _4481_/A2 _4473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold346 _7023_/Q hold346/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold368 _5854_/Z _7187_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4396_ _5385_/A1 _4385_/Z _4922_/A3 _4424_/B _5002_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3416_ _7305_/Q _3415_/Z _3416_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7184_ _7184_/D _7256_/RN _7184_/CLK _7184_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6204_ _6198_/Z _6201_/Z _6204_/A3 _6204_/A4 _6204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold379 _5707_/Z _7057_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3347_ _7177_/Q _3732_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_98_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _6127_/Z _6134_/Z _6447_/B1 _6168_/C _6136_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6066_ _7023_/Q _6068_/A4 _6211_/B1 _6991_/Q _6067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1002 _6868_/Q _3965_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XTAP_3219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _5017_/A1 _5197_/C _5019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_456 _4073__11/I _6709_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_467 net813_467/I _6698_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_489 net813_489/I _6676_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_478 net813_481/I _6687_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6968_ _6968_/D _7258_/RN _6968_/CLK _6968_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_167_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ _6021_/A2 _6015_/A3 _5984_/A1 _6745_/Q _5919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_50_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6899_ hold18/Z _7238_/RN _6899_/CLK _6899_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold880 _5493_/Z _6867_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold891 _7005_/Q hold891/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_107_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4250_ hold65/Z hold149/Z _4252_/S _4250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ hold291/Z hold757/Z _4181_/S _4181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6822_ _6822_/D _7008_/RN _6822_/CLK _6822_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6753_ _6753_/D _7170_/RN _6753_/CLK _6753_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3965_ _6564_/I0 _3965_/A2 _3965_/B1 _3899_/S _3966_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_188_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5704_ hold576/Z hold91/Z _5709_/S _5704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6684_ _6684_/D _7008_/RN _6684_/CLK _6684_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3896_ _3860_/Z _3869_/Z _3885_/Z _3895_/Z _3896_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ hold20/Z hold27/Z _5637_/S hold28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold110 _5547_/Z _6915_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5566_ hold24/Z _3521_/Z hold42/Z hold6/Z _5574_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4517_ _5165_/A4 _5003_/A2 _4491_/B _5438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7305_ _7305_/D _6657_/Z _7305_/CLK _7305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold132 _5775_/Z _7117_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold121 _6705_/Q hold121/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold143 _7109_/Q hold143/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5497_ _5647_/A1 hold16/Z hold32/Z hold6/Z _5502_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4448_ _3401_/I _5288_/C _4369_/Z _5288_/B _4451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7236_ _7236_/D _7235_/RN _4067_/I1 _7236_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold176 _7326_/I hold176/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold154 _5580_/Z _6944_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold165 _7022_/Q hold165/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold198 _7188_/Q hold198/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold187 _5882_/Z _7212_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_120_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4379_ _4853_/A1 _5464_/A1 _4604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_99_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7167_ _7167_/D _7218_/RN _7167_/CLK _7167_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7098_ _7098_/D _7218_/RN _7098_/CLK _7098_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _7057_/Q _5924_/Z _6168_/C _6127_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_3027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6049_ _6942_/Q _5972_/Z _6021_/Z _6998_/Q _6049_/C _6053_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_58_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_32__1359_ clkbuf_opt_3_0__1359_/Z net663_317/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112__1359_ net513_165/I net813_466/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_95__1359_ clkbuf_4_5_0__1359_/Z net763_422/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_95 net413_95/I _7130_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__21 _4073__9/I _7204_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__10 _4073__7/I _7215_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__32 net413_64/I _7193_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet413_73 net413_73/I _7152_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_84 net413_84/I _7141_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_62 net413_62/I _7163_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__43 _4073__43/I _7182_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3750_ _7007_/Q _3934_/A2 _5638_/A1 _6999_/Q _3916_/B1 _6881_/Q _3751_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3681_ _3527_/Z _3680_/Z _3912_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _5420_/A1 _5420_/A2 _5420_/A3 _4456_/B _5420_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet713_400 net413_56/I _6774_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5351_ _5356_/A1 _5387_/A2 _5356_/B _5351_/C _5352_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput215 _4066_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_133_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput226 _7324_/Z mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_127_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput204 _3374_/ZN mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_57_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput237 _4055_/Z mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5282_ _5281_/C _4467_/B _5399_/A2 _4683_/Z _5283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_99_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput248 _4094_/ZN pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4302_ hold871/Z _4103_/I _4303_/S _4302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput259 _6888_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4233_ _4232_/Z hold827/Z _4245_/S _4233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7021_ _7021_/D _7260_/RN _7021_/CLK _7021_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_141_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _5520_/C _3552_/Z hold235/Z _5821_/A3 _4166_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4095_ _4097_/A1 _4900_/B _6831_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6805_ _6805_/D _6818_/CLK _6805_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6736_ _6736_/D _7256_/RN _6736_/CLK _7316_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4997_ _4546_/Z _4716_/Z _4997_/B _4997_/C _4999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_176_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3948_ input43/Z _4210_/S _4194_/A1 input52/Z _3948_/C1 input61/Z _3949_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ _7087_/Q _3945_/B1 _3952_/A2 _7045_/Q _3950_/C1 _6844_/Q _3880_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6667_ _6667_/D _7238_/RN _6667_/CLK _6667_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6598_ _6598_/A1 _4313_/Z _6598_/B _6599_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_164_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ hold12/Z hold276/Z _5619_/S _5618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5549_ hold227/Z hold356/Z _5556_/S _5549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _6818_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7219_ _7219_/D _7237_/RN _7219_/CLK _7219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_48_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _5130_/B2 _5420_/A3 _4367_/Z _4920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_64_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _5287_/C _4833_/Z _4852_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3802_ _3509_/Z _3540_/Z _3925_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_127_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4782_ _4782_/A1 _4510_/Z _5302_/B _5099_/A1 _5213_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_158_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3733_ _7193_/Q _3909_/A2 _5683_/A1 _7039_/Q _3952_/A2 _7047_/Q _3734_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6521_ _6521_/A1 _6521_/A2 _6521_/A3 _6521_/A4 _6521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6452_ _7074_/Q _6484_/A2 _6484_/A3 _6452_/A4 _6456_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3664_ input17/Z _3913_/A2 _5674_/A1 _7033_/Q _3674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_118_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5403_ _4699_/Z _5403_/A2 _5456_/A2 _5403_/B2 _5403_/C _5404_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_173_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6383_ _6383_/A1 _6383_/A2 _6383_/A3 _6383_/A4 _6383_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3595_ _6995_/Q _3954_/A2 _3927_/A2 _6705_/Q _3596_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5334_ _5334_/A1 _5334_/A2 _5334_/A3 _5334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_170_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5265_ _5265_/A1 _4991_/C _5392_/B _5265_/A4 _5265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_142_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5196_ _5347_/A1 _5437_/A1 _5195_/Z _5347_/A3 _5196_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4216_ _4215_/Z hold815/Z _4228_/S _4216_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7004_ _7004_/D _7008_/RN _7004_/CLK _7004_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_69_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4147_ hold687/Z _4103_/I _4148_/S _4147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _4081_/A1 input86/Z _4079_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_44_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6719_ _6719_/D _7008_/RN _6719_/CLK _6719_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold709 _6726_/Q hold709/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_155_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3380_ _6930_/Q _6473_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_124_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _5343_/A2 _5389_/A2 _5078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_112_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4001_ _4001_/I _6836_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_310 net763_409/I _6915_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_321 net413_72/I _6904_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_343 net813_487/I _6882_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_332 net813_491/I _6893_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _6746_/Q _6744_/Q _5952_/A3 _5952_/B _5955_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_81_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _4467_/B _4407_/Z _4495_/Z _5259_/A1 _4903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_179_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5883_ hold2/Z hold129/Z _5883_/S _5883_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4834_ _4834_/A1 _4834_/A2 _4846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_178_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4765_ _4765_/A1 _5302_/B _4700_/Z _5226_/C _4765_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_140_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3716_ _7130_/Q _3930_/A2 _3925_/A2 input7/Z _5647_/A1 _3904_/A2 _3719_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_53_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6504_ _6789_/Q _6245_/Z _6274_/Z _6851_/Q _6512_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4696_ _5099_/A2 _4695_/Z _4704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_162_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3647_ _3647_/A1 _3625_/Z _3646_/Z _3647_/A4 _6570_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6435_ _7187_/Q _6282_/Z _6299_/Z _7057_/Q hold27/I _6237_/Z _6439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6366_ _6366_/I _6367_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3578_ _3653_/A1 hold320/Z _3617_/A1 hold673/Z _3578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5317_ _5317_/A1 _5454_/A1 _5318_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6297_ _6300_/A2 _6484_/A3 _5943_/S _5942_/S _6297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold14 hold14/I hold14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5248_ _5246_/Z _5248_/A2 _5442_/A2 _5056_/C _5248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold47 hold47/I hold47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold25 hold25/I hold25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_57_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold36 hold36/I hold36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _5240_/B _5343_/A2 _5179_/B _5242_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold58 hold58/I hold58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold69 hold69/I hold69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_84_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_273 net813_492/I _6952_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_262 net613_262/I _6963_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_188_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_295 net613_297/I _6930_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_284 net613_284/I _6941_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4550_ _4454_/Z _5269_/A2 _5368_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4481_ _4481_/A1 _4481_/A2 _4486_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3501_ _3499_/I _3305_/I hold54/Z _3501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
Xhold517 _5554_/Z _6921_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold506 _6934_/Q hold506/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3432_ _3432_/I _7299_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold528 _5844_/Z _7178_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold539 _6958_/Q hold539/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6220_ _6217_/Z _6220_/A2 _6220_/A3 _6220_/A4 _6220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3363_ _7055_/Q _3363_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6151_ _7148_/Q _5987_/Z _6015_/Z _7010_/Q _6152_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5102_ _4586_/Z _4817_/Z _5103_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ _7169_/Q _6006_/Z _6014_/Z _6959_/Q _6084_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3294_ _7300_/Q _4081_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _5035_/A4 _5032_/Z _5388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6984_ _6984_/D _7258_/RN _6984_/CLK _6984_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_20_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5935_ _6282_/A2 _6279_/A3 _6300_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_80_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _3485_/Z _3507_/Z hold24/Z _5874_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_167_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _5420_/A3 _5287_/B _3402_/I _5269_/A2 _4817_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5797_ hold91/Z hold221/Z _5802_/S _5797_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_11_0__1359_ clkbuf_0__1359_/Z net413_93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4748_ _4510_/Z _5302_/B _5099_/A1 _5226_/C _4748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_31_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4679_ _4670_/Z _5451_/C _4685_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6418_ _6411_/Z _6417_/Z _6418_/B1 _6286_/Z _6555_/C _6419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_122_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6349_ _7200_/Q _6272_/Z _6282_/Z _7184_/Q _6296_/Z _7160_/Q _6356_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xinput104 wb_adr_i[18] _4391_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput126 wb_adr_i[9] _4388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput115 wb_adr_i[28] _4027_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0__1359_ _4072_/ZN clkbuf_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput148 wb_dat_i[28] _6591_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput137 wb_dat_i[18] _6585_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput159 wb_dat_i[9] _6582_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3981_ _3981_/A1 _3981_/A2 _3981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5720_ hold227/Z hold641/Z _5727_/S _5720_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ hold504/Z hold65/Z _5655_/S _5651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4602_ _4524_/Z _5399_/A2 _4554_/Z _5364_/B _5285_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5582_ hold45/Z hold12/Z _5583_/S hold46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _4736_/A3 _4690_/C _4713_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7321_ _7321_/I _7321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7252_ _7252_/D _7256_/RN _7258_/CLK _7252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold314 _7101_/Q hold314/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold303 _5637_/Z _6995_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold325 _7193_/Q hold325/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold358 _6922_/Q hold358/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4464_ _4456_/B _5051_/S _4460_/B _4436_/B _4464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold336 _6931_/Q hold336/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold347 _5669_/Z _7023_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold369 _7040_/Q hold369/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6203_ _6724_/Q _5984_/Z _6000_/Z _6728_/Q _6710_/Q _6006_/Z _6204_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4395_ _4580_/C _4489_/A1 _4483_/B _5002_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3415_ _7304_/Q _7303_/Q _3415_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_98_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7183_ _7183_/D _7008_/RN _7183_/CLK _7183_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3346_ _7185_/Q _3346_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _6134_/A1 _6134_/A2 _6134_/A3 _6133_/Z _6134_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_113_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6065_ _7243_/Q _6065_/I1 _6558_/S _7243_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold1003 _6875_/Q _3611_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _5438_/C _4551_/Z _4586_/Z _5003_/Z _5016_/B2 _5197_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_85_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_457 net413_74/I _6708_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _6967_/D _7260_/RN _6967_/CLK _6967_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet813_479 net813_487/I _6686_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet813_468 net413_63/I _6697_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5918_ _6745_/Q _5917_/Z _5913_/I _6021_/A2 _7228_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_107_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6898_ _6898_/D _7238_/RN _6898_/CLK hold39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5849_ hold227/Z hold653/Z _5856_/S _5849_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold881 _6693_/Q hold881/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold870 _4148_/Z _6697_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold892 _5649_/Z _7005_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55__1359_ net663_324/I net463_110/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_135__1359_ clkbuf_4_1_0__1359_/Z net813_481/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _4103_/I hold715/Z _4181_/S _4180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6821_ _6821_/D _7008_/RN _6821_/CLK _6821_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6752_ _6752_/D _7260_/RN _6752_/CLK _7311_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3964_ _3898_/S _3899_/S _3965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ hold975/Z hold291/Z _5709_/S _5703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6683_ _6683_/D _7008_/RN _6683_/CLK _6683_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3895_ _3895_/A1 _3889_/Z _3895_/A3 _3894_/Z _3895_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_31_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5634_ hold48/Z hold88/Z _5637_/S hold89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7304_ _7304_/D _6656_/Z _7304_/CLK _7304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5565_ hold2/Z hold336/Z _5565_/S _5565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold100 _5799_/Z _7138_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4516_ _5003_/A2 _4561_/A2 _5389_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_176_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold122 _4157_/Z _6705_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold133 _7165_/Q hold133/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold144 _5766_/Z _7109_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold111 _6783_/Q hold111/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5496_ hold291/Z _6877_/Q _5496_/S _5496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4447_ _5420_/A2 _4853_/A1 _5270_/A1 _4501_/B _4504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_171_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7235_ _7235_/D _7235_/RN _4067_/I1 _7235_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold177 _5543_/Z _6911_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold155 _7137_/Q hold155/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold166 _5668_/Z _7022_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold199 _5855_/Z _7188_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold188 _7327_/I hold188/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7166_ _7166_/D _7218_/RN _7166_/CLK _7166_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4378_ _5281_/C _5464_/A1 _4648_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_101_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6117_ _7073_/Q _7231_/Q _6210_/C _6117_/A4 _6128_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ _7234_/Q _5942_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_7097_ _7097_/D _7218_/RN _7097_/CLK _7097_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6048_ _5925_/Z _6048_/A2 _6048_/B _6048_/C _6049_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_37_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_52 net413_68/I _7173_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__22 _4073__22/I _7203_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073__11 _4073__11/I _7214_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_74 net413_74/I _7151_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_85 net413_89/I _7140_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_63 net413_63/I _7162_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_96 net413_96/I _7129_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__33 net413_80/I _7192_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__44 _4073__46/I _7181_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3680_ _3489_/I _3492_/Z _3497_/I hold673/Z _3680_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet713_401 net763_431/I _6773_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput216 _7315_/Z mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5350_ _5350_/A1 _5350_/A2 _5350_/A3 _5350_/A4 _5350_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput205 _3373_/ZN mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput238 _4048_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput227 _7325_/Z mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5281_ _5288_/A1 _5281_/A2 _5281_/B _5281_/C _5369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput249 _4074_/Z pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4301_ _4301_/A1 hold32/Z _4303_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4232_ hold811/Z hold291/Z _4244_/S _4232_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7020_ _7020_/D _7260_/RN _7020_/CLK _7020_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_96_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ hold957/Z hold291/Z _4163_/S _4163_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4094_ _4094_/I _4094_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_167_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ _5083_/C _4997_/C _4716_/Z _4422_/Z _5341_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6804_ _6804_/D _7265_/CLK _6804_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6735_ _6735_/D _7256_/RN _6735_/CLK _7315_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3947_ _7094_/Q _3947_/A2 _3947_/B1 _6716_/Q _3949_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_165_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6666_ _6666_/D _7238_/RN _6666_/CLK _6666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3878_ _6904_/Q _5532_/A1 _3935_/B1 _6850_/Q _3885_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6597_ _6834_/Q _6597_/A2 _6597_/B1 _6835_/Q _6836_/Q _6597_/C2 _6598_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5617_ hold20/Z hold29/Z _5619_/S hold30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ _3485_/Z _3542_/Z _6652_/A2 hold24/Z _5556_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_132_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5479_ _5479_/A1 _5479_/A2 _5479_/A3 _5479_/A4 _5479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7218_ _7218_/D _7218_/RN _7218_/CLK _7218_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7149_ _7149_/D _7256_/RN _7149_/CLK _7149_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_63_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _5287_/C _4817_/Z _5106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3801_ _3509_/Z _3653_/Z _3928_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_159_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4781_ _4781_/A1 _5121_/A1 _5456_/B _5122_/B _4790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6520_ _6710_/Q _5948_/Z _6292_/Z _6722_/Q _6521_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_186_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3732_ _3732_/A1 _5857_/A3 _5839_/A3 _3552_/Z _3732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_13_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _7212_/Q _6256_/Z _6464_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_9_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _3663_/A1 _3663_/A2 _3663_/A3 _3663_/A4 _3663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6382_ _7039_/Q _6275_/Z _6300_/Z _7105_/Q _6383_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5402_ _5480_/A1 _5480_/A2 _5406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5333_ _4761_/I _5481_/B1 _5334_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3594_ _6963_/Q _3957_/A2 _3927_/C2 input33/Z _5575_/A1 _6947_/Q _3596_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_170_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5264_ _5264_/A1 _5412_/A3 _5264_/A3 _5263_/Z _5265_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_88_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5195_ _5350_/A1 _5350_/A3 _5195_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_141_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4215_ hold781/Z hold291/Z _4227_/S _4215_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7003_ _7003_/D _7258_/RN _7003_/CLK _7003_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_84_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ _4146_/A1 hold32/Z _4148_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_110_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4077_ _4077_/I _4077_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4979_ _4419_/Z _4973_/Z _4979_/B _4979_/C _4986_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6718_ _6718_/D _7008_/RN _6718_/CLK _6718_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6649_ _7235_/RN _6653_/A2 _6649_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_164_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4000_ _6836_/Q _4097_/A1 _6831_/Q _4001_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_111_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet663_311 net763_406/I _6914_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_322 net663_322/I _6903_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_344 net813_455/I _6881_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_333 net813_499/I _6892_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0__1359_ clkbuf_0__1359_/Z _4073__49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5951_ _7225_/Q _7226_/Q _5951_/A3 _6746_/Q _5952_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_92_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _4436_/B _4494_/Z _5323_/B _4902_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5882_ hold12/Z hold186/Z _5883_/S _5882_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _4422_/Z _4530_/I _4878_/A2 _4483_/B _4833_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_140_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4764_ _4765_/A1 _5302_/B _4764_/A3 _4692_/C _4764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_53_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _7258_/Q _6503_/I1 _6558_/S _7258_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3715_ _3715_/A1 _3715_/A2 _3715_/A3 _3715_/A4 _3715_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_119_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4695_ _4736_/A3 _4467_/B _4736_/A1 _4695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6434_ _6434_/A1 _6434_/A2 _6434_/A3 _6434_/A4 _6434_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3646_ _3646_/A1 _3630_/Z _3646_/A3 _3645_/Z _3646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6365_ _6744_/Q _7252_/Q _6365_/B _6366_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_115_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3577_ _3512_/Z _3537_/Z _3947_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_142_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _7235_/Q _7234_/Q _6484_/A2 _6484_/A3 _6296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ _5316_/A1 _5316_/A2 _5315_/Z _4772_/Z _5316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_170_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5247_ _5246_/Z _5442_/A2 _5056_/C _4496_/Z _5247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold15 hold15/I hold15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold37 hold37/I hold37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold26 hold26/I hold26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5178_ _5180_/A3 _5180_/A2 _5211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold48 hold48/I hold48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_69_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold59 hold59/I hold59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_28_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _4103_/I hold941/Z _4136_/S _4129_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_263 net613_263/I _6962_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_252 net613_268/I _6973_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_274 net613_279/I _6951_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_285 net813_492/I _6940_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet613_296 net663_330/I _6929_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3500_ _3500_/I0 _3500_/I1 hold54/Z _3500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_183_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _4463_/Z _4468_/Z _4786_/A2 _4786_/A3 _4808_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold507 _5569_/Z _6934_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold518 _7014_/Q hold518/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_13_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3431_ _6734_/Q _3434_/B _7299_/Q _3432_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold529 _7039_/Q hold529/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3362_ _7063_/Q _3362_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _7092_/Q _6002_/Z _6003_/Z _7164_/Q _6152_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_98_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5101_ _5303_/A1 _5460_/A1 _5101_/A3 _5303_/A2 _5101_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_98_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3293_ _7301_/Q _3428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6081_ _7113_/Q _5984_/Z _5997_/Z _7097_/Q _7071_/Q _5980_/Z _6084_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_98_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _4397_/Z _4411_/Z _5328_/A1 _5387_/A1 _5032_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6983_ _6983_/D _7258_/RN _6983_/CLK _6983_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_53_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _5934_/I _7232_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ hold2/Z hold382/Z _5865_/S _5865_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _5287_/B _4673_/Z _5132_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5796_ hold291/Z hold833/Z _5802_/S _5796_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4747_ _4747_/A1 _4747_/A2 _5231_/C _4751_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_31_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4678_ _4997_/C _4673_/Z _4675_/Z _5451_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3629_ _7124_/Q _3956_/A2 _3927_/B1 _7066_/Q _3630_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6417_ _6554_/A1 _6417_/A2 _6417_/A3 _6417_/A4 _6417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6348_ _7136_/Q _6253_/Z _6293_/Z _7152_/Q _6348_/C _6356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_143_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput127 wb_cyc_i _4032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput116 wb_adr_i[29] _4031_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput105 wb_adr_i[19] _4391_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6279_ _6452_/A4 _6285_/A2 _6279_/A3 _7237_/Q _6279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_131_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput149 wb_dat_i[29] _6594_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput138 wb_dat_i[19] _6588_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_15__1359_ clkbuf_4_2_0__1359_/Z net813_473/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78__1359_ clkbuf_opt_1_0__1359_/Z net413_57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ _6733_/Q _3972_/Z _6659_/Q _3981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_90_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5650_ hold566/Z hold91/Z _5655_/S _5650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4601_ _4601_/A1 _4595_/Z _4599_/Z _4600_/Z _4601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_148_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5581_ hold35/Z hold20/Z _5583_/S hold36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4532_ _5420_/A2 _4456_/B _5051_/S _3401_/I _5414_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7320_ _7320_/I _7320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7251_ _7251_/D _7256_/RN _7258_/CLK _7251_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4463_ _4460_/B _4481_/A2 _4463_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xhold315 _5757_/Z _7101_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold326 _5861_/Z _7193_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold304 _6676_/Q hold304/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3414_ _6733_/Q _3413_/Z _3442_/B _3988_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_172_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold359 _5555_/Z _6922_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold337 _5565_/Z _6931_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold348 _7162_/Q hold348/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6202_ _6799_/Q _5958_/Z _5969_/Z _7296_/Q _6726_/Q _5994_/I _6204_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4394_ _4427_/A3 _4481_/A1 _4922_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ _7182_/D _7218_/RN _7182_/CLK _7182_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3345_ _7193_/Q _3345_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _6133_/A1 _6133_/A2 _6133_/A3 _6133_/A4 _6133_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold1004 _6731_/Q _4023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_112_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6064_ _6064_/I _6065_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _5013_/Z _5350_/A2 _5017_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_458 net413_59/I _6707_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _6966_/D _7238_/RN _6966_/CLK _6966_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_26_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet813_469 net813_469/I _6696_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5917_ _7228_/Q _7227_/Q _5917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6897_ hold92/Z _7238_/RN _6897_/CLK _6897_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _3485_/Z _3521_/Z hold24/Z _5856_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_10_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5779_ hold91/Z hold550/Z _5784_/S _5779_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold882 _4142_/Z _6693_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold871 _6809_/Q hold871/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold860 _4172_/Z _6715_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold893 _6906_/Q hold893/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2__1359_ net763_436/I net763_421/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6820_ _6820_/D _7008_/RN _6820_/CLK _6820_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _6751_/D _7260_/RN _6751_/CLK _7310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3963_ _3915_/Z _3919_/Z _3963_/A3 _3962_/Z _6564_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5702_ hold624/Z hold227/Z _5709_/S _5702_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6682_ _6682_/D _7008_/RN _6682_/CLK _6682_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3894_ _3894_/A1 _3894_/A2 _3894_/A3 _3894_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5633_ hold65/Z hold339/Z _5637_/S _5633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5564_ hold12/Z hold293/Z _5565_/S _5564_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7303_ _7303_/D _6655_/Z _7305_/CLK _7303_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4515_ _5002_/A3 _5002_/A4 _5083_/B _4561_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_89_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold101 _6951_/Q hold101/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold123 _7133_/Q hold123/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold134 _5829_/Z _7165_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold112 _4269_/Z _6783_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5495_ _4103_/I _6876_/Q _5496_/S _5495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7234_ _7234_/D _7235_/RN _4067_/I1 _7234_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4446_ _4441_/B _5281_/C _4467_/B _4501_/B _5287_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_132_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold145 _7173_/Q hold145/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold156 _5798_/Z _7137_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold167 _6966_/Q hold167/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4377_ _3401_/I _3402_/I _4456_/B _5051_/S _5464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_61__1359_ net513_170/I net763_415/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold178 _7325_/I hold178/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold189 _5544_/Z _6912_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7165_ _7165_/D _7256_/RN _7165_/CLK _7165_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_leaf_141__1359_ clkbuf_4_1_0__1359_/Z net813_470/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3328_ _7235_/Q _5943_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_113_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _6116_/A1 _5991_/Z _6132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ _7096_/D _7256_/RN _7096_/CLK _7096_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6047_ _7144_/Q _5987_/Z _6015_/Z _7006_/Q _6047_/C _6048_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_27_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6949_ _6949_/D _7260_/RN _6949_/CLK _6949_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_179_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold690 _4327_/Z _6824_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__12 net413_60/I _7213_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_53 net413_93/I _7172_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__23 net413_57/I _7202_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_64 net413_64/I _7161_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_86 net413_89/I _7139_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_75 net413_75/I _7150_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_97 net413_97/I _7128_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__45 _4073__46/I _7180_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__34 _4073__7/I _7191_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput217 _7316_/Z mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput206 _3372_/ZN mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput239 _4047_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5280_ _5372_/A1 _5055_/Z _5284_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xoutput228 _7326_/Z mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4300_ _6571_/I0 _6808_/Q _4300_/S _6808_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4231_ _4230_/Z hold779/Z _4245_/S _4231_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4162_ hold831/Z _4103_/I _4163_/S _4162_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4093_ _7299_/Q _7170_/RN _4094_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ _4892_/B _4716_/Z _5428_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6803_ _6803_/D _6818_/CLK _6803_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _6734_/D _6625_/Z _7305_/CLK _6734_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3946_ _6720_/Q _3946_/A2 _4161_/A1 _6708_/Q _6674_/Q _3546_/Z _3949_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_182_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6665_ _6665_/D _6620_/Z _7305_/CLK _6665_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_17_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3877_ _7005_/Q _3934_/A2 _3916_/B1 _6879_/Q _3885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6596_ _6596_/I0 _7275_/Q _6602_/S _7275_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5616_ hold48/Z hold464/Z _5619_/S _5616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5547_ hold2/Z hold109/Z _5547_/S _5547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5478_ _4614_/Z _4683_/Z _5302_/B _4700_/Z _5230_/B _5479_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_4429_ _5083_/C _4422_/Z _5340_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7217_ _7217_/D _7237_/RN _7217_/CLK _7217_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_7148_ _7148_/D _7237_/RN _7148_/CLK _7148_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7079_ _7079_/D _7008_/RN _7079_/CLK _7079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xnet463_150 net813_461/I _7075_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4780_ _4716_/Z _4778_/Z _5122_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3800_ _3509_/Z _3680_/Z _3928_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_33_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ input14/Z _3913_/A2 _3758_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6450_ _7256_/Q _6450_/I1 _6558_/S _7256_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3662_ _7131_/Q _3930_/A2 _3901_/A2 _6985_/Q _3663_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6381_ _7097_/Q _6250_/Z _6290_/Z _7081_/Q _6302_/Z _7089_/Q _6383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5401_ _4694_/Z _4703_/Z _5401_/B _5401_/C _5480_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3593_ _6939_/Q _3910_/A2 _3901_/A2 _6987_/Q _3596_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_62_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5332_ _5444_/A2 _5327_/Z _5482_/A1 _5332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_161_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5263_ _4997_/B _5263_/A2 _4716_/Z _5263_/A4 _5263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_141_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _4555_/C _5205_/A1 _5194_/B1 _5346_/A2 _5350_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_96_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7002_ hold13/Z _7238_/RN _7002_/CLK _7002_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4214_ _4213_/Z hold813/Z _4228_/S _4214_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4145_ hold925/Z hold291/Z _4145_/S _4145_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ _7299_/Q input88/Z _4077_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ _5258_/A2 _4977_/Z _4979_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_138_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3929_ _3926_/Z _3929_/A2 _3929_/A3 _3929_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6717_ _6717_/D _7170_/RN _6717_/CLK _6717_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6648_ _7235_/RN _6653_/A2 _6648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6579_ _6834_/Q _6579_/A2 _6579_/B1 _6835_/Q _6836_/Q _6579_/C2 _6580_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_166_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_312 net763_409/I _6913_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_323 net413_66/I _6902_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_334 net813_491/I _6891_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_345 net813_455/I _6880_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ _5950_/A1 _5950_/A2 _5950_/B1 _6302_/A4 _7237_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_25_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _4700_/Z _4716_/Z _5442_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_179_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5881_ hold20/Z hold342/Z _5883_/S _5881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4832_ _5287_/B _4683_/Z _5281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4763_ _4765_/A1 _5302_/B _5226_/C _5403_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_119_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6502_ _6502_/I _6503_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4694_ _5302_/B _4778_/A4 _4468_/Z _5099_/A2 _4694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_14_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3714_ hold93/I _5665_/A1 _3923_/C1 hold95/I _3714_/C _3715_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _7073_/Q _6248_/Z _6297_/Z _6703_/Q _6433_/C _6434_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3645_ _3638_/Z _3642_/Z _3645_/A3 _3645_/A4 _3645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6364_ _6357_/Z _6363_/Z _6364_/B1 _6286_/Z _6555_/C _6365_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3576_ _3521_/Z _3529_/Z _5638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5315_ _5315_/A1 _5315_/A2 _4683_/Z _5302_/B _5315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6295_ _6295_/I _6298_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5246_ _5258_/B2 _5343_/A2 _5389_/A2 _5255_/A2 _5246_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold16 hold16/I hold16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold27 hold27/I hold27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold38 hold38/I hold38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5177_ _4414_/Z _4878_/Z _5180_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold49 hold49/I hold49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4128_ _5520_/C _3533_/Z _5513_/A3 _5839_/A3 _4136_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_28_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4059_ _6753_/Q input77/Z _4059_/S _4059_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_253 _4073__50/I _6972_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_264 net613_288/I _6961_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet613_286 net413_76/I _6939_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_297 net613_297/I _6928_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_275 net613_275/I _6950_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold508 _7046_/Q hold508/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold519 _7098_/Q hold519/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3430_ _7300_/Q _7283_/Q _3430_/S _7300_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3361_ _7071_/Q _3361_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5100_ _5100_/A1 _5312_/A2 _5220_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6080_ _6943_/Q _5972_/Z _6021_/Z _6999_/Q _6085_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_3_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3292_ _7303_/Q _3422_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5031_ _5028_/Z _5354_/A1 _5202_/A3 _5035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_111_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _6982_/D _7258_/RN _6982_/CLK _6982_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_65_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5933_ _5913_/I _6745_/Q _7232_/Q _5934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ hold12/Z hold476/Z _5865_/S _5864_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _5414_/A2 _4764_/Z _5215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5795_ hold227/Z hold354/Z _5802_/S _5795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _4716_/Z _5230_/B _5231_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_162_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4677_ _4673_/Z _4892_/B _5392_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_107_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3628_ input27/Z _3954_/B1 _3925_/A2 input9/Z _3630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6416_ _6944_/Q _6245_/Z _6262_/Z _6968_/Q _7032_/Q _6269_/Z _6417_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_150_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _7038_/Q _6275_/Z _6300_/Z _7104_/Q _6347_/C _6357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3559_ _3523_/Z _3537_/Z _3923_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput117 wb_adr_i[2] _5051_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xinput106 wb_adr_i[1] _3402_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_131_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6278_ _6276_/Z _6277_/Z _6287_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput139 wb_dat_i[1] _3394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput128 wb_dat_i[0] _3393_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _5229_/A1 _5479_/A2 _5234_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ _4524_/Z _5399_/A2 _4546_/Z _5364_/B _4600_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_157_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5580_ hold153/Z hold48/Z _5583_/S _5580_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4531_ _5270_/A1 _4530_/I _5214_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4462_ _4736_/A1 _4736_/A3 _4778_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold316 _7097_/Q hold316/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold305 _4122_/Z _6676_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7250_ _7250_/D _7260_/RN _7260_/CLK _7250_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3413_ _3412_/Z _3409_/Z _6732_/Q _3413_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_144_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold327 _7011_/Q hold327/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold338 _6967_/Q hold338/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6201_ _6201_/A1 _6201_/A2 _6201_/A3 _6201_/A4 _6201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold349 _5826_/Z _7162_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4393_ _4385_/Z _4387_/Z _4390_/Z _4489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7181_ _7181_/D _7237_/RN _7181_/CLK _7181_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3344_ _6926_/Q _6364_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ hold73/I _5994_/I _6132_/B _6133_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold1005 _7298_/Q _3433_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_140_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6063_ _6555_/C _7242_/Q _6063_/B _6064_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _4555_/C _5439_/A1 _5349_/A1 _5439_/B2 _5350_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6965_ _6965_/D _7218_/RN _6965_/CLK _6965_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xnet813_459 net413_63/I _6706_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5916_ _7228_/Q _7227_/Q _6210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_21__1359_ _4073__7/I _4073__50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6896_ _6896_/D _7260_/RN _6896_/CLK _6896_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_84__1359_ net413_62/I net513_153/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_101__1359_ clkbuf_4_5_0__1359_/Z net613_284/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_167_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ hold2/Z hold388/Z _5847_/S _5847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5778_ hold291/Z hold843/Z _5784_/S _5778_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4729_ _4765_/A1 _5302_/B _5099_/A2 _4700_/Z _4729_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold872 _4302_/Z _6809_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold861 _6851_/Q hold861/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold850 _4151_/Z _6699_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold883 _6707_/Q hold883/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold894 _5537_/Z _6906_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_27_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _6750_/D _7238_/RN _6750_/CLK _7309_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ _5701_/A1 hold32/Z _5709_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_32_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ _3938_/Z _3944_/Z _3949_/Z _3961_/Z _3962_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_189_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _6681_/D _7238_/RN _6681_/CLK _6681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3893_ _7151_/Q _3916_/A2 _5536_/A1 _6907_/Q _3894_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_176_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5632_ hold91/Z hold205/Z _5637_/S _5632_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5563_ hold20/Z hold375/Z _5565_/S _5563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7302_ _7302_/D _6654_/Z _7304_/CLK _7302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4514_ _4414_/Z _4421_/Z _4452_/Z _4810_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_145_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold124 _5793_/Z _7133_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_145_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold135 _7189_/Q hold135/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold113 _7205_/Q hold113/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5494_ hold42/Z _3515_/Z hold24/Z hold273/Z _5494_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold102 _5588_/Z _6951_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4445_ _4853_/A1 _4501_/B _5309_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7233_ _7233_/D _7237_/RN _4067_/I1 _7233_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold157 _7328_/I hold157/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold146 _5838_/Z _7173_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold168 _6681_/Q hold168/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4376_ _3401_/I _3402_/I _4456_/B _5051_/S _4376_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_160_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold179 _5542_/Z _6910_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7164_ _7164_/D _7237_/RN _7164_/CLK _7164_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3327_ _7232_/Q _6279_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_113_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ hold80/I _6211_/A2 _6211_/B1 hold27/I _6116_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_113_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7095_ _7095_/D _7218_/RN _7095_/CLK _7095_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _7160_/Q _7231_/Q _6211_/A2 _6117_/A4 _6047_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6948_ _6948_/D _7258_/RN _6948_/CLK _6948_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_168_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _6879_/D input75/Z _6879_/CLK _6879_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold680 _5577_/Z _6941_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold691 _6716_/Q hold691/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_77_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__13 net413_60/I _7212_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_76 net413_76/I _7149_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_65 net413_65/I _7160_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_54 net413_54/I _7171_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__24 net413_80/I _7201_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__46 _4073__46/I _7179_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_98 net413_99/I _7127_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__35 net413_74/I _7190_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet413_87 net413_89/I _7138_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput207 _3371_/ZN mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput218 _7317_/Z mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput229 _7327_/Z mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_127_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4230_ hold356/Z _4102_/Z _4244_/S _4230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4161_ _4161_/A1 hold32/Z _4163_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_68_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _4092_/I _4092_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6802_ _6802_/D _6818_/CLK _6802_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4994_ _5083_/C _4997_/C _4546_/Z _4422_/Z _4994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6733_ _6733_/D _6624_/Z _7305_/CLK _6733_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3945_ _7174_/Q _3945_/A2 _3945_/B1 _7086_/Q _6682_/Q _3945_/C2 _3949_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_189_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _6664_/D _6619_/Z _7304_/CLK _6664_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_17_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ hold65/Z hold69/Z _5619_/S hold70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3876_ _3873_/Z _3876_/A2 _3876_/A3 _3876_/A4 _3876_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6595_ _6595_/A1 _4313_/Z _6595_/B _6596_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_20_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5546_ hold12/Z hold584/Z _5547_/S _5546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5477_ _5352_/Z _5390_/Z _5437_/Z _5476_/Z _5477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_155_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4428_ _4427_/Z _4402_/B _4373_/Z _4428_/B2 _5337_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_133_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7216_ _7216_/D _7237_/RN _7216_/CLK _7216_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_105_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7305_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7147_ hold59/Z _7260_/RN _7147_/CLK hold58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4359_ _4359_/A1 hold32/Z _4361_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_48_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7078_ _7078_/D _7008_/RN _7078_/CLK _7078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_24_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _7103_/Q _5967_/Z _5969_/Z _7119_/Q _6030_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_46_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_151 _4073__9/I _7074_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_140 net413_76/I _7085_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3730_ _7071_/Q _3943_/A2 _3945_/B1 _7089_/Q _3757_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_1992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3661_ _7057_/Q _5701_/A1 _3925_/A2 input8/Z _3663_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6380_ _6380_/A1 _6380_/A2 _6380_/A3 _6380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5400_ _5400_/A1 _5400_/A2 _5399_/Z _4729_/Z _5401_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3592_ _3592_/A1 _3592_/A2 _3592_/A3 _3592_/A4 _3592_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5331_ _5331_/I _5482_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5262_ _5340_/A1 _5262_/A2 _5328_/A2 _5442_/A4 _5262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ hold63/Z _7260_/RN _7001_/CLK hold62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5193_ _5193_/A1 _5193_/A2 _5437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ hold719/Z _4103_/I _4225_/S _4213_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4144_ hold867/Z _4103_/I _4145_/S _4144_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4075_ input83/Z _4075_/I1 _7299_/Q _4075_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _5262_/A2 _5343_/A2 _4495_/Z _4497_/Z _4977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_149_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6716_ _6716_/D _7170_/RN _6716_/CLK _6716_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_165_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3928_ _6940_/Q _5575_/A1 _3928_/B1 _6789_/Q _3928_/C1 _6822_/Q _3929_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6647_ _7235_/RN _6653_/A2 _6647_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3859_ _6933_/Q _3910_/A2 _3959_/B1 _6667_/Q _3925_/A2 input35/Z _3860_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6578_ _6578_/A1 _6578_/A2 _6602_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_165_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ hold32/Z hold587/Z _6901_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_118_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_302 net763_418/I _6923_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_324 net663_324/I _6901_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_313 net663_317/I _6912_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_335 net413_91/I _6890_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_346 net813_455/I _6879_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _5343_/B _5255_/A2 _4900_/B _5341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5880_ hold48/Z hold384/Z _5883_/S _5880_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _5214_/A2 _5420_/A1 _5223_/A2 _5291_/C _5276_/A1 _4840_/B1 _4834_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4762_ _5420_/A2 _5270_/A1 _4761_/I _3401_/I _4762_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_187_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6501_ _6555_/C _7257_/Q _6501_/B _6502_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4693_ _5099_/A1 _5099_/A2 _5097_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3713_ _3713_/I _3714_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6432_ _6432_/A1 _6239_/Z _6433_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3644_ _7010_/Q _3934_/A2 _3916_/A2 _7156_/Q _3645_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3575_ _7067_/Q _3927_/B1 _3592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6363_ _6554_/A1 _6363_/A2 _6363_/A3 _6363_/A4 _6363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5314_ _5314_/A1 _5314_/A2 _5314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_6294_ _7142_/Q _6292_/Z _6293_/Z _7150_/Q _6295_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5245_ _4421_/Z _4510_/Z _4666_/Z _4703_/Z _5245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold17 hold17/I hold17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold28 hold28/I hold28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5176_ _5175_/Z _4313_/Z _5184_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold39 hold39/I hold39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_110_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4127_ hold2/Z hold168/Z _4127_/S _4127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4058_ _6755_/Q input67/Z _7302_/Q _4058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_254 net613_254/I _6971_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_265 net813_463/I _6960_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_298 net613_298/I _6927_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_287 net613_287/I _6938_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_276 net413_84/I _6949_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold509 _6982_/Q hold509/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3360_ _6701_/Q _3360_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5030_ _5471_/B2 _5376_/B2 _5002_/Z _5353_/A1 _5202_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_112_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ _6981_/D _7008_/RN _6981_/CLK _6981_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_20_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ _5932_/I _7231_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5863_ hold20/Z hold502/Z _5865_/S _5863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4814_ _5414_/A2 _5287_/B _4876_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5794_ _3507_/Z _3552_/Z _5520_/C _5802_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_166_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _4700_/Z _5230_/B _4747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4676_ _4675_/Z _4501_/B _4472_/B _4524_/Z _4892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_179_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3627_ _7002_/Q _5638_/A1 _3959_/B1 _6672_/Q input32/Z _3927_/C2 _3630_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6415_ _7048_/Q _6241_/Z _6251_/Z _6984_/Q _6268_/Z _6952_/Q _6417_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3558_ _3515_/Z _3552_/Z _3916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6346_ _7096_/Q _6250_/Z _6302_/Z _7088_/Q _6292_/Z _7144_/Q _6357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_163_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput118 wb_adr_i[30] _4035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput107 wb_adr_i[20] _4483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_131_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ _6261_/Z _6265_/Z _6268_/Z _6269_/Z _6277_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_44__1359_ net663_324/I net413_69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3489_ _3489_/I _3653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
Xclkbuf_leaf_124__1359_ net613_261/I _4073__19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput129 wb_dat_i[10] _6585_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5228_ _5287_/C _5302_/B _4784_/Z _5228_/B _5479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5159_ _4422_/Z _4568_/Z _4641_/Z _4483_/B _5160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_56_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4530_ _4530_/I _4860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold306 _6939_/Q hold306/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4461_ _5281_/C _4481_/A2 _4469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold317 _5753_/Z _7097_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3412_ _3451_/I0 _7292_/Q _7293_/Q _3412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_171_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7180_ _7180_/D _7237_/RN _7180_/CLK _7180_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold328 _5655_/Z _7011_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold339 _6991_/Q hold339/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6200_ _6843_/Q _5971_/Z _5981_/Z _6787_/Q _6005_/Z _6849_/Q _6201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4392_ _4385_/Z _4387_/Z _4390_/Z _4392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_113_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _6703_/Q _5965_/Z _5967_/Z _7107_/Q _7171_/Q _6006_/Z _6133_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_112_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _7136_/Q _6051_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold1006 _7295_/Q _3438_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_100_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6062_ _6053_/Z _6061_/Z _6364_/B1 _6168_/C _6555_/C _6063_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _5347_/A1 _5012_/Z _5347_/A4 _5192_/B _5013_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _6964_/D _7008_/RN _6964_/CLK _6964_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5915_ _5945_/A1 _6745_/Q _5941_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6895_ _6895_/D _7260_/RN _6895_/CLK _6895_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5846_ hold12/Z hold474/Z _5847_/S _5846_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ hold227/Z hold406/Z _5784_/S _5777_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4728_ _4765_/A1 _5302_/B _5099_/A2 _4728_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_162_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4659_ _5281_/C _4436_/B _4472_/B _4501_/B _4659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_107_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold873 _6856_/Q hold873/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_66_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold840 _5512_/Z _6890_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold851 _6989_/Q hold851/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold862 _4351_/Z _6851_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6329_ _6329_/A1 _6329_/A2 _6322_/Z _6328_/Z _6329_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold884 _4160_/Z _6707_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold895 _6810_/Q hold895/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90__1359_ net413_62/I net763_423/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3953_/Z _3958_/Z _3961_/A3 _3961_/A4 _3961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_189_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5700_ hold2/Z hold225/Z hold25/Z _7051_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6680_ _6680_/D _7008_/RN _6680_/CLK _6680_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3892_ _7111_/Q _3917_/A2 _3950_/B1 _6725_/Q _3894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ hold291/Z hold851/Z _5637_/S _5631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ hold48/Z hold286/Z _5565_/S _5562_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _7301_/D _6653_/Z _7305_/CLK _7301_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4513_ _4421_/Z _4506_/Z _5180_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7232_ _7232_/D _7237_/RN _4067_/I1 _7232_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold114 _5874_/Z _7205_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5493_ hold291/Z hold879/Z _5493_/S _5493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold125 _6881_/Q hold125/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold103 _6955_/Q hold103/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4444_ _5288_/B _4472_/B _4868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold136 _5856_/Z _7189_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold158 _5545_/Z _6913_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold147 _6936_/Q hold147/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4375_ _3401_/I _3402_/I _5170_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold169 _4127_/Z _6681_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7163_ _7163_/D _7258_/RN _7163_/CLK _7163_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3326_ _7233_/Q _6282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_101_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7094_ _7094_/D _7218_/RN _7094_/CLK _7094_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ hold71/I _5958_/Z _5969_/Z hold76/I _6133_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_101_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _7088_/Q _6002_/Z _6048_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ hold3/Z _7260_/RN _6947_/CLK _6947_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6878_ _6878_/D _7170_/RN _6878_/CLK _6878_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5829_ hold2/Z hold133/Z _5829_/S _5829_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold670 _7058_/Q hold670/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold681 _6785_/Q hold681/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold692 _4174_/Z _6716_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_77 net413_77/I _7148_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet413_66 net413_66/I _7159_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__14 _4073__15/I _7211_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_55 net413_55/I _7170_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__36 net413_97/I _7189_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_99 net413_99/I _7126_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__25 _4073__25/I _7200_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__47 _4073__47/I _7178_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_88 net413_88/I _7137_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput208 _3370_/ZN mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput219 _7318_/Z mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ hold291/Z hold883/Z _4160_/S _4160_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _7300_/Q _7170_/RN _4092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _6801_/D _7265_/CLK _6801_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4993_ _4993_/A1 _4988_/Z _4993_/A3 _4999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_51_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6732_ _6732_/D _6623_/Z _7304_/CLK _6732_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3944_ _3944_/A1 _3944_/A2 _3944_/A3 _3944_/A4 _3944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6663_ _6663_/D _6618_/Z _7305_/CLK _6663_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3875_ _7053_/Q _5701_/A1 _4188_/A1 _6727_/Q _3914_/B1 _6877_/Q _3876_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ hold91/Z hold556/Z _5619_/S _5614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _6834_/Q _6594_/A2 _6594_/B1 _6835_/Q _6836_/Q _6594_/C2 _6595_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_158_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5545_ hold20/Z hold157/Z _5547_/S _5545_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _5476_/A1 _5476_/A2 _5475_/Z _5151_/B _5476_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_117_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4427_ _4374_/Z _4427_/A2 _4427_/A3 _4481_/A1 _4427_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_144_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7215_ _7215_/D _7218_/RN _7215_/CLK _7215_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7146_ _7146_/D _7238_/RN _7146_/CLK _7146_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4358_ hold291/Z hold873/Z _4358_/S _4358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3309_ hold4/Z hold5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_87_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _4289_/A1 hold32/Z _4291_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_7077_ _7077_/D input75/Z _7077_/CLK _7077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6028_ _7151_/Q _5960_/Z _5965_/Z _6699_/Q _6030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_58_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_141 net413_69/I _7084_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet463_130 net413_66/I _7095_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ hold84/I _3910_/A2 _5575_/A1 hold35/I _3663_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3591_ hold9/I _3951_/A2 _3954_/B1 input28/Z _3959_/B1 _6673_/Q _3592_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5330_ _4936_/I _5246_/Z _5445_/B2 _5330_/B2 _5330_/C _5331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_154_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _5261_/I _5264_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4212_ _4227_/S _4194_/Z _6652_/A2 _3519_/Z hold32/Z _4228_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_7000_ _7000_/D _7260_/RN _7000_/CLK _7000_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5192_ _5438_/C _4547_/Z _5192_/B _5192_/C _5193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_68_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ _4143_/A1 hold32/Z _4145_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_83_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4074_ input84/Z input67/Z _7300_/Q _4074_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4976_ _4421_/Z _5263_/A2 _5324_/A1 _5263_/A4 _5337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_52_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6715_ _6715_/D _7170_/RN _6715_/CLK _6715_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3927_ _6698_/Q _3927_/A2 _3927_/B1 _7060_/Q input4/Z _3927_/C2 _3929_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6646_ _7235_/RN _6653_/A2 _6646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3858_ _6699_/Q _3927_/A2 _3902_/A2 _6890_/Q input15/Z _3927_/C2 _3860_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6577_ _6834_/Q _6607_/A2 _6605_/A2 _6835_/Q _6577_/C _6578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3789_ _7006_/Q _3934_/A2 _5528_/S _6897_/Q _3790_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5528_ hold586/Z _4102_/Z _5528_/S _5528_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_14_0__1359_ clkbuf_0__1359_/Z net663_324/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_173_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5459_ _5459_/A1 _5098_/B _5098_/C _5458_/Z _5460_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_105_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7129_ _7129_/D _7237_/RN _7129_/CLK _7129_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8__1359_ net763_436/I net813_475/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_303 net763_415/I _6922_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_314 net663_317/I _6911_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_325 net713_394/I _6900_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_336 net413_91/I _6889_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_347 net813_455/I _6878_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _5287_/B _4586_/Z _4840_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_73_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4761_ _4761_/I _5071_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6500_ _6493_/Z _6499_/Z _6500_/B1 _6286_/Z _6555_/C _6501_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4692_ _4735_/A2 _4764_/A3 _4692_/B _4692_/C _5099_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_53_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3712_ hold88/I _3954_/A2 _3954_/B1 input24/Z _3713_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_14_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6431_ _7131_/Q _6484_/A2 _6533_/A3 _7115_/Q _6432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3643_ _6688_/Q _3945_/C2 _3941_/A2 _7164_/Q _3645_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _6942_/Q _6245_/Z _6273_/Z _6974_/Q _7120_/Q _6288_/Z _6363_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_155_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5313_ _5313_/A1 _5313_/A2 _5313_/A3 _5312_/Z _5314_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3574_ _3521_/Z _3537_/Z _3927_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_154_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6293_ _7235_/Q _7234_/Q _6302_/A3 _6484_/A3 _6293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5244_ _5324_/A1 _5324_/A2 _5324_/C _5250_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_114_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _5175_/A1 _5380_/C _5175_/A3 _5175_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_111_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold29 hold29/I hold29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold18 hold18/I hold18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_96_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4126_ hold12/Z hold258/Z _4127_/S _4126_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4057_ _6756_/Q _4072_/B2 _7301_/Q _4057_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _4959_/A1 _4959_/A2 _4957_/Z _4958_/Z _4963_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_147__1359_ net763_436/I net763_427/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6629_ _7170_/RN _6652_/A2 _6629_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_153_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_255 net613_255/I _6970_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet613_299 net413_57/I _6926_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_266 net613_266/I _6959_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_277 net413_91/I _6948_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_288 net613_288/I _6937_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _6980_/D _7008_/RN _6980_/CLK _6980_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5931_ _5931_/I0 _7231_/Q _5931_/S _5932_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5862_ hold48/Z hold329/Z _5865_/S _5862_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ hold2/Z hold123/Z _5793_/S _5793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4813_ _4422_/Z _4997_/C _4554_/Z _4483_/B _5167_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4744_ _5302_/B _4501_/B _4786_/A2 _5099_/A1 _5230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_175_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4675_ _4424_/B _4026_/B _4026_/C _4402_/B _4675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_135_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3626_ _7188_/Q _3959_/C1 _3923_/C1 _7084_/Q _3951_/C1 _7148_/Q _3646_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6414_ _7008_/Q _6243_/Z _6273_/Z _6976_/Q _6414_/C _6417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3557_ _3523_/Z _3529_/Z _5665_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6345_ _6345_/I _6347_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6276_ _6235_/Z _6237_/Z _6243_/Z _6266_/Z _6276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_102_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput108 wb_adr_i[21] _4402_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3488_ _3487_/Z _6862_/Q hold54/Z _3489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_115_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _5227_/I _5228_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput119 wb_adr_i[31] _4035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _5293_/A1 _5293_/B _5161_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ hold64/Z _7273_/Q hold54/Z hold65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5089_ _4506_/Z _4666_/Z _5341_/C _5265_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_99_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_50__1359_ net413_93/I net413_96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_130__1359_ net513_165/I net463_147/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_183_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold307 _5574_/Z _6939_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4460_ _4454_/Z _4367_/Z _4460_/B _4736_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4391_ _4391_/A1 _4391_/A2 _4391_/A3 _4391_/A4 _4481_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3411_ _7293_/Q _7292_/Q _4042_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_172_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold318 _6861_/Q _3307_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold329 _7194_/Q hold329/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3342_ _7251_/Q _6310_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6130_ hold84/I _5981_/Z _5984_/Z _7115_/Q _6134_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6061_ _6057_/Z _6061_/A2 _6061_/A3 _6061_/A4 _6061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _5350_/A1 _5192_/C _5009_/Z _4576_/C _5012_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold1007 _6731_/Q _3312_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ hold8/Z _7260_/RN _6963_/CLK _6963_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_146_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _6745_/Q _5913_/I _7227_/Q _7227_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6894_ _6894_/D _7170_/RN _6894_/CLK _7307_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5845_ hold20/Z hold498/Z _5847_/S _5845_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5776_ _3521_/Z _3552_/Z _5520_/C _5784_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_148_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4727_ _4727_/A1 _5223_/C _4727_/A3 _5090_/A1 _4733_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_174_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ _4887_/A1 _5315_/A2 _5172_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_4_2_0__1359_ clkbuf_0__1359_/Z clkbuf_4_2_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3609_ _7294_/Q _6732_/Q _3899_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xinput90 spimemio_flash_io2_oeb input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold830 _5733_/Z _7079_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4589_ _4835_/A2 _4454_/Z _5364_/B _4456_/B _4589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_107_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold841 _6706_/Q hold841/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold863 _6722_/Q hold863/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold852 _5631_/Z _6989_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold885 _7099_/Q hold885/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold874 _4358_/Z _6856_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6328_ _6328_/A1 _6328_/A2 _6328_/A3 _6328_/A4 _6328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold896 _4303_/Z _6810_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6259_ _6259_/A1 _6259_/A2 _6259_/A3 _6259_/A4 _6259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_153_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ _7206_/Q _3960_/A2 _3960_/B1 _6718_/Q _3960_/C _3961_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_44_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _6949_/Q _5584_/A1 _3954_/B1 input21/Z _5575_/A1 _6941_/Q _3894_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5630_ hold227/Z hold396/Z _5637_/S _5630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5561_ hold65/Z hold933/Z _5565_/S _5561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4512_ _4421_/Z _4452_/Z _5043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_145_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5492_ _4103_/I hold821/Z _5493_/S _5492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7300_ _7300_/D _6652_/Z _4075_/I1 _7300_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold115 _7067_/Q hold115/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7231_ _7231_/D _7256_/RN _7258_/CLK _7231_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_105_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold126 _5501_/Z _6881_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold104 _5592_/Z _6955_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4443_ _5288_/B _4380_/Z _4580_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_176_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold137 _7093_/Q hold137/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold148 _5571_/Z _6936_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold159 _6984_/Q hold159/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4374_ _5288_/B _4853_/A1 _4884_/A1 _4374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_132_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7162_ _7162_/D _7170_/RN _7162_/CLK _7162_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3325_ _6745_/Q _5950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_112_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7093_ _7093_/D _7237_/RN _7093_/CLK _7093_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6113_ _7245_/Q _6113_/I1 _6558_/S _7245_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6044_ _6210_/A2 _7054_/Q _6048_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6946_ hold46/Z _7238_/RN _6946_/CLK hold45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_26_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _6877_/D _7170_/RN _6877_/CLK _6877_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_168_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5828_ hold12/Z hold484/Z _5829_/S _5828_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5759_ hold919/Z _4103_/I _5766_/S _5759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold671 _5708_/Z _7058_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold660 _7198_/Q hold660/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold682 _4272_/Z _6785_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold693 _6728_/Q hold693/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_76_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_56 net413_56/I _7169_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_67 net413_67/I _7158_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__37 net413_97/I _7188_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__48 _4073__8/I _7177_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__26 _4073__43/I _7199_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__15 _4073__15/I _7210_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_89 net413_89/I _7136_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_78 net413_78/I _7147_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput209 _4063_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_4_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _4097_/A1 _4686_/B _6827_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6800_ _6800_/D input75/Z _6800_/CLK _6800_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_36_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ _5337_/A2 _5130_/B2 _5368_/A1 _5083_/B _5415_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_56_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _6731_/D _6622_/Z _7304_/CLK _6731_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3943_ _7068_/Q _3943_/A2 _5728_/A1 _7076_/Q _4182_/A1 _6722_/Q _3944_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_189_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6662_ _6662_/D _6617_/Z _7304_/CLK _6662_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3874_ _6884_/Q _3912_/B1 _3934_/B1 _6846_/Q _6858_/Q _4359_/A1 _3876_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ hold291/Z hold995/Z _5619_/S _5613_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _6593_/I0 _7274_/Q _6602_/S _7274_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5544_ hold48/Z hold188/Z _5547_/S _5544_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5475_ _5438_/C _4604_/Z _5475_/A3 _4666_/Z _5475_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_173_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4426_ _4721_/A1 _4721_/A2 _5083_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_133_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7214_ _7214_/D _7218_/RN _7214_/CLK _7214_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_7145_ _7145_/D _7237_/RN _7145_/CLK _7145_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4357_ _4103_/I hold835/Z _4358_/S _4357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3308_ hold40/I _5431_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4288_ _6571_/I0 _6798_/Q _4288_/S _6798_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _7076_/D input75/Z _7076_/CLK _7076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_104_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ _6949_/Q _5958_/Z _5994_/I _7135_/Q _6027_/C _6030_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_120 _4073__22/I _7105_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_131 net413_67/I _7094_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_142 net513_200/I _7083_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _6929_/D _7260_/RN _6929_/CLK _6929_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold490 _7056_/Q hold490/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3590_ _7019_/Q _5656_/A1 _3925_/A2 input10/Z _5665_/A1 _7027_/Q _3592_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_142_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5260_ _4700_/Z _4982_/Z _5260_/B _5261_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_126_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4211_ _4210_/Z hold801/Z _4211_/S _4211_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5191_ _4600_/Z _5190_/Z _5191_/A3 _5191_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_123_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4142_ hold291/Z hold881/Z _4142_/S _4142_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4975_ _4975_/A1 _4975_/A2 _4975_/A3 _4979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_177_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3926_ _3926_/A1 _3926_/A2 _3926_/A3 _3926_/A4 _3926_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6714_ _6714_/D _7170_/RN _6714_/CLK _6714_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6645_ _7235_/RN _6653_/A2 _6645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3857_ _6838_/Q _3923_/B1 _3960_/B1 _6719_/Q _3860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6576_ _6832_/Q _6608_/I1 _6606_/A2 _6836_/Q _6578_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3788_ _7104_/Q _5758_/A1 _3947_/A2 _7096_/Q _3941_/B1 _7168_/Q _3790_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_30_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _6900_/Q hold291/Z hold17/Z _5527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _4539_/I _4683_/Z _5302_/B _4460_/B _5458_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4409_ _4407_/Z _4390_/Z _4485_/A2 _5385_/A1 _4412_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5389_ _5389_/A1 _5389_/A2 _5389_/B _5389_/C _5390_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_114_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7128_ _7128_/D _7237_/RN _7128_/CLK _7128_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_119_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_107__1359_ net613_261/I net813_463/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7059_ _7059_/D _7237_/RN _7059_/CLK _7059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_8_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_315 net663_317/I _6910_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_304 _4073__22/I _6921_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_326 net763_425/I _6899_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_348 net813_455/I _6877_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_337 net813_483/I _6888_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4760_ _5324_/A1 _4436_/B _4495_/Z _4759_/Z _4761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4691_ _4786_/A2 _4692_/B _4692_/C _4691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_53_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3711_ _7016_/Q _5656_/A1 _3924_/A2 _6968_/Q _3927_/A2 _6702_/Q _3715_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3642_ _3642_/A1 _3642_/A2 _3642_/A3 _3642_/A4 _3642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6430_ _7203_/Q _6272_/Z _6275_/Z _7041_/Q _6293_/Z hold82/I _6434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6361_ _7046_/Q _6241_/Z _6251_/Z _6982_/Q _6268_/Z _6950_/Q _6363_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_60_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _5312_/A1 _5312_/A2 _5376_/B2 _5312_/A4 _5312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3573_ _3523_/Z _3552_/Z _3951_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_170_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6292_ _7235_/Q _7234_/Q _6484_/A3 _6533_/A3 _6292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5243_ _5243_/A1 _4890_/I _5324_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold19 hold19/I hold19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5174_ _5392_/B _4893_/Z _4991_/C _5175_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_111_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ hold20/Z hold263/Z _4127_/S _4125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ _6757_/Q input58/Z _7302_/Q _4056_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _5258_/B2 _5442_/A2 _5248_/A2 _4958_/A4 _4958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_61_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4889_ _4997_/C _4700_/Z _4890_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3909_ _7190_/Q _3909_/A2 _3915_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6628_ _7170_/RN _6652_/A2 _6628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _6833_/D _6830_/Q _6826_/Q _6833_/Q _6559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_118_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_256 net613_256/I _6969_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_267 _4073__15/I _6958_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_289 net813_492/I _6936_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_278 net613_279/I _6947_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10__1359_ clkbuf_4_2_0__1359_/Z net413_56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_73__1359_ net513_167/I net563_239/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5930_ _5924_/Z _6210_/A2 _6201_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5861_ hold65/Z hold325/Z _5865_/S _5861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5792_ hold12/Z hold717/Z _5793_/S _5792_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4812_ _4812_/A1 _4812_/A2 _5179_/B _4812_/B _5000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_61_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4743_ _4743_/A1 _4740_/Z _4741_/Z _5111_/C _4747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4674_ _4424_/B _4422_/Z _5172_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6413_ _6413_/I _6414_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3625_ _3625_/A1 _3625_/A2 _3625_/A3 _3866_/B _3625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3556_ _3525_/Z _3529_/Z _5701_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6344_ _7062_/Q _6257_/Z _6299_/Z _7054_/Q _6345_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_142_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6275_ _7235_/Q _7234_/Q _6484_/A2 _6533_/A2 _6275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_88_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput109 wb_adr_i[22] _4026_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3487_ _6658_/Q _7305_/Q _6733_/Q _3487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5226_ _4716_/Z _5310_/A2 _5226_/B _5226_/C _5227_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_69_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5157_ _5157_/A1 _5423_/A1 _5161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5088_ _5340_/C _5417_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ hold91/Z hold298/Z _4118_/S _4108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4039_ _6730_/Q _3464_/Z _6734_/Q _4040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_112_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold308 _7149_/Q hold308/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4390_ _4391_/A1 _4391_/A2 _4391_/A3 _4391_/A4 _4390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3410_ _6732_/Q _3409_/Z _3991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_125_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold319 hold319/I hold319/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3341_ _6925_/Q _6336_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_3_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _6974_/Q _5964_/Z _5984_/Z _7112_/Q _6061_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1008 _7294_/Q _3433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5011_ _5389_/C _5011_/A2 _5002_/Z _5194_/B1 _5350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6962_ _6962_/D _7256_/RN _6962_/CLK _6962_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_93_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5913_ _5913_/I _5952_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6893_ _6893_/D _7170_/RN _6893_/CLK _6893_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ hold48/Z hold527/Z _5847_/S _5844_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5775_ hold2/Z hold131/Z _5775_/S _5775_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4726_ _4703_/Z _5222_/A1 _5090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_163_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4657_ _4657_/A1 _4654_/Z _4657_/A3 _4656_/Z _4664_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_135_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold820 _4203_/Z _6738_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput91 spimemio_flash_io3_do input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3608_ _3589_/Z _3596_/Z _3607_/Z _6571_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xinput80 spi_sck input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xnet513_200 net513_200/I _7025_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4588_ _4546_/Z _5364_/B _5205_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_150_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold831 _6708_/Q hold831/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6327_ _7021_/Q _6235_/Z _6262_/Z _6965_/Q _6327_/C _6328_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold842 _4159_/Z _6706_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold853 _6822_/Q hold853/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold864 _4183_/Z _6722_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold886 _5755_/Z _7099_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3539_ _3509_/Z _3525_/Z _3954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold897 _6823_/Q hold897/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold875 _7076_/Q hold875/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_88_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6258_ _7206_/Q _6256_/Z _6257_/Z _7060_/Q _6259_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5209_ _5438_/B _4397_/Z _5209_/A3 _4666_/Z _5209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_131_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _6690_/Q _5985_/Z _5999_/Z _6847_/Q _6822_/Q _5964_/Z _6193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_57_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _7135_/Q _3951_/A2 _3924_/B1 _6821_/Q _3951_/C1 _7143_/Q _3895_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_43_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ hold91/Z hold442/Z _5565_/S _5560_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4511_ _5129_/A3 _5343_/B _4835_/A2 _3402_/I _4511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5491_ _3485_/Z _5857_/A2 hold235/Z _5520_/C _5493_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4442_ _4380_/Z _4579_/A2 _4607_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold116 _5718_/Z _7067_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7230_ _7230_/D _7256_/RN _7260_/CLK _7230_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold105 _7146_/Q hold105/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold127 _7059_/Q hold127/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold138 _5748_/Z _7093_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold149 _6766_/Q hold149/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4373_ _4501_/B _5288_/C _4369_/Z _4373_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_125_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _7161_/D _7218_/RN _7161_/CLK _7161_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3324_ _6744_/Q _5957_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_7092_ _7092_/D _7237_/RN _7092_/CLK _7092_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6112_ _6555_/C _6109_/Z _6112_/A3 _6112_/B _6113_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_86_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _7022_/Q _6211_/A2 _6211_/B1 _6990_/Q _6051_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_152_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ hold36/Z _7238_/RN _6945_/CLK hold35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _6876_/D _7170_/RN _6876_/CLK _6876_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ hold20/Z hold651/Z _5829_/S _5827_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5758_ _5758_/A1 hold32/Z _5766_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_6_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4709_ _5459_/A1 _5098_/B _4705_/Z _4709_/A4 _4709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_136_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ hold365/Z hold20/Z _5691_/S _5689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold672 _6859_/Q _3305_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_78_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold661 _5867_/Z _7198_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold650 _5764_/Z _7107_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold694 _4192_/Z _6728_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold683 _6849_/Q hold683/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_68 net413_68/I _7157_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_57 net413_57/I _7168_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__16 _4073__8/I _7209_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__27 _4073__27/I _7198_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4073__38 net413_73/I _7187_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_79 net413_79/I _7146_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__49 _4073__49/I _7176_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6730_ _6730_/D _6621_/Z _7304_/CLK _6730_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4991_ _5340_/A1 _5370_/B _4991_/B _4991_/C _4993_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_1_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3942_ _3907_/Z _3942_/A2 _7036_/Q _5683_/A1 _3942_/C1 _6853_/Q _3944_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_44_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ _6661_/D _6616_/Z _7304_/CLK _6661_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_90_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3873_ _3873_/A1 _3873_/A2 _3873_/A3 _3873_/A4 _3873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6592_ _6592_/A1 _4313_/Z _6592_/B _6593_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_177_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5612_ hold227/Z hold633/Z _5619_/S _5612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5543_ hold65/Z hold176/Z _5547_/S _5543_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5474_ hold5/I _5299_/C _5466_/Z _5473_/Z _5474_/C _6864_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_132_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4425_ _4483_/B _4373_/Z _4485_/A2 _4390_/Z _4721_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7213_ _7213_/D _7256_/RN _7213_/CLK _7213_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_132_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4356_ _3485_/Z hold674/Z _5520_/C _4358_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7144_ _7144_/D _7258_/RN _7144_/CLK _7144_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3307_ _3307_/I hold319/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _7075_/D _7235_/RN _7075_/CLK _7075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_140_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4287_ _6570_/I0 _6797_/Q _4288_/S _6797_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6026_ _6026_/A1 _6026_/A2 _6026_/A3 _6026_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_55_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_110 net463_110/I _7115_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_132 net413_69/I _7093_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_121 _4073__15/I _7104_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_143 net613_262/I _7082_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _6928_/D _7256_/RN _6928_/CLK _6928_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6859_ _6859_/D _7279_/RN _7278_/CLK _6859_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold480 _7186_/Q hold480/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold491 _5706_/Z _7056_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4210_ hold214/Z hold2/Z _4210_/S _4210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5190_ _5464_/A1 _5190_/A2 _5438_/C _5435_/A2 _5190_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_141_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ _4103_/I hold837/Z _4142_/S _4141_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4072_ hold54/I _4072_/A2 _4072_/B1 _4072_/B2 _4072_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_84_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4974_ _5359_/A1 _4973_/Z _4975_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3925_ input34/Z _3925_/A2 _3925_/B1 _6824_/Q _6839_/Q _3925_/C2 _3926_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6713_ _6713_/D input75/Z _6713_/CLK _6713_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6644_ _7235_/RN _6657_/A2 _6644_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _7013_/Q _5656_/A1 _5638_/A1 _6997_/Q _5665_/A1 _7021_/Q _3860_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6575_ _6575_/A1 _6575_/A2 _6606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3787_ _7192_/Q _3909_/A2 _4210_/S input45/Z _4227_/S input58/Z _3795_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_30_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5526_ _6899_/Q hold12/Z hold17/Z hold18/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ _5457_/A1 _5457_/A2 _5316_/Z _5457_/A4 _5457_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4408_ _4719_/A2 _4489_/A1 _4428_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5388_ _5388_/A1 _5202_/Z _5354_/Z _5388_/A4 _5388_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_120_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7127_ _7127_/D _7237_/RN _7127_/CLK _7127_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4339_ _4103_/I hold711/Z _4340_/S _4339_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _7058_/D _7256_/RN _7058_/CLK _7058_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _6009_/A1 _6009_/A2 _6009_/A3 _6008_/Z _6010_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_28_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_305 net763_415/I _6920_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_316 net763_406/I _6909_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet663_349 net813_455/I _6876_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_338 net813_487/I _6887_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_327 net763_425/I _6898_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ _6976_/Q _3923_/A2 _3910_/A2 _6936_/Q _3956_/A2 _7122_/Q _3715_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4690_ _4736_/A1 _4736_/A3 _4690_/B _4690_/C _5099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xclkbuf_leaf_33__1359_ clkbuf_4_10_0__1359_/Z _4073__8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3641_ _6704_/Q _3927_/A2 _3924_/A2 _6970_/Q _3642_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_128_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3572_ _3529_/Z _3542_/Z _3952_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6360_ _6966_/Q _6262_/Z _6269_/Z _7030_/Q _6360_/C _6363_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xclkbuf_leaf_113__1359_ net513_165/I net413_91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_96__1359_ clkbuf_4_5_0__1359_/Z net613_256/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5311_ _5308_/Z _5479_/A3 _5318_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ _7190_/Q _6285_/Z _6290_/Z _7078_/Q _6307_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ _4812_/B _5242_/A2 _5242_/A3 _4810_/B _5242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5173_ _4424_/B _4422_/Z _5269_/A2 _4997_/C _5173_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_102_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ hold48/Z hold418/Z _4127_/S _4124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4055_ _6766_/Q input81/Z _4055_/S _4055_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ _5389_/A2 _5442_/A2 _5248_/A2 _4958_/A4 _4957_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4888_ _5263_/A2 _4700_/Z _5445_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3908_ _5821_/A3 _3533_/Z hold235/I _3942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_137_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3839_ _3485_/Z _3680_/Z _3922_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6627_ _7170_/RN _6652_/A2 _6627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_118_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6558_ _7260_/Q _6558_/I1 _6558_/S _7260_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6489_ _6489_/I _6490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ hold392/Z hold20/Z _5509_/S _5509_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_268 net613_268/I _6957_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet613_279 net613_279/I _6946_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_257 net813_463/I _6968_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5860_ hold91/Z hold614/Z _5865_/S _5860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _5094_/C _5312_/A2 _5137_/B1 _5220_/B2 _5179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_179_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5791_ hold20/Z hold200/Z _5793_/S _5791_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4742_ _5302_/B _4695_/Z _4703_/Z _5226_/C _5111_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4673_ _5420_/A3 _5129_/A3 _5051_/S _3402_/I _4673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3624_ _7058_/Q _5701_/A1 _5674_/A1 _7034_/Q _3952_/A2 _7050_/Q _3625_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6412_ hold93/I _6235_/Z _6265_/Z _7000_/Q _6288_/Z _7122_/Q _6413_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_179_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ _7080_/Q _6290_/Z _6357_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3555_ _3507_/Z _3552_/Z _3951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3486_ _7305_/Q _6733_/Q _3987_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_143_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6274_ _7234_/Q _6282_/A1 _6302_/A3 _5943_/S _6274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_89_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _4728_/Z _5310_/A2 _5225_/B _5310_/C _5229_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_116_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _5356_/A1 _5403_/B2 _5156_/B _5423_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4107_ hold90/Z _7272_/Q hold54/Z hold91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5087_ _5087_/A1 _4982_/Z _5340_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _4038_/A1 _6561_/B2 _6826_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_112_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5989_ _7142_/Q _5987_/Z _5988_/Z _6980_/Q _6009_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_178_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 _3352_/ZN mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_2_0__1359_ clkbuf_4_10_0__1359_/Z clkbuf_opt_2_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold309 _5811_/Z _7149_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _4421_/Z _5438_/C _5435_/A2 _4606_/Z _5192_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_113_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1009 _7282_/Q _3466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_94_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ hold87/Z _7260_/RN _6961_/CLK hold86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _6743_/Q _6745_/Q _5913_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_59_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6892_ _6892_/D _7238_/RN _6892_/CLK _6892_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ hold65/Z hold558/Z _5847_/S _5843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5774_ hold12/Z hold456/Z _5775_/S _5774_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4725_ _4510_/Z _5325_/B _4727_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ _5420_/A3 _4374_/Z _5165_/A4 _5209_/A3 _4656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4587_ _4454_/Z _5269_/A2 _5364_/B _4586_/Z _4587_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold810 _4241_/Z _6760_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3607_ _3601_/Z _3607_/A2 _3606_/Z _3607_/A4 _3607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput70 mgmt_gpio_in[7] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold821 _6866_/Q hold821/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_66_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_201 net413_78/I _7024_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput81 spi_sdo input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput92 spimemio_flash_io3_oeb input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3538_ _3505_/Z _3537_/Z _3943_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold832 _4162_/Z _6708_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6326_ _7079_/Q _6290_/Z _6302_/Z _7087_/Q _6326_/C _6328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold854 _4324_/Z _6822_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold843 _7119_/Q hold843/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_88_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold898 _4325_/Z _6823_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold865 _6712_/Q hold865/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold887 _6847_/Q hold887/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold876 _5729_/Z _7076_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3469_ _3991_/A1 _3469_/A2 _7280_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6257_ _6484_/A3 _6282_/A2 _7232_/Q _6452_/A4 _6257_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_107_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _5206_/Z _4662_/B _5433_/A1 _5208_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_88_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6188_ _6857_/Q _5924_/Z _6201_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5139_ _4376_/Z _5139_/A2 _5139_/A3 _5291_/C _5139_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_123_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _5490_/A1 _5299_/C _5466_/Z _5489_/Z _5490_/C _6865_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_129_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _5420_/A2 _4456_/B _5051_/S _3401_/I _4510_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_89_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4441_ _5420_/A3 _5315_/A1 _4884_/A1 _4441_/B _4579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_145_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold117 _7075_/Q hold117/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold106 _5808_/Z _7146_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold128 _5709_/Z _7059_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7160_ _7160_/D _7256_/RN _7160_/CLK _7160_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold139 _7170_/Q hold139/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4372_ _4853_/A1 _4884_/A1 _4759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6111_ _6555_/C _7244_/Q _6112_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_98_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3323_ _6832_/Q _4096_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _7091_/D _7258_/RN _7091_/CLK _7091_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_85_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6042_ _7168_/Q _6006_/Z _6053_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6944_ _6944_/D _7238_/RN _6944_/CLK _6944_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6875_ _6875_/D _6633_/Z _4075_/I1 _6875_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_33_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5826_ hold48/Z hold348/Z _5829_/S _5826_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5757_ hold2/Z hold314/Z _5757_/S _5757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _4708_/A1 _5312_/A2 _5312_/A1 _5094_/C _4709_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5688_ hold369/Z hold48/Z _5691_/S _5688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4639_ _4639_/A1 _5039_/A4 _4638_/Z _4644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_135_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold640 _5741_/Z _7086_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold662 _6710_/Q hold662/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold651 _7163_/Q hold651/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7289_ _7289_/D _6643_/Z _4072_/B2 hold11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6309_ _6554_/A1 _6924_/Q _6310_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold673 _3500_/Z hold673/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold695 _6787_/Q hold695/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold684 _4348_/Z _6849_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_134_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_58 net413_74/I _7167_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__17 _4073__9/I _7208_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__28 _4073__5/I _7197_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_69 net413_69/I _7156_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__39 _4073__39/I _7186_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _4551_/Z _4892_/B _4991_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_90_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ _7158_/Q _3941_/A2 _3941_/B1 _7166_/Q _3941_/C _3944_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6660_ _6660_/D _6615_/Z _7304_/CLK _6660_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_177_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3872_ _6675_/Q _3546_/Z _3945_/C2 _6683_/Q _3873_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6591_ _6834_/Q _6591_/A2 _6591_/B1 _6835_/Q _6836_/Q _6591_/C2 _6592_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_158_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5611_ _3509_/Z hold24/Z _5821_/A3 _5857_/A3 _5619_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_31_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5542_ hold91/Z hold178/Z _5547_/S _5542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5473_ _5469_/Z _5489_/A2 _5472_/Z _5473_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_117_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4424_ _4374_/Z _4489_/A1 _4424_/B _4721_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_172_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7212_ _7212_/D _7237_/RN _7212_/CLK _7212_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4355_ hold291/Z hold735/Z _4355_/S _4355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7143_ _7143_/D _7008_/RN _7143_/CLK _7143_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3306_ _6860_/Q _5185_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7074_ _7074_/D _7237_/RN _7074_/CLK _7074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_58_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _6569_/I0 _6796_/Q _4288_/S _6796_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6025_ _7053_/Q _5924_/Z _6002_/Z _7087_/Q _6168_/C _6026_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_133 net413_77/I _7092_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_111 net413_99/I _7114_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_122 net813_473/I _7103_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_144 net663_322/I _7081_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _6927_/D _7237_/RN _6927_/CLK _6927_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_50_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6858_ _6858_/D _7170_/RN _6858_/CLK _6858_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5809_ hold20/Z hold58/Z _5811_/S hold59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6789_ _6789_/D _7008_/RN _6789_/CLK _6789_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_129_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold481 _5853_/Z _7186_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_8_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold470 _6879_/Q hold470/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold492 _7048_/Q hold492/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_77_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4140_ _3485_/Z _5857_/A2 _5513_/A3 _5520_/C _4142_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_150_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4071_ _3994_/Z hold54/I _4072_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_136__1359_ clkbuf_4_1_0__1359_/Z net813_483/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4973_ _5324_/A1 _5263_/A4 _4718_/B _5072_/A4 _4973_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_51_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _6712_/D input75/Z _6712_/CLK _6712_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3924_ _6964_/Q _3924_/A2 _3924_/B1 _6820_/Q _3926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6643_ _7235_/RN _6657_/A2 _6643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3855_ _3855_/A1 _3855_/A2 _3855_/A3 _3855_/A4 _3855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6574_ _6575_/A2 _6574_/A2 _6605_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_118_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3786_ _3786_/A1 _3786_/A2 _3786_/A3 _3786_/A4 _3786_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_106_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5525_ hold39/Z hold20/Z hold17/Z _6898_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5456_ _5456_/A1 _5456_/A2 _5456_/B _5457_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4407_ _4402_/B _4483_/B _4407_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_145_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5387_ _5387_/A1 _5387_/A2 _5387_/B _5388_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_132_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7126_ _7126_/D _7218_/RN _7126_/CLK _7126_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4338_ _3529_/Z _5520_/C hold235/Z _5857_/A2 _4340_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_115_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4269_ hold111/Z hold12/Z _4270_/S _4269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7057_ _7057_/D _7258_/RN _7057_/CLK _7057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6008_ _6008_/A1 _6008_/A2 _6008_/A3 _6008_/A4 _6008_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_46_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_306 net763_415/I _6919_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet663_317 net663_317/I _6908_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet663_328 net713_394/I _6897_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_339 net813_487/I _6886_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _6962_/Q _3957_/A2 _3901_/A2 _6986_/Q _3642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_127_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ _3542_/Z _3552_/Z _3941_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _6484_/A3 _5943_/S _7234_/Q _6533_/A3 _6290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5310_ _4728_/Z _5310_/A2 _5310_/B _5310_/C _5479_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_6_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _5321_/A1 _5241_/A2 _5451_/B _5242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_69_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _5172_/A1 _5368_/A1 _5172_/B _5172_/C _5380_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_114_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ hold65/Z hold300/Z _4127_/S _4123_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4054_ _6764_/Q input78/Z _4055_/S _4054_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4956_ _5359_/A1 _4761_/I _4959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4887_ _4887_/A1 _5315_/A2 _4554_/Z _4675_/Z _4887_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3907_ _7300_/Q _7283_/Q _6893_/Q _3907_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_20_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3838_ _3485_/Z _3617_/Z _3920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6626_ _7170_/RN _6652_/A2 _6626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_153_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _6557_/I _6558_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3769_ _7038_/Q _5683_/A1 _5674_/A1 _7030_/Q _3912_/B1 _6885_/Q _3773_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5508_ hold552/Z hold48/Z _5509_/S _5508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6488_ _7149_/Q _6292_/Z _6300_/Z _7109_/Q _6489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _5439_/A1 _5468_/A1 _5439_/B1 _5439_/B2 _5439_/C _5440_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_126_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7109_ _7109_/D _7256_/RN _7109_/CLK _7109_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_258 net613_258/I _6967_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_269 net813_467/I _6956_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _4997_/C _4675_/Z _4683_/Z _4810_/B _4812_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_2280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5790_ hold48/Z hold216/Z _5793_/S _5790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4741_ _4510_/Z _5302_/B _4695_/Z _5226_/C _4741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _5269_/A2 _4530_/I _5291_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_174_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3623_ _7108_/Q _5758_/A1 _5683_/A1 _7042_/Q _6930_/Q _3935_/A2 _3625_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6411_ _6401_/Z _6408_/Z _6411_/A3 _6411_/A4 _6411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6342_ _7070_/Q _6484_/A2 _6484_/A3 _6452_/A4 _6348_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3554_ _3505_/Z _3552_/Z _3930_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_131_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6273_ _6484_/A2 _5943_/S _7234_/Q _6533_/A2 _6273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3485_ _3473_/Z hold6/Z hold41/Z _3484_/Z _3485_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_115_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5224_ _5224_/A1 _5224_/A2 _5401_/B _5400_/A2 _5225_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _5275_/B _5153_/Z _5157_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5086_ _5086_/A1 _5412_/A1 _5412_/A2 _5260_/B _5182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_110_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4106_ hold291/Z hold845/Z _4118_/S _4106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4037_ _4036_/I _6826_/Q _6561_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_71_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _7228_/Q _7227_/Q _6002_/A2 _6210_/A2 _5988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4939_ _4939_/A1 _5061_/B _4937_/Z _4938_/Z _4939_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_36_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _6608_/Z _6833_/Q _6830_/Q _4313_/Z _6610_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_123_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput180 _3361_/ZN mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput191 _3351_/ZN mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6960_ _6960_/D _7258_/RN _6960_/CLK _6960_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_38_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ _5911_/A1 _5901_/B _5911_/B _7226_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_98_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6891_ _6891_/D _7170_/RN _6891_/CLK _6891_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5842_ hold91/Z hold969/Z _5847_/S _5842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5773_ hold20/Z hold219/Z _5775_/S _5773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4724_ _5442_/A2 _4500_/Z _5072_/A4 _5248_/A2 _5325_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_166_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4655_ _5043_/A2 _5043_/B _4657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_148_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _5288_/B _5281_/C _4436_/B _4472_/B _4586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold811 _6917_/Q hold811/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput71 mgmt_gpio_in[8] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3606_ _3606_/A1 _3606_/A2 _3606_/A3 _3606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold800 _5514_/Z _6891_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput82 spi_sdoenb input82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_150_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3537_ _3477_/Z hold41/Z _3484_/Z _3473_/Z _3537_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold822 _5492_/Z _6866_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6325_ _6325_/I _6326_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold855 _6718_/Q hold855/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold833 _7135_/Q hold833/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold844 _5778_/Z _7119_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput93 trap _3339_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_171_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold866 _4168_/Z _6712_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold888 _4345_/Z _6847_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold877 _7296_/Q hold877/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3468_ _7295_/Q hold22/Z _3469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6256_ _6282_/A1 _5943_/S _7234_/Q _6533_/A3 _6256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold899 _6723_/Q hold899/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3399_ _3399_/I _6598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5207_ _4662_/B _5433_/A1 _5362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_130_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6187_ _6187_/A1 _5991_/Z _6192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5138_ _5138_/A1 _5287_/B _5148_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5069_ _4761_/I _5078_/A2 _5070_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4440_ _4436_/B _4648_/A1 _4472_/B _4604_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_176_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold107 _7064_/Q hold107/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_176_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold118 _5727_/Z _7075_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold129 _7213_/Q hold129/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_125_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _3402_/I _4456_/B _5051_/S _4460_/B _4497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_171_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ _6201_/A3 _6928_/Q _6112_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3322_ _6746_/Q _4005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_99_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7090_ _7090_/D _7258_/RN _7090_/CLK _7090_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _7242_/Q _6041_/I1 _6558_/S _7242_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ hold66/Z _7238_/RN _6943_/CLK _6943_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6874_ _6874_/D _6632_/Z _4075_/I1 _6874_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5825_ hold65/Z hold323/Z _5829_/S _5825_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ hold12/Z hold493/Z _5757_/S _5756_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ hold529/Z hold65/Z _5691_/S _5687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4707_ _5420_/A3 _5269_/A2 _4708_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4638_ _4436_/B _4638_/A2 _5356_/C _5356_/A1 _4638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_118_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold630 _5888_/Z _7217_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4569_ _5364_/B _4568_/Z _5356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_78_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold641 _7068_/Q hold641/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap360 _7008_/RN _7238_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold663 _4165_/Z _6710_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold652 _5827_/Z _7163_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7288_ _7288_/D _6642_/Z _4072_/B2 hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _6554_/A1 _6307_/Z _6271_/Z _6308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold674 _3560_/Z hold674/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold696 _4275_/Z _6787_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold685 _6714_/Q hold685/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6239_ _5943_/S _6285_/A2 _7237_/Q _7234_/Q _6239_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_94_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_59 net413_59/I _7166_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__29 _4073__46/I _7196_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__18 _4073__43/I _7207_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3940_ _3940_/I _3941_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_182_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _6697_/Q _4146_/A1 _3936_/B1 _6691_/Q _3873_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6590_ _6590_/I0 _7273_/Q _6602_/S _7273_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5610_ hold2/Z hold218/Z hold43/Z _6971_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ hold291/Z hold797/Z _5547_/S _5541_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_16__1359_ clkbuf_4_2_0__1359_/Z net413_59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5472_ _5472_/A1 _5472_/A2 _4841_/B _5472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_117_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79__1359_ net513_167/I net413_65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7211_ _7211_/D _7256_/RN _7211_/CLK _7211_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4423_ _4373_/Z _4385_/Z _4922_/A3 _4423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_160_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7142_ _7142_/D _7008_/RN _7142_/CLK _7142_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4354_ _4103_/I hold668/Z _4355_/S _4354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7073_ _7073_/D _7235_/RN _7073_/CLK _7073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3305_ _3305_/I _3500_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4285_ _6568_/I0 _6795_/Q _4288_/S _6795_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6024_ _6981_/Q _5988_/Z _6015_/Z _7005_/Q _6024_/C _6026_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_58_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_112 net413_96/I _7113_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_123 net413_59/I _7102_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_134 net513_153/I _7091_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_145 net613_262/I _7080_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _6926_/D _7256_/RN _6926_/CLK _6926_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6857_ _6857_/D _7170_/RN _6857_/CLK _6857_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_13_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5808_ hold48/Z hold105/Z _5811_/S _5808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6788_ _6788_/D _7170_/RN _6788_/CLK _6788_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5739_ hold2/Z hold310/Z _5739_/S _5739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold471 _5499_/Z _6879_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold460 _6968_/Q hold460/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold482 _6769_/Q hold482/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold493 _7100_/Q hold493/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7304_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _7240_/Q _6896_/Q _6900_/Q _4070_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_3__1359_ net763_436/I net763_449/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4972_ _4496_/Z _5262_/A2 _5323_/B _4495_/Z _4972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_17_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6711_ _6711_/D _7170_/RN _6711_/CLK _6711_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3923_ _6972_/Q _3923_/A2 _3923_/B1 _6837_/Q _3923_/C1 _7078_/Q _3926_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_189_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _7235_/RN _6657_/A2 _6642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3854_ _7191_/Q _3909_/A2 _4210_/S input44/Z _3854_/C _3855_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_177_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6573_ _6575_/A2 _6573_/A2 _6607_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3785_ _6934_/Q _3910_/A2 _3959_/C1 _7184_/Q _3785_/C _3786_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _6897_/Q hold91/Z hold17/Z hold92/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5455_ _5455_/I _5485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_106_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4406_ _4402_/B _4483_/B _4719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_160_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5386_ _5386_/A1 _5432_/A1 _5386_/A3 _5434_/A1 _5386_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_160_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7125_ _7125_/D _7258_/RN _7125_/CLK _7125_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_119_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4337_ hold291/Z hold765/Z _4337_/S _4337_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4268_ hold37/Z hold20/Z _4270_/S hold38/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7056_ _7056_/D _7256_/RN _7056_/CLK _7056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6007_ _7036_/Q _6005_/Z _6006_/Z _7166_/Q _6008_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4199_ _4198_/Z hold805/Z _4211_/S _4199_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _6909_/D _7218_/RN _6909_/CLK _7324_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62__1359_ net513_170/I net763_418/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_142__1359_ clkbuf_4_1_0__1359_/Z net413_75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold290 _7284_/Q hold290/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_49_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_307 net763_418/I _6918_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_329 net763_423/I _6896_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_318 net713_369/I _6907_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3570_ _3521_/Z _3552_/Z _3956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_161_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5240_ _5368_/A1 _5389_/A2 _5240_/B _5451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_115_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5171_ _5169_/Z _5170_/Z _5175_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4122_ hold91/Z hold304/Z _4127_/S _4122_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4053_ _6763_/Q input80/Z _4055_/S _4053_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _4419_/Z _4951_/Z _4955_/B _5068_/B _4959_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3906_ _3485_/Z _3578_/Z _3920_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _4880_/Z _4886_/A2 _4884_/Z _4885_/Z _4886_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _7235_/RN _6653_/A2 _6625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3837_ input47/Z _4227_/S _3855_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_165_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3768_ _3527_/Z _3540_/Z _5532_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6556_ _6555_/C _7259_/Q _6556_/B _6557_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_173_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5507_ hold427/Z hold65/Z _5509_/S _5507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6487_ _7101_/Q _6250_/Z _6299_/Z _7059_/Q _6995_/Q _6237_/Z _6492_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_105_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3699_ _6887_/Q _3912_/B1 _3916_/B1 _6882_/Q _3701_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_4_5_0__1359_ clkbuf_0__1359_/Z clkbuf_4_5_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_161_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ _4568_/Z _4666_/Z _5438_/B _5438_/C _5439_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xoutput340 _6818_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5369_ _5287_/B _5369_/A2 _5369_/B _5369_/C _5421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_59_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _7108_/D _7256_/RN _7108_/CLK _7108_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7039_ _7039_/D _7237_/RN _7039_/CLK _7039_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet613_259 net763_425/I _6966_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ _5302_/B _4695_/Z _4716_/Z _5226_/C _4740_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _4530_/I _5051_/S _5137_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_179_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3622_ _7180_/Q _3945_/A2 _3913_/A2 input18/Z _3941_/B1 _7172_/Q _3647_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6410_ _7146_/Q _6292_/Z _6300_/Z _7106_/Q hold95/I _6290_/Z _6411_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6341_ _6934_/Q _6263_/Z _6266_/Z _7014_/Q _6355_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_155_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _3525_/Z _3552_/Z _3945_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3484_ _4317_/A1 _3483_/Z _3484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_131_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _6300_/A2 _6285_/A2 _7237_/Q _6452_/A4 _6272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5223_ _5094_/B _5223_/A2 _5223_/B _5223_/C _5400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_88_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _4568_/Z _4624_/Z _5376_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4105_ hold290/Z hold362/Z hold54/Z _4105_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5085_ _4987_/Z _5085_/A2 _5260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4036_ _4036_/I _4045_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _7231_/Q _7230_/Q _7229_/Q _6210_/B _5987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_80_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4938_ _4998_/A2 _5389_/A2 _5056_/C _5442_/A2 _4938_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4869_ _4869_/A1 _4866_/Z _4867_/Z _4868_/Z _4872_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6608_ _6608_/I0 _6608_/I1 _6832_/Q _6608_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6539_ _6729_/Q _6247_/Z _6297_/Z _7077_/Q _6547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_133_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput170 _4089_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput181 _3360_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput192 _3350_/ZN mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5910_ _6746_/Q _4006_/Z _5910_/B _5910_/C _5911_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_35_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _6890_/D _7238_/RN _6890_/CLK _6890_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_146_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ hold291/Z hold991/Z _5847_/S _5841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ hold48/Z hold620/Z _5775_/S _5772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4723_ _4495_/Z _4436_/B _5248_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_187_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ _4467_/B _5315_/A2 _4589_/Z _4460_/B _4654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4585_ _4887_/A1 _5399_/A2 _5276_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold812 _5550_/Z _6917_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput72 mgmt_gpio_in[9] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold801 _7322_/I hold801/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3605_ _7085_/Q _3923_/C1 _3956_/A2 _7125_/Q _3606_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold823 _7317_/I hold823/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput83 spimemio_flash_clk input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6324_ _7143_/Q _6292_/Z _6300_/Z _7103_/Q _6325_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold834 _5796_/Z _7135_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold845 _6667_/Q hold845/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3536_ _3533_/Z _3535_/Z _3927_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput94 uart_enabled _4059_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6255_ _7134_/Q _6253_/Z _6254_/Z _7174_/Q _6259_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold856 _4177_/Z _6718_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold867 _6694_/Q hold867/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold889 _6799_/Q hold889/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold878 _6612_/Z _7296_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ _3467_/I _7282_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5206_ _5189_/Z _5203_/Z _5357_/A2 _5440_/A1 _5206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3398_ _3398_/I _6595_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6186_ _6845_/Q _6211_/A2 _6211_/B1 _6837_/Q _6187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5137_ _5276_/C _5137_/A2 _5137_/B1 _5279_/A2 _5370_/B _5138_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_84_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _4700_/Z _4761_/I _5068_/B _5334_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_42_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4019_ _4006_/Z _4019_/A2 _4014_/Z _4019_/B _6745_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_123_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold108 _5715_/Z _7064_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4370_ _3402_/I _4456_/B _5051_/S _4884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_176_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold119 _7221_/Q hold119/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3321_ _7226_/Q _5911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_99_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6040_ _6040_/I _6041_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6942_ _6942_/D _7238_/RN _6942_/CLK _6942_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xclkbuf_leaf_119__1359_ net613_261/I net563_217/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6873_ _6873_/D _6631_/Z _4075_/I1 _6873_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_179_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5824_ hold91/Z hold606/Z _5829_/S _5824_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5755_ hold20/Z hold885/Z _5757_/S _5755_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4706_ _4765_/A1 _4782_/A1 _5302_/B _5218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5686_ hold588/Z hold91/Z _5691_/S _5686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4637_ _4565_/Z _5293_/B _5039_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_148_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold620 _7114_/Q hold620/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4568_ _5129_/A3 _4835_/A2 _3401_/I _3402_/I _4568_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold653 _7182_/Q hold653/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold642 _5720_/Z _7068_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold631 _7004_/Q hold631/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap361 input75/Z _7008_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_2_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _4759_/A2 _4759_/A3 _4718_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_171_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7287_ _7287_/D _6641_/Z _4072_/B2 hold47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3519_ _3653_/A1 hold673/Z hold320/Z _3497_/I _3519_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_89_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _6307_/A1 _6307_/A2 _6307_/A3 _6306_/Z _6307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold697 _6949_/Q hold697/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold664 _6883_/Q hold664/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold675 _4341_/Z _4343_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold686 _4171_/Z _6714_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6238_ _7020_/Q _6235_/Z _6237_/Z _6988_/Q _6260_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6169_ _6169_/A1 _6169_/A2 _6169_/A3 _6169_/A4 _6169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__19 _4073__19/I _7206_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3870_ _7103_/Q _5758_/A1 _3947_/A2 _7095_/Q _3873_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_16_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ hold227/Z hold246/Z _5547_/S _5540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ _5471_/A1 _5291_/C _4555_/C _5471_/B2 _5472_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4422_ _4402_/B _4026_/B _4026_/C _4422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_145_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7210_ _7210_/D _7256_/RN _7210_/CLK _7210_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ hold10/Z _7238_/RN _7141_/CLK hold9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4353_ _3529_/Z _5520_/C hold235/Z _5821_/A3 _4355_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3304_ _6733_/Q _4041_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_4284_ _6567_/I0 _6794_/Q _4288_/S _6794_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7072_ _7072_/D _7258_/RN _7072_/CLK _7072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6023_ _6941_/Q _5972_/Z _6021_/Z _6997_/Q _6026_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_67_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_124 net613_287/I _7101_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_113 _4073__41/I _7112_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_102 net513_200/I _7123_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_135 net513_153/I _7090_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_146 net463_147/I _7079_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6925_ _6925_/D _7218_/RN _6925_/CLK _6925_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6856_ _6856_/D _7218_/RN _6856_/CLK _6856_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_167_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3999_ _3999_/I _6835_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5807_ hold65/Z hold533/Z _5811_/S _5807_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6787_ _6787_/D _7170_/RN _6787_/CLK _6787_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ hold12/Z hold211/Z _5739_/S _5738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ hold346/Z hold65/Z _5673_/S _5669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold472 _6878_/Q hold472/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold450 _6689_/Q hold450/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold461 _6960_/Q hold461/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold483 _4254_/Z _6769_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_145_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold494 _5756_/Z _7100_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22__1359_ _4073__7/I _4073__43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_102__1359_ clkbuf_4_5_0__1359_/Z net613_275/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_85__1359_ net513_167/I net413_81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4971_ _5464_/A1 _4905_/Z _4975_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _6855_/Q _3922_/A2 _3922_/B1 _6692_/Q _3922_/C _3963_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6710_ _6710_/D _7170_/RN _6710_/CLK _6710_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_32_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _7235_/RN _6657_/A2 _6641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3853_ _3853_/I _3854_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _6575_/A2 _6572_/A2 _6608_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_118_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _3784_/I _3785_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ hold408/Z hold65/Z hold17/Z _6896_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5454_ _5454_/A1 _5454_/A2 _5454_/A3 _5453_/Z _5455_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4405_ _4489_/B _4483_/B _4722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5385_ _5385_/A1 _5389_/C _5439_/B1 _5393_/A1 _5385_/C _5434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7124_ _7124_/D _7258_/RN _7124_/CLK _7124_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4336_ _4103_/I hold713/Z _4337_/S _4336_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7055_ _7055_/D _7256_/RN _7055_/CLK _7055_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4267_ _6781_/Q hold48/Z _4270_/S hold49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4198_ _6770_/Q hold291/Z _4210_/S _4198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6006_ _7231_/Q _7228_/Q _7227_/Q _6068_/A4 _6006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_28_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _6908_/D _7218_/RN _6908_/CLK _7323_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6839_ _6839_/D _7008_/RN _6839_/CLK _6839_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold280 _5636_/Z _6994_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_46_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold291 hold363/Z hold291/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_46_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_308 net763_418/I _6917_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_319 net813_470/I _6906_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _5172_/B _5170_/A2 _5170_/A3 _5172_/C _5170_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4121_ hold291/Z hold847/Z _4127_/S _4121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _4052_/I _4052_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _5464_/A1 _5324_/A1 _4759_/Z _5263_/A4 _5068_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_91_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3905_ _7307_/I _3904_/Z _3944_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_177_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _4887_/A1 _5315_/A2 _4551_/Z _4675_/Z _4885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _7235_/RN _6653_/A2 _6624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_119_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3836_ _3515_/Z _3533_/Z _3914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3767_ _6700_/Q _3927_/A2 _3786_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6555_ _6548_/Z _6554_/Z _6555_/B1 _6286_/Z _6555_/C _6556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ hold454/Z hold91/Z _5509_/S _5506_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6486_ _6486_/A1 _6486_/A2 _6486_/A3 _6486_/A4 _6486_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_106_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3698_ _7056_/Q _5701_/A1 _5674_/A1 _7032_/Q _3952_/A2 _7048_/Q _3701_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5437_ _5437_/A1 _5437_/A2 _5436_/Z _5437_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput330 _7265_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput341 _6801_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5368_ _5368_/A1 _5276_/C _5368_/B _5368_/C _5369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_120_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ _4318_/Z _6833_/Q _6832_/Q _4313_/Z _6819_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5299_ _5210_/Z _5396_/A1 _5267_/Z _5298_/Z _5299_/C _5300_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_7107_ _7107_/D _7256_/RN _7107_/CLK _7107_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_7038_ _7038_/D _7256_/RN _7038_/CLK _7038_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_101_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4670_ _4670_/A1 _4667_/Z _4669_/Z _4670_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_119_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3621_ hold45/I _5575_/A1 _3642_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_30_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3552_ _3473_/Z _3552_/A2 _3484_/Z _3477_/Z _3552_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6340_ _7176_/Q _6254_/Z _6355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_127_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3483_ _6662_/Q _6661_/Q _6733_/Q _3483_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6271_ _6260_/Z _6271_/A2 _6271_/A3 _6271_/A4 _6271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_170_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5222_ _5222_/A1 _5310_/A2 _5223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5153_ _5150_/Z _5487_/A2 _5153_/A3 _5289_/A3 _5153_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_111_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4104_ hold227/Z hold420/Z _4118_/S _4104_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5084_ _5359_/A1 _4982_/Z _5085_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4035_ _4034_/Z _4035_/A2 _4035_/A3 _4035_/A4 _4036_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_110_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _7110_/Q _5984_/Z _5985_/Z _7060_/Q _6009_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4937_ _4998_/A2 _5328_/A1 _5056_/C _5442_/A2 _4937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_24_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _4868_/A1 _4524_/Z _5287_/B _4683_/Z _4868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_20 _4250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _4900_/B _6607_/A2 _6610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3819_ _3552_/Z hold674/Z _4182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4799_ _4422_/Z _4534_/Z _4568_/Z _5312_/A1 _4799_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_118_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _6723_/Q _6292_/Z _6299_/Z _6858_/Q _6548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_4_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _7010_/Q _6243_/Z _6269_/Z _7034_/Q _6469_/C _6472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_134_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput182 _4064_/Z mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput193 _3377_/ZN mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput171 _4065_/Z mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_130_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ hold227/Z hold645/Z _5847_/S _5840_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5771_ hold65/Z hold525/Z _5775_/S _5771_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ _5083_/C _4722_/A2 _4923_/A2 _5083_/B _5324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_159_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4653_ _4653_/A1 _5040_/C _4653_/A3 _5041_/B _4657_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_147_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ _4584_/A1 _4584_/A2 _5349_/B _4591_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_174_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold802 _4211_/Z _6742_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3604_ _7149_/Q _3951_/C1 _5638_/A1 _7003_/Q _3606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput73 pad_flash_io0_di input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput95 wb_adr_i[0] _3401_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold824 _4201_/Z _6737_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput84 spimemio_flash_csb input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3535_ hold320/Z _3617_/A1 hold673/Z _3489_/I _3535_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold835 _6855_/Q hold835/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6323_ _7095_/Q _6250_/Z _6257_/Z _7061_/Q _6275_/Z _7037_/Q _6328_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold813 _6747_/Q hold813/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold846 _4106_/Z _6667_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3466_ _3465_/Z _3466_/A2 input58/Z _3430_/S _3467_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6254_ _7237_/Q _6533_/A3 _6452_/A4 _6285_/A2 _6254_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold879 _6867_/Q hold879/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold868 _4144_/Z _6694_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold857 _6964_/Q hold857/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5205_ _5205_/A1 _5468_/A1 _5205_/B1 _5356_/C _5205_/C _5440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_88_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3397_ _3397_/I _6592_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_69_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _7248_/Q _6185_/I1 _6558_/S _7248_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5136_ _5287_/C _4570_/Z _4598_/Z _4784_/Z _5374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_69_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _4951_/Z _5078_/A2 _5070_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_45_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ _6743_/Q _6901_/Q _4019_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_25_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5969_ _7231_/Q _6211_/B1 _6021_/A2 _7227_/Q _5969_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_12_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold109 _7330_/I hold109/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3320_ _7224_/Q _5954_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_153_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _6941_/D _7260_/RN _6941_/CLK _6941_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_19_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _6872_/D _6630_/Z _4075_/I1 _6872_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_5823_ hold291/Z hold947/Z _5829_/S _5823_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ hold48/Z hold519/Z _5757_/S _5754_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4705_ _5220_/B2 _4536_/Z _4491_/B _4705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5685_ hold977/Z hold291/Z _5691_/S _5685_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4636_ _4636_/A1 _5034_/B _4635_/Z _4639_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_148_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold610 _7050_/Q hold610/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold621 _5772_/Z _7114_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_162_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4567_ _5270_/A1 _4454_/Z _5389_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_104_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold654 _5849_/Z _7182_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold643 _7110_/Q hold643/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6306_ _6306_/A1 _6306_/A2 _6306_/A3 _6306_/A4 _6306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold632 _5648_/Z _7004_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7286_ _7286_/D _6640_/Z _4072_/B2 hold64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4498_ _4494_/Z _4496_/Z _4998_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3518_ _3617_/A1 _3501_/Z _5513_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold665 _5504_/Z _6883_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold676 _4342_/Z _6845_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold687 _6696_/Q hold687/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3449_ _7292_/Q _3449_/A2 _3450_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _7235_/Q _6533_/A2 _6533_/A3 _5942_/S _6237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold698 _5586_/Z _6949_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6168_ _7059_/Q _5924_/Z _6015_/Z _7011_/Q _6168_/C _6169_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_76_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _4773_/Z _4874_/C _5238_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6099_ hold99/I _5994_/I _6015_/Z _7008_/Q _6944_/Q _5972_/Z _6101_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_2837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_45__1359_ net663_324/I net413_60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_125__1359_ net613_261/I net563_221/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5470_ _5470_/A1 _5372_/Z _5470_/A3 _5489_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_9_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _5420_/A3 _5420_/A2 _4456_/B _5051_/S _4421_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_32_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7140_ hold53/Z _7260_/RN _7140_/CLK hold52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4352_ hold291/Z hold905/Z _4352_/S _4352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7071_ _7071_/D _7235_/RN _7071_/CLK _7071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3303_ hold54/Z _4317_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4283_ _6566_/I0 _6793_/Q _4288_/S _6793_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6022_ _7079_/Q _5996_/Z _6005_/Z _7037_/Q _6965_/Q _5979_/Z _6031_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_58_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_125 _4073__6/I _7100_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_114 net413_99/I _7111_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_103 net813_463/I _7122_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_136 net663_322/I _7089_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_147 net463_147/I _7078_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6924_ _6924_/D _7237_/RN _6924_/CLK _6924_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_81_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6855_ _6855_/D _7218_/RN _6855_/CLK _6855_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3998_ _6835_/Q _4097_/A1 _6829_/Q _3999_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5806_ hold91/Z hold602/Z _5811_/S _5806_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6786_ _6786_/D _7170_/RN _6786_/CLK _6786_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5737_ hold20/Z hold78/Z _5739_/S hold79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ hold165/Z hold91/Z _5673_/S _5668_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4619_ _4565_/Z _4614_/Z _5029_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_117_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5599_ hold20/Z hold86/Z hold7/Z hold87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold440 _7042_/Q hold440/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold451 _4136_/Z _6689_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold462 _7122_/Q hold462/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold484 _7164_/Q hold484/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7269_ _7269_/D _7269_/CLK _7269_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold473 _5498_/Z _6878_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold495 _7008_/Q hold495/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_77_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _4970_/A1 _4967_/Z _4968_/Z _4969_/Z _4975_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_189_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ _3921_/I _3922_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6640_ _7235_/RN _6657_/A2 _6640_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3852_ _7215_/Q _3912_/A2 _3922_/A2 _6856_/Q _3853_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_60_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6571_ _6571_/I0 _7269_/Q _6571_/S _7269_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3783_ _7022_/Q _5665_/A1 _3959_/B1 _6668_/Q _3923_/C1 _7080_/Q _3784_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_30_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5522_ hold413/Z hold48/Z hold17/Z _6895_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5453_ _5126_/I _5452_/Z _5129_/Z _5453_/A4 _5453_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4404_ _4424_/B _4402_/B _4922_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_172_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5384_ _6577_/C _5267_/Z _5382_/Z _5384_/B _6862_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_132_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4335_ _5520_/C _3529_/Z _5513_/A3 _5857_/A2 _4337_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7123_ hold77/Z _7260_/RN _7123_/CLK hold76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_119_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4266_ hold67/Z hold65/Z _4270_/S hold68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7054_ _7054_/D _7256_/RN _7054_/CLK _7054_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xclkbuf_leaf_91__1359_ net413_62/I net663_330/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _4196_/Z hold803/Z _4211_/S _4197_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6005_ _7230_/Q _7229_/Q _6117_/A4 _6210_/A2 _6005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_28_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6907_ _6907_/D _7170_/RN _6907_/CLK _6907_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _6838_/D _7008_/RN _6838_/CLK _6838_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6769_ _6769_/D _7256_/RN _6769_/CLK _6769_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold270 _4112_/Z _6670_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold281 _7018_/Q hold281/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_49_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold292 _5496_/Z _6877_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_120_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet663_309 net763_419/I _6916_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _4103_/I hold791/Z _4127_/S _4120_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4051_ _7201_/Q input82/Z _4055_/S _4052_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4953_ _4953_/A1 _5065_/B _4953_/A3 _4955_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_149_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3904_ _3489_/I _3904_/A2 hold320/Z _3904_/A4 _3904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_33_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6623_ _7235_/RN _6653_/A2 _6623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4884_ _4884_/A1 _4659_/Z _4675_/Z _3401_/I _4884_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3835_ _3485_/Z _3560_/Z _3922_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3766_ input26/Z _3927_/C2 _3794_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6554_ _6554_/A1 _6554_/A2 _6554_/A3 _6553_/Z _6554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6485_ _7117_/Q _6240_/Z _6297_/Z _6705_/Q _6485_/C _6486_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5505_ hold771/Z hold291/Z _5509_/S _5505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5436_ _4576_/C _5472_/A2 _5009_/Z _5435_/Z _5436_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3697_ _6944_/Q _5575_/A1 _3707_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput331 _7266_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput342 _6802_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput320 _6793_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5367_ _4568_/Z _4586_/Z _5368_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_120_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4318_ _4316_/Z _4318_/A2 _6833_/D _6828_/Q _4318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5298_ _5296_/Z _5382_/A3 _5173_/Z _5464_/B _5298_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7106_ _7106_/D _7256_/RN _7106_/CLK _7106_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4249_ hold91/Z hold182/Z _4252_/S _4249_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _7037_/D _7218_/RN _7037_/CLK _7037_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_74_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3620_ hold50/I _5584_/A1 _3630_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_128_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3551_ _3525_/Z _3537_/Z _3917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_183_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3482_ _4041_/B1 _6662_/Q _3975_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_115_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6270_ _6948_/Q _6268_/Z _6269_/Z _7028_/Q _6271_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_102_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ _5221_/I _5401_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_44_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5152_ _5364_/B _4614_/Z _4784_/Z _4624_/Z _4570_/Z _5153_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_97_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _4103_/I _5520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5083_ _4977_/Z _4981_/Z _5083_/B _5083_/C _5337_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_56_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ _4033_/Z _4034_/A2 _4388_/A2 _4388_/A1 _4034_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_38_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _7231_/Q _6210_/C _6021_/A2 _7227_/Q _5985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4936_ _4936_/I _5410_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_21_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _5269_/A2 _4530_/I _5287_/B _5293_/B _4867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_21 hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_10 _5505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6606_ _4686_/B _6606_/A2 _6610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3818_ _3535_/Z _3552_/Z _3960_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4798_ _4568_/Z _4793_/Z _5452_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6537_ _6717_/Q _6250_/Z _6290_/Z _6709_/Q _6302_/Z _6713_/Q _6548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3749_ _7129_/Q _3930_/A2 _5758_/A1 _7105_/Q _3941_/B1 _7169_/Q _3751_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_137_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _6468_/I _6469_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5419_ _5419_/A1 _5419_/A2 _5418_/Z _5431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6399_ _7218_/Q _6274_/Z _6285_/Z _7194_/Q _7178_/Q _6254_/Z _6401_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet713_390 net763_423/I _6784_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput194 _3349_/ZN mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput183 _3359_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput172 _3369_/ZN mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ hold91/Z hold604/Z _5775_/S _5770_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _4721_/A1 _4721_/A2 _4721_/B _5323_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_148_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4652_ _4436_/B _5139_/A2 _5471_/B2 _5281_/C _5041_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_30_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3603_ _7117_/Q _3917_/A2 _5758_/A1 _7109_/Q _5674_/A1 _7035_/Q _3606_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4583_ _4570_/Z _5016_/B2 _5349_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_163_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold803 _7315_/I hold803/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput96 wb_adr_i[10] input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput85 spimemio_flash_io0_do input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3534_ _3497_/I _3501_/Z hold235/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold825 _6902_/Q hold825/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6322_ _6322_/A1 _6322_/A2 _6322_/A3 _6322_/A4 _6322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold836 _4357_/Z _6855_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold814 _4214_/Z _6747_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput74 pad_flash_io1_di _3337_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3465_ _3464_/Z _3442_/B _3465_/A3 _3465_/A4 _3465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_143_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _7236_/Q _6300_/A2 _6533_/A4 _6302_/A4 _6253_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_107_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold847 _6675_/Q hold847/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold858 _5603_/Z _6964_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold869 _6697_/Q hold869/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5204_ _5346_/A2 _5387_/A1 _5403_/B2 _5205_/A1 _5204_/C _5357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_103_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9__1359_ clkbuf_4_2_0__1359_/Z net413_67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3396_ _3396_/I _6589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6184_ _6555_/C _6181_/Z _6184_/A3 _6184_/B _6185_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5135_ _4589_/Z _4817_/Z _5287_/C _5487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_97_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _4944_/Z _5078_/A2 _5066_/B _5481_/C _5070_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4017_ _4006_/Z _4019_/A2 _4020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _6014_/A2 _7229_/Q _6211_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4919_ _5343_/A1 _4496_/Z _5056_/C _5442_/A2 _4927_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5899_ _5910_/B _5899_/I1 _7223_/Q _7223_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_68__1359_ net513_175/I net763_419/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6940_ _6940_/D _7258_/RN _6940_/CLK _6940_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_75_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6871_ _6871_/D _6629_/Z _4075_/I1 _6871_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_179_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5822_ _4103_/I hold929/Z _5829_/S _5822_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ hold65/Z hold316/Z _5757_/S _5753_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4704_ _4687_/Z _4704_/A2 _5255_/A2 _5092_/A1 _5098_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_72_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5684_ hold927/Z _4103_/I _5691_/S _5684_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _4868_/A1 _4524_/Z _4546_/Z _5364_/B _4635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_136_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4566_ _4422_/Z _5278_/C _4554_/Z _4483_/B _4576_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_116_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold600 _6768_/Q hold600/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold611 _7044_/Q hold611/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap352 _5364_/B _5287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_143_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold622 _7209_/Q hold622/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3517_ _3489_/I _3492_/Z _5839_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold644 _5768_/Z _7110_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold633 _6972_/Q hold633/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6305_ _7198_/Q _6272_/Z _6275_/Z _7036_/Q _6306_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4497_ _4436_/B _4497_/A2 _4497_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_7285_ _7285_/D _6639_/Z _4072_/B2 hold90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold677 _7312_/I hold677/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold655 _7013_/Q hold655/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold666 _7060_/Q hold666/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold688 _4147_/Z _6696_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3448_ _3448_/I _7293_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6236_ _5943_/S _7234_/Q _6533_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_131_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold699 _6857_/Q hold699/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_134_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6167_ _6947_/Q _5972_/Z _6021_/Z _7003_/Q _6169_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _6929_/Q _6447_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5118_ _5115_/Z _5117_/Z _5118_/A3 _5215_/C _5118_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_94_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _7090_/Q _6002_/Z _6019_/Z _7048_/Q _6098_/C _6101_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5049_ _5049_/A1 _5210_/A4 _5180_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_72_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4420_ _5170_/A2 _4836_/A4 _5258_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4351_ _4103_/I hold861/Z _4352_/S _4351_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3302_ hold31/Z _6608_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7070_ _7070_/D _7235_/RN _7070_/CLK _7070_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_141_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4282_ _6565_/I0 _6792_/Q _4288_/S _6792_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ _6211_/B1 _6021_/A2 _6210_/A2 _7227_/Q _6021_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_95_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_104 _4073__49/I _7121_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_115 _4073__47/I _7110_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_126 _4073__49/I _7099_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_137 _4073__25/I _7088_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_148 _4073__3/I _7077_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6923_ _6923_/D _7256_/RN _6923_/CLK _6923_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6854_ _6854_/D _7170_/RN _6854_/CLK _6854_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3997_ _3997_/I _6834_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6785_ _6785_/D _7170_/RN _6785_/CLK _6785_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5805_ hold291/Z hold973/Z _5811_/S _5805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_131__1359_ net513_165/I net713_373/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5736_ hold48/Z hold95/Z _5739_/S hold96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ hold647/Z hold291/Z _5673_/S _5667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _4618_/A1 _5151_/B _4616_/Z _4617_/Z _4622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_135_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ hold48/Z hold461/Z hold7/Z _6960_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold452 _6771_/Q hold452/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4549_ _5288_/B _4467_/B _4460_/B _4472_/B _4549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_150_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold430 _5788_/Z _7128_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold441 _5690_/Z _7042_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold463 _5781_/Z _7122_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold485 _5828_/Z _7164_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold474 _7180_/Q hold474/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7268_ _7268_/D _7269_/CLK _7268_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold496 _5652_/Z _7008_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6219_ _6844_/Q _5971_/Z _5981_/Z _6788_/Q _6005_/Z _6850_/Q _6220_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_135_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7199_ _7199_/D _7218_/RN _7199_/CLK _7199_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_38_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ input71/Z _4244_/S _3920_/B1 _6866_/Q _6902_/Q _3920_/C2 _3921_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_17_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ _7159_/Q _3941_/A2 _3912_/C1 _6707_/Q _4170_/A1 _6715_/Q _3855_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_158_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6570_ _6570_/I0 _7268_/Q _6571_/S _7268_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3782_ _7014_/Q _5656_/A1 _5638_/A1 _6998_/Q _3951_/C1 _7144_/Q _3786_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_185_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5521_ hold16/Z _5521_/A2 hold55/I hold6/Z hold17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_74_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5452_ _4791_/Z _5452_/A2 _5452_/A3 _4801_/Z _5452_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4403_ _4424_/B _4402_/B _4923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5383_ _6862_/Q _6577_/C _5212_/Z _5320_/Z _5383_/C _5384_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_160_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7122_ _7122_/D _7258_/RN _7122_/CLK _7122_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4334_ hold291/Z hold738/Z _4334_/S _6840_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _7053_/D _7008_/RN _7053_/CLK _7053_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4265_ hold97/Z hold91/Z _4270_/S hold98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6004_ _7086_/Q _6002_/Z _6003_/Z _7158_/Q _6008_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4196_ hold482/Z _4102_/Z _4210_/S _4196_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _6906_/D _7170_/RN _6906_/CLK _6906_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6837_ _6837_/D _7008_/RN _6837_/CLK _6837_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_148_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _6768_/D _7218_/RN _6768_/CLK _6768_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5719_ _5857_/A2 _5857_/A3 _3537_/Z hold24/Z _5727_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6699_ _6699_/D _7258_/RN _6699_/CLK _6699_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_163_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold271 _6659_/Q hold271/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold260 _6671_/Q hold260/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold293 _6930_/Q hold293/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold282 _6669_/Q hold282/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_10_0__1359_ clkbuf_0__1359_/Z clkbuf_4_10_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_74_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4050_ _4050_/I0 input90/Z _4050_/S _4050_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _5359_/A1 _4951_/Z _4953_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_149_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4883_ _4881_/Z _4882_/Z _4886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3903_ _3903_/A1 _5821_/A3 _5513_/A3 _3533_/Z _3903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_32_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6622_ _7235_/RN _6653_/A2 _6622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3834_ _3485_/Z _3535_/Z _3956_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3765_ _7046_/Q _3952_/A2 _3916_/B1 _6880_/Q _3790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6553_ _6553_/A1 _6553_/A2 _6553_/A3 _6553_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_173_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6484_ _7133_/Q _6484_/A2 _6484_/A3 _6533_/A4 _6485_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_118_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5504_ hold664/Z _4103_/I _5509_/S _5504_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3696_ _7008_/Q _3934_/A2 _3701_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5435_ _5438_/C _5435_/A2 _5475_/A3 _4666_/Z _5435_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput310 _7261_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput332 _7267_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput321 _6794_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5366_ _5366_/A1 _5366_/A2 _5365_/Z _5469_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_114_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4317_ _4317_/A1 _6826_/Q _4318_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5297_ _4882_/Z _5170_/Z _5382_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7105_ _7105_/D _7237_/RN _7105_/CLK _7105_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7036_ _7036_/D _7218_/RN _7036_/CLK _7036_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4248_ hold291/Z hold743/Z _4252_/S _4248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4179_ _5821_/A3 hold235/Z _3537_/Z _5520_/C _4181_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_71_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet763_450 net413_63/I _6715_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3550_ _3485_/Z _3507_/Z _3955_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_182_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3481_ hold41/Z _3552_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_5220_ _4694_/Z _5310_/A2 _5220_/B1 _5220_/B2 _5221_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_142_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5151_ _5287_/C _5364_/B _4784_/Z _5151_/B _5487_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_96_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4102_ input58/Z hold226/Z hold54/Z _4102_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5082_ _4980_/Z _5081_/Z _5412_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4033_ _4028_/Z _4030_/Z _4026_/B _4026_/C _4033_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_99_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5984_ _5984_/A1 _6210_/B _7231_/Q _7230_/Q _5984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_36_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _5442_/A2 _4497_/Z _4495_/Z _5056_/C _4936_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_21_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4866_ _4868_/A1 _4524_/Z _5414_/A2 _5287_/B _4866_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_22 _7111_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_11 _5518_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ _4415_/B _6605_/A2 _6610_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4797_ _4791_/Z _5452_/A2 _5453_/A4 _4797_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3817_ _3527_/Z _3542_/Z _5536_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3748_ _6677_/Q _3546_/Z _3947_/A2 _7097_/Q _6896_/Q _5528_/S _3758_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6536_ _6691_/Q _6257_/Z _6275_/Z _6850_/Q _6300_/Z _6721_/Q _6548_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_137_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ _5857_/A2 _5513_/A3 _5503_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6467_ _7026_/Q _6235_/Z _6262_/Z _6970_/Q _6265_/Z _7002_/Q _6468_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_161_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _5418_/A1 _5418_/A2 _5417_/Z _5418_/A4 _5418_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6398_ _7098_/Q _6250_/Z _6302_/Z _7090_/Q _6401_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet713_380 net813_481/I _6810_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5349_ _5349_/A1 _5387_/A2 _5349_/B _5350_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput195 _3348_/ZN mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput173 _3368_/ZN mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput184 _3358_/ZN mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_391 net763_444/I _6783_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7019_ _7019_/D _7258_/RN _7019_/CLK _7019_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_46_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28__1359_ net613_298/I net763_430/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_79_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_108__1359_ clkbuf_4_5_0__1359_/Z net413_79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4720_ _5083_/C _5083_/B _5259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_159_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4651_ _4467_/B _4460_/B _4501_/B _4472_/B _4651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3602_ _7213_/Q _3960_/A2 _3955_/A2 _7205_/Q _6955_/Q _5584_/A1 _3607_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _4638_/A2 _5345_/A2 _4438_/B _4467_/B _5016_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput97 wb_adr_i[11] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold804 _4197_/Z _6735_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_115_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3533_ hold15/Z _3477_/Z hold41/Z _3484_/Z _3533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold815 _6748_/Q hold815/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput86 spimemio_flash_io0_oeb input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6321_ _7069_/Q _6248_/Z _6297_/Z _6699_/Q _6321_/C _6322_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold826 _5531_/Z _6902_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold837 _6692_/Q hold837/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput75 porb input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
X_3464_ _7283_/Q _6665_/Q _6664_/Q _6663_/Q _3464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold859 _6715_/Q hold859/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6252_ _7094_/Q _6250_/Z _6251_/Z _6980_/Q _6259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold848 _4121_/Z _6675_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5203_ _5199_/Z _5354_/A2 _5202_/Z _5203_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_103_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6183_ _6555_/C _7247_/Q _6184_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3395_ _3395_/I _6586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5134_ _5293_/A1 _4624_/Z _5275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5065_ _4699_/Z _5252_/B _5065_/B _5481_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_85_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _6744_/Q _5896_/I0 _4019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_72_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _7231_/Q _7228_/Q _7227_/Q _6002_/A2 _5967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_52_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _4927_/A1 _4927_/A2 _5444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_40_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ _5901_/B _5899_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ _4598_/Z _4681_/Z _4849_/B _5373_/B _4852_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_21_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6519_ _6716_/Q _6250_/Z _6293_/Z _6718_/Q _6521_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_4_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6870_ _6870_/D _6628_/Z _4075_/I1 _6870_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_179_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5821_ _5520_/C _3552_/Z _5821_/A3 _5857_/A3 _5829_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_34_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5752_ hold91/Z hold596/Z _5757_/S _5752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ _5420_/A2 _5129_/A3 _4835_/A2 _3401_/I _4703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_176_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5683_ _5683_/A1 hold32/Z _5691_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_30_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _4868_/A1 _4524_/Z _4551_/Z _5364_/B _5034_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_129_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4565_ _5364_/B _5051_/S _4456_/B _4454_/Z _4565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold612 _6935_/Q hold612/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold601 _4252_/Z _6768_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap353 _7237_/RN _7235_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_128_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold623 _5879_/Z _7209_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3516_ _3485_/Z _3515_/Z _3912_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold645 _7174_/Q hold645/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold634 _5612_/Z _6972_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6304_ _7166_/Q _5948_/Z _6273_/Z _6972_/Q _6306_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4496_ _4467_/B _4497_/A2 _4496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_7284_ _7284_/D _6638_/Z _4072_/B2 _7284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold678 _4228_/Z _6754_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold656 _6997_/Q hold656/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold667 _5711_/Z _7060_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3447_ _7293_/Q _3449_/A2 _3447_/B1 _7292_/Q _3448_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_6235_ _7235_/Q _7234_/Q _6533_/A2 _6533_/A3 _6235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold689 _6824_/Q hold689/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6166_ _6987_/Q _5988_/Z _6019_/Z _7051_/Q _6169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11__1359_ clkbuf_4_2_0__1359_/Z net413_64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3378_ _6928_/Q _6418_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5117_ _5117_/A1 _5117_/A2 _5117_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6097_ _6097_/I _6098_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5048_ _5395_/A1 _4991_/C _5210_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _6999_/D _7260_/RN _6999_/CLK _6999_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_185_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ _3485_/Z _3535_/Z _5520_/C _4352_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3301_ _6663_/Q _3971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_153_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4281_ _6564_/I0 _6791_/Q _4288_/S _6791_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6020_ _6933_/Q _5981_/Z _6019_/Z _7045_/Q _6037_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_140_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_116 net413_68/I _7109_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_105 net613_266/I _7120_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_127 _4073__47/I _7098_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_138 _4073__50/I _7087_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_149 _4073__3/I _7076_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6922_ _6922_/D _7256_/RN _6922_/CLK _6922_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ _6853_/D _7170_/RN _6853_/CLK _6853_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5804_ hold227/Z hold635/Z _5811_/S _5804_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3996_ _6834_/Q _4097_/A1 _6828_/Q _3997_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_149_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6784_ _6784_/D _7260_/RN _6784_/CLK _6784_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5735_ hold65/Z hold560/Z _5739_/S _5735_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5666_ hold231/Z hold227/Z _5673_/S _5666_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4617_ _4422_/Z _4546_/Z _4614_/Z _4483_/B _4617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_108_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5597_ hold65/Z hold426/Z hold7/Z _6959_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold420 _6666_/Q hold420/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold453 _4256_/Z _6771_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4548_ _4441_/B _5281_/C _4436_/B _4501_/B _4555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_104_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_8_0__1359_ clkbuf_0__1359_/Z net613_298/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold442 _6926_/Q hold442/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold431 _6980_/Q hold431/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_145_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold475 _5846_/Z _7180_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4479_ _4786_/A1 _4786_/A2 _4786_/A3 _5094_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold486 _7092_/Q hold486/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7267_ _7267_/D _7269_/CLK _7267_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold464 _6976_/Q hold464/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold497 _7032_/Q hold497/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6218_ _6790_/Q _5972_/Z _6021_/Z _6840_/Q _6220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_98_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7198_ _7198_/D _7218_/RN _7198_/CLK _7198_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_180_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6149_ _6986_/Q _5988_/Z _5996_/Z _7084_/Q _6152_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_79_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ _7069_/Q _3943_/A2 _4244_/S input72/Z _4161_/A1 _6709_/Q _3855_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3781_ _6974_/Q _3923_/A2 _3957_/A2 _6958_/Q _3956_/A2 _7120_/Q _3786_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_60_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5520_ hold321/Z _5520_/A2 _5520_/B _5520_/C hold322/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_185_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5451_ _4492_/Z _4536_/Z _5451_/B _5451_/C _5454_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_67_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4402_ _4580_/C _4489_/A1 _4402_/B _4412_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5382_ _5379_/Z _5464_/B _5382_/A3 _5382_/A4 _5382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_132_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7121_ _7121_/D _7218_/RN _7121_/CLK _7121_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4333_ hold227/Z _6839_/Q _4334_/S _4333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4264_ hold781/Z hold291/Z _4270_/S _4264_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7052_ _7052_/D _7008_/RN _7052_/CLK _7052_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6003_ _6015_/A3 _6211_/A2 _7231_/Q _7228_/Q _6003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4195_ _4210_/S _4194_/Z _6652_/A2 _3540_/Z hold32/Z _4211_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_95_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6905_ _6905_/D _7237_/RN _6905_/CLK _6905_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6836_ _6836_/D _7279_/RN _7279_/CLK _6836_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _6767_/D _7218_/RN _6767_/CLK _6767_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3979_ _3978_/Z _6661_/Q _3988_/S _6661_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5718_ hold2/Z hold115/Z _5718_/S _5718_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6698_ _6698_/D _7258_/RN _6698_/CLK _6698_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_164_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ hold891/Z hold291/Z _5655_/S _5649_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7319_ _7319_/I _7319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold261 _4114_/Z _6671_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold250 _6892_/Q hold250/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold272 _3476_/I hold272/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold294 _5564_/Z _6930_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold283 _4110_/Z _6669_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_46_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4951_ _4407_/Z _5259_/A1 _4759_/Z _5263_/A4 _4951_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_36_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4882_ _4367_/Z _4555_/B _5172_/B _5172_/C _4882_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_51_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3902_ _6889_/Q _3902_/A2 _3960_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_189_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ _7235_/RN _6653_/A2 _6621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3833_ _3529_/Z _3578_/Z _3936_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3764_ _6676_/Q _3546_/Z _3776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6552_ _6848_/Q _6269_/Z _6273_/Z _6823_/Q _6553_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6483_ _7205_/Q _6272_/Z _6296_/Z _7165_/Q _7067_/Q _6257_/Z _6486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5503_ hold16/Z _5503_/A2 hold32/Z hold6/Z _5509_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3695_ _7106_/Q _5758_/A1 _3719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5434_ _5434_/A1 _5434_/A2 _5432_/Z _5433_/Z _5441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xoutput300 _3990_/I serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_69_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput311 _6811_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput322 _6812_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput333 _6813_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5365_ _5468_/B1 _5288_/B _4441_/B _4363_/Z _5365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_113_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ _7104_/D _7256_/RN _7104_/CLK _7104_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4316_ _6830_/Q _6829_/Q _6831_/Q _4316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_141_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5296_ _5271_/Z _5296_/A2 _5295_/Z _5467_/B _5296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_101_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7035_ _7035_/D _7258_/RN _7035_/CLK _7035_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_75_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4247_ _4103_/I hold701/Z _4252_/S _4247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4178_ hold291/Z hold903/Z _4178_/S _4178_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6819_ _6819_/D _7279_/RN _7279_/CLK hold54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_24_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_440 net413_55/I _6725_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_451 net813_469/I _6714_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3480_ _3479_/Z hold40/Z hold54/I hold41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_127_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5150_ _5374_/A2 _5148_/Z _5374_/A1 _5487_/A1 _5150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5081_ _5340_/A1 _5262_/A2 _5343_/A2 _5442_/A4 _5081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ _3533_/Z _5520_/C hold235/Z _5839_/A3 _4118_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4032_ _4032_/A1 _4032_/A2 _4031_/Z _4035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_96_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5983_ _7231_/Q _5983_/A2 _5983_/B _5983_/C _6010_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4934_ _5464_/A1 _5325_/B _5061_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_178_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4865_ _4865_/A1 _4865_/A2 _5156_/B _4869_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_23 _7161_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_12 _5537_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6604_ _4316_/Z _6604_/A2 _6833_/D _6828_/Q _7278_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_123_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4796_ _4793_/Z _5394_/A2 _5453_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3816_ _3521_/Z _3527_/Z _3902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3747_ _3747_/A1 _3747_/A2 _3747_/A3 _3747_/A4 _3747_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6535_ _6856_/Q _6256_/Z _6546_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_21_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6466_ _6466_/A1 _6466_/A2 _6466_/A3 _6465_/Z _6466_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_106_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3678_ input31/Z _3927_/C2 _3951_/A2 hold73/I _3686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5417_ _5417_/A1 _5417_/A2 _5263_/Z _5417_/A4 _5417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_133_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6397_ _7186_/Q _6282_/Z _6299_/Z _7056_/Q hold88/I _6237_/Z _6401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet713_370 net713_385/I _6840_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_381 net813_453/I _6809_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5348_ _5348_/I _5437_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput174 _3367_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput185 _3357_/ZN mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet713_392 net713_394/I _6782_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput196 _3732_/A1 mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5279_ _5288_/A1 _5279_/A2 _4555_/C _5439_/A1 _5279_/C _5284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_88_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _7018_/D _7258_/RN _7018_/CLK _7018_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_47_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4650_ _4441_/B _5288_/B _5281_/C _4436_/B _4650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3601_ _3601_/A1 _3601_/A2 _3601_/A3 _3601_/A4 _3601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4581_ _4557_/Z _5435_/A2 _5349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6320_ _6320_/A1 _6239_/Z _6321_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput98 wb_adr_i[12] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_183_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput65 mgmt_gpio_in[36] _7333_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold805 _7316_/I hold805/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold827 _6756_/Q hold827/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput87 spimemio_flash_io1_do _7332_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold816 _4216_/Z _6748_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3532_ hold42/Z hold273/Z _3904_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput76 qspi_enabled _4050_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3463_ _7283_/Q _3462_/Z _3463_/S _7283_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6251_ _6300_/A2 _5943_/S _7234_/Q _6533_/A2 _6251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold838 _4141_/Z _6692_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold849 _6699_/Q hold849/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5202_ _4626_/Z _5201_/Z _5202_/A3 _5202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_131_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6182_ _6201_/A3 _6931_/Q _6184_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3394_ _3394_/I _6583_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5133_ _5165_/A2 _5287_/B _5288_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_57_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5064_ _5064_/A1 _5410_/B _5063_/I _5064_/A4 _5066_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _5957_/S _3990_/I _5953_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _6972_/Q _5964_/Z _5965_/Z _6698_/Q _5974_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4917_ _5328_/A1 _5056_/C _5442_/A2 _5442_/A4 _4927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5897_ _6744_/Q _3990_/I _5901_/A1 _5950_/A1 _5901_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_33_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4848_ _4853_/A1 _5414_/A2 _5287_/B _4501_/B _5373_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_34__1359_ clkbuf_4_10_0__1359_/Z net413_72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_114__1359_ net513_165/I net813_499/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4779_ _4700_/Z _4778_/Z _5456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_97__1359_ clkbuf_4_5_0__1359_/Z net763_425/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6518_ _6824_/Q _6251_/Z _6256_/Z _6855_/Q _6521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_10_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6449_ _6449_/I _6450_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5820_ hold2/Z hold141/Z _5820_/S _5820_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ hold291/Z hold953/Z _5757_/S _5751_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4702_ _4884_/A1 _3401_/I _5255_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5682_ hold204/Z hold2/Z hold33/Z _7035_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4633_ _4633_/A1 _5035_/A4 _5387_/B _4636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_175_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _4554_/Z _5364_/B _5439_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_116_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold602 _7144_/Q hold602/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap343 _6653_/A2 _6657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_7283_ _7283_/D _6637_/Z _7305_/CLK _7283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold613 _5570_/Z _6935_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3515_ _3653_/A1 _3492_/Z _3497_/I _3501_/Z _3515_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xmax_cap354 _7218_/RN _7237_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold624 _7052_/Q hold624/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6303_ _7214_/Q _6274_/Z _6302_/Z _7086_/Q _6306_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold635 _7142_/Q hold635/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4495_ _4460_/B _4884_/A1 _4495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_144_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6234_ _7233_/Q _7232_/Q _6533_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_131_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold646 _5840_/Z _7174_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold679 _6941_/Q hold679/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold657 _5640_/Z _6997_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold668 _6853_/Q hold668/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3446_ _3449_/A2 _3450_/A1 _3447_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_170_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6165_ _7019_/Q _5971_/Z _6005_/Z _7043_/Q _6169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_69_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3377_ _6943_/Q _3377_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5116_ _5117_/A1 _5117_/A2 _5316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _7146_/Q _5987_/Z _6003_/Z _7162_/Q _6097_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5047_ _5047_/A1 _5360_/B _5049_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6998_ _6998_/D _7260_/RN _6998_/CLK _6998_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_14_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ _6282_/A1 _5948_/Z _5950_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80__1359_ net513_167/I _4073__25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3300_ _6664_/Q _3465_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_126_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _6831_/Q _7279_/RN _4288_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_4_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_106 net713_373/I _7119_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_117 net413_60/I _7108_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_128 net413_64/I _7097_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_139 _4073__51/I _7086_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6921_ _6921_/D _7237_/RN _6921_/CLK _6921_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_94_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _6852_/D input75/Z _6852_/CLK _6852_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5803_ _3523_/Z _3552_/Z hold24/Z _5811_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_50_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3995_ _3994_/Z _3995_/A2 _4097_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6783_ _6783_/D _7170_/RN _6783_/CLK _6783_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5734_ hold91/Z hold194/Z _5739_/S _5734_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5665_ _5665_/A1 hold32/Z _5673_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_163_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4616_ _4422_/Z _4551_/Z _4614_/Z _4483_/B _4616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_117_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ hold91/Z hold539/Z hold7/Z _6958_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold410 _5643_/Z _7000_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _5278_/C _4878_/A2 _3401_/I _3402_/I _4547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_150_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold443 _5560_/Z _6926_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold454 _6885_/Q hold454/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold421 _4104_/Z _6666_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold432 _5621_/Z _6980_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold487 _5747_/Z _7092_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold476 _7196_/Q hold476/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4478_ _4786_/A2 _4786_/A3 _4782_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7266_ _7266_/D _7269_/CLK _7266_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold465 _5616_/Z _6976_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3429_ _3971_/A1 _6730_/Q _6665_/Q _6664_/Q _3430_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_132_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7197_ _7197_/D _7237_/RN _7197_/CLK _7197_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold498 _7179_/Q hold498/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6217_ _6217_/A1 _6217_/A2 _6217_/A3 _6217_/A4 _6217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6148_ _6970_/Q _5979_/Z _5999_/Z _7034_/Q _6152_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6079_ _7129_/Q _6000_/Z _6019_/Z _7047_/Q _6967_/Q _5979_/Z _6085_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_46_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3780_ _7208_/Q _3960_/A2 _3955_/A2 _7200_/Q _3796_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _5450_/I _5463_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ _4412_/A1 _4399_/Z _5083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_173_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5381_ _5381_/I _5382_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7120_ _7120_/D _7258_/RN _7120_/CLK _7120_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4332_ _3509_/Z _5839_/A3 hold235/Z _5520_/C _4332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7051_ _7051_/D _7256_/RN _7051_/CLK _7051_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4263_ hold719/Z _4103_/I _4270_/S _4263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6002_ _7231_/Q _6002_/A2 _6021_/A2 _7227_/Q _6002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4194_ _4194_/A1 _3994_/Z _4194_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_94_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6904_ _6904_/D _7237_/RN _6904_/CLK _6904_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_39_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6835_ _6835_/D _7279_/RN _7279_/CLK _6835_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_51_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3978_ _3977_/Z _6660_/Q _6733_/Q _3978_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6766_ _6766_/D _7170_/RN _6766_/CLK _6766_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5717_ hold12/Z hold170/Z _5718_/S _5717_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4072_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6697_ _6697_/D _7170_/RN _6697_/CLK _6697_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5648_ hold631/Z hold227/Z _5655_/S _5648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5579_ _6943_/Q hold65/Z _5583_/S hold66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7318_ _7318_/I _7318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold240 _7216_/Q hold240/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold251 _5516_/Z _6892_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold262 _7012_/Q hold262/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold273 _3477_/Z hold273/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold295 _6962_/Q hold295/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold284 _6880_/Q hold284/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7249_ _7249_/D _7260_/RN _7260_/CLK _7249_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_46_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4950_ _5442_/A2 _4495_/Z _4496_/Z _4958_/A4 _5252_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_91_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4881_ _5104_/A1 _4555_/B _4650_/Z _5172_/C _4881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3901_ _6980_/Q _3901_/A2 _3926_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_33_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6620_ _7235_/RN _6653_/A2 _6620_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3832_ _3519_/Z _3529_/Z _4359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6551_ _6790_/Q _6245_/Z _6288_/Z _7297_/Q _6553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3763_ input54/Z _4194_/A1 _3795_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_119_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5502_ hold422/Z hold48/Z _5502_/S _5502_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6482_ _7075_/Q _6248_/Z _6253_/Z hold9/I _7157_/Q _6293_/Z _6486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_9_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3694_ _7064_/Q _3927_/B1 _3715_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5433_ _5433_/A1 _5433_/A2 _5433_/A3 _4662_/B _5433_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput301 _3683_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5364_ _5414_/A2 _4551_/Z _5364_/B _5468_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_133_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput334 _7268_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput323 _6795_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput312 _6803_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _6834_/Q _6835_/Q _6836_/Q _6832_/Q _5299_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7103_ _7103_/D _7218_/RN _7103_/CLK _7103_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_0_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _5295_/A1 _4501_/B _4472_/B _5315_/A1 _5295_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_102_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7034_ _7034_/D _7258_/RN _7034_/CLK _7034_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4246_ _3485_/Z _5821_/A3 _5513_/A3 _5520_/C _4252_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_95_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4177_ _4103_/I hold855/Z _4178_/S _4177_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _6818_/D _6818_/CLK _6818_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_430 net763_430/I _6740_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6749_ _6749_/D _7238_/RN _6749_/CLK _7308_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet763_441 net763_449/I _6724_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_167_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5080_ _4977_/Z _4981_/Z _5083_/B _5080_/C _5412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4100_ hold22/Z hold31/Z hold54/Z hold55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_116_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4031_ _4031_/A1 _4031_/A2 _4031_/A3 _4031_/A4 _4031_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5982_ _6964_/Q _5979_/Z _5981_/Z _6932_/Q _5980_/Z _7068_/Q _5983_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4933_ _4933_/A1 _4930_/Z _4933_/A3 _4933_/A4 _4939_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_80_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_13 hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4864_ _4624_/Z _4844_/Z _5156_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_61_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _5299_/C _6833_/Q _6826_/Q _6603_/A4 _6604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4795_ _5328_/A1 _4699_/Z _5394_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_24 _7193_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3815_ _3552_/Z _3617_/Z _4188_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_146_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3746_ _7185_/Q _3959_/C1 _3901_/A2 _6983_/Q _3747_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6534_ _6727_/Q _6253_/Z _6296_/Z _6715_/Q _6542_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ _6465_/A1 _6465_/A2 _6465_/A3 _6464_/Z _6465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5416_ _5416_/I _5417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3677_ input49/Z _4210_/S _5521_/A2 _3904_/A2 _3947_/A2 _7099_/Q _3687_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_161_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_371 net813_489/I _6839_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6396_ _7064_/Q _6257_/Z _6408_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xnet713_360 net813_475/I _6850_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5347_ _5347_/A1 _5347_/A2 _5347_/A3 _5347_/A4 _5348_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xoutput175 _3366_/ZN mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput186 _3356_/ZN mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet713_382 net813_453/I _6800_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_393 net763_422/I _6781_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput197 _3346_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5278_ _4554_/Z _4683_/Z _5287_/B _5278_/C _5279_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_87_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4229_ _4244_/S _4194_/Z _6652_/A2 _3542_/Z hold32/Z _4245_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_102_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7017_ _7017_/D _7260_/RN _7017_/CLK _7017_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_leaf_57__1359_ net663_324/I net513_163/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_137__1359_ clkbuf_4_1_0__1359_/Z net813_453/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _4604_/A2 _4604_/A3 _4580_/B _4580_/C _5435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_128_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3600_ _7181_/Q _3945_/A2 _3945_/B1 _7093_/Q _3601_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3531_ _3505_/Z _3529_/Z _3934_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 mgmt_gpio_in[37] _7334_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold817 _6770_/Q hold817/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold806 _4199_/Z _6736_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold828 _4233_/Z _6756_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput88 spimemio_flash_io1_oeb input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput77 ser_tx input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput99 wb_adr_i[13] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3462_ _3465_/A3 _6665_/Q input58/Z _3462_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_143_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6250_ _7236_/Q _6484_/A2 _6311_/A3 _6302_/A4 _6250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold839 _6890_/Q hold839/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3393_ _3393_/I _6580_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5201_ _5464_/A1 _5438_/C _4557_/Z _4604_/Z _5201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6181_ _6169_/Z _6181_/A2 _6181_/A3 _6180_/Z _6181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_69_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5132_ _5205_/A1 _5132_/A2 _5293_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_97_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _5063_/I _5330_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4014_ _7237_/Q _6484_/A2 _6311_/A3 _6285_/A2 _4014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_92_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ _7231_/Q _7228_/Q _7227_/Q _6210_/C _5965_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_34_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4916_ _5324_/A1 _5263_/A4 _5056_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5896_ _5896_/I0 _6746_/Q _5957_/S _5910_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4847_ _4530_/I _5399_/A2 _5104_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_178_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4778_ _4468_/Z _4782_/A1 _5302_/B _4778_/A4 _4778_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3729_ _7201_/Q _3955_/A2 _3747_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6517_ _6706_/Q _6254_/Z _6273_/Z _6822_/Q _6521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _6744_/Q _7255_/Q _6448_/B _6449_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_106_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6379_ _7137_/Q _6253_/Z _6297_/Z _6701_/Q _6380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_121_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40__1359_ net413_93/I _4073__6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5750_ _4103_/I hold917/Z _5757_/S _5750_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4701_ _4687_/Z _5097_/A1 _4699_/Z _5092_/A1 _5459_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5681_ hold439/Z hold12/Z hold33/Z _7034_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4632_ _4441_/B _4501_/B _4460_/B _4436_/B _5293_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_30_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ _4402_/B _4483_/B _4026_/B _4026_/C _5364_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_128_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold603 _5806_/Z _7144_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4494_ _5281_/C _4884_/A1 _4494_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xmax_cap344 _4064_/S _6653_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7282_ _7282_/D _6636_/Z _7305_/CLK _7282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6302_ _7236_/Q _6311_/A3 _6302_/A3 _6302_/A4 _6302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold614 _7192_/Q hold614/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3514_ _6979_/Q _3923_/A2 _3592_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold625 _5702_/Z _7052_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold636 _5804_/Z _7142_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3445_ _3452_/S _7291_/Q _3450_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6233_ _7236_/Q _7237_/Q _6533_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold658 _6924_/Q hold658/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap355 _7170_/RN _7218_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold669 _4354_/Z _6853_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold647 _7021_/Q hold647/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_98_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6164_ _7027_/Q _6211_/A2 _6211_/B1 _6995_/Q _6176_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3376_ _6951_/Q _3376_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5115_ _5113_/Z _5403_/C _5233_/A1 _5156_/B _5115_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_85_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _6968_/Q _5979_/Z _5996_/Z hold95/I _6095_/C _6101_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5046_ _5044_/Z _5433_/A1 _5047_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_2819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6997_ _6997_/D _7260_/RN _6997_/CLK _6997_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _7235_/Q _7234_/Q _6300_/A2 _6484_/A3 _5948_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_129_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5879_ hold65/Z hold622/Z _5883_/S _5879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_107 net463_147/I _7118_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_129 net413_65/I _7096_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_118 net413_62/I _7107_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6920_ _6920_/D _7258_/RN _6920_/CLK _6920_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _6851_/D input75/Z _6851_/CLK _6851_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5802_ hold2/Z hold9/Z _5802_/S hold10/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3994_ _3994_/A1 _6902_/Q input67/Z _3994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6782_ hold38/Z _7238_/RN _6782_/CLK hold37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5733_ hold291/Z hold829/Z _5739_/S _5733_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5664_ hold213/Z hold2/Z hold56/Z _7019_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4615_ _4422_/Z _4568_/Z _4614_/Z _4483_/B _5151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5595_ hold291/Z hold988/Z hold7/Z _6957_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold411 _6920_/Q hold411/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_135_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4546_ _4835_/A2 _4456_/B _3402_/I _3401_/I _4546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_117_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7334_ _7334_/I _7334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold400 _7171_/Q hold400/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold444 _6938_/Q hold444/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold433 _7106_/Q hold433/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold422 _6882_/Q hold422/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold477 _5864_/Z _7196_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4477_ _4692_/B _4692_/C _4786_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_89_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7265_ _7265_/D _7265_/CLK _7265_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold455 _5506_/Z _6885_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold466 _6702_/Q hold466/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3428_ _3427_/Z _6734_/Q _3428_/A3 _3428_/B _7301_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xhold499 _5845_/Z _7179_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7196_ _7196_/D _7237_/RN _7196_/CLK _7196_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold488 _7148_/Q hold488/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6216_ _6723_/Q _5987_/Z _6015_/Z _6842_/Q _6217_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_48_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3359_ _7081_/Q _3359_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6147_ _6147_/A1 _6147_/A2 _6147_/A3 _6147_/A4 _6147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_58_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6078_ _6078_/A1 _6078_/A2 _6078_/A3 _6078_/A4 _6078_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_85_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5029_ _5353_/A1 _5439_/B2 _5029_/B _5354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4400_ _4412_/A1 _4399_/Z _4491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_157_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ _4568_/Z _4892_/B _4821_/Z _4675_/Z _5380_/C _5381_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_153_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4331_ hold291/Z hold747/Z _4331_/S _4331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7050_ _7050_/D _7256_/RN _7050_/CLK _7050_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4262_ _4227_/S _3994_/Z hold32/Z _4270_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_86_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _7028_/Q _5999_/Z _6000_/Z _7126_/Q _6008_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_67_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ hold961/Z hold291/Z _4193_/S _4193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6903_ _6903_/D _7237_/RN _6903_/CLK _6903_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_51_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _6834_/D _7279_/RN _7279_/CLK _6834_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_90_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3977_ _6661_/Q _3973_/Z _3977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6765_ _6765_/D _7218_/RN _6765_/CLK _7331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5716_ hold20/Z hold60/Z _5718_/S hold61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6696_ _6696_/D _7170_/RN _6696_/CLK _6696_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_163_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ _5647_/A1 hold32/Z hold16/Z hold273/Z _5655_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5578_ hold161/Z hold91/Z _5583_/S _5578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7317_ _7317_/I _7317_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold252 _6701_/Q hold252/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_145_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold241 _5887_/Z _7216_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4529_ _5420_/A2 _3401_/I _4530_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold230 _4278_/Z _6789_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold296 _6774_/Q hold296/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold274 _5494_/Z _5496_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold285 _5500_/Z _6880_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold263 _6679_/Q hold263/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7248_ _7248_/D _7260_/RN _7260_/CLK _7248_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_172_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7179_ _7179_/D _7237_/RN _7179_/CLK _7179_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7238__362 _7238_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_3169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4880_ _4880_/A1 _4877_/Z _4879_/Z _5167_/B _4880_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3900_ _6728_/Q _4191_/A1 _3919_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_178_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3831_ _3537_/Z _3578_/Z _6611_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_177_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ _6854_/Q _6241_/Z _6251_/Z _6825_/Q _6268_/Z _6800_/Q _6553_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3762_ _3761_/Z hold998/Z _3899_/S _6871_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5501_ hold125/Z hold65/Z _5502_/S _5501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ _7213_/Q _6256_/Z _6263_/Z _6939_/Q _6493_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3693_ _7000_/Q _5638_/A1 _3724_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5432_ _5432_/A1 _5189_/Z _5209_/Z _4985_/Z _5432_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5363_ _5363_/A1 _5342_/I _5363_/B1 _5396_/A1 _5383_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_127_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput335 _7269_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput324 _6796_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput313 _6804_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput302 _3619_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4314_ _4313_/Z _6832_/Q _6577_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_142_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _7102_/D _7218_/RN _7102_/CLK _7102_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5294_ _5294_/A1 _5366_/A2 _5296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4245_ _4244_/Z hold769/Z _4245_/S _4245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7033_ hold34/Z _7260_/RN _7033_/CLK _7033_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_171_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _3535_/Z _3552_/Z _5520_/C _4178_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_28_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _6817_/D _6818_/CLK _6817_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6748_ _6748_/D _7258_/RN _6748_/CLK _6748_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet763_431 net763_431/I _6739_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_420 net763_420/I _6754_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_442 net413_75/I _6723_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_17__1359_ clkbuf_4_2_0__1359_/Z net513_189/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6679_ _6679_/D _7008_/RN _6679_/CLK _6679_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_164_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_174_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _4386_/A3 _4386_/A4 _4391_/A1 _4391_/A2 _4030_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_37_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5981_ _6210_/C _6021_/A2 _6210_/A2 _7227_/Q _5981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4932_ _5258_/B2 _5056_/C _5442_/A2 _5248_/A2 _4933_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_80_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6602_ _6602_/I0 _7277_/Q _6602_/S _7277_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4863_ _4624_/Z _4833_/Z _4865_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_14 _6951_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_25 user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4794_ _4673_/Z _4793_/Z _5452_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3814_ _6729_/Q _4191_/A1 _3876_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_158_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3745_ _7209_/Q _3960_/A2 _5665_/A1 _7023_/Q _3747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6533_ _6838_/Q _6533_/A2 _6533_/A3 _6533_/A4 _6540_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6464_ _6464_/A1 _6464_/A2 _6464_/A3 _6464_/A4 _6464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_107_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ _4703_/Z _4982_/Z _5415_/B1 _5083_/C _5416_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_134_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3676_ _7115_/Q _3917_/A2 _5683_/A1 _7041_/Q _3687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6395_ _7254_/Q _6395_/I1 _6558_/S _7254_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet713_372 net713_373/I _6838_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_361 net763_449/I _6849_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5346_ _5393_/A2 _5346_/A2 _5346_/B _5347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput176 _3365_/ZN mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_394 net713_394/I _6780_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_383 net713_383/I _6799_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput198 _3345_/ZN mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput187 _3355_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5277_ _5277_/I _5421_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ _4227_/Z hold677/Z _4228_/S _4228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7016_ hold57/Z _7260_/RN _7016_/CLK _7016_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_130_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4159_ _4103_/I hold841/Z _4160_/S _4159_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_4__1359_ net763_436/I net413_55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3530_ _3507_/Z _3529_/Z _5656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_7_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold818 _4255_/Z _6770_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_156_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold807 _6757_/Q hold807/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_115_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput89 spimemio_flash_io2_do input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput78 spi_csb input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_182_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3461_ _6665_/Q _6663_/Q _6730_/Q _3463_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_143_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63__1359_ net513_170/I net763_417/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_143__1359_ clkbuf_4_1_0__1359_/Z net813_487/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold829 _7079_/Q hold829/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5200_ _5205_/A1 _5291_/B _5200_/B1 _5346_/A2 _5200_/C _5354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_112_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _6180_/A1 _6180_/A2 _6180_/A3 _6180_/A4 _6180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3392_ _6891_/Q _3903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _5172_/A1 _5291_/A2 _5165_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_123_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ _4699_/Z _5330_/B2 _5062_/B _5063_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_112_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4013_ _5942_/S _7235_/Q _6311_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_111_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5964_ _6117_/A4 _6014_/A2 _6210_/A2 _7229_/Q _5964_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4915_ _4496_/Z _4495_/Z _5263_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5895_ _6746_/Q _6744_/Q _5901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_61_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4846_ _4846_/A1 _4846_/A2 _5090_/A2 _4849_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_21_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4777_ _4782_/A1 _5099_/A1 _5456_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6516_ _6512_/Z _6516_/A2 _6516_/A3 _6516_/A4 _6516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3728_ input46/Z _4210_/S _3739_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3659_ _7091_/Q _3945_/B1 _3927_/B1 hold60/I _3663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6447_ _6440_/Z _6446_/Z _6447_/B1 _6286_/Z _6555_/C _6448_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _7071_/Q _6248_/Z _6293_/Z _7153_/Q _6380_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5329_ _5359_/A1 _4716_/Z _5445_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_103_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4700_ _5420_/A2 _5129_/A3 _5051_/S _3401_/I _4700_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ _7033_/Q hold20/Z hold33/Z hold34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4631_ _4868_/A1 _4524_/Z _5403_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_72_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4562_ _4422_/Z _4483_/B _5291_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_183_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7281_ _7281_/D _6635_/Z _7305_/CLK _7281_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
Xhold615 _5860_/Z _7192_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4493_ _4808_/A2 _4492_/Z _5240_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3513_ _3509_/Z _3512_/Z _3923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold604 _7112_/Q hold604/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6301_ _7052_/Q _6299_/Z _6300_/Z _7102_/Q _6306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold626 _7028_/Q hold626/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3444_ _3442_/B _3452_/S _3449_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold659 _5558_/Z _6924_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap345 _4064_/S _6652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold637 _7206_/Q hold637/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap356 input75/Z _7170_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold648 _5667_/Z _7021_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6232_ _7250_/Q _6232_/I1 _6558_/S _7250_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ _7125_/Q _5969_/Z _6176_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3375_ _6959_/Q _3375_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _4762_/Z _4867_/Z _5403_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_85_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _6094_/I _6095_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5045_ _5214_/A2 _5389_/A1 _5172_/B _5045_/C _5433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_97_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6996_ _6996_/D _7260_/RN _6996_/CLK _6996_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5947_ _6285_/A2 _7237_/Q _6484_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_129_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ hold91/Z hold242/Z _5883_/S _5878_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4829_ _4673_/Z _4683_/Z _5276_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_21_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_13_0__1359_ clkbuf_0__1359_/Z net513_175/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_72_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold1 hold1/I hold1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_95_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_108 net463_110/I _7117_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_119 net413_73/I _7106_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _6850_/D _7170_/RN _6850_/CLK _6850_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ hold12/Z hold52/Z _5802_/S hold53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ hold49/Z _7260_/RN _6781_/CLK _6781_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3993_ _3994_/A1 _6902_/Q input67/Z _4064_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_50_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5732_ hold227/Z hold404/Z _5739_/S _5732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5663_ hold281/Z hold12/Z hold56/Z _7018_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4614_ _4441_/B _4467_/B _4460_/B _4501_/B _4614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5594_ hold227/Z hold394/Z hold7/Z _5594_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4545_ _4454_/Z _4878_/A2 _5172_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7333_ _7333_/I _7333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold401 _5836_/Z _7171_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold412 _5553_/Z _6920_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold445 _5573_/Z _6938_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold434 _5763_/Z _7106_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold423 _5502_/Z _6882_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold478 _6772_/Q hold478/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold456 _7116_/Q hold456/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4476_ _4853_/A1 _4481_/A2 _5288_/B _4692_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_104_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7264_ _7264_/D _7265_/CLK _7264_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold467 _4154_/Z _6702_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3427_ _6733_/Q _6732_/Q _6730_/Q _3427_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_131_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold489 _5810_/Z _7148_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7195_ _7195_/D _7237_/RN _7195_/CLK _7195_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6215_ _6713_/Q _6002_/Z _6003_/Z _6715_/Q _6217_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3358_ _7089_/Q _3358_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6146_ _7124_/Q _5969_/Z _6146_/B _6147_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6077_ _7055_/Q _5924_/Z _5988_/Z _6983_/Q _6168_/C _6078_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_57_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _5023_/Z _5476_/A1 _5027_/I _5028_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_2617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6979_ _6979_/D _7258_/RN _6979_/CLK _6979_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_41_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold990 _5787_/Z _7127_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_135_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4330_ hold227/Z hold244/Z _4331_/S _4330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ hold2/Z hold214/Z _4261_/S _4261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6000_ _6015_/A3 _6211_/B1 _7231_/Q _7228_/Q _6000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_140_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4192_ hold693/Z _4103_/I _4193_/S _4192_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6902_ _6902_/D _7218_/RN _6902_/CLK _6902_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_70_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _6833_/D _7279_/RN _7278_/CLK _6833_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_63_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ _3975_/Z _6662_/Q _3988_/S _6662_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _6764_/D _7170_/RN _6764_/CLK _6764_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5715_ hold48/Z hold107/Z _5718_/S _5715_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6695_ _6695_/D input75/Z _6695_/CLK _6695_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_148_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5646_ hold207/Z hold2/Z _5646_/S _5646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold220 _5773_/Z _7115_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_129_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5577_ hold679/Z hold291/Z _5583_/S _5577_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7316_ _7316_/I _7316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold253 _4153_/Z _6701_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4528_ _5359_/A1 _4524_/Z _4472_/B _4501_/B _4528_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold242 _7208_/Q hold242/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold231 _7020_/Q hold231/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ _4555_/B _5270_/A1 _5281_/C _4459_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7247_ _7247_/D _7258_/RN _7258_/CLK _7247_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold286 _6928_/Q hold286/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold275 _5495_/Z _6876_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold264 _4125_/Z _6679_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold297 _4259_/Z _6774_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_86_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7178_ _7178_/D _7218_/RN _7178_/CLK _7178_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_3104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ hold29/I _5964_/Z _6014_/Z hold86/I _6000_/Z _7131_/Q _6134_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_3137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3830_ _3529_/Z _3540_/Z _3942_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_189_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3761_ _6567_/I0 _6870_/Q _3898_/S _3761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5500_ hold284/Z hold91/Z _5502_/S _5500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6480_ _7221_/Q _6274_/Z _6285_/Z _7197_/Q _7181_/Q _6254_/Z _6493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3692_ _3505_/Z _3527_/Z _3916_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_173_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _5431_/A1 _5299_/C _5431_/B _5431_/C _6863_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _5362_/A1 _5362_/A2 _5362_/A3 _5363_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_160_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput314 _6805_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput325 _6797_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput303 _4070_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4313_ _6834_/Q _6835_/Q _6836_/Q _4313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7101_ _7101_/D _7256_/RN _7101_/CLK _7101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_5_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput336 _6814_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5293_ _5293_/A1 _5295_/A1 _5293_/B _5366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_102_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7032_ _7032_/D _7258_/RN _7032_/CLK _7032_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_141_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4244_ hold288/Z hold2/Z _4244_/S _4244_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ hold291/Z hold755/Z _4175_/S _4175_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6816_ _6816_/D _7265_/CLK _6816_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6747_ _6747_/D _7170_/RN _6747_/CLK _6747_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet763_432 net763_435/I _6738_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet763_421 net763_421/I _6753_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_410 net763_421/I _6764_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3959_ _7012_/Q _5656_/A1 _3959_/B1 _6666_/Q _3959_/C1 _7182_/Q _3961_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_167_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _6678_/D input75/Z _6678_/CLK _6678_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet763_443 net413_75/I _6722_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5629_ _3509_/Z _5520_/C _5839_/A3 _5857_/A3 _5637_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_152_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1_0__1359_ clkbuf_0__1359_/Z clkbuf_4_1_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _6015_/A3 _6210_/C _7231_/Q _7228_/Q _5980_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_92_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_23__1359_ _4073__49/I net613_268/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_103__1359_ clkbuf_4_5_0__1359_/Z net413_84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _5389_/A2 _5056_/C _5442_/A2 _5248_/A2 _4933_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_86__1359_ net513_175/I net563_222/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4862_ _4862_/A1 _4859_/Z _4861_/Z _4819_/Z _4865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6601_ _6601_/A1 _4313_/Z _6601_/B _6602_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_177_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3813_ _3552_/Z _3680_/Z _4191_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_36_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4793_ _4534_/Z _5312_/A1 _4491_/B _4402_/B _4793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_26 user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_15 _6951_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3744_ _6959_/Q _3957_/A2 _3927_/A2 _6701_/Q _3747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6532_ _6697_/Q _6282_/Z _6542_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_118_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _6938_/Q _6263_/Z _6266_/Z _7018_/Q _6464_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3675_ _7179_/Q _3945_/A2 _5758_/A1 _7107_/Q _3687_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ _4997_/B _5414_/A2 _4659_/Z _5414_/B _5418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_127_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ _6394_/I _6395_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet713_362 net713_383/I _6848_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5345_ _5389_/C _5345_/A2 _5356_/B _5389_/A2 _5346_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput177 _3364_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_395 net763_425/I _6779_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_373 net713_373/I _6837_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_384 net713_385/I _6790_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput199 _4052_/ZN mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput188 _3354_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5276_ _5276_/A1 _5276_/A2 _5291_/C _5276_/C _5277_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_99_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4227_ hold256/Z hold2/Z _4227_/S _4227_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7015_ _7015_/D _7238_/RN _7015_/CLK hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_68_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _5520_/C _3552_/Z _5513_/A3 _5839_/A3 _4160_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_55_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _6907_/Q input39/Z _4089_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_102_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold819 _7318_/I hold819/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_156_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold808 _4235_/Z _6757_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_122_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput68 mgmt_gpio_in[5] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput79 spi_enabled _4055_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3460_ hold290/Z input58/Z _3460_/S _7284_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3391_ _7222_/Q _5894_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ _5240_/B _5328_/A2 _5130_/B1 _5130_/B2 _5321_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5061_ _4699_/Z _4936_/I _5061_/B _5410_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_97_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4012_ _6302_/A4 _7236_/Q _6282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ _6021_/A2 _7227_/Q _6117_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_25_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4914_ _4497_/Z _4494_/Z _5442_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_52_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ _5894_/A1 _5894_/A2 _5894_/A3 _4019_/B _6746_/Q _7222_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_178_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _4596_/Z _4817_/Z _5090_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _4703_/Z _5236_/B _5121_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_165_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3727_ _3726_/Z _6872_/Q _3899_/S _6872_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6515_ _6845_/Q _6235_/Z _6237_/Z _6837_/Q _6516_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3658_ hold58/I _3951_/C1 _3924_/A2 _6969_/Q input25/Z _3954_/B1 _3688_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6446_ _6554_/A1 _6446_/A2 _6446_/A3 _6446_/A4 _6446_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_164_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6377_ _7201_/Q _6272_/Z _6282_/Z _7185_/Q _6296_/Z _7161_/Q _6384_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3589_ _3589_/A1 _3589_/A2 _3589_/A3 _3589_/A4 _3589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5328_ _5328_/A1 _5328_/A2 _5481_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_161_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ _5259_/A1 _5259_/A2 _5337_/A2 _5449_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_130_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4630_ _4367_/Z _4555_/B _5291_/C _5387_/A1 _5387_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_72_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4561_ _4556_/Z _4561_/A2 _5003_/A2 _4561_/B _4584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _7234_/Q _6300_/A2 _6484_/A3 _5943_/S _6300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7280_ _7280_/D _6634_/Z _7305_/CLK hold22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_155_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4492_ _4402_/B _4026_/B _4026_/C _5312_/A1 _4492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_143_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold616 _6767_/Q hold616/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3512_ _3653_/A1 _3617_/A1 _3501_/Z _3492_/Z _3512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold605 _5770_/Z _7112_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold627 _6932_/Q hold627/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3443_ _3438_/S _3440_/S _3443_/A3 _3443_/A4 _3452_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xmax_cap346 _4225_/S _4227_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold638 _5876_/Z _7206_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap357 _7008_/RN _7256_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold649 _7107_/Q hold649/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6231_ _6231_/I _6232_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6162_ _7247_/Q _6162_/I1 _6558_/S _7247_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5113_ _5113_/A1 _5113_/A2 _5313_/A1 _5313_/A3 _5113_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3374_ _6967_/Q _3374_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _7000_/Q _6021_/Z _6090_/Z _5924_/Z _6094_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5044_ _5044_/A1 _5386_/A1 _5044_/A3 _5432_/A1 _5044_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_38_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _6995_/D _7256_/RN _6995_/CLK _6995_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5946_ _5950_/B1 _5945_/B _7236_/Q _7236_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5877_ hold291/Z hold943/Z _5883_/S _5877_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _5287_/B _4586_/Z _4784_/Z _4598_/Z _5414_/A2 _5421_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_4759_ _4501_/B _4759_/A2 _4759_/A3 _4759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_181_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6429_ hold73/I _6253_/Z _6296_/Z _7163_/Q _6434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_175_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold2 hold2/I hold2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_66_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_109 net413_96/I _7116_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3992_ _7298_/Q hold22/I _3995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_90_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5800_ hold20/Z hold73/Z _5802_/S hold74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6780_ hold68/Z _7238_/RN _6780_/CLK hold67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ _3523_/Z _3537_/Z hold24/Z _5739_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_95_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ hold377/Z hold20/Z hold56/Z _7017_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4613_ _5288_/B _5281_/C _4436_/B _4472_/B _5291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_129_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5593_ hold24/I _3523_/Z hold42/I hold6/Z hold7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold402 _7070_/Q hold402/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4544_ _4454_/Z _4456_/B _5276_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_8_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _7332_/I _7332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7263_ _7263_/D _7269_/CLK _7263_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold424 _7202_/Q hold424/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold435 _7154_/Q hold435/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold413 _6895_/Q hold413/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold457 _5774_/Z _7116_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4475_ _5288_/C _4454_/Z _4367_/Z _4501_/B _4692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold468 _7220_/Q hold468/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold446 _7124_/Q hold446/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6214_ _6825_/Q _5988_/Z _6019_/Z _6854_/Q _6217_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3426_ _6733_/Q _6732_/Q _6730_/Q _3434_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold479 _4257_/Z _6772_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7194_ _7194_/D _7218_/RN _7194_/CLK _7194_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3357_ _7097_/Q _3357_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6145_ hold50/I _5958_/Z _5994_/I hold52/I _6147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6076_ _7089_/Q _6002_/Z _6015_/Z _7007_/Q _6076_/C _6078_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_97_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _5027_/I _5200_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6978_ _6978_/D _7258_/RN _6978_/CLK _6978_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_167_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _5925_/Z _7231_/Q _6168_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_55_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold980 _7111_/Q hold980/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold991 _7175_/Q hold991/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4260_ hold12/Z hold594/Z _4261_/S _4260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ _4191_/A1 hold32/Z _4193_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_121_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6901_ _6901_/D _7235_/RN _6901_/CLK _6901_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_78_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _6832_/D _7279_/RN _7279_/CLK _6832_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_165_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3975_ _3483_/Z _3975_/I1 _3975_/S _3975_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6763_ _6763_/D _7170_/RN _6763_/CLK _6763_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5714_ hold65/Z hold248/Z _5718_/S _5714_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _6694_/D input75/Z _6694_/CLK _6694_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_31_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _7002_/Q hold12/Z _5646_/S hold13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold210 _5673_/Z _7027_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5576_ hold390/Z hold227/Z _5583_/S _5576_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4527_ _5359_/A1 _4997_/C _5243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7315_ _7315_/I _7315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold243 _5878_/Z _7208_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold221 _7136_/Q hold221/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold232 _5666_/Z _7020_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold254 _7071_/Q hold254/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4458_ _4467_/A1 _4555_/B _4736_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold287 _5562_/Z _6928_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7246_ _7246_/D _7256_/RN _7260_/CLK _7246_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_85_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold276 _6978_/Q hold276/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold265 _7026_/Q hold265/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3409_ _6665_/Q _6664_/Q _6663_/Q _3409_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_172_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7177_ _7177_/D _7237_/RN _7177_/CLK _7177_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold298 _6668_/Q hold298/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4389_ _4427_/A2 _4427_/A3 _4485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6128_ hold60/I _5985_/Z _5997_/Z _7099_/Q _6128_/C _6134_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ _7030_/Q _5999_/Z _6014_/Z _6958_/Q _6000_/Z _7128_/Q _6061_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_3149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_190 net763_426/I _7035_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _3760_/A1 _3739_/Z _3759_/Z _6567_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_60_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _5268_/Z _5430_/A2 _5428_/Z _5429_/Z _5431_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3691_ _3690_/Z hold997/Z _3899_/S _6873_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5361_ _5361_/A1 _5209_/Z _5362_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput304 _4069_/Z serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput315 _6806_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput326 _6798_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_46__1359_ net663_324/I _4073__9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5292_ _5423_/A2 _5292_/A2 _5292_/A3 _5292_/A4 _5294_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7100_ _7100_/D _7237_/RN _7100_/CLK _7100_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_leaf_126__1359_ _4073__7/I _4073__27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput337 _6815_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _6571_/I0 _6818_/Q _4312_/S _6818_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4243_ _4242_/Z hold777/Z _4245_/S _4243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7031_ _7031_/D _7258_/RN _7031_/CLK _7031_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _4103_/I hold691/Z _4175_/S _4174_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _6815_/D _6818_/CLK _6815_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6746_ _6746_/D _7235_/RN _4067_/I1 _6746_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_50_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_433 net763_434/I _6737_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet763_411 net763_444/I _6763_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3958_ _3958_/A1 _3958_/A2 _3958_/A3 _3958_/A4 _3958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet763_422 net763_422/I _6752_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6677_ _6677_/D _7008_/RN _6677_/CLK _6677_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xnet763_444 net763_444/I _6721_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3889_ _3889_/A1 _3889_/A2 _3889_/A3 _3889_/A4 _3889_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_164_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5628_ hold2/Z hold223/Z _5628_/S _5628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ hold291/Z hold951/Z _5565_/S _5559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _7229_/D _7256_/RN _7258_/CLK _7229_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_101_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4930_ _5129_/A3 _5325_/B _5051_/S _5170_/A2 _4930_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_75_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4861_ _4887_/A1 _4868_/A1 _5414_/A2 _5287_/B _4861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_75_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6600_ _6834_/Q _6600_/A2 _6600_/B1 _6835_/Q _6836_/Q _6600_/C2 _6601_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_178_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3812_ _3552_/Z _3578_/Z _4146_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_162_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_27 _7279_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ _4492_/Z _4534_/Z _5129_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_16 pad_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3743_ _7063_/Q _3927_/B1 _3924_/A2 _6967_/Q _3743_/C _3759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6531_ _6821_/Q _6262_/Z _6554_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_185_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6462_ _7172_/Q _5948_/Z _6261_/Z _6962_/Q _6464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3674_ _3674_/A1 _3674_/A2 _3674_/A3 _3673_/Z _3674_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5413_ _5448_/A1 _5483_/A1 _5412_/Z _5414_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6393_ _6744_/Q _7253_/Q _6393_/B _6394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_118_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5344_ _5438_/C _4666_/Z _5387_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_363 net713_383/I _6847_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_352 net763_439/I _6858_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_396 net763_426/I _6778_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput167 _4087_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet713_374 net713_385/I _6825_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_385 net713_385/I _6789_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput178 _3363_/ZN mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput189 _3353_/ZN mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5275_ _5376_/B2 _5468_/A2 _5275_/B _5423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_87_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7014_ _7014_/D _7258_/RN _7014_/CLK _7014_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4226_ _4225_/Z hold592/Z _4228_/S _4226_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4157_ hold2/Z hold121/Z _4157_/S _4157_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4088_ _6906_/Q input70/Z _4088_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_37_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6729_ _6729_/D _7170_/RN _6729_/CLK _6729_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_183_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92__1359_ net413_62/I net613_266/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold809 _6760_/Q hold809/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput69 mgmt_gpio_in[6] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3390_ _7241_/Q _6011_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _5058_/Z _5060_/A2 _4928_/Z _5060_/A4 _5064_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_123_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _6282_/A2 _7232_/Q _6484_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_84_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _5984_/A1 _7230_/Q _6002_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_52_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _4376_/Z _5442_/A2 _4909_/Z _4927_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_18_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ _5945_/A1 _6746_/Q _5894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4844_ _5287_/B _4456_/B _4530_/I _5051_/S _4844_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4775_ _4775_/A1 _4772_/Z _4773_/Z _4774_/Z _4781_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_20_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3726_ _4309_/I0 _6871_/Q _3898_/S _3726_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6514_ _6787_/Q _6263_/Z _6266_/Z _6843_/Q _6516_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3657_ _3657_/A1 _3657_/A2 _3657_/A3 _3657_/A4 _3657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6445_ _7049_/Q _6241_/Z _6268_/Z hold71/I _6256_/Z _7211_/Q _6446_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6376_ _7113_/Q _6240_/Z _6376_/B _6384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3588_ _7133_/Q _3930_/A2 _3941_/B1 _7173_/Q _3588_/C _3589_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5327_ _4928_/Z _5326_/Z _5327_/A3 _5327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_138_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5258_ _4890_/I _5258_/A2 _4972_/Z _5258_/B2 _5258_/C _5412_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_180_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5189_ _5386_/A1 _5386_/A3 _5189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4209_ _4208_/Z hold783/Z _4211_/S _4209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4560_ _5002_/A3 _5002_/A4 _5083_/B _5393_/B1 _4561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_129_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _4491_/A1 _4491_/A2 _4491_/B _5312_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold617 _4251_/Z _6767_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3511_ hold320/Z _3489_/I _5821_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold606 _7160_/Q hold606/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3442_ _3991_/A1 _4042_/A3 _6733_/Q _3442_/B _3443_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xmax_cap347 _5323_/B _5442_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_143_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6230_ _6555_/C _7249_/Q _6230_/B _6231_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold639 _7086_/Q hold639/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap358 _7238_/RN _7260_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold628 _5567_/Z _6932_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ _6161_/I _6162_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3373_ hold69/I _3373_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5112_ _4614_/Z _5302_/B _4784_/Z _5230_/B _4716_/Z _5113_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_69_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6092_ _6092_/A1 _5991_/Z _6102_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _5385_/A1 _5043_/A2 _5043_/B _5432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_111_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0_wbbd_sck _7278_/Q clkbuf_0_wbbd_sck/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6994_ _6994_/D _7258_/RN _6994_/CLK _6994_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5945_ _5945_/A1 _6745_/Q _5945_/B _5950_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_40_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ hold227/Z hold637/Z _5883_/S _5876_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4827_ _4586_/Z _4784_/Z _5223_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _5072_/A4 _4500_/Z _4958_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_181_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4689_ _4687_/Z _5092_/A1 _5302_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3709_ _7210_/Q _3960_/A2 _3955_/A2 _7202_/Q _7186_/Q _3959_/C1 _3724_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _7009_/Q _6243_/Z _6269_/Z _7033_/Q _6440_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_175_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6359_ _6359_/I _6360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold3 hold3/I hold3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_12_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3991_ _3991_/A1 _3412_/Z _3442_/B _3409_/Z _6730_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_16_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5730_ hold907/Z hold291/Z _5730_/S _5730_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ _7016_/Q hold48/Z hold56/Z hold57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4612_ _4612_/A1 _4612_/A2 _5025_/B _4618_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_148_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5592_ hold103/Z hold2/Z _5592_/S _5592_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _5129_/A3 _5051_/S _4878_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_144_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7331_ _7331_/I _7331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold403 _5722_/Z _7070_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold425 _5871_/Z _7202_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7262_ _7262_/D _7265_/CLK _7262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold436 _5817_/Z _7154_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold414 _7072_/Q hold414/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4474_ _5288_/C _4454_/Z _4367_/Z _4501_/B _4474_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold458 _6919_/Q hold458/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold469 _5891_/Z _7220_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold447 _5783_/Z _7124_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6213_ _6821_/Q _5979_/Z _5996_/Z _6709_/Q _6217_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3425_ _3425_/I0 _7302_/Q _3425_/S _7302_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _7193_/D _7218_/RN _7193_/CLK _7193_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_174_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3356_ _7105_/Q _3356_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6144_ _7066_/Q _5985_/Z _6000_/Z _7132_/Q _6144_/C _6147_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_58_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ hold75/I _5971_/Z _6003_/Z _7161_/Q _6078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xload_slew350 _4102_/Z _4103_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _5471_/B2 _5291_/B _5002_/Z _5200_/B1 _5027_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6977_ hold30/Z _7260_/RN _6977_/CLK hold29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5928_ _7231_/Q _5941_/A1 _5931_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ hold291/Z hold993/Z _5865_/S _5859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold981 _5769_/Z _7111_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold970 _5842_/Z _7176_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold992 _5841_/Z _7175_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_62_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_250 net613_256/I _6975_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ hold733/Z hold291/Z _4190_/S _4190_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6900_ _6900_/D _7238_/RN _6900_/CLK _6900_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_6831_ _6831_/D _7279_/RN _7279_/CLK _6831_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_91_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69__1359_ net513_175/I net613_263/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ _6661_/Q _6660_/Q _6659_/Q _3972_/Z _3975_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_165_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ _6762_/D _7256_/RN _6762_/CLK _6762_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_189_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5713_ hold91/Z hold386/Z _5718_/S _5713_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6693_ _6693_/D _7218_/RN _6693_/CLK _6693_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_137_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5644_ hold62/Z hold20/Z _5646_/S hold63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7314_ _7314_/I _7314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold200 _7131_/Q hold200/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold211 _7084_/Q hold211/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5575_ _5575_/A1 hold32/Z _5583_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4526_ _4472_/B _4501_/B _4460_/B _4436_/B _4997_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold233 _6860_/Q hold233/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold244 _6837_/Q hold244/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold222 _5797_/Z _7136_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold255 _5723_/Z _7071_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4457_ _4456_/B _5051_/S _4460_/B _4467_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_116_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _7245_/D _7256_/RN _7258_/CLK _7245_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold277 _5618_/Z _6978_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold266 _5672_/Z _7026_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold288 _6923_/Q hold288/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3408_ _4436_/B _4467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
X_7176_ _7176_/D _7008_/RN _7176_/CLK _7176_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_59_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold299 _4108_/Z _6668_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4388_ _4388_/A1 _4388_/A2 input97/Z input96/Z _4427_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_59_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _6127_/A1 _6124_/Z _6127_/A3 _6127_/A4 _6127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_112_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3339_ _3339_/I _3932_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _7062_/Q _5985_/Z _5997_/Z _7096_/Q _6061_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_65_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _5438_/C _5359_/A1 _5435_/A2 _5475_/A3 _5009_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_191 net563_239/I _7034_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_180 _4073__50/I _7045_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_188_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3690_ _6569_/I0 _6872_/Q _3898_/S _3690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _5045_/C _5393_/B1 _5360_/B _5360_/C _5361_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_154_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput316 _6807_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput305 _4086_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5291_ _4542_/Z _5291_/A2 _5291_/B _5291_/C _5377_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput327 _7262_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4311_ _6570_/I0 _6817_/Q _4312_/S _6817_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput338 _6816_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4242_ hold358/Z hold12/Z _4244_/S _4242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7030_ _7030_/D _7260_/RN _7030_/CLK _7030_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_113_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_1_0__1359_ _4073__49/I clkbuf_opt_1_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _5821_/A3 _5513_/A3 _3537_/Z _5520_/C _4175_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_45_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _6814_/D _6818_/CLK _6814_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6745_ _6745_/D _7235_/RN _4067_/I1 _6745_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3957_ _6956_/Q _3957_/A2 _4289_/A1 _6799_/Q _3958_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet763_412 net763_417/I _6762_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_423 net763_423/I _6751_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_434 net763_434/I _6736_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6676_ _6676_/D _7008_/RN _6676_/CLK _6676_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3888_ _6989_/Q _3954_/A2 _3956_/A2 _7119_/Q _3889_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet763_445 net763_445/I _6720_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5627_ hold12/Z hold437/Z _5628_/S _5627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5558_ hold227/Z hold658/Z _5565_/S _5558_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _5087_/A1 _5051_/S _5343_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5489_ _5489_/A1 _5489_/A2 _5472_/Z _5489_/A4 _5489_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_132_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7228_ _7228_/D _7256_/RN _7258_/CLK _7228_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_120_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7159_ _7159_/D _7218_/RN _7159_/CLK _7159_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52__1359_ net663_324/I net813_464/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_132__1359_ net513_165/I net813_488/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _5104_/A1 _4860_/A2 _5291_/C _5291_/B _5376_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_82_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3811_ _3509_/Z _3578_/Z _3925_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_17 user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4791_ _5312_/A2 _5214_/A2 _5456_/A1 _5220_/B2 _4791_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ _7259_/Q _6529_/Z _6558_/S _7259_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3742_ _3742_/I _3743_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _7220_/Q _6274_/Z _6285_/Z _7196_/Q _7180_/Q _6254_/Z _6464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3673_ _3673_/A1 _3673_/A2 _3673_/A3 _3673_/A4 _3673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5412_ _5412_/A1 _5412_/A2 _5412_/A3 _4984_/B _5412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6392_ _6385_/Z _6391_/Z _6392_/B1 _6286_/Z _6744_/Q _6393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _5343_/A1 _5343_/A2 _5343_/B _5418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xnet713_353 net763_439/I _6857_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput168 _7307_/Z irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet713_375 net813_489/I _6824_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_386 net413_55/I _6788_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_364 net763_421/I _6846_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput179 _3362_/ZN mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5274_ _5370_/A1 _5312_/A4 _5291_/C _5295_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_102_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_397 net763_427/I _6777_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7013_ _7013_/D _7260_/RN _7013_/CLK _7013_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4225_ hold111/Z hold12/Z _4225_/S _4225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4156_ hold12/Z hold180/Z _4157_/S _4156_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ input1/Z input36/Z _4087_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_70_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _5340_/A1 _5262_/A2 _5328_/A2 _5248_/A2 _4991_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_51_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6728_ _6728_/D _7170_/RN _6728_/CLK _6728_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_178_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _6659_/D _6614_/Z _7305_/CLK _6659_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_164_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _4010_/I _6744_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _6948_/Q _5958_/Z _5960_/Z _7150_/Q _5974_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4912_ _5464_/A1 _5443_/A1 _5193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5892_ hold2/Z hold119/Z _5892_/S _5892_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4843_ _5287_/B _4784_/Z _5231_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_61_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4774_ _4782_/A1 _4510_/Z _5302_/B _4695_/Z _4774_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_146_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3725_ _3708_/Z _3724_/Z _3725_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6513_ _6809_/Q _6261_/Z _6268_/Z _6799_/Q _6265_/Z _6839_/Q _6516_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6444_ _7219_/Q _6274_/Z _6285_/Z _7195_/Q _7179_/Q _6254_/Z _6446_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_106_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3656_ _6679_/Q _3546_/Z _3945_/C2 _6687_/Q _3657_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6375_ _7129_/Q _6484_/A2 _6484_/A3 _6533_/A4 _6376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3587_ _3587_/I _3588_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5326_ _5246_/Z _5442_/A4 _5442_/A2 _5056_/C _5326_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _5257_/A1 _5246_/Z _5257_/B _5257_/C _5264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_142_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4208_ hold594/Z hold12/Z _4210_/S _4208_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _5243_/A1 _5043_/B _5205_/A1 _4650_/Z _5386_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_95_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4139_ hold291/Z hold761/Z _4139_/S _4139_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3510_ _3507_/Z _3509_/Z _5584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4490_ _4491_/A1 _4491_/A2 _5092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold618 _6773_/Q hold618/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold607 _5824_/Z _7160_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3441_ _6664_/Q _6663_/Q _6730_/Q _6665_/Q _3443_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_171_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold629 _7217_/Q hold629/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap348 _6068_/A4 _6211_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xmax_cap359 _7238_/RN _7258_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_6160_ _6555_/C _7246_/Q _6160_/B _6161_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3372_ _6983_/Q _3372_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5111_ _4614_/Z _4817_/Z _5111_/B _5111_/C _5113_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ hold93/I _6211_/A2 _6211_/B1 hold88/I _6092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _5385_/A1 _5389_/C _5439_/B1 _5393_/A1 _5044_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_111_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ hold28/Z _7260_/RN _6993_/CLK hold27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5944_ _6745_/Q _7235_/Q _7234_/Q _6300_/A2 _5945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_41_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ _3485_/Z _3523_/Z hold24/Z _5883_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_167_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4826_ _4826_/A1 _5370_/B _4826_/A3 _4826_/B _4834_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_139_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4757_ _4757_/I _4766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4688_ _5083_/B _5092_/A1 _5312_/A1 _5094_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_88_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ _3701_/Z _3708_/A2 _3708_/A3 _3707_/Z _3708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3639_ hold52/I _3951_/A2 _5665_/A1 _7026_/Q _7018_/Q _5656_/A1 _3642_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6427_ hold35/I _6245_/Z _6288_/Z hold76/I _6440_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_115_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6358_ _7022_/Q _6235_/Z _6243_/Z _7006_/Q _6265_/Z _6998_/Q _6359_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _4699_/Z _5309_/A2 _5456_/A2 _5309_/B2 _5309_/C _5310_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_68_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6289_ _7182_/Q _6282_/Z _6288_/Z _7118_/Q _6307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_124_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold4 hold4/I hold4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_79_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3990_ _3990_/I _5896_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_90_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ hold75/Z hold65/Z hold56/Z _7015_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _5287_/C _4565_/Z _5025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5591_ hold50/Z hold12/Z _5592_/S hold51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _5420_/A2 _5129_/A3 _5051_/S _4542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7330_ _7330_/I _7330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7261_ _7261_/D _7279_/RN _7278_/CLK _7261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4473_ _4472_/B _4473_/A2 _4481_/A2 _4853_/A1 _4786_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xhold404 _7078_/Q hold404/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold426 _6959_/Q hold426/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold415 _5724_/Z _7072_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3424_ _3465_/A4 _3465_/A3 _3971_/A1 _3442_/B _3425_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_144_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold459 _5552_/Z _6919_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold448 _6918_/Q hold448/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold437 _6986_/Q hold437/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6212_ _6212_/A1 _5991_/Z _6226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7192_ _7192_/D _7237_/RN _7192_/CLK _7192_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_98_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_29__1359_ net613_298/I net763_431/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_109__1359_ clkbuf_4_5_0__1359_/Z net413_89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3355_ _7113_/Q _3355_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6143_ _6143_/I _6144_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew351 _6744_/Q _6555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_112_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6074_ _7081_/Q _5996_/Z _6005_/Z _7039_/Q _6078_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_86_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _5439_/B2 _5200_/B1 _5025_/B _5476_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_100_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6976_ _6976_/D _7258_/RN _6976_/CLK _6976_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5927_ _5919_/Z _6014_/A2 _5941_/A1 _5925_/Z _5950_/A1 _7230_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_80_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _4103_/I hold913/Z _5865_/S _5858_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5789_ hold65/Z hold521/Z _5793_/S _5789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4809_ _4809_/A1 _4805_/Z _4807_/Z _4808_/Z _4812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold982 _7069_/Q hold982/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold971 _6965_/Q hold971/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold960 _5712_/Z _7061_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_135_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold993 _7191_/Q hold993/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_95_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_240 net763_422/I _6985_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_251 net613_266/I _6974_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6830_ _6833_/Q _7279_/RN _7279_/CLK _6830_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_36_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _6761_/D _7256_/RN _6761_/CLK _6761_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _6660_/Q _6659_/Q _3972_/Z _3973_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_149_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5712_ hold291/Z hold959/Z _5718_/S _5712_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6692_ _6692_/D _7218_/RN _6692_/CLK _6692_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_148_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5643_ hold409/Z hold48/Z _5646_/S _5643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5574_ hold2/Z hold306/Z _5574_/S _5574_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold201 _5791_/Z _7131_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7313_ _7313_/I _7313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4525_ _5315_/A2 _4524_/Z _5130_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_102_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold234 _3496_/Z _3497_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold212 _5738_/Z _7084_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold223 _6987_/Q hold223/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4456_ _3401_/I _3402_/I _4456_/B _5051_/S _4481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_7244_ _7244_/D _7258_/RN _7260_/CLK _7244_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold267 _7010_/Q hold267/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold278 _6970_/Q hold278/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold245 _4330_/Z _6837_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold256 _6784_/Q hold256/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4387_ _4388_/A1 _4388_/A2 input97/Z input96/Z _4387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3407_ _4460_/B _5281_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
Xhold289 _5556_/Z _6923_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_98_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7175_ _7175_/D _7218_/RN _7175_/CLK _7175_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_105_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3338_ _6927_/Q _6392_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ hold78/I _5996_/Z _5999_/Z _7033_/Q _6969_/Q _5979_/Z _6127_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_112_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6057_ _6057_/A1 _6057_/A2 _6057_/A3 _6057_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_22_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _5438_/C _5359_/A1 _5439_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_2417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6959_ _6959_/D _7260_/RN _6959_/CLK _6959_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_139_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_170 net513_170/I _7055_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold790 _4207_/Z _6740_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_12__1359_ clkbuf_4_2_0__1359_/Z net413_66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet513_192 net763_422/I _7033_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_181 net413_54/I _7044_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_75__1359_ net663_324/I net413_68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4075_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_185_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput306 _4081_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput317 _6808_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5290_ _4422_/Z _4554_/Z _4614_/Z _4483_/B _5290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xoutput339 _6817_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput328 _7263_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4310_ _6569_/I0 _6816_/Q _4312_/S _6816_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4241_ _4240_/Z hold809/Z _4245_/S _4241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4172_ hold859/Z hold291/Z _4172_/S _4172_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6813_ _6813_/D _6818_/CLK _6813_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6744_ _6744_/D _7256_/RN _4067_/I1 _6744_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3956_ _7118_/Q _3956_/A2 _3956_/B1 _6712_/Q _3956_/C1 _6851_/Q _3958_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet763_402 net763_434/I _6772_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_413 net763_415/I _6761_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _6675_/D input75/Z _6675_/CLK _6675_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xnet763_424 net763_425/I _6750_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_435 net763_435/I _6735_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_446 net813_483/I _6719_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3887_ _6840_/Q _3925_/C2 _3956_/C1 _6852_/Q _3889_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5626_ hold20/Z _6985_/Q _5628_/S hold21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5557_ _5520_/C _3527_/Z _5839_/A3 _5857_/A3 _5565_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4508_ _4698_/B _5087_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_145_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _5374_/Z _5487_/Z _5489_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7227_ _7227_/D _7235_/RN _4067_/I1 _7227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4439_ _4363_/Z _4369_/Z _4472_/B _4759_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_132_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7158_ _7158_/D _7170_/RN _7158_/CLK _7158_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_7089_ _7089_/D _7237_/RN _7089_/CLK _7089_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _6101_/Z _6106_/Z _6109_/A3 _6109_/A4 _6109_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_47_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4790_ _4790_/A1 _5213_/C _4787_/Z _4789_/Z _4803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_60_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _3509_/Z hold674/Z _4301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3741_ _7081_/Q _3923_/C1 _5575_/A1 _6943_/Q _3925_/A2 input6/Z _3742_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_60_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_18 _4226_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6460_ _6994_/Q _6237_/Z _6247_/Z _7132_/Q _6460_/C _6465_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3672_ _7073_/Q _3943_/A2 _3941_/A2 _7163_/Q _3673_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5411_ _5248_/Z _5327_/Z _5411_/A3 _5483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6391_ _6554_/A1 _6391_/A2 _6391_/A3 _6390_/Z _6391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_63_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5342_ _5342_/I _5418_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet713_354 net813_473/I _6856_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet713_376 net813_481/I _6823_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_387 net413_55/I _6787_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_365 net763_421/I _6845_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5273_ _4554_/Z _4683_/Z _5287_/B _5468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_88_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet713_398 net413_56/I _6776_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7012_ _7012_/D _7260_/RN _7012_/CLK _7012_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xoutput169 _4088_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _4223_/Z hold540/Z _4228_/S _4224_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4155_ hold20/Z hold184/Z _4157_/S _4155_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4086_ _4055_/S input63/Z _4086_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_102_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4988_ _5083_/C _4568_/Z _4659_/Z _4422_/Z _4988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_23_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6727_ _6727_/D _7170_/RN _6727_/CLK _6727_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3939_ _6696_/Q _4146_/A1 _4359_/A1 _6857_/Q _3939_/C1 _6710_/Q _3940_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6658_ _6658_/D _4098_/Z _7305_/CLK _6658_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_127_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ hold12/Z hold278/Z hold43/Z _6970_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6589_ _6589_/A1 _4313_/Z _6589_/B _6590_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_164_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _7231_/Q _6068_/A4 _6021_/A2 _7227_/Q _5960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_65_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4911_ _5464_/A1 _4903_/Z _5205_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5891_ hold12/Z hold468/Z _5892_/S _5891_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4842_ _5104_/A1 _4860_/A2 _4555_/C _5291_/C _4842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_60_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4773_ _4782_/A1 _5302_/B _4695_/Z _4716_/Z _4773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_187_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3724_ _3715_/Z _3724_/A2 _3724_/A3 _3723_/Z _3724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6512_ _6512_/A1 _6512_/A2 _6512_/A3 _6511_/Z _6512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _7219_/Q _3912_/A2 _3948_/C1 _7334_/I _3657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6443_ hold80/I _6235_/Z _6261_/Z hold86/I _6443_/C _6446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_173_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6374_ _7209_/Q _6256_/Z _6263_/Z _6935_/Q _6385_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3586_ _6931_/Q _3935_/A2 _3943_/A2 _7075_/Q _7157_/Q _3916_/A2 _3587_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_161_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5325_ _4716_/Z _5394_/A2 _5325_/B _5327_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_115_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5256_ _5262_/A2 _4902_/Z _5246_/Z _5257_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_88_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ _4206_/Z hold789/Z _4211_/S _4207_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5187_ _5392_/B _5339_/A4 _5417_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _4103_/I hold707/Z _4139_/S _4138_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4069_ _7238_/Q _6897_/Q _6900_/Q _4069_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold608 _7184_/Q hold608/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3440_ input58/Z _3440_/I1 _3440_/S _7294_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold619 _4258_/Z _6773_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3371_ _6991_/Q _3371_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5110_ _4614_/Z _4817_/Z _5111_/C _5479_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_88_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _6210_/A2 _7056_/Q _6090_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_5041_ _5439_/B1 _5002_/Z _5041_/B _5386_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ hold89/Z _7260_/RN _6992_/CLK hold88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_179_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5943_ _5943_/I0 _5940_/Z _5943_/S _7235_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ hold2/Z hold113/Z _5874_/S _5874_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4825_ _4539_/I _4683_/Z _4826_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4756_ _4510_/Z _4752_/Z _4757_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_161_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _5083_/B _4687_/A2 _4687_/A3 _4687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_3707_ _3707_/A1 _3707_/A2 _3707_/A3 _3707_/A4 _3707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3638_ _3638_/A1 _3638_/A2 _3638_/A3 _3638_/A4 _3638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6426_ _6969_/Q _6262_/Z _6266_/Z _7017_/Q _6426_/C _6440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3569_ _3515_/Z _3529_/Z _5674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6357_ _6357_/A1 _6357_/A2 _6356_/Z _6357_/A4 _6357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5308_ _5303_/Z _5308_/A2 _5221_/I _5480_/A1 _5308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_130_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _7236_/Q _6302_/A3 _6533_/A4 _6302_/A4 _6288_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _5238_/Z _4801_/Z _5453_/A4 _5452_/A2 _5241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_102_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold5 hold5/I hold5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_94_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ _5287_/C _4589_/Z _4612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5590_ hold71/Z hold20/Z _5592_/S hold72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4541_ _5278_/C _5279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_4472_ _4464_/Z _4454_/Z _4472_/B _4764_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold416 _7090_/Q hold416/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold427 _6886_/Q hold427/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold405 _5732_/Z _7078_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7260_ _7260_/D _7260_/RN _7260_/CLK _7260_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3423_ _3422_/Z _7303_/Q _3988_/S _7303_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold449 _5551_/Z _6918_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold438 _5627_/Z _6986_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7191_ _7191_/D _7218_/RN _7191_/CLK _7191_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6211_ _6846_/Q _6211_/A2 _6211_/B1 _6838_/Q _6212_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_135_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6142_ _6978_/Q _5964_/Z _5981_/Z _6938_/Q _6014_/Z _6962_/Q _6143_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_48_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3354_ _7121_/Q _3354_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6073_ _6073_/A1 _6073_/A2 _6073_/A3 _6073_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _4604_/Z _5475_/A3 _5200_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ hold70/Z _7260_/RN _6975_/CLK hold69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_5926_ _5950_/A1 _5925_/Z _5931_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5857_ _3485_/Z _5857_/A2 _5857_/A3 _5520_/C _5865_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_55_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5788_ hold91/Z hold429/Z _5793_/S _5788_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4808_ _4422_/Z _4808_/A2 _5312_/A1 _4666_/Z _4808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _4739_/A1 _5106_/A1 _4738_/Z _4743_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_147_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _7170_/Q _5948_/Z _6261_/Z _6960_/Q _6266_/Z _7016_/Q _6411_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_89_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold950 _5814_/Z _7151_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold972 _7029_/Q hold972/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold961 _6729_/Q hold961/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold994 _5859_/Z _7191_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold983 _5721_/Z _7069_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_4_0__1359_ clkbuf_0__1359_/Z net513_165/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_35__1359_ clkbuf_4_10_0__1359_/Z _4073__22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_115__1359_ net513_165/I net563_245/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_98__1359_ clkbuf_4_5_0__1359_/Z net713_394/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_185_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_230 net563_239/I _6995_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_241 net813_466/I _6984_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6760_ _6760_/D _7237_/RN _6760_/CLK _6760_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _7305_/Q _7304_/Q _7303_/Q _6658_/Q _3972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_149_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ hold227/Z hold666/Z _5718_/S _5711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6691_ _6691_/D _7170_/RN _6691_/CLK _6691_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_176_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5642_ hold344/Z hold65/Z _5646_/S _5642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ hold12/Z hold444/Z _5574_/S _5573_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold202 _7156_/Q hold202/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4524_ _4460_/B _4436_/B _4524_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_7312_ _7312_/I _7312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold224 _5628_/Z _6987_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold213 _7019_/Q hold213/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold235 hold235/I hold235/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4455_ _4555_/B _5270_/A1 _5170_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold246 _7323_/I hold246/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold268 _5654_/Z _7010_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7243_ _7243_/D _7260_/RN _7260_/CLK _7243_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold257 _4270_/Z _6784_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4386_ input99/Z input98/Z _4386_/A3 _4386_/A4 _4427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ _4501_/B _5288_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_132_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7174_ _7174_/D _7218_/RN _7174_/CLK _7174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold279 _6994_/Q hold279/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_113_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ _3337_/I _4082_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6125_ hold35/I _5972_/Z _6021_/Z hold62/I _6127_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_100_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _7070_/Q _5980_/Z _6005_/Z _7038_/Q _6057_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _5435_/A2 _5475_/A3 _5194_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6958_ _6958_/D _7256_/RN _6958_/CLK _6958_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_53_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5909_ _7226_/Q _5908_/Z _5910_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6889_ _6889_/D _7238_/RN _6889_/CLK _6889_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_22_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold780 _4231_/Z _6755_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold791 _6674_/Q hold791/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_160 net613_262/I _7065_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_182 net613_294/I _7043_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_171 net413_57/I _7054_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_193 net563_217/I _7032_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput307 _4082_/ZN spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput329 _7264_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput318 _6791_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ hold516/Z hold20/Z _4244_/S _4240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4171_ hold685/Z _4103_/I _4172_/S _4171_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _6812_/D _7265_/CLK _6812_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _6743_/D _7235_/RN _4067_/I1 _6743_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_91_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3955_ _7198_/Q _3955_/A2 _3955_/B1 _6847_/Q _3958_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet763_403 net763_435/I _6771_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_414 net413_72/I _6760_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ _6674_/D input75/Z _6674_/CLK _6674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_149_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_447 net813_483/I _6718_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5625_ hold48/Z hold159/Z _5628_/S _5625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3886_ _6790_/Q _3928_/B1 _4289_/A1 _6800_/Q _6810_/Q _4301_/A1 _3889_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet763_425 net763_425/I _6749_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_436 net763_436/I _6729_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_81__1359_ net513_167/I _4073__41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5556_ hold2/Z hold288/Z _5556_/S _5556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4507_ _5420_/A3 _5129_/A3 _3402_/I _4698_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5487_ _5487_/A1 _5487_/A2 _5487_/A3 _5487_/A4 _5487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4438_ _4648_/A1 _4648_/A2 _4438_/B _4438_/C _5190_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_172_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7226_ _7226_/D _7235_/RN _4067_/I1 _7226_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4369_ _3402_/I _4456_/B _5051_/S _4369_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7157_ _7157_/D _7256_/RN _7157_/CLK _7157_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7088_ _7088_/D _7256_/RN _7088_/CLK _7088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _7154_/Q _5960_/Z _5964_/Z _6976_/Q _5981_/Z _6936_/Q _6109_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_47_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _6555_/C _7241_/Q _6039_/B _6040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3740_ _6935_/Q _3910_/A2 _3927_/C2 input29/Z _3954_/A2 _6991_/Q _3759_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA_19 _4247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3671_ hold29/I _3923_/A2 _5665_/A1 hold80/I _3673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5410_ _5410_/A1 _5481_/B1 _5410_/B _5411_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_127_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6390_ _6390_/A1 _6390_/A2 _6390_/A3 _6390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_9_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5341_ _4997_/B _4878_/Z _5341_/B _5341_/C _5342_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_126_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet713_355 net813_473/I _6855_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_377 net813_481/I _6822_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_366 net763_445/I _6844_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5272_ _5165_/Z _5270_/Z _4877_/Z _5425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7011_ _7011_/D _7258_/RN _7011_/CLK _7011_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet713_399 net763_430/I _6775_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_388 net813_469/I _6786_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4223_ hold37/Z hold20/Z _4227_/S _4223_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4154_ hold48/Z hold466/Z _4157_/S _4154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4085_ _4059_/S input68/Z _4085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_102_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4987_ _4367_/Z _5340_/A1 _4555_/B _5172_/B _4987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6726_ _6726_/D _7170_/RN _6726_/CLK _6726_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3938_ _3929_/Z _3938_/A2 _3938_/A3 _3937_/Z _3938_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_176_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6657_ _7235_/RN _6657_/A2 _6657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3869_ _3869_/A1 _3869_/A2 _3869_/A3 _3868_/Z _3869_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6588_ _6834_/Q _6588_/A2 _6588_/B1 _6835_/Q _6836_/Q _6588_/C2 _6589_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5608_ hold20/Z _6969_/Q hold43/Z hold44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5539_ _3485_/Z _5857_/A3 _5821_/A3 _5520_/C _5547_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_132_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _7209_/D _7237_/RN _7209_/CLK _7209_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_154_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4910_ _5442_/A2 _4909_/Z _5443_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5890_ hold20/Z hold500/Z _5892_/S _5890_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _5287_/B _4836_/Z _4841_/B _4841_/C _4846_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_178_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _4782_/A1 _5302_/B _4695_/Z _4700_/Z _4772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_158_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3723_ _3719_/Z _3723_/A2 _3723_/A3 _3723_/A4 _3723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6511_ _6511_/A1 _6511_/A2 _6511_/A3 _6511_/A4 _6511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3654_ _3485_/Z _3653_/Z _3948_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6442_ _6442_/I _6443_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _7217_/Q _6274_/Z _6285_/Z _7193_/Q _7177_/Q _6254_/Z _6385_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3585_ _7221_/Q _3912_/A2 _3959_/C1 _7189_/Q _3589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_170_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5324_ _5324_/A1 _5324_/A2 _5324_/B _5324_/C _5444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_138_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5255_ _5258_/B2 _5255_/A2 _5051_/Z _5255_/B _5446_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_142_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4206_ hold296/Z hold20/Z _4210_/S _4206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _4506_/Z _4700_/Z _5339_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4137_ _3529_/Z _5520_/C hold235/Z _5839_/A3 _4139_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4068_ _6760_/Q _3339_/I _6905_/Q _4068_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6709_ _6709_/D _7218_/RN _6709_/CLK _6709_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_165_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold609 _5851_/Z _7184_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_109_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3370_ _6999_/Q _3370_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _5439_/B1 _5439_/B2 _5040_/B _5040_/C _5044_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _6991_/D _7258_/RN _6991_/CLK _6991_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_65_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5942_ _5943_/I0 _5936_/Z _5942_/S _7234_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5873_ hold12/Z hold174/Z _5874_/S _5873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _4997_/C _4703_/Z _5370_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4755_ _4755_/A1 _5313_/A2 _5233_/A1 _4766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_159_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3706_ _6952_/Q _5584_/A1 _3951_/C1 _7146_/Q _3707_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_175_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _5240_/B _5214_/A2 _4686_/B _4812_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_134_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3637_ input59/Z _4194_/A1 _3917_/A2 _7116_/Q _5528_/S _3619_/Z _3638_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6425_ _6425_/I _6426_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3568_ _3512_/Z _3552_/Z _3941_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6356_ _6356_/A1 _6356_/A2 _6356_/A3 _6355_/Z _6356_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5307_ _4586_/Z _4683_/Z _5302_/B _5307_/B _5480_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_88_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6287_ _6287_/A1 _6287_/A2 _6287_/A3 _6554_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3499_ _3499_/I _3500_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _5238_/A1 _5454_/A1 _5238_/A3 _5238_/A4 _5238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_64_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _5169_/A1 _5425_/A1 _5425_/A3 _5169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_56_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold6 hold6/I hold6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_87_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_138__1359_ clkbuf_4_1_0__1359_/Z net713_383/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _4441_/B _4501_/B _4460_/B _4436_/B _5278_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_129_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _4853_/A1 _4481_/A2 _4735_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold417 _5745_/Z _7090_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold406 _7118_/Q hold406/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3422_ _3422_/I0 input58/Z _6733_/Q _3422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold439 _7034_/Q hold439/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7190_ _7190_/D _7218_/RN _7190_/CLK _7190_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6210_ _6858_/Q _6210_/A2 _6210_/B _6210_/C _6220_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold428 _5507_/Z _6886_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_87_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6141_ _6141_/A1 _5991_/Z _6146_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_48_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3353_ _7129_/Q _3353_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _7121_/Q _5969_/Z _6072_/B _6073_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _5019_/Z _5020_/Z _5023_/A3 _5285_/B _5023_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6974_ _6974_/D _7260_/RN _6974_/CLK _6974_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_53_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ _7228_/Q _7227_/Q _7230_/Q _7229_/Q _5925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_80_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ hold2/Z hold135/Z _5856_/S _5856_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _4422_/Z _4534_/Z _5312_/A1 _5414_/A2 _4807_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_182_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5787_ hold291/Z hold989/Z _5793_/S _5787_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4738_ _4699_/Z _5309_/A2 _4738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4669_ _4397_/Z _5209_/A3 _4997_/C _5464_/A1 _4669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_162_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold940 _5813_/Z _7150_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6408_ _6408_/A1 _6408_/A2 _6408_/A3 _6408_/A4 _6408_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_122_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold951 _6925_/Q hold951/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold962 _4193_/Z _6729_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold973 _7143_/Q hold973/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6339_ _7252_/Q _6339_/I1 _6558_/S _7252_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold995 _6973_/Q hold995/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold984 _7087_/Q hold984/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_62_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_231 net613_258/I _6994_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_220 net613_261/I _7005_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet563_242 net613_254/I _6983_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3971_ _3971_/A1 _3434_/B _6663_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ _3521_/Z _3537_/Z hold24/Z _5718_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_90_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6690_ _6690_/D _7170_/RN _6690_/CLK _6690_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_86_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ hold568/Z hold91/Z _5646_/S _5641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ hold20/Z hold84/Z _5574_/S hold85/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4523_ _4460_/B _4436_/B _5139_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7311_ _7311_/I _7311_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold203 _5819_/Z _7156_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold225 _7051_/Q hold225/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_102_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold214 _6776_/Q hold214/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7242_ _7242_/D _7258_/RN _7260_/CLK _7242_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold247 _5540_/Z _6908_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4454_ _3401_/I _3402_/I _4454_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_104_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold236 _4332_/Z _4334_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold258 _6680_/Q hold258/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold269 _6670_/Q hold269/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4385_ input99/Z input98/Z _4386_/A3 _4386_/A4 _4385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3405_ _4472_/B _4441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_7173_ _7173_/D _7256_/RN _7173_/CLK _7173_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3336_ _7209_/Q _4050_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _6124_/A1 _6124_/A2 _6124_/A3 _6124_/A4 _6124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6055_ _7014_/Q _5971_/Z _5979_/Z _6966_/Q _5996_/Z _7080_/Q _6057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _5389_/C _5170_/A2 _5170_/A3 _5130_/B2 _5347_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41__1359_ net413_93/I _4073__46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _6957_/D _7237_/RN _6957_/CLK _6957_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ _7223_/Q _7224_/Q _7225_/Q _5908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_139_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6888_ _6888_/D _7008_/RN _6888_/CLK _6888_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5839_ hold24/Z _3552_/Z _5839_/A3 _5857_/A3 _5847_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_22_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold770 _4245_/Z _6762_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_122_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold781 _6778_/Q hold781/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_161 net413_79/I _7064_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_183 net413_76/I _7042_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_194 net763_426/I _7031_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_172 _4073__19/I _7053_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold792 _4120_/Z _6674_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_49_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput308 _7333_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput319 _6792_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ _4170_/A1 hold32/Z _4172_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_171_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6811_ _6811_/D _7265_/CLK _6811_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _6742_/D _7218_/RN _6742_/CLK _7322_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3954_ _6988_/Q _3954_/A2 _3954_/B1 input20/Z _4301_/A1 _6809_/Q _3958_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet763_404 net763_434/I _6770_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_415 net763_415/I _6759_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6673_ _6673_/D _7238_/RN _6673_/CLK _6673_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3885_ _3876_/Z _3885_/A2 _3885_/A3 _3884_/Z _3885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_426 net763_426/I _6748_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5624_ hold65/Z hold350/Z _5628_/S _5624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet763_437 net413_55/I _6728_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_448 net763_449/I _6717_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ hold12/Z hold358/Z _5556_/S _5555_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4506_ _4997_/B _4494_/Z _4496_/Z _5263_/A2 _4506_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5486_ _4616_/Z _4855_/C _5487_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_133_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4437_ _4438_/B _4438_/C _4648_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7225_ _7225_/D _7235_/RN _4067_/I1 _7225_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_160_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7156_ _7156_/D _7237_/RN _7156_/CLK _7156_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4368_ _4456_/B _5051_/S _5270_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6107_ _7064_/Q _5985_/Z _5997_/Z _7098_/Q _7170_/Q _6006_/Z _6109_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3319_ _7223_/Q _5900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7087_ _7087_/D _7218_/RN _7087_/CLK _7087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_58_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _6570_/I0 _6807_/Q _4300_/S _6807_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6038_ _6031_/Z _6037_/Z _6336_/B1 _6168_/C _6555_/C _6039_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_67_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3670_ _6703_/Q _3927_/A2 _3952_/A2 _7049_/Q _3673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5340_ _5340_/A1 _5370_/B _5340_/B _5340_/C _5363_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_127_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ _5165_/Z _5270_/Z _4877_/Z _5271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xnet713_378 net713_379/I _6821_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_356 net763_421/I _6854_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_367 net763_445/I _6843_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7010_ _7010_/D _7258_/RN _7010_/CLK _7010_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_389 net813_469/I _6785_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4222_ _4221_/Z hold793/Z _4228_/S _4222_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4153_ hold65/Z hold252/Z _4157_/S _4153_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4084_ _4084_/I0 _4084_/I1 _6732_/Q _7281_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4986_ _4986_/A1 _4980_/Z _4986_/A3 _4993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_177_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6725_ _6725_/D _7170_/RN _6725_/CLK _6725_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3937_ _3937_/A1 _3937_/A2 _3937_/A3 _3903_/Z _3937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6656_ _7235_/RN _6657_/A2 _6656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3868_ _3868_/A1 _3868_/A2 _3868_/A3 _3868_/A4 _3868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6587_ _6587_/I0 _7272_/Q _6602_/S _7272_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5607_ hold48/Z hold460/Z hold43/Z _6968_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3799_ _3798_/Z _3799_/I1 _3899_/S _6870_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5538_ hold751/Z hold291/Z _5538_/S _5538_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5469_ _5469_/A1 _5423_/Z _5469_/A3 _5469_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_133_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7208_ _7208_/D _7237_/RN _7208_/CLK _7208_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7139_ hold74/Z _7260_/RN _7139_/CLK hold73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_100_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4840_ _5281_/B _5132_/A2 _4840_/B1 _5214_/A2 _4841_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_60_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _4467_/B _4463_/Z _4782_/A1 _5302_/B _5236_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_14_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ _6841_/Q _6243_/Z _6288_/Z _7296_/Q _6511_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_33_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3722_ _7194_/Q _3909_/A2 _3948_/C1 _7333_/I _4225_/S _4075_/I1 _3723_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_158_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3653_ _3653_/A1 _3492_/Z _3497_/I hold673/Z _3653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6441_ _6985_/Q _6251_/Z _6273_/Z hold29/I _6265_/Z hold62/I _6442_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6372_ _7169_/Q _5948_/Z _6261_/Z _6959_/Q _6266_/Z hold75/I _6385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5323_ _5323_/A1 _4920_/Z _5322_/Z _5323_/B _5324_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_155_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3584_ _7197_/Q _3909_/A2 _4227_/S input70/Z _4194_/A1 input60/Z _3589_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5254_ _4761_/I _5245_/Z _5254_/B _5254_/C _5257_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_102_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ _5185_/A1 _5185_/A2 _6577_/C _5185_/B2 _6860_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ _4204_/Z hold785/Z _4211_/S _4205_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4136_ hold2/Z hold450/Z _4136_/S _4136_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4067_ _6761_/Q _4067_/I1 _6903_/Q _4067_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _4718_/B _4903_/Z _5072_/A4 _4421_/Z _4969_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_184_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6708_ _6708_/D _7218_/RN _6708_/CLK _6708_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_22_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _7235_/RN _6657_/A2 _6639_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_138_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_300 _4073__51/I _6925_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18__1359_ _4073__7/I _4073__51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_184_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6990_ _6990_/D _7238_/RN _6990_/CLK _6990_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5941_ _5941_/A1 _5940_/Z _5943_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5872_ hold20/Z hold514/Z _5874_/S _5872_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _5270_/A1 _4454_/Z _4997_/C _4554_/Z _4659_/Z _4826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_21_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4754_ _4716_/Z _4752_/Z _5233_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_105_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3705_ _6960_/Q _3957_/A2 _3959_/B1 _6670_/Q _3707_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4685_ _4685_/A1 _4685_/A2 _5180_/A3 _5211_/C _5001_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_146_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3636_ _7196_/Q _3909_/A2 _4227_/S input69/Z _3945_/B1 _7092_/Q _3638_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6424_ _7171_/Q _5948_/Z _6263_/Z hold84/I _6425_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_108_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3567_ _3512_/Z _3529_/Z _5683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6355_ _6355_/A1 _6355_/A2 _6355_/A3 _6355_/A4 _6355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6286_ _6287_/A1 _6287_/A2 _6287_/A3 _6286_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_89_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5306_ _5306_/I _5307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3498_ _7303_/Q input58/Z _6733_/Q _3499_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5237_ _5238_/A1 _5238_/A4 _5457_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _4454_/Z _4997_/C _4820_/Z _4456_/B _5425_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_112_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _5099_/A1 _5099_/A2 _4716_/Z _4784_/Z _4549_/Z _5100_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_83_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4119_ _5520_/C _3533_/Z _5839_/A3 _5857_/A3 _4127_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_17_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_1__f__1062_ clkbuf_0__1062_/Z _6568_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_180_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold7 hold7/I hold7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_48_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_5__1359_ net763_436/I net763_439/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _4463_/Z _4468_/Z _4765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold418 _6678_/Q hold418/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold407 _5777_/Z _7118_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3421_ _3421_/A1 _3421_/A2 _7304_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xhold429 _7128_/Q hold429/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_125_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3352_ _7137_/Q _3352_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6140_ _7026_/Q _6211_/A2 _6211_/B1 _6994_/Q _6141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6071_ _7153_/Q _5960_/Z _5965_/Z _6701_/Q _5981_/Z _6935_/Q _6073_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_58_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _5198_/C _5023_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _6973_/D _7237_/RN _6973_/CLK _6973_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_0_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5924_ _6021_/A2 _6015_/A3 _6014_/A2 _5984_/A1 _5924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5855_ hold12/Z hold198/Z _5856_/S _5855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _4492_/Z _4536_/Z _5319_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5786_ hold227/Z hold767/Z _5793_/S _5786_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4737_ _5226_/C _5226_/B _5309_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4668_ _4411_/Z _5343_/A1 _5393_/A2 _5165_/A4 _5360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_64__1359_ net513_170/I net413_76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_144__1359_ net763_436/I net813_455/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold930 _5822_/Z _7158_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3619_ _7260_/Q _6899_/Q _6900_/Q _3619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6407_ _7072_/Q _6248_/Z _6293_/Z _7154_/Q _6407_/C _6408_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4599_ _5129_/A3 _4598_/Z _5051_/S _4454_/Z _4599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold963 _7183_/Q hold963/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold952 _5559_/Z _6925_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold941 _6682_/Q hold941/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6338_ _6338_/I _6339_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold996 _5613_/Z _6973_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold985 _5742_/Z _7087_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold974 _5805_/Z _7143_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6269_ _7235_/Q _7234_/Q _6302_/A3 _6533_/A2 _6269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_48_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet563_221 net563_221/I _7004_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_210 net763_425/I _7015_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_172_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet563_243 net763_420/I _6982_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_232 net763_422/I _6993_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3970_ _3967_/Z _3970_/A2 _6664_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_189_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ hold656/Z hold291/Z _5646_/S _5640_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5571_ hold48/Z hold147/Z _5574_/S _5571_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _4441_/B _5288_/B _5315_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_129_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7310_ _7310_/I _7310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold226 _7270_/Q hold226/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4453_ _3401_/I _3402_/I _4555_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7241_ _7241_/D _7256_/RN _7258_/CLK _7241_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold204 _7035_/Q hold204/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold215 _4261_/Z _6776_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold248 _7063_/Q hold248/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3404_ _5051_/S _4835_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_116_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold237 _4333_/Z _6839_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold259 _4126_/Z _6680_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4384_ _4376_/Z _4381_/Z _4580_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7172_ _7172_/D _7237_/RN _7172_/CLK _7172_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3335_ _7217_/Q _4049_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ hold58/I _5987_/Z _6015_/Z _7009_/Q _6124_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_100_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6054_ _6934_/Q _5981_/Z _5988_/Z _6982_/Q _7046_/Q _6019_/Z _6057_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_58_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _5043_/A2 _5389_/C _5393_/B1 _5043_/B _5347_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_105_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3340__1 _3340__1/I _6603_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _6956_/D _7258_/RN _6956_/CLK _6956_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_42_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5907_ _5906_/Z _5904_/B _7225_/Q _7225_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6887_ _6887_/D input75/Z _6887_/CLK _6887_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_22_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ hold2/Z hold145/Z _5838_/S _5838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5769_ hold291/Z hold980/Z _5775_/S _5769_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold782 _4264_/Z _6778_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold771 _6884_/Q hold771/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold760 _4349_/Z _6850_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_162 net813_464/I _7063_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_173 net563_221/I _7052_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_195 net763_420/I _7030_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold793 _7310_/I hold793/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_184 net613_266/I _7041_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput309 _7334_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6810_ _6810_/D _7008_/RN _6810_/CLK _6810_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6741_ _6741_/D _7218_/RN _6741_/CLK _7321_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_16_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3953_ _3953_/A1 _3953_/A2 _3953_/A3 _3953_/A4 _3953_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_189_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet763_405 net763_415/I _6769_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3884_ _3884_/A1 _3884_/A2 _3884_/A3 _3884_/A4 _3884_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_52_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _6672_/D _7238_/RN _6672_/CLK _6672_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xnet763_416 net763_418/I _6758_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5623_ hold91/Z hold509/Z _5628_/S _5623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet763_427 net763_427/I _6747_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_438 net763_439/I _6727_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_449 net763_449/I _6716_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5554_ hold20/Z hold516/Z _5556_/S _5554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4505_ _5340_/A1 _4495_/Z _4497_/Z _5262_/A2 _5343_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_145_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5485_ _5480_/Z _5485_/A2 _5485_/B _5490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4436_ _5281_/C _5464_/A1 _4436_/B _4438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7224_ _7224_/D _7235_/RN _4067_/I1 _7224_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_117_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4367_ _4456_/B _5051_/S _4367_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_116_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7155_ hold83/Z _7260_/RN _7155_/CLK hold82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3318_ _6743_/Q _5945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_100_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6106_ _6106_/A1 _6106_/A2 _6106_/A3 _6106_/A4 _6106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7086_ _7086_/D _7218_/RN _7086_/CLK _7086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_58_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _6569_/I0 _6806_/Q _4300_/S _6806_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6037_ _6037_/A1 _6037_/A2 _6037_/A3 _6037_/A4 _6037_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_27_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6939_ _6939_/D _7256_/RN _6939_/CLK _6939_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold590 _7088_/Q hold590/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5270_ _5270_/A1 _4454_/Z _4997_/C _4820_/Z _5270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_5_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet713_368 net713_369/I _6842_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_357 net763_421/I _6853_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_379 net713_379/I _6820_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4221_ _6781_/Q hold48/Z _4227_/S _4221_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4152_ hold91/Z hold537/Z _4157_/S _4152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4083_ _6734_/Q _6731_/Q _4084_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4985_ _4397_/Z _5209_/A3 _4659_/Z _4703_/Z _4985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_63_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6724_ _6724_/D _7170_/RN _6724_/CLK _6724_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3936_ _7028_/Q _5674_/A1 _3936_/B1 _6690_/Q _3937_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_32_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6655_ _7235_/RN _6657_/A2 _6655_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3867_ _7079_/Q _3923_/C1 _3956_/B1 _6713_/Q _3867_/C _3868_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6586_ _6586_/A1 _4313_/Z _6586_/B _6587_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_178_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5606_ hold65/Z hold338/Z hold43/Z _6967_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3798_ _6566_/I0 _6869_/Q _3898_/S _3798_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5537_ hold893/Z _4103_/I _5538_/S _5537_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _5468_/A1 _5468_/A2 _5468_/B1 _4650_/Z _5468_/C _5469_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_105_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ _7207_/D _7218_/RN _7207_/CLK _7207_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4419_ _5420_/A3 _5420_/A2 _4456_/B _4419_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_132_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5399_ _4524_/Z _5399_/A2 _4683_/Z _5302_/B _5399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_87_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7138_ _7138_/D _7238_/RN _7138_/CLK hold99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_143_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7069_ _7069_/D _7218_/RN _7069_/CLK _7069_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _4770_/A1 _5118_/A3 _4770_/A3 _5117_/A1 _4775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_174_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _6678_/Q _3546_/Z _3916_/A2 _7154_/Q _7170_/Q _3941_/B1 _3723_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3652_ input68/Z _4227_/S _4244_/S input40/Z _3657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6440_ _6440_/A1 _6440_/A2 _6440_/A3 _6439_/Z _6440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _7063_/Q _6257_/Z _6299_/Z _7055_/Q _6383_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3583_ _6971_/Q _3924_/A2 _3607_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_61_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5322_ _4436_/B _4494_/Z _5328_/A2 _5056_/C _5322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _5254_/C _5334_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5184_ _6834_/Q _5182_/Z _5184_/B _5184_/C _5185_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4204_ hold618/Z hold48/Z _4210_/S _4204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ hold12/Z hold511/Z _4136_/S _4135_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ _6762_/Q user_clock _6904_/Q _4066_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ _4903_/Z _5072_/A4 _4718_/B _4666_/Z _4968_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_51_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4899_ _6577_/C _4899_/A2 _5000_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6707_ _6707_/D _7218_/RN _6707_/CLK _6707_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3919_ _3919_/A1 _3919_/A2 _3919_/A3 _3919_/A4 _3919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6638_ _7235_/RN _6657_/A2 _6638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_164_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _6569_/I0 _7267_/Q _6571_/S _7267_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_301 net413_72/I _6924_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__2 _4073__3/I _7297_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _6745_/Q _7233_/Q _7232_/Q _7234_/Q _5940_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5871_ hold48/Z hold424/Z _5874_/S _5871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4822_ _4554_/Z _4659_/Z _4820_/Z _5364_/B _4826_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_33_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4753_ _4700_/Z _4752_/Z _5313_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ hold99/I _3951_/A2 _3901_/A2 _6984_/Q input30/Z _3927_/C2 _3707_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_175_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4684_ _4414_/Z _4452_/Z _4666_/Z _4892_/B _4683_/Z _4685_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_119_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6423_ _7099_/Q _6250_/Z _6439_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_174_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3635_ input50/Z _4210_/S _3947_/A2 _7100_/Q _3638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6354_ _7168_/Q _5948_/Z _6261_/Z _6958_/Q _6355_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3566_ _3507_/Z _3533_/Z _3954_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6285_ _6484_/A2 _6285_/A2 _7237_/Q _6452_/A4 _6285_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5305_ _4586_/Z _4673_/Z _5302_/B _5305_/B _5306_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3497_ _3497_/I _3617_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_130_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5236_ _4510_/Z _5414_/A2 _5236_/B _5238_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_124_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _4546_/Z _4651_/Z _4675_/Z _5167_/B _5425_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_97_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ _5098_/A1 _5302_/B _5098_/B _5098_/C _5101_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_57_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4118_ hold2/Z hold163/Z _4118_/S _4118_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4049_ _4049_/I0 input92/Z _4050_/S _4049_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_24__1359_ net613_298/I net413_99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_84_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104__1359_ clkbuf_4_5_0__1359_/Z net613_262/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_87__1359_ net513_175/I net613_255/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold8 hold8/I hold8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_181_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold408 _6896_/Q hold408/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3420_ _3988_/S _3422_/I0 _3421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_172_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold419 _4124_/Z _6678_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3351_ _7145_/Q _3351_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6070_ _6951_/Q _5958_/Z _5967_/Z _7105_/Q _7137_/Q _5994_/I _6073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _4604_/Z _4606_/Z _5003_/Z _5021_/B _5198_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _6972_/D _7218_/RN _6972_/CLK _6972_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_19_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5923_ _7230_/Q _7229_/Q _6210_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_94_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5854_ hold20/Z hold367/Z _5856_/S _5854_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _4835_/A2 _4492_/Z _4534_/Z _4681_/Z _4805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5785_ _5520_/C _3552_/Z _5857_/A3 _5857_/A2 _5793_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_148_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _4736_/A1 _5302_/B _4736_/A3 _4467_/B _5226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4667_ _4414_/Z _5038_/A1 _4557_/Z _4666_/Z _4667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_135_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold931 _6904_/Q hold931/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3618_ _3527_/Z _3617_/Z _5528_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold920 _5759_/Z _7102_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6406_ _6406_/I _6407_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6337_ _6744_/Q _7251_/Q _6337_/B _6338_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4598_ _5287_/B _4460_/B _5399_/A2 _4436_/B _4598_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_116_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold964 _5850_/Z _7183_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold953 _7095_/Q hold953/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold942 _4129_/Z _6682_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3549_ _3485_/Z _3512_/Z _4194_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold986 _7199_/Q hold986/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold975 _7053_/Q hold975/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold997 _6873_/Q hold997/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6268_ _7233_/Q _7232_/Q _6533_/A2 _6452_/A4 _6268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_135_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _5303_/A1 _5303_/A3 _5224_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ _6789_/Q _5972_/Z _6021_/Z _6839_/Q _6201_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_84_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_222 net563_222/I _7003_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_211 net563_222/I _7014_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_233 net613_279/I _6992_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_244 net813_467/I _6981_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70__1359_ net513_175/I net763_426/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ hold65/Z hold612/Z _5574_/S _5570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ _4472_/B _4501_/B _5139_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4452_ _5038_/A1 _4648_/B _4638_/A2 _4452_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7240_ _7240_/D _7256_/RN _4067_/I1 _7240_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold216 _7130_/Q hold216/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold205 _6990_/Q hold205/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold249 _5714_/Z _7063_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3403_ _4456_/B _5129_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xhold227 _4102_/Z hold227/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold238 _6672_/Q hold238/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4383_ _5464_/A1 _4383_/A2 _5385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_171_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _7171_/D _7258_/RN _7171_/CLK _7171_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3334_ _3334_/I _4029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _7091_/Q _6002_/Z _6003_/Z _7163_/Q _6124_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_140_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6053_ _6053_/A1 _6053_/A2 _6053_/A3 _6053_/A4 _6053_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _5368_/A1 _5420_/A1 _5002_/Z _5389_/B _5191_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6955_ _6955_/D _7260_/RN _6955_/CLK _6955_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5906_ _7223_/Q _7224_/Q _5910_/B _5906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6886_ _6886_/D input75/Z _6886_/CLK _6886_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5837_ hold12/Z hold721/Z _5838_/S _5837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ hold227/Z hold643/Z _5775_/S _5768_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4719_ _5083_/B _4719_/A2 _4721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_175_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5699_ hold12/Z hold610/Z hold25/Z _7050_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_152 net513_163/I _7073_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold750 _5889_/Z _7218_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold772 _5505_/Z _6884_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold761 _6691_/Q hold761/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_157_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_163 net513_163/I _7062_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_174 net613_263/I _7051_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold783 _7321_/I hold783/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_77_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_185 net513_189/I _7040_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold794 _4222_/Z _6751_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_162_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_196 net563_221/I _7029_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _6740_/D _7218_/RN _6740_/CLK _7320_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3952_ _7044_/Q _3952_/A2 _5638_/A1 _6996_/Q _6948_/Q _5584_/A1 _3953_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet763_406 net763_406/I _6768_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3883_ input53/Z _4194_/A1 _3948_/C1 input62/Z _3941_/B1 _7167_/Q _3884_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6671_ _6671_/D _7238_/RN _6671_/CLK _6671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_31_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet763_417 net763_417/I _6757_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_428 net763_431/I _6742_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5622_ hold291/Z hold773/Z _5628_/S _5622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet763_439 net763_439/I _6726_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5553_ hold48/Z hold411/Z _5556_/S _5553_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4504_ _4759_/A2 _4759_/A3 _4504_/B _4504_/C _5263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_145_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5484_ _5483_/Z _5450_/I _5477_/Z _5441_/B _5485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_133_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4435_ _5281_/C _5270_/A1 _5170_/A2 _4436_/B _4438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7223_ _7223_/D _7235_/RN _4067_/I1 _7223_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4366_ _4472_/B _4460_/B _4436_/B _4853_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7154_ _7154_/D input75/Z _7154_/CLK _7154_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3317_ _6836_/Q _4686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_141_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6105_ _7114_/Q _5984_/Z _6000_/Z _7130_/Q _6106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_59_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7085_ _7085_/D _7256_/RN _7085_/CLK _7085_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4297_ _6568_/I0 _6805_/Q _4300_/S _6805_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _6973_/Q _5964_/Z _5984_/Z _7111_/Q _6036_/C _6037_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6938_ _6938_/D _7256_/RN _6938_/CLK _6938_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _6869_/D _6627_/Z _4075_/I1 _6869_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_22_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold580 _7309_/I hold580/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_173_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold591 _5743_/Z _7088_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_358 net813_483/I _6852_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_369 net713_369/I _6841_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4220_ _4219_/Z hold580/Z _4228_/S _4220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4151_ hold291/Z hold849/Z _4157_/S _4151_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _4082_/A1 _7299_/Q _4082_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4984_ _4700_/Z _4982_/Z _4984_/B _4986_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6723_ _6723_/D input75/Z _6723_/CLK _6723_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3935_ _6924_/Q _3935_/A2 _3935_/B1 _6849_/Q _3937_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_189_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _7235_/RN _4064_/S _6654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_108_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3866_ _3866_/A1 _3537_/Z _3617_/Z _3866_/B _3867_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5605_ hold91/Z hold167/Z hold43/Z _6966_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6585_ _6834_/Q _6585_/A2 _6585_/B1 _6835_/Q _6836_/Q _6585_/C2 _6586_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3797_ _3776_/Z _3797_/A2 _3797_/A3 _3796_/Z _6566_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_118_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5536_ _5536_/A1 hold32/Z _5538_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_172_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _4570_/Z _4651_/Z _5467_/B _5467_/C _5468_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_117_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4418_ _5170_/A2 _4456_/B _5343_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_160_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ _7206_/D _7008_/RN _7206_/CLK _7206_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5398_ _5391_/Z _5398_/A2 _5419_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7137_ _7137_/D _7238_/RN _7137_/CLK _7137_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4349_ hold291/Z hold759/Z _4349_/S _4349_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7068_ _7068_/D _7218_/RN _7068_/CLK _7068_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_115_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _7228_/Q _7227_/Q _6211_/A2 _6210_/A2 _6019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _7114_/Q _3917_/A2 _3947_/A2 _7098_/Q _3945_/A2 _7178_/Q _3723_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_187_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3651_ _7187_/Q _3959_/C1 _3960_/A2 _7211_/Q _3657_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6370_ _6991_/Q _6237_/Z _6380_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3582_ _3509_/Z _3515_/Z _3924_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_161_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5321_ _5321_/A1 _5212_/Z _5454_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5252_ _5343_/A1 _5343_/A2 _5255_/A2 _5252_/B _5254_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_115_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ _4202_/Z hold819/Z _4211_/S _4203_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5183_ _5181_/Z _4686_/B _5299_/C _5184_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_68_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ hold20/Z hold531/Z _4136_/S _4134_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _6392_/B1 input2/Z input1/Z _4065_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4967_ _4903_/Z _5072_/A4 _4718_/B _5359_/A1 _4967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4898_ _3401_/I _4893_/Z _4898_/B _4898_/C _4899_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6706_ _6706_/D _7170_/RN _6706_/CLK _6706_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3918_ input36/Z _4225_/S _4143_/A1 _6694_/Q _3919_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_165_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6637_ _7235_/RN _6657_/A2 _6637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3849_ _7175_/Q _3945_/A2 _3939_/C1 _6711_/Q _3897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _6568_/I0 _7266_/Q _6571_/S _7266_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_47__1359_ net663_324/I net413_97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ _7307_/I hold321/Z _5520_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_173_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6499_ _6554_/A1 _6499_/A2 _6499_/A3 _6498_/Z _6499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__3 _4073__3/I _7296_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0__1359_ clkbuf_0__1359_/Z net413_62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_129_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ hold65/Z hold535/Z _5874_/S _5870_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ _4554_/Z _4472_/B _4887_/A1 _4501_/B _4821_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4752_ _5302_/B _4436_/B _4463_/Z _5226_/C _4752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4683_ _5420_/A3 _4835_/A2 _4456_/B _3402_/I _4683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3703_ input48/Z _4210_/S _4244_/S input39/Z _3708_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3634_ _7220_/Q _3912_/A2 _4244_/S input41/Z _3930_/A2 _7132_/Q _3638_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_88_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6422_ hold60/I _6257_/Z _6434_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_175_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _7208_/Q _6256_/Z _6285_/Z _7192_/Q _6274_/Z _7216_/Q _6355_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3565_ _3509_/Z _3542_/Z _3901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3496_ _3495_/Z hold233/Z hold54/Z _3496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6284_ _6281_/Z _6283_/Z _6251_/Z _6273_/Z _6287_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ _4683_/Z _5302_/B _5456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_130_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5235_ _5316_/A2 _5234_/Z _5238_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_69_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5166_ _5166_/A1 _5467_/B _5166_/A3 _5165_/Z _5169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_96_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4117_ hold1/Z _7277_/Q hold54/I hold2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_151_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5097_ _5097_/A1 _5328_/A2 _5368_/B _3401_/I _5098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_110_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4048_ _6767_/Q input89/Z _4050_/S _4048_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ _6211_/A2 _6021_/A2 _6210_/A2 _7227_/Q _5999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_166_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput290 _6685_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_94_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 hold9/I hold9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_47_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold409 _7000_/Q hold409/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_174_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3350_ _7153_/Q _3350_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_30__1359_ net613_298/I net763_406/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_110__1359_ net513_165/I net413_88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_93__1359_ clkbuf_4_5_0__1359_/Z net513_200/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5020_ _5438_/C _5359_/A1 _4604_/Z _4606_/Z _5020_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_97_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6971_ _6971_/D _7258_/RN _6971_/CLK _6971_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ _5922_/I _7229_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5853_ hold48/Z hold480/Z _5856_/S _5853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _4681_/Z _4793_/Z _5319_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5784_ hold2/Z hold312/Z _5784_/S _5784_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _4501_/B _4735_/A2 _4764_/A3 _5226_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_174_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _5420_/A3 _5420_/A2 _4835_/A2 _4456_/B _4666_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4597_ _5287_/B _4596_/Z _5420_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3617_ _3617_/A1 hold673/Z _3489_/I _3492_/Z _3617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold921 _7166_/Q hold921/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold910 _6613_/Z _7297_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6405_ hold99/I _6253_/Z _6297_/Z _6702_/Q _6406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold932 _5534_/Z _6904_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold943 _7207_/Q hold943/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3548_ _3519_/Z _3533_/Z _3945_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6336_ _6329_/Z _6335_/Z _6336_/B1 _6286_/Z _6555_/C _6337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold954 _5751_/Z _7095_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold987 _5868_/Z _7199_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold976 _5703_/Z _7053_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold998 _6871_/Q hold998/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold965 _6683_/Q hold965/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3479_ _6659_/Q _6658_/Q _6733_/Q _3479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _6996_/Q _6265_/Z _6266_/Z _7012_/Q _6271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5218_ _4673_/Z _4700_/Z _5218_/B _5303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_97_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _6198_/A1 _6198_/A2 _6198_/A3 _6198_/A4 _6198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5149_ _5165_/A2 _4598_/Z _5374_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_212 net613_256/I _7013_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_234 net613_255/I _6991_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_223 net713_394/I _7002_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_245 net563_245/I _6980_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_153_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _4835_/A2 _4456_/B _3402_/I _3401_/I _5359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_11_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _4604_/A2 _4604_/A3 _4451_/B _4451_/C _5038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold217 _5790_/Z _7130_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold206 _5632_/Z _6990_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3402_ _3402_/I _5420_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xhold239 _4116_/Z _6672_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7170_ _7170_/D _7170_/RN _7170_/CLK _7170_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold228 _5639_/Z _6996_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4382_ _4472_/B _4501_/B _4460_/B _4436_/B _4383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _6985_/Q _5988_/Z _6019_/Z _7049_/Q _6124_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3333_ _4483_/B _4424_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_112_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6052_ _6950_/Q _5958_/Z _5967_/Z _7104_/Q _6052_/C _6053_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _5165_/A4 _5003_/A2 _4421_/Z _4491_/B _5003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_67_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0__1062_ _3725_/ZN clkbuf_0__1062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6954_ hold51/Z _7238_/RN _6954_/CLK hold50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_26_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5905_ _5905_/I _7224_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _6885_/D input75/Z _6885_/CLK _6885_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5836_ hold20/Z hold400/Z _5838_/S _5836_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5767_ _5857_/A3 _5839_/A3 _3537_/Z _5520_/C _5775_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_50_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4718_ _4504_/B _4504_/C _4718_/B _5056_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_108_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5698_ hold20/Z _7049_/Q hold25/Z hold26/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4649_ _4570_/Z _5438_/B _4653_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_89_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold740 _4328_/Z _6825_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold751 _6907_/Q hold751/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold773 _6981_/Q hold773/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold762 _4139_/Z _6691_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7299_ _7299_/D _6651_/Z _7304_/CLK _7299_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold795 _7314_/I hold795/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_186 _4073__5/I _7039_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_175 net513_175/I _7050_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold784 _4209_/Z _6741_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6319_ _7127_/Q _6484_/A2 _6533_/A3 _7111_/Q _6320_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet513_164 net413_57/I _7061_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_153 net513_153/I _7072_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_197 _4073__39/I _7028_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3951_ _7134_/Q _3951_/A2 _5665_/A1 _7020_/Q _3951_/C1 _7142_/Q _3953_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_177_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3882_ _6925_/Q _3935_/A2 _3933_/B1 _6786_/Q _3942_/C1 _6854_/Q _3884_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6670_ _6670_/D _7238_/RN _6670_/CLK _6670_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_31_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_418 net763_418/I _6756_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_407 net763_431/I _6767_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_429 net763_431/I _6741_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ hold227/Z hold431/Z _5628_/S _5621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5552_ hold65/Z hold458/Z _5556_/S _5552_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4503_ _4718_/B _5072_/A4 _5262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5483_ _5483_/A1 _5483_/A2 _5483_/A3 _5483_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7222_ _7222_/D _7235_/RN _4067_/I1 _7222_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4434_ _4467_/B _4460_/B _4887_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_132_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4365_ _4472_/B _4460_/B _4436_/B _5288_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_160_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7153_ _7153_/D _7237_/RN _7153_/CLK _7153_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3316_ _6835_/Q _4415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_141_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7084_ _7084_/D _7237_/RN _7084_/CLK _7084_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6104_ _7106_/Q _5967_/Z _5980_/Z _7072_/Q _5969_/Z _7122_/Q _6106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_140_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6035_ _6035_/I _6036_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _6567_/I0 _6804_/Q _4300_/S _6804_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6937_ hold85/Z _7260_/RN _6937_/CLK hold84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6868_ _6868_/D _6626_/Z _4075_/I1 _6868_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_167_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5819_ hold12/Z hold202/Z _5820_/S _5819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6799_ _6799_/D input75/Z _6799_/CLK _6799_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_136_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold570 _6685_/Q hold570/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold581 _4220_/Z _6750_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold592 _6753_/Q hold592/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_65_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet713_359 net813_453/I _6851_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150_ hold227/Z hold398/Z _4157_/S _4150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4081_ _4081_/A1 input73/Z _4081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_49_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4983_ _5083_/C _4659_/Z _4703_/Z _4422_/Z _4984_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_51_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6722_ _6722_/D input75/Z _6722_/CLK _6722_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3934_ _7004_/Q _3934_/A2 _3934_/B1 _6845_/Q _5532_/A1 _6905_/Q _3937_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6653_ _7235_/RN _6653_/A2 _6653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_176_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3865_ _6900_/Q _5528_/S _6611_/A1 _7297_/Q _3868_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_149_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5604_ hold291/Z hold971/Z hold43/Z _6965_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6584_ _6584_/I0 _7271_/Q _6602_/S _7271_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3796_ _3796_/A1 _3796_/A2 _3786_/Z _3795_/Z _3796_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5535_ hold935/Z _4102_/Z _5535_/S _5535_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5466_ _5425_/Z _5428_/Z _5429_/Z _5465_/Z _5466_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4417_ _5129_/A3 _4835_/A2 _4836_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_133_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7205_ _7205_/D _7237_/RN _7205_/CLK _7205_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5397_ _5433_/A2 _5433_/A3 _5434_/A2 _5209_/Z _5398_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_114_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7136_ _7136_/D _7260_/RN _7136_/CLK _7136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_28_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4348_ _4103_/I hold683/Z _4349_/S _4348_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7067_ _7067_/D _7235_/RN _7067_/CLK _7067_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4279_ hold291/Z hold741/Z _4279_/S _4279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _7143_/Q _7231_/Q _6210_/B _6068_/A4 _6024_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3650_ _7195_/Q _3909_/A2 _4194_/A1 input57/Z _3955_/A2 _7203_/Q _3689_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3581_ _3523_/Z _3533_/Z _3925_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5320_ _5320_/A1 _5319_/Z _5452_/A2 _5453_/A4 _5320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5251_ _5330_/B2 _5246_/Z _5251_/B _5254_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_170_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4202_ hold478/Z hold65/Z _4210_/S _4202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5182_ _5182_/A1 _5340_/C _5265_/A4 _4511_/Z _5182_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_142_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4133_ hold48/Z hold544/Z _4136_/S _4133_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4064_ _6392_/B1 _7281_/Q _4064_/S _4064_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4966_ _4966_/A1 _4966_/A2 _5073_/B _4970_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6705_ _6705_/D _7237_/RN _6705_/CLK _6705_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_40_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4897_ _6834_/Q _6835_/Q _6836_/Q _4897_/A4 _4898_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3917_ _7110_/Q _3917_/A2 _6611_/A1 _7296_/Q _3919_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _7235_/RN _4064_/S _6636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3848_ _7127_/Q _3930_/A2 _3920_/B1 _6867_/Q _3922_/B1 _6693_/Q _3897_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3779_ _6982_/Q _3901_/A2 _3927_/B1 _7062_/Q _3796_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6567_ _6567_/I0 _7265_/Q _6571_/S _7265_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5518_ _4103_/I hold703/Z _5518_/S _5518_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _6498_/A1 _6498_/A2 _6498_/A3 _6498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5449_ _5449_/A1 _5342_/I _5416_/I _5449_/A4 _5450_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_133_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7119_ _7119_/D _7008_/RN _7119_/CLK _7119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_28_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/Z _4072_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__4 _4073__9/I _7221_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _4489_/B _4483_/B _4026_/B _4026_/C _4820_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_53__1359_ net663_324/I net813_461/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_133__1359_ net513_165/I net813_489/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _4751_/A1 _4748_/Z _4750_/Z _4755_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_187_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4682_ _4530_/I _4878_/A2 _5312_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3702_ _7218_/Q _3912_/A2 _4194_/A1 input56/Z _3941_/A2 _7162_/Q _3708_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_147_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6421_ _7255_/Q _6421_/I1 _6558_/S _7255_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3633_ _6978_/Q _3923_/A2 _3960_/A2 _7212_/Q _3633_/C _3646_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_175_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3564_ _3515_/Z _3537_/Z _3945_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6352_ _6990_/Q _6237_/Z _6240_/Z _7112_/Q _6352_/C _6356_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3495_ _7304_/Q _7303_/Q _6733_/Q _3495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6283_ _6241_/Z _6275_/Z _6282_/Z _6283_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_115_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5303_ _5303_/A1 _5303_/A2 _5303_/A3 _5303_/A4 _5303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_130_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5234_ _5234_/A1 _5314_/A1 _5404_/A1 _5234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5165_ _5209_/A3 _5165_/A2 _4651_/Z _5165_/A4 _5165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_130_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4116_ hold12/Z hold238/Z _4118_/S _4116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _4539_/I _5287_/B _4673_/Z _4460_/B _5098_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_83_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4047_ _6768_/Q input91/Z _4050_/S _4047_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _7078_/Q _5996_/Z _5997_/Z _7094_/Q _6008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_185_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4949_ _5464_/A1 _4944_/Z _5065_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _7235_/RN _6653_/A2 _6619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_138_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput280 _6668_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput291 _6686_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _6970_/D _7258_/RN _6970_/CLK _6970_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_66_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5921_ _5920_/Z _6745_/Q _7229_/Q _5913_/I _5922_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_53_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5852_ hold65/Z hold523/Z _5856_/S _5852_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _4803_/A1 _4797_/Z _4803_/B _4809_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5783_ hold12/Z hold446/Z _5784_/S _5783_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4734_ _4703_/Z _4728_/Z _5106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_148_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _5170_/A2 _4878_/A2 _5389_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4596_ _5288_/B _4460_/B _4436_/B _4472_/B _4596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold911 _7121_/Q hold911/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3616_ _5857_/A2 hold235/I _5521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold922 _5831_/Z _7166_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold900 _4184_/Z _6723_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6404_ _7202_/Q _6272_/Z _6275_/Z _7040_/Q _6296_/Z _7162_/Q _6408_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_150_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold933 _6927_/Q hold933/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3547_ _3485_/Z _3523_/Z _3960_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold944 _5877_/Z _7207_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6335_ _6554_/A1 _6335_/A2 _6335_/A3 _6335_/A4 _6335_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold955 _7103_/Q hold955/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold988 _6957_/Q hold988/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold977 _7037_/Q hold977/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold966 _4130_/Z _6683_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3478_ _3478_/I0 hold5/Z hold54/I hold6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6266_ _6300_/A2 _6533_/A4 _6285_/A2 _6302_/A4 _6266_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_88_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold999 _6874_/Q hold999/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5217_ _5460_/A1 _5460_/A4 _5224_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6197_ _6722_/Q _5987_/Z _6015_/Z _6841_/Q _6198_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5148_ _5147_/Z _5139_/Z _5148_/A3 _5470_/A3 _5148_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5079_ _5079_/A1 _5258_/C _5086_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_151_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_202 net613_258/I _7023_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_213 net413_78/I _7012_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_246 net563_246/I _6979_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet563_235 net613_284/I _6990_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_224 net413_78/I _7001_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_153_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4450_ _4607_/A1 _4451_/B _4451_/C _5356_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_129_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold207 _7003_/Q hold207/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4381_ _4472_/B _4501_/B _4460_/B _4436_/B _4381_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3401_ _3401_/I _5420_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_116_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold218 _6971_/Q hold218/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold229 _6789_/Q hold229/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3332_ _4402_/B _4489_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_6120_ _7017_/Q _5971_/Z _6005_/Z _7041_/Q _6124_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_140_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _6051_/A1 _6051_/A2 _6051_/B1 _5991_/Z _6052_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_5002_ _4411_/Z _5258_/B2 _5002_/A3 _5002_/A4 _5002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_67_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ hold72/Z _7238_/RN _6953_/CLK hold71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ _7224_/Q _5903_/Z _5904_/B _5905_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6884_ _6884_/D input75/Z _6884_/CLK _6884_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_22_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ hold48/Z hold139/Z _5838_/S _5835_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5766_ hold143/Z hold2/Z _5766_/S _5766_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4717_ _5222_/A1 _4716_/Z _5223_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5697_ hold48/Z hold492/Z hold25/Z _7048_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4648_ _4648_/A1 _4648_/A2 _4648_/B _5356_/C _5438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_135_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold730 _4276_/Z _6788_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_30_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4579_ _4380_/Z _4579_/A2 _4451_/B _4451_/C _5345_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold741 _6790_/Q hold741/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold752 _5538_/Z _6907_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold763 _6844_/Q hold763/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7298_ _7298_/D _6650_/Z _7305_/CLK _7298_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_157_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_154 net513_163/I _7071_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold796 _4239_/Z _6759_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_118_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold785 _7319_/I hold785/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6318_ _7199_/Q _6272_/Z _6293_/Z _7151_/Q _6318_/C _6322_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold774 _5622_/Z _6981_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_165 net513_165/I _7060_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_176 net763_422/I _7049_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_187 _4073__25/I _7038_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_198 net613_255/I _7027_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6249_ _7126_/Q _6247_/Z _6248_/Z _7068_/Q _6259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_57_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold90 hold90/I hold90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_48_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ _6726_/Q _4188_/A1 _3950_/B1 _6724_/Q _3950_/C1 _6843_/Q _3953_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_35_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3881_ _7037_/Q _5683_/A1 _5674_/A1 _7029_/Q _3881_/C _3884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xnet763_419 net763_419/I _6755_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5620_ hold24/Z _3542_/Z hold42/Z hold6/Z _5628_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet763_408 net763_444/I _6766_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5551_ hold91/Z hold448/Z _5556_/S _5551_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4502_ _4504_/B _4504_/C _5072_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_145_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5482_ _5482_/A1 _5482_/A2 _5483_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7221_ _7221_/D _7237_/RN _7221_/CLK _7221_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4433_ _4648_/A1 _4648_/A2 _4638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4364_ _4460_/B _4436_/B _5315_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7152_ _7152_/D _7256_/RN _7152_/CLK _7152_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3315_ _6834_/Q _4900_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_4295_ _6566_/I0 _6803_/Q _4300_/S _6803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7083_ hold79/Z _7260_/RN _7083_/CLK hold78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6103_ _6702_/Q _5965_/Z _6014_/Z _6960_/Q _6106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_112_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6034_ _7029_/Q _5999_/Z _6014_/Z _6957_/Q _6000_/Z _7127_/Q _6035_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_132_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _6936_/D _7238_/RN _6936_/CLK _6936_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _6867_/D _7218_/RN _6867_/CLK _6867_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6798_ _6798_/D _7265_/CLK _6798_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5818_ hold20/Z hold82/Z _5820_/S hold83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5749_ _5857_/A3 _5821_/A3 _3537_/Z _5520_/C _5757_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_157_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold560 _7081_/Q hold560/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold571 _4132_/Z _6685_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold593 _4226_/Z _6753_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold582 _7308_/I hold582/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ input85/Z input58/Z _7300_/Q _4080_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4982_ _4997_/B _4495_/Z _5263_/A2 _4436_/B _4982_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_63_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3933_ _7222_/Q _5528_/S _3933_/B1 _6785_/Q _3933_/C _3938_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6721_ _6721_/D _7170_/RN _6721_/CLK _6721_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3864_ _6723_/Q _4182_/A1 _3946_/A2 _6721_/Q input12/Z _3913_/A2 _3868_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6652_ _7170_/RN _6652_/A2 _6652_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ _4102_/Z hold857/Z hold43/Z _5603_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6583_ _6583_/A1 _4313_/Z _6583_/B _6584_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_176_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ _3795_/A1 _3790_/Z _3794_/Z _3795_/A4 _3795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ hold931/Z hold291/Z _5535_/S _5534_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5465_ _5465_/A1 _5170_/Z _4882_/Z _4881_/Z _5465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7204_ _7204_/D _7237_/RN _7204_/CLK _7204_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4416_ _4456_/B _5051_/S _5104_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ _5396_/A1 _5395_/Z _5434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7135_ _7135_/D _7238_/RN _7135_/CLK _7135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_98_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4347_ _5520_/C _3529_/Z _5513_/A3 _5821_/A3 _4349_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7066_ _7066_/D _7235_/RN _7066_/CLK _7066_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4278_ hold227/Z hold229/Z _4279_/S _4278_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6017_ _7167_/Q _6006_/Z _6030_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_2006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/Z _3340__1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6919_ _6919_/D _7258_/RN _6919_/CLK _6919_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold390 _6940_/Q hold390/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3580_ _3505_/Z _3509_/Z _5575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_142_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5250_ _5250_/A1 _5247_/Z _5248_/Z _5250_/A4 _5251_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_142_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4201_ _4200_/Z hold823/Z _4211_/S _4201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_13__1359_ clkbuf_4_2_0__1359_/Z net413_74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5181_ _5127_/Z _5181_/A2 _5321_/A1 _5242_/A3 _5181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_76__1359_ net513_167/I net613_287/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_69_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4132_ hold65/Z hold570/Z _4136_/S _4132_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4063_ _6747_/Q input3/Z input1/Z _4063_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _5464_/A1 _4908_/Z _5073_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6704_ _6704_/D _7235_/RN _6704_/CLK _6704_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3916_ _7150_/Q _3916_/A2 _3916_/B1 _6878_/Q _4274_/A1 _6787_/Q _3919_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_33_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4896_ _4554_/Z _4892_/B _4897_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6635_ _7235_/RN _4064_/S _6635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3847_ _3552_/Z _3653_/Z _4170_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3778_ input37/Z _4244_/S _3948_/C1 input63/Z _3797_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6566_ _6566_/I0 _7264_/Q _6571_/S _7264_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5517_ _5821_/A3 _3533_/Z hold235/Z _5520_/C _5518_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_161_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6497_ _7035_/Q _6269_/Z _6273_/Z _6979_/Q _6498_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5448_ _5448_/A1 _5483_/A2 _5448_/A3 _5463_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_154_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5379_ _5469_/A1 _5379_/A2 _5377_/Z _5379_/A4 _5379_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_120_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _7118_/D _7008_/RN _7118_/CLK _7118_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_102_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ hold26/Z _7260_/RN _7049_/CLK _7049_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_47_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__5 _4073__5/I _7220_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _5302_/B _5099_/A1 _4703_/Z _5226_/C _4750_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_61_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0__1359_ net763_436/I net763_444/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4681_ _5420_/A3 _3402_/I _4456_/B _4681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3701_ _3701_/A1 _3701_/A2 _3701_/A3 _3701_/A4 _3701_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6420_ _6420_/I _6421_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3632_ _3632_/I _3633_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6351_ _6351_/I _6352_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5302_ _4536_/Z _5283_/B _5302_/B _5303_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_108_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3563_ _3537_/Z _3542_/Z _5758_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6282_ _6282_/A1 _6282_/A2 _7232_/Q _6452_/A4 _6282_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3494_ _3653_/A1 hold320/Z _5857_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_88_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ _5233_/A1 _4757_/I _5156_/B _5233_/A4 _5404_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5164_ _5315_/A1 _5315_/A2 _5287_/B _4784_/Z _5467_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4115_ hold11/Z _7276_/Q hold54/I hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_110_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _5278_/C _5302_/B _4784_/Z _4716_/Z _4697_/Z _5460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_68_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _4046_/I _6832_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _7231_/Q _6117_/A4 _6014_/A2 _7229_/Q _5997_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_12_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4948_ _4948_/A1 _4945_/Z _4946_/Z _4947_/Z _4953_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_178_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ _5315_/A2 _4524_/Z _4546_/Z _4820_/Z _4879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_71_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6618_ _7235_/RN _6657_/A2 _6618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_166_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _6846_/Q _6235_/Z _6243_/Z _6842_/Q _6265_/Z _6840_/Q _6554_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xoutput270 _6885_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput281 _6669_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput292 _6687_/Q pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_75_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _7229_/Q _6210_/B _5920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ hold91/Z hold608/Z _5856_/S _5851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _5453_/A4 _5420_/A3 _5456_/A1 _5130_/B1 _5129_/A2 _5389_/A1 _4803_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_21_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ hold20/Z hold76/Z _5784_/S hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4733_ _4733_/A1 _4729_/Z _4731_/Z _4732_/Z _4739_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_187_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _4664_/A1 _4664_/A2 _4663_/Z _4670_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6403_ _7114_/Q _6240_/Z _6403_/B _6408_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_174_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4595_ _5190_/A2 _5364_/B _4568_/Z _5435_/A2 _4595_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_128_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3615_ _5857_/A2 _5857_/A3 hold42/I _3477_/Z _3866_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold912 _5780_/Z _7121_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold901 _6800_/Q hold901/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_31_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold934 _5561_/Z _6927_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3546_ _3489_/I _3492_/Z _3904_/A4 _3904_/A2 _3546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold945 _7167_/Q hold945/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6334_ _7045_/Q _6241_/Z _6268_/Z _6949_/Q _6274_/Z _7215_/Q _6335_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold923 _6848_/Q hold923/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6265_ _6302_/A3 _6533_/A4 _6285_/A2 _6302_/A4 _6265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold989 _7127_/Q hold989/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold967 _7214_/Q hold967/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold956 _5760_/Z _7103_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold978 _5685_/Z _7037_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_142_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3477_ hold272/Z hold4/Z hold54/Z _3477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5216_ _4697_/Z _5310_/A2 _5460_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6196_ _6712_/Q _6002_/Z _6003_/Z _6714_/Q _6198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5147_ _4842_/Z _5147_/A2 _5147_/A3 _5147_/A4 _5147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_111_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5078_ _5324_/A1 _5078_/A2 _5263_/A4 _5263_/A2 _5337_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_72_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4029_ _4029_/A1 _4029_/A2 _4391_/A3 _4391_/A4 _4031_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_38_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet563_203 net613_256/I _7022_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_214 net563_246/I _7011_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_247 net613_255/I _6978_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_236 net563_245/I _6989_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_225 net563_225/I _7000_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold208 _5646_/Z _7003_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4380_ _4853_/A1 _5270_/A1 _5170_/A2 _4380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3400_ _3400_/I _6601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold219 _7115_/Q hold219/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3331_ _7237_/Q _6302_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_98_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6050_ _7152_/Q _5960_/Z _5965_/Z _6700_/Q _5969_/Z _7120_/Q _6053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _5000_/Z _5001_/A2 _5001_/B _6859_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_100_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6952_ _6952_/D _7238_/RN _6952_/CLK _6952_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5903_ _5901_/B _5902_/Z _7223_/Q _5903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_81_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6883_ _6883_/D input75/Z _6883_/CLK _6883_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5834_ hold65/Z hold352/Z _5838_/S _5834_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ hold190/Z hold12/Z _5766_/S _5765_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4716_ _5420_/A2 _4835_/A2 _4456_/B _3401_/I _4716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5696_ hold65/Z hold341/Z hold25/Z _7047_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4647_ _5038_/A1 _5475_/A3 _5439_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold720 _4263_/Z _6777_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4578_ _5464_/A1 _5438_/C _5346_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _7135_/Q _6253_/Z _6296_/Z _7159_/Q _6322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold742 _4279_/Z _6790_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold764 _4340_/Z _6844_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold731 _6858_/Q hold731/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold753 _6786_/Q hold753/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_155 net813_461/I _7070_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_166 net413_95/I _7059_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold797 _7324_/I hold797/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3529_ hold6/Z _3552_/A2 _3484_/Z hold15/Z _3529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold786 _4205_/Z _6739_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold775 _6821_/Q hold775/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7297_ _7297_/D input75/Z _7297_/CLK _7297_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet513_177 net563_217/I _7048_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6248_ _7236_/Q _6484_/A2 _6452_/A4 _6302_/A4 _6248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet513_199 net763_420/I _7026_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_188 _4073__7/I _7037_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6179_ _7117_/Q _5984_/Z _5997_/Z _7101_/Q _7075_/Q _5980_/Z _6180_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_130_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold91 hold91/I hold91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold80 hold80/I hold80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_36_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3880_ _3880_/I _3881_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_409 net763_409/I _6765_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ hold291/Z hold811/Z _5556_/S _5550_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4501_ _4853_/A1 _4884_/A1 _4501_/B _4504_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5481_ _4944_/Z _5245_/Z _5481_/B1 _4951_/Z _5481_/C _5482_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_129_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4432_ _4460_/B _4376_/Z _4648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7220_ _7220_/D _7237_/RN _7220_/CLK _7220_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_145_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4363_ _4460_/B _4436_/B _4363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_116_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7151_ _7151_/D _7218_/RN _7151_/CLK _7151_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_112_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3314_ _6950_/Q _3994_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_59_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7082_ hold96/Z _7260_/RN _7082_/CLK hold95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6102_ _6952_/Q _5958_/Z _5999_/Z _7032_/Q _6102_/C _6106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4294_ _6565_/I0 _6802_/Q _4300_/S _6802_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6033_ _7061_/Q _5985_/Z _5997_/Z _7095_/Q _6037_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_100_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6935_ _6935_/D _7237_/RN _6935_/CLK _6935_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _6866_/D _7218_/RN _6866_/CLK _6866_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_22_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6797_ _6797_/D _7265_/CLK _6797_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5817_ hold48/Z hold435/Z _5820_/S _5817_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5748_ hold2/Z hold137/Z _5748_/S _5748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ hold497/Z hold48/Z hold33/Z _7032_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold561 _5735_/Z _7081_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold572 _7152_/Q hold572/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold550 _7120_/Q hold550/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold594 _6775_/Q hold594/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold583 _4218_/Z _6749_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _5262_/A2 _5255_/A2 _4495_/Z _4497_/Z _4981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_51_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3932_ _3932_/A1 _3533_/Z _3542_/Z _3932_/B _3933_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_6720_ _6720_/D _7170_/RN _6720_/CLK _6720_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_176_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _7235_/RN _4064_/S _6651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_108_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36__1359_ clkbuf_4_10_0__1359_/Z net663_322/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3863_ _6973_/Q _3923_/A2 _3959_/C1 _7183_/Q _3869_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_116__1359_ net513_165/I net813_467/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6582_ _6834_/Q _6582_/A2 _6582_/B1 _6835_/Q _6836_/Q _6582_/C2 _6583_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5602_ hold24/Z _3515_/Z hold42/Z hold6/Z hold43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_99__1359_ clkbuf_4_5_0__1359_/Z net613_279/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5533_ hold548/Z hold91/Z _5535_/S _5533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3794_ _3794_/A1 _3794_/A2 _3794_/A3 _3794_/A4 _3794_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5464_ _5464_/A1 _4659_/Z _4675_/Z _5464_/B _5465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_117_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4415_ _5385_/A1 _5045_/C _4415_/B _5211_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5395_ _5395_/A1 _4991_/C _5428_/A2 _5395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7203_ _7203_/D _7237_/RN _7203_/CLK _7203_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_154_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7134_ _7134_/D _7258_/RN _7134_/CLK _7134_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4346_ hold291/Z hold923/Z _4346_/S _4346_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7065_ hold61/Z _7260_/RN _7065_/CLK hold60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4277_ _3509_/Z _5520_/C _5513_/A3 _5857_/A2 _4279_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6016_ _7013_/Q _5971_/Z _6031_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_2007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _6918_/D _7258_/RN _6918_/CLK _6918_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _6849_/D _7170_/RN _6849_/CLK _6849_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_167_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold380 _6889_/Q hold380/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold391 _5576_/Z _6940_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_120_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_490 net813_491/I _6675_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_187_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ hold452/Z hold91/Z _4210_/S _4200_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5180_ _5180_/A1 _5180_/A2 _5180_/A3 _5211_/C _5185_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_111_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0__1359_ clkbuf_0__1359_/Z net513_167/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_3_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4131_ hold91/Z hold578/Z _4136_/S _4131_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _4061_/Z _3337_/I _7299_/Q _4062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _4421_/Z _4908_/Z _4966_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_184_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6703_ _6703_/D _7235_/RN _6703_/CLK _6703_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_20_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3915_ _3915_/A1 _3915_/A2 _3915_/A3 _3915_/A4 _3915_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4895_ _4886_/Z _4887_/Z _4891_/Z _4895_/A4 _4898_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6634_ _7235_/RN _6653_/A2 _6634_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3846_ _3540_/Z _3552_/Z _3939_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_158_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3777_ _7176_/Q _3945_/A2 _5532_/A1 _6903_/Q _3797_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6565_ _6565_/I0 _7263_/Q _6571_/S _7263_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _6947_/Q _6245_/Z _6288_/Z _7125_/Q _6498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5516_ hold227/Z hold250/Z _5516_/S _5516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5447_ _5447_/A1 _5447_/A2 _5448_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _5425_/A2 _5425_/A3 _5379_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7117_ _7117_/D _7237_/RN _7117_/CLK _7117_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4329_ _3509_/Z _5839_/A3 _5513_/A3 _5520_/C _4331_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_86_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7048_ _7048_/D _7258_/RN _7048_/CLK _7048_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_170_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4073__6 _4073__6/I _7219_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_82__1359_ net413_62/I _4073__15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_183_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3700_ _6686_/Q _3945_/C2 _5683_/A1 _7040_/Q _3701_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_175_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4680_ _4414_/Z _4452_/Z _4666_/Z _5395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_119_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _6938_/Q _3910_/A2 _3954_/A2 _6994_/Q _7204_/Q _3955_/A2 _3632_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6350_ _7128_/Q _6247_/Z _6297_/Z _6700_/Q _6351_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3562_ _3507_/Z _3537_/Z _3927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_128_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5301_ _5301_/I _6861_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6281_ _6484_/A3 _6256_/Z _6272_/Z _6274_/Z _6281_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3493_ _3493_/I0 hold319/Z hold54/Z _3493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5232_ _5414_/A2 _4752_/Z _5233_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5163_ _5356_/A1 _4650_/Z _5231_/A2 _5468_/A1 _5166_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_111_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4114_ hold20/Z hold260/Z _4118_/S _4114_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5094_ _5328_/A1 _5389_/A1 _5094_/B _5094_/C _5347_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_68_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4045_ _6832_/Q _4097_/A1 _4045_/B1 _6826_/Q _4046_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_37_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _7231_/Q _6210_/B _6014_/A2 _7229_/Q _5996_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_80_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _5072_/A4 _4903_/Z _4421_/Z _4500_/Z _4947_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_33_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _4997_/C _4878_/A2 _3401_/I _3402_/I _4878_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_138_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6617_ _7235_/RN _6657_/A2 _6617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3829_ _3537_/Z hold674/Z _4161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _6548_/A1 _6548_/A2 _6548_/A3 _6547_/Z _6548_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _7189_/Q _6282_/Z _6492_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_106_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput271 _6682_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput260 _6891_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput282 _6683_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput293 _6688_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5850_ hold291/Z hold963/Z _5856_/S _5850_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _5312_/A2 _5312_/A4 _5456_/A1 _5220_/B2 _4801_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_15_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ hold48/Z hold462/Z _5784_/S _5781_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4732_ _4765_/A1 _4510_/Z _5302_/B _5099_/A2 _4732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4663_ _4411_/Z _5214_/A2 _5172_/B _5165_/A4 _4663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6402_ _7130_/Q _6484_/A2 _6484_/A3 _6533_/A4 _6403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3614_ _3505_/Z _3533_/Z _3770_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4594_ _5190_/A2 _5435_/A2 _5389_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold913 _7190_/Q hold913/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold902 _4291_/Z _6800_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_155_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold935 _6905_/Q hold935/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold946 _5832_/Z _7167_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6333_ _7207_/Q _6256_/Z _6261_/Z _6957_/Q _6285_/Z _7191_/Q _6335_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3545_ _3485_/Z _3521_/Z _3959_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold924 _4346_/Z _6848_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3476_ _3476_/I _3478_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold968 _5885_/Z _7214_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold979 _7045_/Q hold979/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold957 _6709_/Q hold957/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _6956_/Q _6261_/Z _6263_/Z _6932_/Q _6262_/Z _6964_/Q _6271_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_170_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _4698_/B _5403_/A2 _5215_/B _5215_/C _5316_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6195_ _6824_/Q _5988_/Z _6019_/Z _6853_/Q _6198_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5146_ _4546_/Z _5364_/B _4586_/Z _4598_/Z _4568_/Z _5147_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_97_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ _4973_/Z _5078_/A2 _5258_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4028_ input97/Z input96/Z input99/Z input98/Z _4028_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_84_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ _6002_/A2 _6021_/A2 _6210_/A2 _7227_/Q _5979_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_139_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_204 net763_422/I _7021_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_154_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_215 net763_426/I _7010_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_226 net613_258/I _6999_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_237 net813_467/I _6988_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_248 net763_422/I _6977_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold209 _7027_/Q hold209/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3330_ _7236_/Q _6285_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_4_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _5000_/A1 _5000_/A2 _5000_/A3 _5000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_0_0__1359_ clkbuf_0__1359_/Z net763_436/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_121_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _6951_/D _7238_/RN _6951_/CLK _6951_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_5902_ _5911_/A1 _6746_/Q _7225_/Q _5902_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_53_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6882_ _6882_/D input75/Z _6882_/CLK _6882_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5833_ hold91/Z hold564/Z _5838_/S _5833_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5764_ hold649/Z hold20/Z _5766_/S _5764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4715_ _4835_/A2 _5087_/A1 _5328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5695_ hold91/Z hold508/Z hold25/Z _7046_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4646_ _4648_/A1 _4648_/A2 _4648_/B _5475_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4577_ _5002_/A3 _5002_/A4 _5083_/B _5003_/A2 _5043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold721 _7172_/Q hold721/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold710 _4189_/Z _6726_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _7167_/Q _5948_/Z _6245_/Z _6941_/Q _6263_/Z _6933_/Q _6329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold754 _4273_/Z _6786_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold743 _6764_/Q hold743/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold732 _4361_/Z _6858_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_157_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold787 _7313_/I hold787/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet513_167 net513_167/I _7058_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3528_ _3525_/Z _3527_/Z _3935_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet513_156 _4073__50/I _7069_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold776 _4322_/Z _6821_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold765 _6842_/Q hold765/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7296_ _7296_/D input75/Z _7296_/CLK _7296_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3459_ hold90/Z hold290/Z _3460_/S _7285_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6247_ _7236_/Q _6484_/A2 _6533_/A4 _6302_/A4 _6247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet513_178 net763_419/I _7047_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold798 _5541_/Z _6909_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_77_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_189 net513_189/I _7036_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _7157_/Q _5960_/Z _5965_/Z _6705_/Q _6006_/Z _7173_/Q _6180_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5129_ _5420_/A2 _5129_/A2 _5129_/A3 _3401_/I _5129_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_97_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold81 hold81/I hold81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold70 hold70/I hold70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold92 hold92/I hold92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_152_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4500_ _4759_/A2 _4759_/A3 _4500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_145_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5480_ _5480_/A1 _5480_/A2 _5480_/A3 _5479_/Z _5480_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4431_ _4414_/Z _4421_/Z _5393_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_6_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_1 _4121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4362_ _5299_/C _6859_/Q _5001_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7150_ _7150_/D input75/Z _7150_/CLK _7150_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3313_ _6830_/Q _4038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7081_ _7081_/D _7237_/RN _7081_/CLK _7081_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6101_ _6101_/A1 _6101_/A2 _6101_/A3 _6101_/A4 _6101_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4293_ _6564_/I0 _6801_/Q _4300_/S _6801_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_59__1359_ net513_170/I net763_434/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ _7069_/Q _5980_/Z _6003_/Z _7159_/Q _6037_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_139__1359_ clkbuf_4_1_0__1359_/Z _4073__3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6934_ _6934_/D _7258_/RN _6934_/CLK _6934_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6865_ _6865_/D _7279_/RN _7278_/CLK hold14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5816_ hold65/Z hold542/Z _5820_/S _5816_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6796_ _6796_/D _7265_/CLK _6796_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5747_ hold12/Z hold486/Z _5748_/S _5747_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5678_ hold331/Z hold65/Z hold33/Z _7031_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4629_ _5190_/A2 _4604_/Z _5387_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold562 _7105_/Q hold562/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold551 _5779_/Z _7120_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold540 _7311_/I hold540/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7279_ _7279_/D _7279_/RN _7279_/CLK hold31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold584 _7329_/I hold584/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold595 _4260_/Z _6775_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold573 _5815_/Z _7152_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput160 wb_rstn_i _7279_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_36_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4980_ _4998_/A2 _5262_/A2 _5255_/A2 _5442_/A2 _4980_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet413_100 net563_239/I _7125_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3931_ _7052_/Q _5701_/A1 _5536_/A1 _6906_/Q _3932_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_16_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6650_ _7235_/RN _6657_/A2 _6650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3862_ _6957_/Q _3957_/A2 _3928_/C1 _6823_/Q _3925_/B1 _6825_/Q _3869_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_31_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6581_ _6581_/I0 _7270_/Q _6602_/S _7270_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5601_ hold2/Z _6963_/Q hold7/Z hold8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5532_ _5532_/A1 hold32/Z _5535_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3793_ _7136_/Q _3951_/A2 _3924_/A2 _6966_/Q _3794_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_31_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ _5463_/A1 _5463_/A2 _5485_/A2 _5463_/B2 _5463_/C _5474_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_8_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4414_ _4397_/Z _4491_/B _5003_/A2 _4414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5394_ _4892_/B _5394_/A2 _5428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7202_ _7202_/D _7256_/RN _7202_/CLK _7202_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_7133_ _7133_/D _7237_/RN _7133_/CLK _7133_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4345_ _4103_/I hold887/Z _4346_/S _4345_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _7064_/D _7238_/RN _7064_/CLK _7064_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4276_ hold729/Z hold291/Z _4276_/S _4276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6015_ _7228_/Q _6211_/B1 _6015_/A3 _6210_/A2 _6015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_100_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6917_ _6917_/D _7258_/RN _6917_/CLK _6917_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6848_ _6848_/D input75/Z _6848_/CLK _6848_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6779_ hold98/Z _7238_/RN _6779_/CLK hold97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_164_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold370 _5688_/Z _7040_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold381 _5511_/Z _6889_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold392 _6888_/Q hold392/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_leaf_42__1359_ net413_93/I net413_77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_480 net813_481/I _6685_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_491 net813_491/I _6674_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4130_ hold291/Z hold965/Z _4136_/S _4130_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4061_ _4060_/Z input38/Z _7301_/Q _4061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4963_ _4963_/A1 _4960_/Z _4961_/Z _4962_/Z _4966_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_184_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6702_ _6702_/D _7238_/RN _6702_/CLK _6702_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3914_ _7102_/Q _5758_/A1 _3914_/B1 _6876_/Q _3915_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_189_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4894_ _4894_/A1 _4893_/Z _4895_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6633_ _7170_/RN _6652_/A2 _6633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ _7061_/Q _3927_/B1 _3955_/B1 _6848_/Q _3895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3776_ _3773_/Z _3776_/A2 _3776_/A3 _3776_/A4 _3776_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6564_ _6564_/I0 _7262_/Q _6571_/S _7262_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _7051_/Q _6241_/Z _6251_/Z _6987_/Q _6268_/Z _6955_/Q _6498_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5515_ _3485_/Z _5857_/A3 _5839_/A3 _5520_/C _5516_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_172_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _5446_/A1 _5446_/A2 _5447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_146_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _5377_/A1 _5290_/Z _5377_/A3 _5377_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_114_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7116_ _7116_/D _7237_/RN _7116_/CLK _7116_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4328_ hold291/Z hold739/Z _4328_/S _4328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7047_ _7047_/D _7258_/RN _7047_/CLK _7047_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4259_ hold20/Z hold296/Z _4261_/S _4259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__7 _4073__7/I _7218_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3630_ _3630_/A1 _3630_/A2 _3630_/A3 _3630_/A4 _3630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3561_ _3533_/Z _3560_/Z _3913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _5242_/Z _5266_/Z _5300_/A3 _5299_/C _6861_/Q _5301_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_115_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6280_ _6245_/Z _6262_/Z _6263_/Z _6279_/Z _6287_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3492_ _3491_/I _3307_/I hold54/Z _3492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_103_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5231_ _5291_/B _5231_/A2 _5231_/B _5231_/C _5314_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_45_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _5165_/A2 _5287_/B _5315_/A2 _5315_/A1 _5467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4113_ hold19/Z _7275_/Q hold54/I hold20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5093_ _5359_/A1 _4568_/Z _5218_/B _5303_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _4044_/I _6732_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _7052_/Q _5924_/Z _5994_/I _7134_/Q _5995_/C _6009_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_24_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _4500_/Z _4903_/Z _5072_/A4 _4666_/Z _4946_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_149_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4877_ _4651_/Z _4483_/B _4422_/Z _4683_/Z _4877_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_71_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6616_ _7235_/RN _6657_/A2 _6616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3828_ _3535_/Z _3537_/Z _3956_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6547_ _6547_/A1 _6547_/A2 _6542_/Z _6546_/Z _6547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_152_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3759_ _3759_/A1 _3759_/A2 _3747_/Z _3758_/Z _3759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_165_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6478_ _7043_/Q _6275_/Z _6486_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5429_ _4898_/C _4991_/C _5392_/B _4893_/Z _5429_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput250 _4092_/ZN pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput261 _6877_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput272 _6676_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput294 _6689_/Q pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput283 _6670_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew349 hold24/Z _5520_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_78_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4800_ _4675_/Z _4683_/Z _5130_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ hold65/Z hold911/Z _5784_/S _5780_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4731_ _4765_/A1 _5302_/B _5099_/A2 _4716_/Z _4731_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _5464_/A1 _4414_/Z _4659_/Z _4662_/B _4664_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_147_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3613_ _7074_/Q _3943_/A2 _3647_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_70_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6401_ _6401_/A1 _6401_/A2 _6401_/A3 _6401_/A4 _6401_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _4593_/A1 _5018_/B _4601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold903 _6719_/Q hold903/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_31_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3544_ input51/Z _4210_/S _4244_/S input42/Z _3589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_127_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold936 _5535_/Z _6905_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold914 _5858_/Z _7190_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6332_ _6981_/Q _6251_/Z _6254_/Z _7175_/Q _6332_/C _6335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold925 _6695_/Q hold925/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3475_ _6660_/Q hold271/Z _6733_/Q _3476_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6263_ _7232_/Q _6533_/A2 _6452_/A4 _6282_/A2 _6263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_131_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold969 _7176_/Q hold969/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold947 _7159_/Q hold947/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold958 _4163_/Z _6709_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5214_ _5343_/A2 _5214_/A2 _5310_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6194_ _6820_/Q _5979_/Z _5996_/Z _6708_/Q _6198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5145_ _4570_/Z _5145_/A2 _4878_/Z _5287_/B _4820_/Z _4821_/Z _5147_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_111_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5076_ _5464_/A1 _4905_/Z _4973_/Z _4700_/Z _5076_/C _5079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_84_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4027_ _4027_/A1 _4027_/A2 _4031_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ _5924_/Z _5975_/Z _5976_/Z _5977_/Z _5983_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_25_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _4929_/A1 _4928_/Z _4929_/A3 _4933_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_60_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_238 net613_254/I _6987_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_227 net763_423/I _6998_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_205 net613_256/I _7020_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_216 net563_225/I _7009_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_249 net813_463/I _6976_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6950_ _6950_/D _7238_/RN _6950_/CLK _6950_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5901_ _5901_/A1 _5951_/A3 _5901_/B _5904_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_93_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6881_ _6881_/D input75/Z _6881_/CLK _6881_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5832_ hold291/Z hold945/Z _5838_/S _5832_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5763_ hold433/Z hold48/Z _5766_/S _5763_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4714_ _4709_/Z _4711_/Z _5305_/B _4714_/A4 _4727_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_19__1359_ _4073__7/I _4073__47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5694_ hold291/Z hold979/Z hold25/Z _7045_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4645_ _4565_/Z _4641_/Z _5040_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4576_ _4549_/Z _4570_/Z _5192_/B _4576_/C _4584_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_162_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold711 _6843_/Q hold711/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold700 _4360_/Z _6857_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold722 _5837_/Z _7172_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3527_ _3552_/A2 _3484_/Z hold15/Z _3477_/Z _3527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6315_ _7183_/Q _6282_/Z _6322_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold744 _4248_/Z _6764_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold755 _6717_/Q hold755/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold733 _6727_/Q hold733/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7295_ _7295_/D _6649_/Z _7304_/CLK _7295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold777 _6761_/Q hold777/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold788 _4237_/Z _6758_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_157 _4073__51/I _7068_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_168 net663_330/I _7057_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold766 _4337_/Z _6842_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3458_ hold64/Z hold90/Z _3460_/S _7286_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet513_179 net763_420/I _7046_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold799 _6891_/Q hold799/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6246_ _7004_/Q _6243_/Z _6245_/Z _6940_/Q _6260_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3389_ _7229_/Q _5984_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_97_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _7109_/Q _5967_/Z _6177_/B _6180_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5128_ _5453_/A4 _5319_/A3 _5181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _4700_/Z _5325_/B _5060_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold60 hold60/I hold60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold82 hold82/I hold82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold71 hold71/I hold71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_75_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold93 hold93/I hold93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_91_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4430_ _4402_/B _4026_/B _4026_/C _5083_/C _4997_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_144_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_2 _4124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4361_ hold731/Z hold291/Z _4361_/S _4361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6100_ _7016_/Q _5971_/Z _5988_/Z _6984_/Q _6005_/Z _7040_/Q _6101_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3312_ _3312_/I _3428_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ _6828_/Q _7279_/RN _4300_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7080_ _7080_/D _7260_/RN _7080_/CLK _7080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_98_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ _6031_/A1 _6026_/Z _6030_/Z _6031_/A4 _6031_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_100_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_6__1359_ net763_436/I net813_469/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6933_ _6933_/D _7238_/RN _6933_/CLK _6933_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _6864_/D _7279_/RN _7278_/CLK hold4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5815_ hold91/Z hold572/Z _5820_/S _5815_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6795_ _6795_/D _7269_/CLK _6795_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5746_ hold20/Z hold373/Z _5748_/S _5746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5677_ hold513/Z hold91/Z hold33/Z _7030_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4628_ _4565_/Z _4624_/Z _5035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_163_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold530 _5687_/Z _7039_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4559_ _5464_/A1 _4997_/C _5393_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold563 _5762_/Z _7105_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold552 _6887_/Q hold552/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold541 _4224_/Z _6752_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7278_ _7278_/D _7279_/RN _7278_/CLK _7278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold585 _5546_/Z _6914_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold596 _7096_/Q hold596/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold574 _6820_/Q hold574/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6229_ _6220_/Z _6228_/Z _6555_/B1 _6168_/C _6555_/C _6230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_103_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_65__1359_ net513_175/I net613_297/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_145__1359_ net763_436/I net713_369/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput161 wb_sel_i[0] _6572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput150 wb_dat_i[2] _3395_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_163_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_101 net413_81/I _7124_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ _7126_/Q _3930_/A2 _3930_/B1 _6841_/Q _4170_/A1 _6714_/Q _3938_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_177_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3861_ _7207_/Q _3960_/A2 _3955_/A2 _7199_/Q _3924_/A2 _6965_/Q _3869_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6580_ _6580_/A1 _4313_/Z _6580_/B _6581_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_108_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ hold12/Z hold295/Z hold7/Z _6962_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3792_ _6990_/Q _3954_/A2 _3954_/B1 input22/Z _3794_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_31_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5531_ _4103_/I hold825/Z _5531_/S _5531_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7201_ _7201_/D _7237_/RN _7201_/CLK _7201_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5462_ _5404_/Z _5457_/Z _5461_/I _5463_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5393_ _5393_/A1 _5393_/A2 _5393_/B1 _5045_/C _5433_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4413_ _5209_/A3 _4397_/Z _5045_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7132_ _7132_/D _7237_/RN _7132_/CLK _7132_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _3529_/Z _3535_/Z _5520_/C _4346_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_28_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ _7063_/D _7235_/RN _7063_/CLK _7063_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_140_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _6210_/B _6014_/A2 _6210_/A2 _7229_/Q _6014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_87_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4275_ hold695/Z _4103_/I _4276_/S _4275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6916_ _6916_/D _7258_/RN _6916_/CLK _6916_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6847_ _6847_/D input75/Z _6847_/CLK _6847_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_161_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _6778_/D _7258_/RN _6778_/CLK _6778_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5729_ hold875/Z _4103_/I _5730_/S _5729_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold360 _6948_/Q hold360/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold371 _7009_/Q hold371/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold382 _7197_/Q hold382/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold393 _5509_/Z _6888_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_481 net813_481/I _6684_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_492 net813_492/I _6673_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_470 net813_470/I _6695_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4060_ _6748_/Q _6875_/Q _4064_/S _4060_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4962_ _4500_/Z _4906_/Z _5072_/A4 _4666_/Z _4962_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_64_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6701_ _6701_/D _7235_/RN _6701_/CLK _6701_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4893_ _5139_/A2 _5139_/A3 _4542_/Z _5172_/C _4893_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3913_ input11/Z _3913_/A2 _3913_/B1 _6892_/Q _3915_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3844_ _3529_/Z _3535_/Z _3955_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6632_ _7170_/RN _6652_/A2 _6632_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6563_ _6833_/D _7279_/RN _6571_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3775_ _7112_/Q _3917_/A2 _3913_/A2 input13/Z _3916_/A2 _7152_/Q _3776_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_118_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6494_ _7027_/Q _6235_/Z _6243_/Z _7011_/Q _6265_/Z _7003_/Q _6499_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5514_ _4103_/I hold799/Z _5514_/S _5514_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5445_ _4376_/Z _5255_/B _4972_/Z _5445_/B2 _5056_/B _5445_/C2 _5446_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_145_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5376_ _5291_/C _5376_/A2 _5468_/B1 _5376_/B2 _5376_/C _5377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7115_ _7115_/D _7237_/RN _7115_/CLK _7115_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4327_ _4103_/I hold689/Z _4328_/S _4327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4258_ hold48/Z hold618/Z _4261_/S _4258_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _7046_/D _7260_/RN _7046_/CLK _7046_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4189_ hold709/Z _4103_/I _4190_/S _4189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__8 _4073__8/I _7217_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold190 _7108_/Q hold190/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3560_ hold320/Z _3497_/I hold673/Z _3489_/I _3560_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_183_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3491_ _3491_/I _3493_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5230_ _4510_/Z _5414_/A2 _5230_/B _5231_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_170_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5161_ _5161_/A1 _5161_/A2 _5366_/A1 _5166_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_123_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _5092_/A1 _4705_/Z _5218_/B _4784_/Z _5303_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_84_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4112_ hold48/Z hold269/Z _4118_/S _4112_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4043_ _4043_/A1 _6732_/Q _6733_/Q _3409_/Z _4044_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_56_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5994_ _5994_/I _6051_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4945_ _4500_/Z _4903_/Z _5072_/A4 _5359_/A1 _4945_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _4650_/Z _4876_/A2 _4876_/B _4876_/C _4880_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6615_ _7235_/RN _6653_/A2 _6615_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3827_ _3537_/Z _3540_/Z _3946_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3758_ _3758_/A1 _3751_/Z _3757_/Z _3758_/A4 _3758_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6546_ _6546_/A1 _6546_/A2 _6546_/A3 _6546_/A4 _6546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6477_ _6971_/Q _6262_/Z _6499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3689_ _3689_/A1 _3657_/Z _3688_/Z _6569_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_161_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5428_ _5381_/I _5428_/A2 _6577_/C _5428_/A4 _5428_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xoutput251 _4080_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput240 _7309_/Z mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput262 _6878_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5359_ _5359_/A1 _4892_/B _5360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_87_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput273 _6677_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput295 _6674_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput284 _6671_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _7029_/D _7008_/RN _7029_/CLK _7029_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_101_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4730_ _4716_/Z _4728_/Z _5105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _4414_/Z _5038_/A1 _5359_/A1 _4557_/Z _4662_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6400_ _7210_/Q _6256_/Z _6263_/Z _6936_/Q _6401_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3612_ _6680_/Q _3546_/Z _3625_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_162_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4592_ _4565_/Z _4586_/Z _5018_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_156_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6331_ _6331_/I _6332_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold904 _4178_/Z _6719_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold937 _7215_/Q hold937/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3543_ _3485_/Z _3542_/Z _4244_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_7_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold926 _4145_/Z _6695_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold915 _6713_/Q hold915/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3474_ _4041_/B1 _6660_/Q _3981_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_142_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6262_ _6302_/A3 _5943_/S _7234_/Q _6533_/A2 _6262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold948 _5823_/Z _7159_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold959 _7061_/Q hold959/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5213_ _4673_/Z _5124_/B _5213_/B _5213_/C _5454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_9_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6193_ _6193_/A1 _6193_/A2 _6193_/A3 _6193_/A4 _6193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5144_ _4555_/C _5276_/C _5145_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5075_ _5255_/B _5051_/Z _5075_/B _5076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_85_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4026_ _4402_/B _4483_/B _4026_/B _4026_/C _4412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_37_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _6996_/Q _6211_/B1 _6021_/A2 _7227_/Q _5977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4928_ _4376_/Z _5056_/C _5442_/A2 _5442_/A4 _4928_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_100_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ _4614_/Z _5051_/S _5287_/B _4681_/Z _4859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet563_206 net563_222/I _7019_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_228 net613_256/I _6997_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_217 net563_217/I _7008_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_239 net563_239/I _6986_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _6529_/I0 _7258_/Q _6555_/C _6529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5900_ _5900_/A1 _5954_/A3 _5951_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_75_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6880_ _6880_/D _7170_/RN _6880_/CLK _6880_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_34_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5831_ _4103_/I hold921/Z _5838_/S _5831_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5762_ hold562/Z hold65/Z _5766_/S _5762_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4713_ _4713_/A1 _5094_/B _4691_/Z _4699_/Z _5305_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ hold227/Z hold611/Z hold25/Z _7044_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4644_ _4644_/A1 _5038_/B _4643_/Z _4653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4575_ _5281_/C _4539_/I _4551_/Z _5364_/B _5192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_129_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold701 _6763_/Q hold701/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold712 _4339_/Z _6843_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7294_ _7294_/D _6648_/Z _7305_/CLK _7294_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold723 _7055_/Q hold723/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3526_ _3552_/A2 _3484_/Z hold15/Z hold16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6314_ _7053_/Q _6299_/Z _6328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold745 _6725_/Q hold745/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold734 _4190_/Z _6727_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_157_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_158 net513_163/I _7067_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold778 _4243_/Z _6761_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6245_ _7233_/Q _6533_/A2 _6452_/A4 _6279_/A3 _6245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold767 _7126_/Q hold767/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold756 _4175_/Z _6717_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3457_ hold47/Z hold64/Z _3460_/S _7287_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold789 _7320_/I hold789/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_169 _4073__39/I _7056_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3388_ _7230_/Q _6014_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_6176_ _5991_/Z _6176_/A2 _6176_/B _6176_/C _6177_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_5127_ _5127_/A1 _5457_/A1 _5213_/B _5127_/A4 _5127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_85_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ _5058_/A1 _5055_/Z _5193_/A2 _5058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XTAP_2928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4009_ _4009_/A1 _6744_/Q _6745_/Q _4010_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 hold50/I hold50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_152_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold83 hold83/I hold83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold61 hold61/I hold61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold72 hold72/I hold72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_leaf_105__1359_ clkbuf_4_5_0__1359_/Z net613_288/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_88__1359_ net513_175/I net613_258/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold94 hold94/I hold94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_16_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_3 _4133_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ hold699/Z _4103_/I _4361_/S _4360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3311_ _6730_/Q _3442_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_141_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ hold901/Z hold291/Z _4291_/S _4291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6030_ _6030_/A1 _6030_/A2 _6030_/A3 _6030_/A4 _6030_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_3_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6932_ _6932_/D _7008_/RN _6932_/CLK _6932_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_35_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _6863_/D _7279_/RN _7278_/CLK hold40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5814_ hold291/Z hold949/Z _5820_/S _5814_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6794_ _6794_/D _7265_/CLK _6794_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5745_ hold48/Z hold416/Z _5748_/S _5745_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5676_ hold972/Z hold291/Z hold33/Z _7029_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4627_ _4627_/A1 _4625_/Z _4626_/Z _4633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_135_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold520 _5754_/Z _7098_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4558_ _5038_/A1 _4557_/Z _5393_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold542 _7153_/Q hold542/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold553 _5508_/Z _6887_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold531 _6687_/Q hold531/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7277_ _7277_/D _7279_/RN _7279_/CLK _7277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold586 _6901_/Q hold586/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4489_ _4489_/A1 _4692_/B _4489_/B _4491_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3509_ hold6/Z hold41/Z _3484_/Z hold15/Z _3509_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold597 _5752_/Z _7096_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold564 _7168_/Q hold564/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold575 _4321_/Z _6820_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6228_ _6228_/A1 _6228_/A2 _6228_/A3 _6227_/Z _6228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_44_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6159_ _6147_/Z _6158_/Z _6473_/B1 _6168_/C _6555_/C _6160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_100_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput162 wb_sel_i[1] _6574_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput151 wb_dat_i[30] _6597_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput140 wb_dat_i[20] _6591_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _3860_/A1 _3860_/A2 _3860_/A3 _3860_/A4 _3860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3791_ _6950_/Q _5584_/A1 _5575_/A1 _6942_/Q _3925_/A2 input5/Z _3794_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5530_ _3485_/Z _5839_/A3 hold235/Z _5520_/C _5531_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_157_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5461_ _5461_/I _5480_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_172_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4412_ _4412_/A1 _4399_/Z _4412_/B _4412_/C _5209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_7200_ _7200_/D _7256_/RN _7200_/CLK _7200_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_68_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5392_ _5051_/S _5360_/B _5392_/B _5433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7131_ _7131_/D _7237_/RN _7131_/CLK _7131_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ hold291/Z hold737/Z _4343_/S _6846_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7062_ _7062_/D _7235_/RN _7062_/CLK _7062_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_141_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _4274_/A1 hold32/Z _4276_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_101_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _6013_/A1 _5991_/Z _6027_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6915_ _6915_/D _7218_/RN _6915_/CLK _7330_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_71__1359_ net513_175/I net613_254/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _6846_/D _7170_/RN _6846_/CLK _6846_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_51_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6777_ _6777_/D _7170_/RN _6777_/CLK _6777_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3989_ _7239_/Q _6895_/Q _6900_/Q _3990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_22_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5728_ _5728_/A1 hold32/Z _5730_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_176_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5659_ hold518/Z hold91/Z hold56/Z _7014_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ _7329_/I _7329_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold350 _6983_/Q hold350/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold361 _5585_/Z _6948_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold383 _5865_/Z _7197_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold394 _6956_/Q hold394/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold372 _5653_/Z _7009_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_460 net813_461/I _6705_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_493 net413_88/I _6672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_482 net813_487/I _6683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_471 net413_75/I _6694_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _4500_/Z _4906_/Z _5072_/A4 _5359_/A1 _4961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_92_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4892_ _4551_/Z _4716_/Z _4892_/B _4894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6700_ _6700_/D _7256_/RN _6700_/CLK _6700_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3912_ _7214_/Q _3912_/A2 _3912_/B1 _6883_/Q _3912_/C1 _6706_/Q _3915_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_33_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3843_ _3529_/Z _3617_/Z _3950_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6631_ _7170_/RN _6652_/A2 _6631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_32_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6562_ _6562_/I _7261_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3774_ _6926_/Q _3935_/A2 _3945_/C2 _6684_/Q _5701_/A1 _7054_/Q _3776_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _6493_/A1 _6493_/A2 _6486_/Z _6492_/Z _6493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5513_ _5520_/C _3533_/Z _5513_/A3 _5821_/A3 _5514_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_172_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ _5444_/A1 _5444_/A2 _5442_/Z _5444_/A4 _5483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_172_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5375_ _5421_/A2 _5470_/A1 _5372_/Z _5374_/Z _5379_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_102_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7114_ _7114_/D _7237_/RN _7114_/CLK _7114_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4326_ _3509_/Z _5821_/A3 hold235/Z _5520_/C _4328_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4257_ hold65/Z hold478/Z _4261_/S _4257_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7045_ _7045_/D _7218_/RN _7045_/CLK _7045_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4188_ _4188_/A1 hold32/Z _4190_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_28_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6829_ _6829_/D _7279_/RN _7279_/CLK _6829_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4073__9 _4073__9/I _7216_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold180 _6704_/Q hold180/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_151_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold191 _5765_/Z _7108_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3490_ _7305_/Q _7304_/Q _6733_/Q _3491_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5160_ _5287_/B _5293_/B _4784_/Z _5160_/B _5366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4111_ hold47/Z _7274_/Q hold54/I hold48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5091_ _4586_/Z _5302_/B _4784_/Z _4716_/Z _5222_/A1 _5103_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_4042_ _7291_/Q _3409_/Z _4042_/A3 _4043_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_97_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5993_ _7231_/Q _7228_/Q _7227_/Q _6211_/B1 _5994_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_25_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4944_ _4467_/B _4495_/Z _5324_/A1 _4759_/Z _4944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4875_ _4651_/Z _4817_/Z _4876_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6614_ _7235_/RN _6657_/A2 _6614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3826_ _3529_/Z _3560_/Z _3934_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3757_ _3757_/A1 _3757_/A2 _3757_/A3 _3757_/A4 _3757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6545_ _6788_/Q _6263_/Z _6266_/Z _6844_/Q _6546_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6476_ _7257_/Q _6476_/I1 _6558_/S _7257_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3688_ _3688_/A1 _3663_/Z _3674_/Z _3687_/Z _3688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput230 _7328_/Z mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5427_ _5427_/A1 _5425_/Z _5426_/Z _4881_/Z _5430_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_133_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput252 _4079_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput241 _7310_/Z mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5358_ _5432_/A1 _5189_/Z _5355_/Z _5357_/Z _5362_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput263 _6879_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput274 _6678_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput285 _6672_/Q pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4309_ _4309_/I0 _6815_/Q _4312_/S _6815_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput296 _6675_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5289_ _5029_/B _5289_/A2 _5289_/A3 _5292_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_75_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7028_ _7028_/D _7008_/RN _7028_/CLK _7028_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_47_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4660_ _4376_/Z _4411_/Z _5172_/B _5165_/A4 _5385_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_30_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ _3610_/Z _3611_/I1 _3899_/S _6875_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4591_ _4591_/A1 _4587_/Z _4590_/Z _4593_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_156_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6330_ _7005_/Q _6243_/Z _6269_/Z _7029_/Q _7119_/Q _6288_/Z _6331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_183_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3542_ _3653_/A1 hold320/Z _3497_/I _3501_/Z _3542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold927 _7036_/Q hold927/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_50_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold905 _6852_/Q hold905/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold916 _4169_/Z _6713_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3473_ _3471_/I _5490_/A1 hold54/Z _3473_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6261_ _7234_/Q _6533_/A2 _6533_/A3 _5943_/S _6261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold938 _5886_/Z _7215_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold949 _7151_/Q hold949/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5212_ _5242_/A3 _4810_/B _4812_/B _5212_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6192_ _6718_/Q _5960_/Z _6192_/B _6193_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5143_ _4820_/Z _4821_/Z _4878_/Z _5287_/B _5372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_9_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _5074_/A1 _5408_/C _5072_/Z _5335_/C _5075_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_69_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4025_ _4489_/B _4424_/B _4034_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _6015_/A3 _6211_/B1 _7004_/Q _7228_/Q _5976_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_13_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _4927_/A1 _4927_/A2 _4927_/A3 _4929_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4858_ _4858_/A1 _4858_/A2 _5289_/A2 _4862_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_166_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet563_218 net563_246/I _7007_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_207 net563_222/I _7018_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3809_ _3509_/Z _3617_/Z _4289_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet563_229 net763_422/I _6996_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4789_ _5270_/A1 _4808_/A2 _4530_/I _5302_/B _4789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_146_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ _6516_/Z _6527_/Z _6528_/B1 _6286_/Z _6529_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6459_ _6459_/I _6460_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48__1359_ net413_93/I _4073__5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_128__1359_ net613_261/I net713_379/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5830_ _3542_/Z _3552_/Z _5520_/C _5838_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_61_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5761_ hold546/Z hold91/Z _5766_/S _5761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _4687_/Z _5092_/A1 _4713_/A1 _4691_/Z _5222_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_148_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5692_ _3529_/Z _3542_/Z hold24/Z hold25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_4643_ _5315_/A1 _5315_/A2 _4546_/Z _5364_/B _4643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4574_ _5278_/C _4551_/Z _5370_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold702 _4247_/Z _6763_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7293_ _7293_/D _6647_/Z _7305_/CLK _7293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold724 _5705_/Z _7055_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_128_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3525_ _3653_/A1 hold320/Z _3617_/A1 _3501_/Z _3525_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6313_ _6997_/Q _6265_/Z _6266_/Z _7013_/Q _6329_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold713 _6841_/Q hold713/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold735 _6854_/Q hold735/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold746 _4187_/Z _6725_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet513_159 net813_464/I _7066_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6244_ _7235_/Q _7234_/Q _6452_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold779 _6755_/Q hold779/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_115_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold768 _5786_/Z _7126_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold757 _6721_/Q hold757/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3456_ hold19/Z hold47/Z _3460_/S _7288_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3387_ _7227_/Q _6015_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_85_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6175_ _6955_/Q _5958_/Z _5994_/I hold9/I _6176_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5126_ _5126_/I _5127_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ _5078_/A2 _5443_/A1 _5057_/B _5324_/C _5058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_2918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4008_ _4008_/I _4009_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5959_ _6014_/A2 _5984_/A1 _6068_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_40_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold40 hold40/I hold40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_96_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold73 hold73/I hold73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold62 hold62/I hold62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold51 hold51/I hold51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_63_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold95 hold95/I hold95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold84 hold84/I hold84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_90_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_4 _4181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3310_ hold14/Z _5490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_125_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4290_ hold889/Z _4103_/I _4291_/S _4290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_15_0__1359_ clkbuf_0__1359_/Z net513_170/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_120_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6931_ _6931_/D _7256_/RN _6931_/CLK _6931_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_54_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _6862_/D _7279_/RN _7278_/CLK _6862_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5813_ _4103_/I hold939/Z _5820_/S _5813_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6793_ _6793_/D _7265_/CLK _6793_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5744_ hold65/Z hold554/Z _5748_/S _5744_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ hold626/Z hold227/Z hold33/Z _7028_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4626_ _4887_/A1 _4868_/A1 _4546_/Z _5364_/B _4626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_129_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold510 _5623_/Z _6982_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4557_ _4436_/B _4648_/A1 _4648_/A2 _4557_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xhold521 _7129_/Q hold521/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31__1359_ clkbuf_opt_2_0__1359_/Z net763_409/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold543 _5816_/Z _7153_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold554 _7089_/Q hold554/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_leaf_111__1359_ net513_165/I net813_492/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold532 _4134_/Z _6687_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_leaf_94__1359_ net413_62/I net563_225/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7276_ _7276_/D _7279_/RN _7279_/CLK _7276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4488_ _4392_/Z _4474_/Z _4722_/A2 _4923_/A2 _4491_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold587 _5528_/Z hold587/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3508_ hold15/Z hold41/Z _3484_/Z hold42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xhold576 _7054_/Q hold576/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold565 _5833_/Z _7168_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3439_ _3971_/A1 _3442_/B _6665_/Q _6664_/Q _3440_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold598 _7200_/Q hold598/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6227_ _6227_/A1 _6227_/A2 _6227_/A3 _6227_/A4 _6227_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _6152_/Z _6155_/Z _6158_/A3 _6158_/A4 _6158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _5108_/Z _4853_/Z _4740_/Z _5111_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_85_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6089_ _7244_/Q _6089_/I1 _6558_/S _7244_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput163 wb_sel_i[2] _6573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput152 wb_dat_i[31] _6600_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput141 wb_dat_i[21] _6594_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput130 wb_dat_i[11] _6588_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ _3790_/A1 _3790_/A2 _3790_/A3 _3790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_20_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5460_ _5460_/A1 _5303_/Z _5460_/A3 _5460_/A4 _5461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4411_ _5083_/B _4412_/B _4412_/C _4411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_145_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5391_ _5388_/Z _4985_/Z _5386_/Z _5390_/Z _5391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_160_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7130_ _7130_/D _7237_/RN _7130_/CLK _7130_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_125_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _4103_/I _6845_/Q _4343_/S _4342_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7061_ _7061_/D _7008_/RN _7061_/CLK _7061_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4273_ hold291/Z hold753/Z _4273_/S _4273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _7021_/Q _6068_/A4 _6211_/B1 _6989_/Q _6013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
.ends

