magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 0 108 756
<< properties >>
string FIXED_BBOX 0 -216 216 756
<< end >>
