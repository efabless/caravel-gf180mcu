magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 72 720 252 756
rect 36 684 288 720
rect 0 612 324 684
rect 0 324 108 612
rect 216 324 324 612
rect 0 216 324 324
rect 0 0 108 216
rect 216 0 324 216
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
