magic
tech gf180mcuC
magscale 6 5
timestamp 1654634570
<< metal5 >>
rect 0 720 252 756
rect 0 684 288 720
rect 0 612 324 684
rect 0 432 108 612
rect 216 432 324 612
rect 0 324 324 432
rect 0 144 108 324
rect 216 144 324 324
rect 0 72 324 144
rect 0 36 288 72
rect 0 0 252 36
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
