magic
tech gf180mcuC
magscale 1 10
timestamp 1654613370
<< metal1 >>
rect 967 720 1039 739
rect 2311 720 2383 739
rect 3431 720 3503 739
rect 4775 720 4847 739
rect 5895 720 5967 739
rect 7239 720 7311 739
rect 8359 720 8431 739
rect 9703 720 9775 739
rect 10823 720 10895 739
rect 12167 720 12239 739
rect 967 648 1172 720
rect 2311 648 2516 720
rect 3431 648 3636 720
rect 4775 648 4980 720
rect 5895 648 6100 720
rect 7239 648 7444 720
rect 8359 648 8564 720
rect 9703 648 9908 720
rect 10823 648 11028 720
rect 12167 648 12372 720
rect 1097 587 1172 648
rect 1097 527 1104 587
rect 1164 527 1172 587
rect 1097 394 1172 527
rect 1415 384 1490 608
rect 2441 587 2516 648
rect 2441 527 2448 587
rect 2508 527 2516 587
rect 2441 394 2516 527
rect 2759 384 2834 608
rect 3561 587 3636 648
rect 3561 527 3568 587
rect 3628 527 3636 587
rect 3561 394 3636 527
rect 3879 384 3954 608
rect 4905 394 4980 648
rect 5223 587 5298 608
rect 5223 527 5230 587
rect 5290 527 5298 587
rect 5223 384 5298 527
rect 6025 394 6100 648
rect 6343 587 6418 608
rect 6343 527 6350 587
rect 6410 527 6418 587
rect 6343 384 6418 527
rect 7369 394 7444 648
rect 7687 587 7762 608
rect 7687 527 7694 587
rect 7754 527 7762 587
rect 7687 384 7762 527
rect 8489 394 8564 648
rect 8807 587 8882 608
rect 8807 527 8814 587
rect 8874 527 8882 587
rect 8807 384 8882 527
rect 9833 394 9908 648
rect 10151 587 10226 608
rect 10151 527 10158 587
rect 10218 527 10226 587
rect 10151 384 10226 527
rect 10953 394 11028 648
rect 11271 587 11346 608
rect 11271 527 11278 587
rect 11338 527 11346 587
rect 11271 384 11346 527
rect 12297 394 12372 648
rect 12615 587 12690 608
rect 12615 527 12622 587
rect 12682 527 12690 587
rect 12615 384 12690 527
<< via1 >>
rect 532 1028 1201 1088
rect 6432 1028 7101 1088
rect 12332 1028 13001 1088
rect 1104 527 1164 587
rect 2448 527 2508 587
rect 3568 527 3628 587
rect 5230 527 5290 587
rect 6350 527 6410 587
rect 7694 527 7754 587
rect 8814 527 8874 587
rect 10158 527 10218 587
rect 11278 527 11338 587
rect 12622 527 12682 587
rect 541 249 1210 309
rect 6441 249 7110 309
rect 12341 249 13010 309
<< metal2 >>
rect 519 1088 1215 1099
rect 519 1028 532 1088
rect 1201 1028 1215 1088
rect 519 1016 1215 1028
rect 6420 1088 7115 1099
rect 6420 1028 6432 1088
rect 7101 1028 7115 1088
rect 6420 1016 7115 1028
rect 12320 1088 13015 1099
rect 12320 1028 12332 1088
rect 13001 1028 13015 1088
rect 12320 1016 13015 1028
rect 0 587 1503 589
rect 0 527 1104 587
rect 1164 527 1503 587
rect 0 525 1503 527
rect 1648 587 2847 589
rect 1648 527 2448 587
rect 2508 527 2847 587
rect 1648 525 2847 527
rect 3018 587 3967 589
rect 3018 527 3568 587
rect 3628 527 3967 587
rect 4475 587 5311 589
rect 4475 564 5230 587
rect 3018 525 3967 527
rect 4474 527 5230 564
rect 5290 527 5311 587
rect 4474 525 5311 527
rect 6012 587 6431 589
rect 6012 527 6350 587
rect 6410 527 6431 587
rect 6012 525 6431 527
rect 7356 587 7775 589
rect 7356 527 7694 587
rect 7754 527 7775 587
rect 7356 525 7775 527
rect 8476 587 9114 589
rect 8476 527 8814 587
rect 8874 527 9114 587
rect 8476 525 9114 527
rect 9820 587 10570 589
rect 9820 527 10158 587
rect 10218 527 10570 587
rect 9820 525 10570 527
rect 10940 587 12134 589
rect 10940 527 11278 587
rect 11338 527 12134 587
rect 10940 525 12134 527
rect 12284 587 13590 589
rect 12284 527 12622 587
rect 12682 527 13590 587
rect 12284 525 13590 527
rect 0 5 56 525
rect 1648 322 1712 525
rect 529 309 1222 321
rect 529 249 541 309
rect 1210 249 1222 309
rect 529 238 1222 249
rect 1456 258 1712 322
rect 1456 5 1512 258
rect 3018 0 3074 525
rect 4474 0 4530 525
rect 6038 0 6094 525
rect 6429 309 7122 321
rect 6429 249 6441 309
rect 7110 249 7122 309
rect 6429 238 7122 249
rect 7494 0 7550 525
rect 9058 0 9114 525
rect 10514 0 10570 525
rect 12078 0 12134 525
rect 12329 309 13022 321
rect 12329 249 12341 309
rect 13010 249 13022 309
rect 12329 237 13022 249
rect 13534 0 13590 525
<< via2 >>
rect 532 1028 1201 1088
rect 6432 1028 7101 1088
rect 12332 1028 13001 1088
rect 541 249 1210 309
rect 6441 249 7110 309
rect 12341 249 13010 309
<< metal3 >>
rect 519 1088 1215 1099
rect 519 1028 532 1088
rect 1201 1028 1215 1088
rect 519 1016 1215 1028
rect 6420 1088 7115 1099
rect 6420 1028 6432 1088
rect 7101 1028 7115 1088
rect 6420 1016 7115 1028
rect 12320 1088 13015 1099
rect 12320 1028 12332 1088
rect 13001 1028 13015 1088
rect 12320 1016 13015 1028
rect 529 309 1222 321
rect 529 249 541 309
rect 1210 249 1222 309
rect 529 238 1222 249
rect 6429 309 7122 321
rect 6429 249 6441 309
rect 7110 249 7122 309
rect 6429 238 7122 249
rect 12329 309 13022 321
rect 12329 249 12341 309
rect 13010 249 13022 309
rect 12329 237 13022 249
<< via3 >>
rect 532 1028 1201 1088
rect 6432 1028 7101 1088
rect 12332 1028 13001 1088
rect 541 249 1210 309
rect 6441 249 7110 309
rect 12341 249 13010 309
<< metal4 >>
rect 519 1088 1215 1099
rect 519 1028 532 1088
rect 1201 1028 1215 1088
rect 519 1016 1215 1028
rect 6420 1088 7115 1099
rect 6420 1028 6432 1088
rect 7101 1028 7115 1088
rect 6420 1016 7115 1028
rect 12320 1088 13015 1099
rect 12320 1028 12332 1088
rect 13001 1028 13015 1088
rect 12320 1016 13015 1028
rect 529 309 1222 321
rect 529 249 541 309
rect 1210 249 1222 309
rect 529 238 1222 249
rect 6429 309 7122 321
rect 6429 249 6441 309
rect 7110 249 7122 309
rect 6429 238 7122 249
rect 12329 309 13022 321
rect 12329 249 12341 309
rect 13010 249 13022 309
rect 12329 237 13022 249
<< via4 >>
rect 532 1028 1201 1088
rect 6432 1028 7101 1088
rect 12332 1028 13001 1088
rect 541 249 1210 309
rect 6441 249 7110 309
rect 12341 249 13010 309
<< metal5 >>
rect 351 1088 13247 1235
rect 351 1028 532 1088
rect 1201 1028 6432 1088
rect 7101 1028 12332 1088
rect 13001 1028 13247 1088
rect 351 915 13247 1028
rect 351 309 13247 435
rect 351 249 541 309
rect 1210 249 6441 309
rect 7110 249 12341 309
rect 13010 249 13247 309
rect 351 115 13247 249
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1653775443
transform 1 0 499 0 1 278
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_1
timestamp 1653775443
transform 1 0 12819 0 1 278
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1653775443
transform 1 0 1619 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_2
timestamp 1653775443
transform 1 0 4083 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_4
timestamp 1653775443
transform 1 0 6547 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_6
timestamp 1653775443
transform 1 0 9011 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_8
timestamp 1653775443
transform 1 0 11475 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1653775443
transform 1 0 2963 0 1 278
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_1
timestamp 1653775443
transform 1 0 5427 0 1 278
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_2
timestamp 1653775443
transform 1 0 7891 0 1 278
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_3
timestamp 1653775443
transform 1 0 10355 0 1 278
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1653775443
transform 1 0 723 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_1
timestamp 1653775443
transform 1 0 2067 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_2
timestamp 1653775443
transform 1 0 3187 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_3
timestamp 1653775443
transform 1 0 4531 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_4
timestamp 1653775443
transform 1 0 5651 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_5
timestamp 1653775443
transform 1 0 6995 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_6
timestamp 1653775443
transform 1 0 8115 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_7
timestamp 1653775443
transform 1 0 9459 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_8
timestamp 1653775443
transform 1 0 10579 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_9
timestamp 1653775443
transform 1 0 11923 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1653775443
transform 1 0 1171 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_1
timestamp 1653775443
transform 1 0 2515 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_2
timestamp 1653775443
transform 1 0 3635 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_3
timestamp 1653775443
transform 1 0 4979 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_4
timestamp 1653775443
transform 1 0 6099 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_5
timestamp 1653775443
transform 1 0 7443 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_6
timestamp 1653775443
transform 1 0 8563 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_7
timestamp 1653775443
transform 1 0 9907 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_8
timestamp 1653775443
transform 1 0 11027 0 1 278
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_9
timestamp 1653775443
transform 1 0 12371 0 1 278
box -86 -86 534 870
<< labels >>
flabel metal2 0 5 56 239 0 FreeSans 400 90 0 0 gpio_defaults[0]
port 1 nsew
flabel metal2 1456 5 1512 239 0 FreeSans 400 90 0 0 gpio_defaults[1]
port 2 nsew
flabel metal2 12078 0 12134 234 0 FreeSans 400 90 0 0 gpio_defaults[8]
port 9 nsew
flabel metal2 13534 0 13590 234 0 FreeSans 400 90 0 0 gpio_defaults[9]
port 10 nsew
flabel metal2 3018 0 3074 234 0 FreeSans 400 90 0 0 gpio_defaults[2]
port 3 nsew
flabel metal2 4474 0 4530 234 0 FreeSans 400 90 0 0 gpio_defaults[3]
port 4 nsew
flabel metal2 6038 0 6094 234 0 FreeSans 400 90 0 0 gpio_defaults[4]
port 5 nsew
flabel metal2 7494 0 7550 234 0 FreeSans 400 90 0 0 gpio_defaults[5]
port 6 nsew
flabel metal2 9058 0 9114 234 0 FreeSans 400 90 0 0 gpio_defaults[6]
port 7 nsew
flabel metal2 10514 0 10570 234 0 FreeSans 400 90 0 0 gpio_defaults[7]
port 8 nsew
flabel metal5 351 915 490 1235 0 FreeSans 1600 0 0 0 VDD
port 11 nsew
flabel metal5 351 115 490 435 0 FreeSans 1600 0 0 0 VSS
port 12 nsew
<< end >>
