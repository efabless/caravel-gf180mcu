magic
tech gf180mcuC
magscale 6 5
timestamp 1654634570
<< metal5 >>
rect 0 648 324 756
rect 0 432 108 648
rect 0 324 216 432
rect 0 108 108 324
rect 0 0 324 108
<< properties >>
string FIXED_BBOX 0 0 432 756
<< end >>
