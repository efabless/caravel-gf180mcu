magic
tech gf180mcuC
magscale 1 10
timestamp 1638586442
<< metal5 >>
tri 528 1376 544 1392 se
rect 544 1376 704 1424
tri 704 1376 720 1392 sw
tri 512 1328 528 1344 se
rect 528 1328 720 1376
tri 720 1328 736 1344 sw
tri 256 1296 287 1328 se
tri 287 1312 303 1328 sw
rect 287 1296 319 1312
tri 319 1296 335 1312 sw
rect 512 1296 736 1328
tri 944 1312 960 1328 se
tri 912 1296 928 1312 se
rect 928 1296 960 1312
tri 192 1232 256 1296 se
rect 256 1280 351 1296
tri 351 1280 367 1296 sw
rect 256 1248 383 1280
tri 383 1248 415 1280 sw
tri 463 1264 495 1296 se
rect 495 1264 752 1296
tri 752 1264 784 1296 sw
tri 880 1280 896 1296 se
rect 896 1280 960 1296
tri 415 1248 431 1264 se
rect 431 1248 816 1264
tri 816 1248 832 1264 sw
tri 832 1248 864 1280 se
rect 864 1248 960 1280
rect 256 1232 960 1248
tri 960 1232 1056 1328 sw
tri 192 1200 224 1232 ne
rect 224 1184 1024 1232
tri 1024 1200 1056 1232 nw
tri 224 1136 272 1184 ne
tri 256 1072 272 1088 se
rect 272 1072 976 1184
tri 976 1136 1024 1184 nw
tri 976 1072 992 1088 sw
rect 1254 1084 1307 1095
rect 1382 1084 1435 1095
rect 1499 1084 1574 1095
rect 1617 1084 1691 1095
rect 1830 1084 1905 1095
rect 1958 1084 2011 1095
rect 1243 1073 1318 1084
rect 1371 1073 1446 1084
rect 256 1056 576 1072
tri 576 1056 592 1072 nw
tri 656 1056 672 1072 ne
rect 672 1056 992 1072
tri 224 1008 256 1040 se
rect 256 1008 480 1056
tri 144 992 160 1008 se
rect 160 992 480 1008
rect 96 848 480 992
tri 480 976 560 1056 nw
tri 688 976 768 1056 ne
rect 768 1008 992 1056
rect 1233 1052 1329 1073
tri 992 1008 1024 1040 sw
rect 768 992 1088 1008
tri 1088 992 1104 1008 sw
rect 768 848 1152 992
rect 1233 977 1265 1052
rect 1297 977 1329 1052
rect 1233 956 1329 977
rect 1361 1052 1457 1073
rect 1361 977 1393 1052
rect 1425 977 1457 1052
rect 1361 956 1457 977
rect 1489 1063 1585 1084
rect 1489 1031 1521 1063
rect 1553 1031 1585 1063
rect 1489 1009 1585 1031
rect 1617 1073 1702 1084
rect 1819 1073 1905 1084
rect 1947 1073 2022 1084
rect 1617 1052 1713 1073
rect 1489 999 1574 1009
rect 1489 967 1521 999
rect 1243 945 1318 956
rect 1361 945 1446 956
rect 1489 945 1585 967
rect 1254 935 1307 945
rect 1361 935 1435 945
rect 1499 935 1585 945
rect 1617 935 1649 1052
rect 1681 935 1713 1052
rect 1809 1063 1905 1073
rect 1809 1031 1851 1063
rect 1937 1052 2033 1073
rect 1809 1020 1883 1031
rect 1819 1009 1894 1020
rect 1830 999 1905 1009
rect 1862 967 1905 999
rect 1809 956 1905 967
rect 1937 977 1969 1052
rect 2001 977 2033 1052
rect 1937 956 2033 977
rect 2065 977 2097 1095
rect 2129 977 2161 1095
rect 2065 956 2161 977
rect 2193 1084 2267 1095
rect 2342 1084 2395 1095
rect 2459 1084 2534 1095
rect 2193 1073 2278 1084
rect 2331 1073 2406 1084
rect 2193 1052 2289 1073
rect 1809 945 1894 956
rect 1947 945 2022 956
rect 2075 945 2150 956
rect 1809 935 1883 945
rect 1958 935 2011 945
rect 2086 935 2139 945
rect 2193 935 2225 1052
rect 2257 1031 2289 1052
rect 2321 1052 2417 1073
rect 2321 977 2353 1052
rect 2385 1031 2417 1052
rect 2449 1063 2545 1084
rect 2449 1031 2481 1063
rect 2513 1031 2545 1063
rect 2449 1009 2545 1031
rect 2449 999 2534 1009
rect 2385 977 2417 999
rect 2321 956 2417 977
rect 2449 967 2481 999
rect 2331 945 2406 956
rect 2449 945 2545 967
rect 2342 935 2395 945
rect 2459 935 2545 945
rect 1361 871 1393 935
rect 1809 871 1841 935
rect 1361 860 1435 871
rect 1489 860 1574 871
rect 1617 860 1691 871
rect 1766 860 1841 871
rect 1361 849 1446 860
tri 144 832 160 848 ne
rect 160 832 480 848
tri 208 800 240 832 ne
rect 240 784 480 832
tri 480 784 544 848 sw
rect 240 768 544 784
tri 240 752 256 768 ne
rect 256 752 544 768
rect 256 736 528 752
tri 528 736 544 752 nw
tri 704 784 768 848 se
rect 768 832 1088 848
tri 1088 832 1104 848 nw
rect 768 784 1008 832
tri 1008 800 1040 832 nw
rect 1361 828 1457 849
rect 1489 839 1585 860
rect 704 768 1008 784
rect 704 752 992 768
tri 992 752 1008 768 nw
tri 704 736 720 752 ne
rect 720 736 992 752
tri 256 720 272 736 ne
tri 256 704 272 720 se
rect 272 704 528 736
tri 224 656 256 688 se
rect 256 672 512 704
tri 512 688 528 704 nw
rect 720 704 976 736
tri 976 720 992 736 nw
tri 976 704 992 720 sw
rect 1361 711 1393 828
rect 1425 711 1457 828
rect 1553 807 1585 839
rect 1489 775 1585 807
rect 1489 743 1521 775
rect 1553 743 1585 775
rect 1489 721 1585 743
rect 1499 711 1585 721
rect 1617 849 1702 860
rect 1755 849 1841 860
rect 1617 828 1713 849
rect 1617 711 1649 828
rect 1681 807 1713 828
rect 1745 828 1841 849
rect 1745 753 1777 828
rect 1809 753 1841 828
rect 1745 732 1841 753
rect 1873 753 1905 871
rect 1937 753 1969 871
rect 2001 753 2033 871
rect 2065 860 2150 871
rect 2193 860 2267 871
rect 2331 860 2406 871
rect 2065 839 2161 860
rect 2129 807 2161 839
rect 2075 796 2161 807
rect 1873 732 2033 753
rect 2065 775 2161 796
rect 2065 743 2097 775
rect 2129 743 2161 775
rect 1755 721 1841 732
rect 1883 721 2022 732
rect 2065 721 2161 743
rect 1766 711 1841 721
rect 1894 711 1937 721
rect 1969 711 2011 721
rect 2075 711 2161 721
rect 2193 849 2278 860
rect 2193 828 2289 849
rect 2193 711 2225 828
rect 2257 807 2289 828
rect 2321 839 2417 860
rect 2321 807 2353 839
rect 2385 807 2417 839
rect 2321 775 2417 807
rect 2321 743 2353 775
rect 2321 721 2417 743
rect 2331 711 2417 721
tri 720 688 736 704 ne
rect 256 656 496 672
tri 496 656 512 672 nw
rect 736 672 992 704
tri 736 656 752 672 ne
rect 752 656 992 672
tri 992 656 1024 688 sw
tri 192 608 224 640 se
rect 224 624 496 656
rect 224 608 480 624
tri 480 608 496 624 nw
rect 752 624 1024 656
tri 752 608 768 624 ne
rect 768 608 1024 624
tri 1024 608 1056 640 sw
tri 192 512 288 608 ne
rect 288 592 480 608
rect 288 576 468 592
tri 468 580 480 592 nw
rect 768 592 960 608
tri 768 585 774 592 ne
rect 774 585 960 592
tri 774 580 779 585 ne
rect 288 560 384 576
tri 384 560 400 576 nw
rect 288 544 352 560
tri 352 544 368 560 nw
tri 411 544 443 576 ne
rect 443 564 468 576
rect 443 544 448 564
tri 448 544 468 564 nw
rect 779 576 960 585
rect 779 564 804 576
tri 779 544 800 564 ne
rect 800 544 804 564
tri 804 544 836 576 nw
tri 848 560 864 576 ne
rect 864 560 960 576
tri 880 544 896 560 ne
rect 896 544 960 560
rect 288 512 304 544
tri 304 512 336 544 nw
tri 912 512 944 544 ne
rect 944 512 960 544
tri 960 512 1056 608 nw
<< fillblock >>
rect 66 458 1173 1443
rect 1208 679 2580 1129
<< end >>
