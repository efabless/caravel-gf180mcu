magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 540 216 756
rect 108 432 216 540
<< properties >>
string FIXED_BBOX 0 -216 324 756
<< end >>
