* Simple POR testbench

.include /usr/share/pdk/gf180mcuC/libs.ref/gf180mcu_pr/spice/design.hspice
.lib /usr/share/pdk/gf180mcuC/libs.ref/gf180mcu_pr/spice/sm141064.hspice typical
.lib /usr/share/pdk/gf180mcuC/libs.ref/gf180mcu_pr/spice/sm141064.hspice res_typical
.lib /usr/share/pdk/gf180mcuC/libs.ref/gf180mcu_pr/spice/sm141064.hspice mimcap_typical
.include simple_por.spice

V0 VDD 0 PWL(0 0 100u 5 5m 5)

X0 VDD 0 POR PORB simple_por

.control
tran 1u 75m
plot V(VDD) V(POR) V(PORB)
.endc
