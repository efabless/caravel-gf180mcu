magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< metal1 >>
rect 1101 2992 1587 3292
rect 1249 2492 1384 2992
rect 1604 2871 1656 2883
rect 1604 2685 1656 2697
rect 1436 2599 1448 2651
rect 1542 2599 1554 2651
rect 1094 2171 1494 2185
rect 1094 1999 1310 2171
rect 1478 1999 1494 2171
rect 1094 1985 1494 1999
rect 2580 1980 2780 2180
rect 1222 592 1356 1483
rect 1424 1342 1437 1414
rect 1511 1342 1524 1414
rect 1553 1271 1605 1283
rect 1553 705 1605 717
rect 1111 292 1596 592
<< via1 >>
rect 1604 2697 1656 2871
rect 1448 2599 1542 2651
rect 1310 1999 1478 2171
rect 1607 1995 1775 2167
rect 1437 1342 1511 1414
rect 1553 717 1605 1271
<< metal2 >>
rect 1604 2885 1673 2888
rect 1602 2871 1673 2885
rect 1602 2697 1604 2871
rect 1656 2697 1673 2871
rect 1602 2683 1673 2697
rect 1446 2651 1544 2665
rect 1446 2599 1448 2651
rect 1542 2599 1544 2651
rect 1446 2584 1544 2599
rect 1446 2185 1513 2584
rect 1294 2171 1513 2185
rect 1604 2182 1673 2683
rect 1294 1999 1310 2171
rect 1478 1999 1513 2171
rect 1294 1985 1513 1999
rect 1435 1414 1513 1985
rect 1435 1342 1437 1414
rect 1511 1342 1513 1414
rect 1435 1327 1513 1342
rect 1578 2167 1788 2182
rect 1578 1995 1607 2167
rect 1775 1995 1788 2167
rect 1578 1982 1788 1995
rect 1578 1285 1649 1982
rect 1551 1271 1649 1285
rect 1551 717 1553 1271
rect 1605 717 1649 1271
rect 1551 703 1649 717
use std_inverter  X0
timestamp 1655304105
transform 1 0 1322 0 1 1642
box 265 -1350 1460 1650
use pmos_6p0_GUW2N9  XM2 primitives
timestamp 1655304105
transform 1 0 1474 0 1 1028
box -378 -586 368 586
use nmos_6p0_BUMBUS  XM3 primitives
timestamp 1655304105
transform 1 0 1505 0 1 2760
box -334 -332 334 332
<< labels >>
flabel metal1 1094 1985 1294 2185 0 FreeSans 1280 0 0 0 Vin
port 2 nsew
flabel metal1 1206 3043 1406 3243 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 1268 357 1468 557 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 2580 1980 2780 2180 0 FreeSans 1280 0 0 0 Vout
port 3 nsew
<< end >>
