magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 72 720 216 756
rect 36 684 216 720
rect 0 612 216 684
rect 0 144 108 612
rect 0 72 216 144
rect 36 36 216 72
rect 72 0 216 36
<< properties >>
string FIXED_BBOX 0 -216 324 756
<< end >>
