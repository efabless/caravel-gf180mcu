magic
tech gf180mcuC
magscale 1 10
timestamp 1669052252
<< checkpaint >>
rect -5616 68968 783615 1022000
rect -2000 -2000 783615 68968
<< metal2 >>
rect 104752 943800 104828 944076
rect 104898 943800 104974 944076
rect 105044 943800 105120 944076
rect 105190 943800 105266 944076
rect 116647 943800 116723 944076
rect 116858 943800 116934 944076
rect 117360 943800 117436 944076
rect 117502 943800 117578 944076
rect 117731 943800 117807 944076
rect 118252 943800 118328 944076
rect 159752 943800 159828 944076
rect 159898 943800 159974 944076
rect 160044 943800 160120 944076
rect 160190 943800 160266 944076
rect 171647 943800 171723 944076
rect 171858 943800 171934 944076
rect 172360 943800 172436 944076
rect 172502 943800 172578 944076
rect 172731 943800 172807 944076
rect 173252 943800 173328 944076
rect 214752 943800 214828 944076
rect 214898 943800 214974 944076
rect 215044 943800 215120 944076
rect 215190 943800 215266 944076
rect 226647 943800 226723 944076
rect 226858 943800 226934 944076
rect 227360 943800 227436 944076
rect 227502 943800 227578 944076
rect 227731 943800 227807 944076
rect 228252 943800 228328 944076
rect 269752 943800 269828 944076
rect 269898 943800 269974 944076
rect 270044 943800 270120 944076
rect 270190 943800 270266 944076
rect 281647 943800 281723 944076
rect 281858 943800 281934 944076
rect 282360 943800 282436 944076
rect 282502 943800 282578 944076
rect 282731 943800 282807 944076
rect 283252 943800 283328 944076
rect 324752 943800 324828 944076
rect 324898 943800 324974 944076
rect 325044 943800 325120 944076
rect 325190 943800 325266 944076
rect 336647 943800 336723 944076
rect 336858 943800 336934 944076
rect 337360 943800 337436 944076
rect 337502 943800 337578 944076
rect 337731 943800 337807 944076
rect 338252 943800 338328 944076
rect 434752 943800 434828 944076
rect 434898 943800 434974 944076
rect 435044 943800 435120 944076
rect 435190 943800 435266 944076
rect 446647 943800 446723 944076
rect 446858 943800 446934 944076
rect 447360 943800 447436 944076
rect 447502 943800 447578 944076
rect 447731 943800 447807 944076
rect 448252 943800 448328 944076
rect 489752 943800 489828 944076
rect 489898 943800 489974 944076
rect 490044 943800 490120 944076
rect 490190 943800 490266 944076
rect 501647 943800 501723 944076
rect 501858 943800 501934 944076
rect 502360 943800 502436 944076
rect 502502 943800 502578 944076
rect 502731 943800 502807 944076
rect 503252 943800 503328 944076
rect 544752 943800 544828 944076
rect 544898 943800 544974 944076
rect 545044 943800 545120 944076
rect 545190 943800 545266 944076
rect 556647 943800 556723 944076
rect 556858 943800 556934 944076
rect 557360 943800 557436 944076
rect 557502 943800 557578 944076
rect 557731 943800 557807 944076
rect 558252 943800 558328 944076
rect 654752 943800 654828 944076
rect 654898 943800 654974 944076
rect 655044 943800 655120 944076
rect 655190 943800 655266 944076
rect 666647 943800 666723 944076
rect 666858 943800 666934 944076
rect 667360 943800 667436 944076
rect 667502 943800 667578 944076
rect 667731 943800 667807 944076
rect 668252 943800 668328 944076
rect 705800 920172 706076 920248
rect 705800 920026 706076 920102
rect 705800 919880 706076 919956
rect 705800 919734 706076 919810
rect 69924 919252 70200 919328
rect 69924 918731 70200 918807
rect 69924 918502 70200 918578
rect 69924 918360 70200 918436
rect 69924 917858 70200 917934
rect 69924 917647 70200 917723
rect 705800 908277 706076 908353
rect 705800 908066 706076 908142
rect 705800 907564 706076 907640
rect 705800 907422 706076 907498
rect 705800 907193 706076 907269
rect 705800 906672 706076 906748
rect 69924 906190 70200 906266
rect 69924 906044 70200 906120
rect 69924 905898 70200 905974
rect 69924 905752 70200 905828
rect 705800 834172 706076 834248
rect 705800 834026 706076 834102
rect 705800 833880 706076 833956
rect 705800 833734 706076 833810
rect 705800 822277 706076 822353
rect 705800 822066 706076 822142
rect 705800 821564 706076 821640
rect 705800 821422 706076 821498
rect 705800 821193 706076 821269
rect 705800 820672 706076 820748
rect 69924 755252 70200 755328
rect 69924 754731 70200 754807
rect 69924 754502 70200 754578
rect 69924 754360 70200 754436
rect 69924 753858 70200 753934
rect 69924 753647 70200 753723
rect 705800 748172 706076 748248
rect 705800 748026 706076 748102
rect 705800 747880 706076 747956
rect 705800 747734 706076 747810
rect 69924 742190 70200 742266
rect 69924 742044 70200 742120
rect 69924 741898 70200 741974
rect 69924 741752 70200 741828
rect 705800 736277 706076 736353
rect 705800 736066 706076 736142
rect 705800 735564 706076 735640
rect 705800 735422 706076 735498
rect 705800 735193 706076 735269
rect 705800 734672 706076 734748
rect 69924 714252 70200 714328
rect 69924 713731 70200 713807
rect 69924 713502 70200 713578
rect 69924 713360 70200 713436
rect 69924 712858 70200 712934
rect 69924 712647 70200 712723
rect 705800 705172 706076 705248
rect 705800 705026 706076 705102
rect 705800 704880 706076 704956
rect 705800 704734 706076 704810
rect 69924 701190 70200 701266
rect 69924 701044 70200 701120
rect 69924 700898 70200 700974
rect 69924 700752 70200 700828
rect 705800 693277 706076 693353
rect 705800 693066 706076 693142
rect 705800 692564 706076 692640
rect 705800 692422 706076 692498
rect 705800 692193 706076 692269
rect 705800 691672 706076 691748
rect 69924 673252 70200 673328
rect 69924 672731 70200 672807
rect 69924 672502 70200 672578
rect 69924 672360 70200 672436
rect 69924 671858 70200 671934
rect 69924 671647 70200 671723
rect 705800 662172 706076 662248
rect 705800 662026 706076 662102
rect 705800 661880 706076 661956
rect 705800 661734 706076 661810
rect 69924 660190 70200 660266
rect 69924 660044 70200 660120
rect 69924 659898 70200 659974
rect 69924 659752 70200 659828
rect 705800 650277 706076 650353
rect 705800 650066 706076 650142
rect 705800 649564 706076 649640
rect 705800 649422 706076 649498
rect 705800 649193 706076 649269
rect 705800 648672 706076 648748
rect 69924 632252 70200 632328
rect 69924 631731 70200 631807
rect 69924 631502 70200 631578
rect 69924 631360 70200 631436
rect 69924 630858 70200 630934
rect 69924 630647 70200 630723
rect 69924 619190 70200 619266
rect 705800 619172 706076 619248
rect 69924 619044 70200 619120
rect 705800 619026 706076 619102
rect 69924 618898 70200 618974
rect 705800 618880 706076 618956
rect 69924 618752 70200 618828
rect 705800 618734 706076 618810
rect 705800 607277 706076 607353
rect 705800 607066 706076 607142
rect 705800 606564 706076 606640
rect 705800 606422 706076 606498
rect 705800 606193 706076 606269
rect 705800 605672 706076 605748
rect 69924 591252 70200 591328
rect 69924 590731 70200 590807
rect 69924 590502 70200 590578
rect 69924 590360 70200 590436
rect 69924 589858 70200 589934
rect 69924 589647 70200 589723
rect 69924 578190 70200 578266
rect 69924 578044 70200 578120
rect 69924 577898 70200 577974
rect 69924 577752 70200 577828
rect 705800 576172 706076 576248
rect 705800 576026 706076 576102
rect 705800 575880 706076 575956
rect 705800 575734 706076 575810
rect 705800 564277 706076 564353
rect 705800 564066 706076 564142
rect 705800 563564 706076 563640
rect 705800 563422 706076 563498
rect 705800 563193 706076 563269
rect 705800 562672 706076 562748
rect 69924 550252 70200 550328
rect 69924 549731 70200 549807
rect 69924 549502 70200 549578
rect 69924 549360 70200 549436
rect 69924 548858 70200 548934
rect 69924 548647 70200 548723
rect 69924 537190 70200 537266
rect 69924 537044 70200 537120
rect 69924 536898 70200 536974
rect 69924 536752 70200 536828
rect 705800 533172 706076 533248
rect 705800 533026 706076 533102
rect 705800 532880 706076 532956
rect 705800 532734 706076 532810
rect 705800 521277 706076 521353
rect 705800 521066 706076 521142
rect 705800 520564 706076 520640
rect 705800 520422 706076 520498
rect 705800 520193 706076 520269
rect 705800 519672 706076 519748
rect 69924 509252 70200 509328
rect 69924 508731 70200 508807
rect 69924 508502 70200 508578
rect 69924 508360 70200 508436
rect 69924 507858 70200 507934
rect 69924 507647 70200 507723
rect 69924 496190 70200 496266
rect 69924 496044 70200 496120
rect 69924 495898 70200 495974
rect 69924 495752 70200 495828
rect 69924 386252 70200 386328
rect 69924 385731 70200 385807
rect 69924 385502 70200 385578
rect 69924 385360 70200 385436
rect 69924 384858 70200 384934
rect 69924 384647 70200 384723
rect 69924 373190 70200 373266
rect 69924 373044 70200 373120
rect 69924 372898 70200 372974
rect 69924 372752 70200 372828
rect 705800 361172 706076 361248
rect 705800 361026 706076 361102
rect 705800 360880 706076 360956
rect 705800 360734 706076 360810
rect 705800 349277 706076 349353
rect 705800 349066 706076 349142
rect 705800 348564 706076 348640
rect 705800 348422 706076 348498
rect 705800 348193 706076 348269
rect 705800 347672 706076 347748
rect 69924 345252 70200 345328
rect 69924 344731 70200 344807
rect 69924 344502 70200 344578
rect 69924 344360 70200 344436
rect 69924 343858 70200 343934
rect 69924 343647 70200 343723
rect 69924 332190 70200 332266
rect 69924 332044 70200 332120
rect 69924 331898 70200 331974
rect 69924 331752 70200 331828
rect 705800 318172 706076 318248
rect 705800 318026 706076 318102
rect 705800 317880 706076 317956
rect 705800 317734 706076 317810
rect 705800 306277 706076 306353
rect 705800 306066 706076 306142
rect 705800 305564 706076 305640
rect 705800 305422 706076 305498
rect 705800 305193 706076 305269
rect 705800 304672 706076 304748
rect 69924 304252 70200 304328
rect 69924 303731 70200 303807
rect 69924 303502 70200 303578
rect 69924 303360 70200 303436
rect 69924 302858 70200 302934
rect 69924 302647 70200 302723
rect 69924 291190 70200 291266
rect 69924 291044 70200 291120
rect 69924 290898 70200 290974
rect 69924 290752 70200 290828
rect 705800 275172 706076 275248
rect 705800 275026 706076 275102
rect 705800 274880 706076 274956
rect 705800 274734 706076 274810
rect 69924 263252 70200 263328
rect 705800 263277 706076 263353
rect 705800 263066 706076 263142
rect 69924 262731 70200 262807
rect 69924 262502 70200 262578
rect 705800 262564 706076 262640
rect 69924 262360 70200 262436
rect 705800 262422 706076 262498
rect 705800 262193 706076 262269
rect 69924 261858 70200 261934
rect 69924 261647 70200 261723
rect 705800 261672 706076 261748
rect 69924 250190 70200 250266
rect 69924 250044 70200 250120
rect 69924 249898 70200 249974
rect 69924 249752 70200 249828
rect 705800 232172 706076 232248
rect 705800 232026 706076 232102
rect 705800 231880 706076 231956
rect 705800 231734 706076 231810
rect 69924 222252 70200 222328
rect 69924 221731 70200 221807
rect 69924 221502 70200 221578
rect 69924 221360 70200 221436
rect 69924 220858 70200 220934
rect 69924 220647 70200 220723
rect 705800 220277 706076 220353
rect 705800 220066 706076 220142
rect 705800 219564 706076 219640
rect 705800 219422 706076 219498
rect 705800 219193 706076 219269
rect 705800 218672 706076 218748
rect 69924 209190 70200 209266
rect 69924 209044 70200 209120
rect 69924 208898 70200 208974
rect 69924 208752 70200 208828
rect 705800 189172 706076 189248
rect 705800 189026 706076 189102
rect 705800 188880 706076 188956
rect 705800 188734 706076 188810
rect 69924 181252 70200 181328
rect 69924 180731 70200 180807
rect 69924 180502 70200 180578
rect 69924 180360 70200 180436
rect 69924 179858 70200 179934
rect 69924 179647 70200 179723
rect 705800 177277 706076 177353
rect 705800 177066 706076 177142
rect 705800 176564 706076 176640
rect 705800 176422 706076 176498
rect 705800 176193 706076 176269
rect 705800 175672 706076 175748
rect 69924 168190 70200 168266
rect 69924 168044 70200 168120
rect 69924 167898 70200 167974
rect 69924 167752 70200 167828
rect 705621 146172 706010 146248
rect 705621 146026 706010 146102
rect 705621 145880 706010 145956
rect 705621 145734 706010 145810
rect 705621 134277 706020 134353
rect 705621 134066 706020 134142
rect 705621 133564 706020 133640
rect 705621 133422 706020 133498
rect 705621 133193 706020 133269
rect 705621 132672 706020 132748
rect 705800 103172 706076 103248
rect 705800 103026 706076 103102
rect 705800 102880 706076 102956
rect 705800 102734 706076 102810
rect 705800 91277 706076 91353
rect 705800 91066 706076 91142
rect 705800 90564 706076 90640
rect 705800 90422 706076 90498
rect 705800 90193 706076 90269
rect 705800 89672 706076 89748
rect 161193 69925 161269 70225
rect 162066 69925 162142 70225
rect 174172 69924 174248 70200
rect 216193 70078 216269 70199
rect 216193 70002 217142 70078
rect 216193 69925 216269 70002
rect 217066 69925 217142 70002
rect 229172 69924 229248 70200
rect 325672 70088 325748 70113
rect 325672 70032 325678 70088
rect 325734 70032 325748 70088
rect 325672 69924 325748 70032
rect 326193 69924 326269 70156
rect 326422 70088 326498 70113
rect 326422 70032 326429 70088
rect 326485 70032 326498 70088
rect 326422 69924 326498 70032
rect 326564 70088 326640 70113
rect 326564 70032 326570 70088
rect 326626 70032 326640 70088
rect 326564 69924 326640 70032
rect 327066 70088 327142 70113
rect 327066 70032 327073 70088
rect 327129 70032 327142 70088
rect 327066 69924 327142 70032
rect 327277 70088 327353 70113
rect 338733 70097 338810 70202
rect 327277 70032 327287 70088
rect 327343 70032 327353 70088
rect 327277 69924 327353 70032
rect 338626 70088 338810 70097
rect 338626 70032 338634 70088
rect 338690 70032 338810 70088
rect 338626 70023 338810 70032
rect 338733 69924 338810 70023
rect 338880 69924 338956 70200
rect 339026 69924 339102 70200
rect 380672 70088 380748 70113
rect 380672 70032 380678 70088
rect 380734 70032 380748 70088
rect 380672 70000 380748 70032
rect 381193 70088 381269 70113
rect 381193 70032 381203 70088
rect 381259 70032 381269 70088
rect 381193 70000 381269 70032
rect 381422 70088 381498 70113
rect 381422 70032 381429 70088
rect 381485 70032 381498 70088
rect 381422 70000 381498 70032
rect 381564 70088 381640 70113
rect 381564 70032 381570 70088
rect 381626 70032 381640 70088
rect 381564 70000 381640 70032
rect 382066 70088 382142 70113
rect 382066 70032 382073 70088
rect 382129 70032 382142 70088
rect 382066 70000 382142 70032
rect 382277 70088 382353 70113
rect 393734 70097 393810 70198
rect 382277 70032 382287 70088
rect 382343 70032 382353 70088
rect 382277 70000 382353 70032
rect 393626 70088 393810 70097
rect 393626 70032 393634 70088
rect 393690 70032 393810 70088
rect 393626 70023 393810 70032
rect 393734 69924 393810 70023
rect 393880 69924 393956 70200
rect 394026 69924 394102 70200
rect 435672 70088 435748 70113
rect 435672 70032 435678 70088
rect 435734 70032 435748 70088
rect 435672 70000 435748 70032
rect 436193 70088 436269 70113
rect 436193 70032 436203 70088
rect 436259 70032 436269 70088
rect 436193 70000 436269 70032
rect 436422 70088 436498 70113
rect 436422 70032 436429 70088
rect 436485 70032 436498 70088
rect 436422 70000 436498 70032
rect 436564 70088 436640 70113
rect 436564 70032 436570 70088
rect 436626 70032 436640 70088
rect 436564 70000 436640 70032
rect 437066 70088 437142 70113
rect 437066 70032 437073 70088
rect 437129 70032 437142 70088
rect 437066 70000 437142 70032
rect 437277 69924 437353 70200
rect 448734 70097 448810 70198
rect 448626 70088 448810 70097
rect 448626 70032 448634 70088
rect 448690 70032 448810 70088
rect 448626 70023 448810 70032
rect 448734 69924 448810 70023
rect 448880 69924 448956 70200
rect 449026 69924 449102 70200
rect 449171 70111 449247 70200
rect 449171 70000 449248 70111
rect 490672 70088 490748 70113
rect 490672 70032 490678 70088
rect 490734 70032 490748 70088
rect 490672 70000 490748 70032
rect 491193 70088 491269 70113
rect 491193 70032 491203 70088
rect 491259 70032 491269 70088
rect 491193 70000 491269 70032
rect 491422 70088 491498 70113
rect 491422 70032 491429 70088
rect 491485 70032 491498 70088
rect 491422 70000 491498 70032
rect 491564 70088 491640 70113
rect 491564 70032 491570 70088
rect 491626 70032 491640 70088
rect 491564 70000 491640 70032
rect 492066 70088 492142 70113
rect 492066 70032 492073 70088
rect 492129 70032 492142 70088
rect 492066 70000 492142 70032
rect 449171 69924 449247 70000
rect 492277 69924 492353 70200
rect 503734 70097 503810 70198
rect 503626 70088 503810 70097
rect 503626 70032 503634 70088
rect 503690 70032 503810 70088
rect 503626 70023 503810 70032
rect 503734 69924 503810 70023
rect 503880 69924 503956 70200
rect 504026 69924 504102 70200
rect 504172 69924 504248 70200
rect 545672 69924 545748 70200
rect 546193 69924 546269 70200
rect 546422 69924 546498 70200
rect 546564 69923 546640 70199
rect 547066 69924 547142 70200
rect 547277 69924 547353 70200
rect 558734 69924 558810 70200
rect 558880 69924 558956 70200
rect 559026 69924 559102 70200
rect 559172 69924 559248 70200
<< via2 >>
rect 325678 70032 325734 70088
rect 326429 70032 326485 70088
rect 326570 70032 326626 70088
rect 327073 70032 327129 70088
rect 327287 70032 327343 70088
rect 338634 70032 338690 70088
rect 380678 70032 380734 70088
rect 381203 70032 381259 70088
rect 381429 70032 381485 70088
rect 381570 70032 381626 70088
rect 382073 70032 382129 70088
rect 382287 70032 382343 70088
rect 393634 70032 393690 70088
rect 435678 70032 435734 70088
rect 436203 70032 436259 70088
rect 436429 70032 436485 70088
rect 436570 70032 436626 70088
rect 437073 70032 437129 70088
rect 448634 70032 448690 70088
rect 490678 70032 490734 70088
rect 491203 70032 491259 70088
rect 491429 70032 491485 70088
rect 491570 70032 491626 70088
rect 492073 70032 492129 70088
rect 503634 70032 503690 70088
<< metal3 >>
rect 325655 70032 325678 70088
rect 325734 70032 326429 70088
rect 326485 70032 326570 70088
rect 326626 70032 327073 70088
rect 327129 70032 327287 70088
rect 327343 70032 338634 70088
rect 338690 70032 338706 70088
rect 380655 70032 380678 70088
rect 380734 70032 381203 70088
rect 381259 70032 381429 70088
rect 381485 70032 381570 70088
rect 381626 70032 382073 70088
rect 382129 70032 382287 70088
rect 382343 70032 393634 70088
rect 393690 70032 393710 70088
rect 435655 70032 435678 70088
rect 435734 70032 436203 70088
rect 436259 70032 436429 70088
rect 436485 70032 436570 70088
rect 436626 70032 437073 70088
rect 437129 70032 448634 70088
rect 448690 70032 448709 70088
rect 490655 70032 490678 70088
rect 490734 70032 491203 70088
rect 491259 70032 491429 70088
rect 491485 70032 491570 70088
rect 491626 70032 492073 70088
rect 492129 70032 503634 70088
rect 503690 70032 503723 70088
<< metal5 >>
rect 105500 1001600 117500 1013600
rect 160500 1001600 172500 1013600
rect 215500 1001600 227500 1013600
rect 270500 1001600 282500 1013600
rect 325500 1001600 337500 1013600
rect 380500 1001600 392500 1013600
rect 435500 1001600 447500 1013600
rect 490500 1001600 502500 1013600
rect 545500 1001600 557500 1013600
rect 600500 1001600 612500 1013600
rect 655500 1001600 667500 1013600
rect 400 906500 12400 918500
rect 763600 907500 775600 919500
rect 400 865500 12400 877500
rect 763600 864500 775600 876500
rect 400 824500 12400 836500
rect 763600 821500 775600 833500
rect 400 783500 12400 795500
rect 763600 778500 775600 790500
rect 400 742500 12400 754500
rect 763600 735500 775600 747500
rect 400 701500 12400 713500
rect 763600 692500 775600 704500
rect 400 660500 12400 672500
rect 763600 649500 775600 661500
rect 400 619500 12400 631500
rect 763600 606500 775600 618500
rect 400 578500 12400 590500
rect 763600 563500 775600 575500
rect 400 537500 12400 549500
rect 763600 520500 775600 532500
rect 400 496500 12400 508500
rect 763600 477500 775600 489500
rect 400 455500 12400 467500
rect 763600 434500 775600 446500
rect 400 414500 12400 426500
rect 763600 391500 775600 403500
rect 400 373500 12400 385500
rect 763600 348500 775600 360500
rect 400 332500 12400 344500
rect 763600 305500 775600 317500
rect 400 291500 12400 303500
rect 763600 262500 775600 274500
rect 400 250500 12400 262500
rect 400 209500 12400 221500
rect 763600 219500 775600 231500
rect 400 168500 12400 180500
rect 763600 176500 775600 188500
rect 400 127500 12400 139500
rect 763600 133500 775600 145500
rect 400 86500 12400 98500
rect 763600 90500 775600 102500
rect 106500 400 118500 12400
rect 161500 400 173500 12400
rect 216500 400 228500 12400
rect 271500 400 283500 12400
rect 326500 400 338500 12400
rect 381500 400 393500 12400
rect 436500 400 448500 12400
rect 491500 400 503500 12400
rect 546500 400 558500 12400
rect 601500 400 613500 12400
rect 656500 400 668500 12400
use gf180mcu_fd_io__bi_t  flash_clk_pad $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 1 0 380000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  flash_csb_pad
timestamp 1670211287
transform 1 0 325000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  flash_io0_pad
timestamp 1670211287
transform 1 0 435000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  flash_io1_pad
timestamp 1670211287
transform 1 0 490000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_0 $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 1 0 704000 0 1 0
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_1
timestamp 1670211287
transform -1 0 72000 0 -1 1014000
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_2
timestamp 1670211287
transform 0 1 0 -1 0 943000
box -32 13097 1032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1 $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 1 0 71000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_2
timestamp 1670211287
transform 1 0 73000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_3
timestamp 1670211287
transform 1 0 75000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_4
timestamp 1670211287
transform 1 0 77000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_5
timestamp 1670211287
transform 1 0 79000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_6
timestamp 1670211287
transform 1 0 81000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_7
timestamp 1670211287
transform 1 0 83000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_8
timestamp 1670211287
transform 1 0 85000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_9
timestamp 1670211287
transform 1 0 87000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_10
timestamp 1670211287
transform 1 0 89000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_11
timestamp 1670211287
transform 1 0 91000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_12
timestamp 1670211287
transform 1 0 93000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_13
timestamp 1670211287
transform 1 0 95000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_14
timestamp 1670211287
transform 1 0 97000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_15
timestamp 1670211287
transform 1 0 99000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_16
timestamp 1670211287
transform 1 0 101000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_17
timestamp 1670211287
transform 1 0 103000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_18
timestamp 1670211287
transform 1 0 120000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_19
timestamp 1670211287
transform 1 0 122000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_20
timestamp 1670211287
transform 1 0 124000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_21
timestamp 1670211287
transform 1 0 126000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_22
timestamp 1670211287
transform 1 0 128000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_23
timestamp 1670211287
transform 1 0 130000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_24
timestamp 1670211287
transform 1 0 132000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_25
timestamp 1670211287
transform 1 0 134000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_26
timestamp 1670211287
transform 1 0 136000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_27
timestamp 1670211287
transform 1 0 138000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_28
timestamp 1670211287
transform 1 0 140000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_29
timestamp 1670211287
transform 1 0 142000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_30
timestamp 1670211287
transform 1 0 144000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_31
timestamp 1670211287
transform 1 0 146000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_32
timestamp 1670211287
transform 1 0 148000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_33
timestamp 1670211287
transform 1 0 150000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_34
timestamp 1670211287
transform 1 0 152000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_35
timestamp 1670211287
transform 1 0 154000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_36
timestamp 1670211287
transform 1 0 156000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_37
timestamp 1670211287
transform 1 0 158000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_38
timestamp 1670211287
transform 1 0 175000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_39
timestamp 1670211287
transform 1 0 177000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_40
timestamp 1670211287
transform 1 0 179000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_41
timestamp 1670211287
transform 1 0 181000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_42
timestamp 1670211287
transform 1 0 183000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_43
timestamp 1670211287
transform 1 0 185000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_44
timestamp 1670211287
transform 1 0 187000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_45
timestamp 1670211287
transform 1 0 189000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_46
timestamp 1670211287
transform 1 0 213000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_47
timestamp 1670211287
transform 1 0 211000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_48
timestamp 1670211287
transform 1 0 209000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_49
timestamp 1670211287
transform 1 0 207000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_50
timestamp 1670211287
transform 1 0 205000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_51
timestamp 1670211287
transform 1 0 203000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_52
timestamp 1670211287
transform 1 0 201000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_53
timestamp 1670211287
transform 1 0 199000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_54
timestamp 1670211287
transform 1 0 197000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_55
timestamp 1670211287
transform 1 0 195000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_56
timestamp 1670211287
transform 1 0 193000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_57
timestamp 1670211287
transform 1 0 191000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_58
timestamp 1670211287
transform 1 0 246000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_59
timestamp 1670211287
transform 1 0 230000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_60
timestamp 1670211287
transform 1 0 232000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_61
timestamp 1670211287
transform 1 0 234000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_62
timestamp 1670211287
transform 1 0 236000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_63
timestamp 1670211287
transform 1 0 238000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_64
timestamp 1670211287
transform 1 0 240000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_65
timestamp 1670211287
transform 1 0 242000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_66
timestamp 1670211287
transform 1 0 244000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_67
timestamp 1670211287
transform 1 0 268000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_68
timestamp 1670211287
transform 1 0 266000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_69
timestamp 1670211287
transform 1 0 264000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_70
timestamp 1670211287
transform 1 0 262000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_71
timestamp 1670211287
transform 1 0 260000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_72
timestamp 1670211287
transform 1 0 258000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_73
timestamp 1670211287
transform 1 0 256000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_74
timestamp 1670211287
transform 1 0 254000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_75
timestamp 1670211287
transform 1 0 252000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_76
timestamp 1670211287
transform 1 0 250000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_77
timestamp 1670211287
transform 1 0 248000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_78
timestamp 1670211287
transform 1 0 303000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_79
timestamp 1670211287
transform 1 0 301000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_80
timestamp 1670211287
transform 1 0 285000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_81
timestamp 1670211287
transform 1 0 287000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_82
timestamp 1670211287
transform 1 0 289000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_83
timestamp 1670211287
transform 1 0 291000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_84
timestamp 1670211287
transform 1 0 293000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_85
timestamp 1670211287
transform 1 0 295000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_86
timestamp 1670211287
transform 1 0 297000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_87
timestamp 1670211287
transform 1 0 299000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_88
timestamp 1670211287
transform 1 0 323000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_89
timestamp 1670211287
transform 1 0 321000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_90
timestamp 1670211287
transform 1 0 319000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_91
timestamp 1670211287
transform 1 0 317000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_92
timestamp 1670211287
transform 1 0 315000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_93
timestamp 1670211287
transform 1 0 313000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_94
timestamp 1670211287
transform 1 0 311000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_95
timestamp 1670211287
transform 1 0 309000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_96
timestamp 1670211287
transform 1 0 307000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_97
timestamp 1670211287
transform 1 0 305000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_98
timestamp 1670211287
transform 1 0 360000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_99
timestamp 1670211287
transform 1 0 358000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_100
timestamp 1670211287
transform 1 0 356000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_101
timestamp 1670211287
transform 1 0 340000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_102
timestamp 1670211287
transform 1 0 342000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_103
timestamp 1670211287
transform 1 0 344000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_104
timestamp 1670211287
transform 1 0 346000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_105
timestamp 1670211287
transform 1 0 348000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_106
timestamp 1670211287
transform 1 0 350000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_107
timestamp 1670211287
transform 1 0 352000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_108
timestamp 1670211287
transform 1 0 354000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_109
timestamp 1670211287
transform 1 0 378000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_110
timestamp 1670211287
transform 1 0 376000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_111
timestamp 1670211287
transform 1 0 374000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_112
timestamp 1670211287
transform 1 0 372000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_113
timestamp 1670211287
transform 1 0 370000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_114
timestamp 1670211287
transform 1 0 368000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_115
timestamp 1670211287
transform 1 0 366000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_116
timestamp 1670211287
transform 1 0 364000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_117
timestamp 1670211287
transform 1 0 362000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_118
timestamp 1670211287
transform 1 0 415000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_119
timestamp 1670211287
transform 1 0 413000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_120
timestamp 1670211287
transform 1 0 411000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_121
timestamp 1670211287
transform 1 0 395000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_122
timestamp 1670211287
transform 1 0 397000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_123
timestamp 1670211287
transform 1 0 399000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_124
timestamp 1670211287
transform 1 0 401000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_125
timestamp 1670211287
transform 1 0 403000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_126
timestamp 1670211287
transform 1 0 405000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_127
timestamp 1670211287
transform 1 0 407000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_128
timestamp 1670211287
transform 1 0 409000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_129
timestamp 1670211287
transform 1 0 433000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_130
timestamp 1670211287
transform 1 0 431000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_131
timestamp 1670211287
transform 1 0 429000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_132
timestamp 1670211287
transform 1 0 427000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_133
timestamp 1670211287
transform 1 0 425000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_134
timestamp 1670211287
transform 1 0 423000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_135
timestamp 1670211287
transform 1 0 421000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_136
timestamp 1670211287
transform 1 0 419000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_137
timestamp 1670211287
transform 1 0 417000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_138
timestamp 1670211287
transform 1 0 450000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_139
timestamp 1670211287
transform 1 0 452000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_140
timestamp 1670211287
transform 1 0 454000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_141
timestamp 1670211287
transform 1 0 456000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_142
timestamp 1670211287
transform 1 0 458000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_143
timestamp 1670211287
transform 1 0 460000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_144
timestamp 1670211287
transform 1 0 462000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_145
timestamp 1670211287
transform 1 0 466000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_146
timestamp 1670211287
transform 1 0 464000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_147
timestamp 1670211287
transform 1 0 470000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_148
timestamp 1670211287
transform 1 0 468000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_149
timestamp 1670211287
transform 1 0 474000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_150
timestamp 1670211287
transform 1 0 472000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_151
timestamp 1670211287
transform 1 0 478000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_152
timestamp 1670211287
transform 1 0 476000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_153
timestamp 1670211287
transform 1 0 482000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_154
timestamp 1670211287
transform 1 0 480000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_155
timestamp 1670211287
transform 1 0 486000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_156
timestamp 1670211287
transform 1 0 484000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_157
timestamp 1670211287
transform 1 0 488000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_158
timestamp 1670211287
transform 1 0 505000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_159
timestamp 1670211287
transform 1 0 507000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_160
timestamp 1670211287
transform 1 0 509000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_161
timestamp 1670211287
transform 1 0 511000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_162
timestamp 1670211287
transform 1 0 513000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_163
timestamp 1670211287
transform 1 0 515000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_164
timestamp 1670211287
transform 1 0 517000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_165
timestamp 1670211287
transform 1 0 521000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_166
timestamp 1670211287
transform 1 0 519000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_167
timestamp 1670211287
transform 1 0 525000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_168
timestamp 1670211287
transform 1 0 523000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_169
timestamp 1670211287
transform 1 0 529000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_170
timestamp 1670211287
transform 1 0 527000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_171
timestamp 1670211287
transform 1 0 533000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_172
timestamp 1670211287
transform 1 0 531000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_173
timestamp 1670211287
transform 1 0 537000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_174
timestamp 1670211287
transform 1 0 535000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_175
timestamp 1670211287
transform 1 0 541000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_176
timestamp 1670211287
transform 1 0 539000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_177
timestamp 1670211287
transform 1 0 543000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_178
timestamp 1670211287
transform 1 0 560000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_179
timestamp 1670211287
transform 1 0 562000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_180
timestamp 1670211287
transform 1 0 564000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_181
timestamp 1670211287
transform 1 0 566000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_182
timestamp 1670211287
transform 1 0 568000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_183
timestamp 1670211287
transform 1 0 570000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_184
timestamp 1670211287
transform 1 0 572000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_185
timestamp 1670211287
transform 1 0 576000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_186
timestamp 1670211287
transform 1 0 574000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_187
timestamp 1670211287
transform 1 0 580000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_188
timestamp 1670211287
transform 1 0 578000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_189
timestamp 1670211287
transform 1 0 584000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_190
timestamp 1670211287
transform 1 0 582000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_191
timestamp 1670211287
transform 1 0 588000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_192
timestamp 1670211287
transform 1 0 586000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_193
timestamp 1670211287
transform 1 0 592000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_194
timestamp 1670211287
transform 1 0 590000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_195
timestamp 1670211287
transform 1 0 596000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_196
timestamp 1670211287
transform 1 0 594000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_197
timestamp 1670211287
transform 1 0 598000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_198
timestamp 1670211287
transform 1 0 615000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_199
timestamp 1670211287
transform 1 0 617000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_200
timestamp 1670211287
transform 1 0 619000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_201
timestamp 1670211287
transform 1 0 621000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_202
timestamp 1670211287
transform 1 0 623000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_203
timestamp 1670211287
transform 1 0 625000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_204
timestamp 1670211287
transform 1 0 627000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_205
timestamp 1670211287
transform 1 0 631000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_206
timestamp 1670211287
transform 1 0 629000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_207
timestamp 1670211287
transform 1 0 635000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_208
timestamp 1670211287
transform 1 0 633000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_209
timestamp 1670211287
transform 1 0 639000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_210
timestamp 1670211287
transform 1 0 637000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_211
timestamp 1670211287
transform 1 0 643000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_212
timestamp 1670211287
transform 1 0 641000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_213
timestamp 1670211287
transform 1 0 647000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_214
timestamp 1670211287
transform 1 0 645000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_215
timestamp 1670211287
transform 1 0 651000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_216
timestamp 1670211287
transform 1 0 649000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_217
timestamp 1670211287
transform 1 0 653000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_218
timestamp 1670211287
transform 1 0 670000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_219
timestamp 1670211287
transform 1 0 672000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_220
timestamp 1670211287
transform 1 0 674000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_221
timestamp 1670211287
transform 1 0 676000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_222
timestamp 1670211287
transform 1 0 678000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_223
timestamp 1670211287
transform 1 0 680000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_224
timestamp 1670211287
transform 1 0 682000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_225
timestamp 1670211287
transform 1 0 686000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_226
timestamp 1670211287
transform 1 0 684000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_227
timestamp 1670211287
transform 1 0 690000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_228
timestamp 1670211287
transform 1 0 688000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_229
timestamp 1670211287
transform 1 0 694000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_230
timestamp 1670211287
transform 1 0 692000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_231
timestamp 1670211287
transform 1 0 698000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_232
timestamp 1670211287
transform 1 0 696000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_233
timestamp 1670211287
transform 1 0 702000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_234
timestamp 1670211287
transform 1 0 700000 0 1 0
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_238
timestamp 1670211287
transform 0 -1 776000 1 0 71000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_239
timestamp 1670211287
transform 0 -1 776000 1 0 73000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_240
timestamp 1670211287
transform 0 -1 776000 1 0 75000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_241
timestamp 1670211287
transform 0 -1 776000 1 0 77000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_242
timestamp 1670211287
transform 0 -1 776000 1 0 79000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_243
timestamp 1670211287
transform 0 -1 776000 1 0 81000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_244
timestamp 1670211287
transform 0 -1 776000 1 0 83000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_245
timestamp 1670211287
transform 0 -1 776000 1 0 85000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_246
timestamp 1670211287
transform 0 -1 776000 1 0 87000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_247
timestamp 1670211287
transform 0 -1 776000 1 0 112000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_248
timestamp 1670211287
transform 0 -1 776000 1 0 108000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_249
timestamp 1670211287
transform 0 -1 776000 1 0 110000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_250
timestamp 1670211287
transform 0 -1 776000 1 0 116000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_251
timestamp 1670211287
transform 0 -1 776000 1 0 114000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_252
timestamp 1670211287
transform 0 -1 776000 1 0 120000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_253
timestamp 1670211287
transform 0 -1 776000 1 0 118000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_254
timestamp 1670211287
transform 0 -1 776000 1 0 124000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_255
timestamp 1670211287
transform 0 -1 776000 1 0 122000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_256
timestamp 1670211287
transform 0 -1 776000 1 0 128000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_257
timestamp 1670211287
transform 0 -1 776000 1 0 126000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_258
timestamp 1670211287
transform 0 -1 776000 1 0 130000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_259
timestamp 1670211287
transform 0 -1 776000 1 0 106000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_260
timestamp 1670211287
transform 0 -1 776000 1 0 104000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_261
timestamp 1670211287
transform 0 -1 776000 1 0 147000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_262
timestamp 1670211287
transform 0 -1 776000 1 0 149000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_263
timestamp 1670211287
transform 0 -1 776000 1 0 151000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_264
timestamp 1670211287
transform 0 -1 776000 1 0 153000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_265
timestamp 1670211287
transform 0 -1 776000 1 0 157000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_266
timestamp 1670211287
transform 0 -1 776000 1 0 155000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_267
timestamp 1670211287
transform 0 -1 776000 1 0 161000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_268
timestamp 1670211287
transform 0 -1 776000 1 0 159000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_269
timestamp 1670211287
transform 0 -1 776000 1 0 165000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_270
timestamp 1670211287
transform 0 -1 776000 1 0 163000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_271
timestamp 1670211287
transform 0 -1 776000 1 0 169000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_272
timestamp 1670211287
transform 0 -1 776000 1 0 167000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_273
timestamp 1670211287
transform 0 -1 776000 1 0 173000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_274
timestamp 1670211287
transform 0 -1 776000 1 0 171000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_275
timestamp 1670211287
transform 0 -1 776000 1 0 190000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_276
timestamp 1670211287
transform 0 -1 776000 1 0 192000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_277
timestamp 1670211287
transform 0 -1 776000 1 0 194000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_278
timestamp 1670211287
transform 0 -1 776000 1 0 196000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_279
timestamp 1670211287
transform 0 -1 776000 1 0 200000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_280
timestamp 1670211287
transform 0 -1 776000 1 0 198000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_281
timestamp 1670211287
transform 0 -1 776000 1 0 204000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_282
timestamp 1670211287
transform 0 -1 776000 1 0 202000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_283
timestamp 1670211287
transform 0 -1 776000 1 0 208000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_284
timestamp 1670211287
transform 0 -1 776000 1 0 206000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_285
timestamp 1670211287
transform 0 -1 776000 1 0 212000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_286
timestamp 1670211287
transform 0 -1 776000 1 0 210000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_287
timestamp 1670211287
transform 0 -1 776000 1 0 216000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_288
timestamp 1670211287
transform 0 -1 776000 1 0 214000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_289
timestamp 1670211287
transform 0 -1 776000 1 0 233000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_290
timestamp 1670211287
transform 0 -1 776000 1 0 235000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_291
timestamp 1670211287
transform 0 -1 776000 1 0 237000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_292
timestamp 1670211287
transform 0 -1 776000 1 0 239000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_293
timestamp 1670211287
transform 0 -1 776000 1 0 243000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_294
timestamp 1670211287
transform 0 -1 776000 1 0 241000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_295
timestamp 1670211287
transform 0 -1 776000 1 0 247000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_296
timestamp 1670211287
transform 0 -1 776000 1 0 245000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_297
timestamp 1670211287
transform 0 -1 776000 1 0 251000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_298
timestamp 1670211287
transform 0 -1 776000 1 0 249000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_299
timestamp 1670211287
transform 0 -1 776000 1 0 255000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_300
timestamp 1670211287
transform 0 -1 776000 1 0 253000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_301
timestamp 1670211287
transform 0 -1 776000 1 0 259000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_302
timestamp 1670211287
transform 0 -1 776000 1 0 257000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_303
timestamp 1670211287
transform 0 -1 776000 1 0 276000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_304
timestamp 1670211287
transform 0 -1 776000 1 0 278000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_305
timestamp 1670211287
transform 0 -1 776000 1 0 280000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_306
timestamp 1670211287
transform 0 -1 776000 1 0 282000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_307
timestamp 1670211287
transform 0 -1 776000 1 0 286000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_308
timestamp 1670211287
transform 0 -1 776000 1 0 284000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_309
timestamp 1670211287
transform 0 -1 776000 1 0 290000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_310
timestamp 1670211287
transform 0 -1 776000 1 0 288000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_311
timestamp 1670211287
transform 0 -1 776000 1 0 294000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_312
timestamp 1670211287
transform 0 -1 776000 1 0 292000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_313
timestamp 1670211287
transform 0 -1 776000 1 0 298000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_314
timestamp 1670211287
transform 0 -1 776000 1 0 296000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_315
timestamp 1670211287
transform 0 -1 776000 1 0 302000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_316
timestamp 1670211287
transform 0 -1 776000 1 0 300000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_317
timestamp 1670211287
transform 0 -1 776000 1 0 319000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_318
timestamp 1670211287
transform 0 -1 776000 1 0 321000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_319
timestamp 1670211287
transform 0 -1 776000 1 0 323000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_320
timestamp 1670211287
transform 0 -1 776000 1 0 325000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_321
timestamp 1670211287
transform 0 -1 776000 1 0 329000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_322
timestamp 1670211287
transform 0 -1 776000 1 0 327000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_323
timestamp 1670211287
transform 0 -1 776000 1 0 333000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_324
timestamp 1670211287
transform 0 -1 776000 1 0 331000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_325
timestamp 1670211287
transform 0 -1 776000 1 0 337000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_326
timestamp 1670211287
transform 0 -1 776000 1 0 335000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_327
timestamp 1670211287
transform 0 -1 776000 1 0 341000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_328
timestamp 1670211287
transform 0 -1 776000 1 0 339000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_329
timestamp 1670211287
transform 0 -1 776000 1 0 345000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_330
timestamp 1670211287
transform 0 -1 776000 1 0 343000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_331
timestamp 1670211287
transform 0 -1 776000 1 0 362000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_332
timestamp 1670211287
transform 0 -1 776000 1 0 364000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_333
timestamp 1670211287
transform 0 -1 776000 1 0 366000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_334
timestamp 1670211287
transform 0 -1 776000 1 0 368000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_335
timestamp 1670211287
transform 0 -1 776000 1 0 372000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_336
timestamp 1670211287
transform 0 -1 776000 1 0 370000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_337
timestamp 1670211287
transform 0 -1 776000 1 0 376000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_338
timestamp 1670211287
transform 0 -1 776000 1 0 374000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_339
timestamp 1670211287
transform 0 -1 776000 1 0 380000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_340
timestamp 1670211287
transform 0 -1 776000 1 0 378000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_341
timestamp 1670211287
transform 0 -1 776000 1 0 384000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_342
timestamp 1670211287
transform 0 -1 776000 1 0 382000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_343
timestamp 1670211287
transform 0 -1 776000 1 0 388000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_344
timestamp 1670211287
transform 0 -1 776000 1 0 386000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_345
timestamp 1670211287
transform 0 -1 776000 1 0 405000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_346
timestamp 1670211287
transform 0 -1 776000 1 0 407000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_347
timestamp 1670211287
transform 0 -1 776000 1 0 409000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_348
timestamp 1670211287
transform 0 -1 776000 1 0 411000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_349
timestamp 1670211287
transform 0 -1 776000 1 0 415000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_350
timestamp 1670211287
transform 0 -1 776000 1 0 413000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_351
timestamp 1670211287
transform 0 -1 776000 1 0 419000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_352
timestamp 1670211287
transform 0 -1 776000 1 0 417000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_353
timestamp 1670211287
transform 0 -1 776000 1 0 423000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_354
timestamp 1670211287
transform 0 -1 776000 1 0 421000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_355
timestamp 1670211287
transform 0 -1 776000 1 0 427000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_356
timestamp 1670211287
transform 0 -1 776000 1 0 425000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_357
timestamp 1670211287
transform 0 -1 776000 1 0 431000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_358
timestamp 1670211287
transform 0 -1 776000 1 0 429000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_359
timestamp 1670211287
transform 0 -1 776000 1 0 448000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_360
timestamp 1670211287
transform 0 -1 776000 1 0 450000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_361
timestamp 1670211287
transform 0 -1 776000 1 0 452000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_362
timestamp 1670211287
transform 0 -1 776000 1 0 454000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_363
timestamp 1670211287
transform 0 -1 776000 1 0 458000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_364
timestamp 1670211287
transform 0 -1 776000 1 0 456000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_365
timestamp 1670211287
transform 0 -1 776000 1 0 462000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_366
timestamp 1670211287
transform 0 -1 776000 1 0 460000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_367
timestamp 1670211287
transform 0 -1 776000 1 0 466000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_368
timestamp 1670211287
transform 0 -1 776000 1 0 464000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_369
timestamp 1670211287
transform 0 -1 776000 1 0 470000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_370
timestamp 1670211287
transform 0 -1 776000 1 0 468000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_371
timestamp 1670211287
transform 0 -1 776000 1 0 474000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_372
timestamp 1670211287
transform 0 -1 776000 1 0 472000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_373
timestamp 1670211287
transform 0 -1 776000 1 0 491000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_374
timestamp 1670211287
transform 0 -1 776000 1 0 493000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_375
timestamp 1670211287
transform 0 -1 776000 1 0 495000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_376
timestamp 1670211287
transform 0 -1 776000 1 0 497000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_377
timestamp 1670211287
transform 0 -1 776000 1 0 501000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_378
timestamp 1670211287
transform 0 -1 776000 1 0 499000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_379
timestamp 1670211287
transform 0 -1 776000 1 0 505000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_380
timestamp 1670211287
transform 0 -1 776000 1 0 503000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_381
timestamp 1670211287
transform 0 -1 776000 1 0 509000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_382
timestamp 1670211287
transform 0 -1 776000 1 0 507000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_383
timestamp 1670211287
transform 0 -1 776000 1 0 513000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_384
timestamp 1670211287
transform 0 -1 776000 1 0 511000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_385
timestamp 1670211287
transform 0 -1 776000 1 0 517000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_386
timestamp 1670211287
transform 0 -1 776000 1 0 515000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_387
timestamp 1670211287
transform 0 -1 776000 1 0 534000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_388
timestamp 1670211287
transform 0 -1 776000 1 0 536000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_389
timestamp 1670211287
transform 0 -1 776000 1 0 538000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_390
timestamp 1670211287
transform 0 -1 776000 1 0 540000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_391
timestamp 1670211287
transform 0 -1 776000 1 0 544000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_392
timestamp 1670211287
transform 0 -1 776000 1 0 542000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_393
timestamp 1670211287
transform 0 -1 776000 1 0 548000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_394
timestamp 1670211287
transform 0 -1 776000 1 0 546000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_395
timestamp 1670211287
transform 0 -1 776000 1 0 552000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_396
timestamp 1670211287
transform 0 -1 776000 1 0 550000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_397
timestamp 1670211287
transform 0 -1 776000 1 0 556000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_398
timestamp 1670211287
transform 0 -1 776000 1 0 554000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_399
timestamp 1670211287
transform 0 -1 776000 1 0 560000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_400
timestamp 1670211287
transform 0 -1 776000 1 0 558000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_401
timestamp 1670211287
transform 0 -1 776000 1 0 577000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_402
timestamp 1670211287
transform 0 -1 776000 1 0 579000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_403
timestamp 1670211287
transform 0 -1 776000 1 0 581000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_404
timestamp 1670211287
transform 0 -1 776000 1 0 583000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_405
timestamp 1670211287
transform 0 -1 776000 1 0 587000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_406
timestamp 1670211287
transform 0 -1 776000 1 0 585000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_407
timestamp 1670211287
transform 0 -1 776000 1 0 591000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_408
timestamp 1670211287
transform 0 -1 776000 1 0 589000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_409
timestamp 1670211287
transform 0 -1 776000 1 0 595000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_410
timestamp 1670211287
transform 0 -1 776000 1 0 593000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_411
timestamp 1670211287
transform 0 -1 776000 1 0 599000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_412
timestamp 1670211287
transform 0 -1 776000 1 0 597000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_413
timestamp 1670211287
transform 0 -1 776000 1 0 603000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_414
timestamp 1670211287
transform 0 -1 776000 1 0 601000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_415
timestamp 1670211287
transform 0 -1 776000 1 0 620000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_416
timestamp 1670211287
transform 0 -1 776000 1 0 622000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_417
timestamp 1670211287
transform 0 -1 776000 1 0 624000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_418
timestamp 1670211287
transform 0 -1 776000 1 0 626000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_419
timestamp 1670211287
transform 0 -1 776000 1 0 630000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_420
timestamp 1670211287
transform 0 -1 776000 1 0 628000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_421
timestamp 1670211287
transform 0 -1 776000 1 0 634000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_422
timestamp 1670211287
transform 0 -1 776000 1 0 632000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_423
timestamp 1670211287
transform 0 -1 776000 1 0 638000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_424
timestamp 1670211287
transform 0 -1 776000 1 0 636000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_425
timestamp 1670211287
transform 0 -1 776000 1 0 642000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_426
timestamp 1670211287
transform 0 -1 776000 1 0 640000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_427
timestamp 1670211287
transform 0 -1 776000 1 0 646000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_428
timestamp 1670211287
transform 0 -1 776000 1 0 644000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_429
timestamp 1670211287
transform 0 -1 776000 1 0 663000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_430
timestamp 1670211287
transform 0 -1 776000 1 0 665000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_431
timestamp 1670211287
transform 0 -1 776000 1 0 667000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_432
timestamp 1670211287
transform 0 -1 776000 1 0 669000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_433
timestamp 1670211287
transform 0 -1 776000 1 0 673000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_434
timestamp 1670211287
transform 0 -1 776000 1 0 671000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_435
timestamp 1670211287
transform 0 -1 776000 1 0 677000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_436
timestamp 1670211287
transform 0 -1 776000 1 0 675000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_437
timestamp 1670211287
transform 0 -1 776000 1 0 681000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_438
timestamp 1670211287
transform 0 -1 776000 1 0 679000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_439
timestamp 1670211287
transform 0 -1 776000 1 0 685000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_440
timestamp 1670211287
transform 0 -1 776000 1 0 683000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_441
timestamp 1670211287
transform 0 -1 776000 1 0 689000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_442
timestamp 1670211287
transform 0 -1 776000 1 0 687000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_443
timestamp 1670211287
transform 0 -1 776000 1 0 706000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_444
timestamp 1670211287
transform 0 -1 776000 1 0 708000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_445
timestamp 1670211287
transform 0 -1 776000 1 0 710000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_446
timestamp 1670211287
transform 0 -1 776000 1 0 712000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_447
timestamp 1670211287
transform 0 -1 776000 1 0 716000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_448
timestamp 1670211287
transform 0 -1 776000 1 0 714000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_449
timestamp 1670211287
transform 0 -1 776000 1 0 720000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_450
timestamp 1670211287
transform 0 -1 776000 1 0 718000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_451
timestamp 1670211287
transform 0 -1 776000 1 0 724000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_452
timestamp 1670211287
transform 0 -1 776000 1 0 722000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_453
timestamp 1670211287
transform 0 -1 776000 1 0 728000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_454
timestamp 1670211287
transform 0 -1 776000 1 0 726000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_455
timestamp 1670211287
transform 0 -1 776000 1 0 732000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_456
timestamp 1670211287
transform 0 -1 776000 1 0 730000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_457
timestamp 1670211287
transform 0 -1 776000 1 0 749000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_458
timestamp 1670211287
transform 0 -1 776000 1 0 751000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_459
timestamp 1670211287
transform 0 -1 776000 1 0 753000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_460
timestamp 1670211287
transform 0 -1 776000 1 0 755000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_461
timestamp 1670211287
transform 0 -1 776000 1 0 759000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_462
timestamp 1670211287
transform 0 -1 776000 1 0 757000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_463
timestamp 1670211287
transform 0 -1 776000 1 0 763000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_464
timestamp 1670211287
transform 0 -1 776000 1 0 761000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_465
timestamp 1670211287
transform 0 -1 776000 1 0 767000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_466
timestamp 1670211287
transform 0 -1 776000 1 0 765000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_467
timestamp 1670211287
transform 0 -1 776000 1 0 771000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_468
timestamp 1670211287
transform 0 -1 776000 1 0 769000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_469
timestamp 1670211287
transform 0 -1 776000 1 0 775000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_470
timestamp 1670211287
transform 0 -1 776000 1 0 773000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_471
timestamp 1670211287
transform 0 -1 776000 1 0 792000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_472
timestamp 1670211287
transform 0 -1 776000 1 0 794000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_473
timestamp 1670211287
transform 0 -1 776000 1 0 796000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_474
timestamp 1670211287
transform 0 -1 776000 1 0 798000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_475
timestamp 1670211287
transform 0 -1 776000 1 0 802000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_476
timestamp 1670211287
transform 0 -1 776000 1 0 800000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_477
timestamp 1670211287
transform 0 -1 776000 1 0 806000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_478
timestamp 1670211287
transform 0 -1 776000 1 0 804000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_479
timestamp 1670211287
transform 0 -1 776000 1 0 810000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_480
timestamp 1670211287
transform 0 -1 776000 1 0 808000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_481
timestamp 1670211287
transform 0 -1 776000 1 0 814000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_482
timestamp 1670211287
transform 0 -1 776000 1 0 812000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_483
timestamp 1670211287
transform 0 -1 776000 1 0 818000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_484
timestamp 1670211287
transform 0 -1 776000 1 0 816000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_485
timestamp 1670211287
transform 0 -1 776000 1 0 835000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_486
timestamp 1670211287
transform 0 -1 776000 1 0 837000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_487
timestamp 1670211287
transform 0 -1 776000 1 0 839000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_488
timestamp 1670211287
transform 0 -1 776000 1 0 841000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_489
timestamp 1670211287
transform 0 -1 776000 1 0 845000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_490
timestamp 1670211287
transform 0 -1 776000 1 0 843000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_491
timestamp 1670211287
transform 0 -1 776000 1 0 849000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_492
timestamp 1670211287
transform 0 -1 776000 1 0 847000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_493
timestamp 1670211287
transform 0 -1 776000 1 0 853000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_494
timestamp 1670211287
transform 0 -1 776000 1 0 851000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_495
timestamp 1670211287
transform 0 -1 776000 1 0 857000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_496
timestamp 1670211287
transform 0 -1 776000 1 0 855000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_497
timestamp 1670211287
transform 0 -1 776000 1 0 861000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_498
timestamp 1670211287
transform 0 -1 776000 1 0 859000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_499
timestamp 1670211287
transform 0 -1 776000 1 0 878000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_500
timestamp 1670211287
transform 0 -1 776000 1 0 880000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_501
timestamp 1670211287
transform 0 -1 776000 1 0 882000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_502
timestamp 1670211287
transform 0 -1 776000 1 0 884000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_503
timestamp 1670211287
transform 0 -1 776000 1 0 888000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_504
timestamp 1670211287
transform 0 -1 776000 1 0 886000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_505
timestamp 1670211287
transform 0 -1 776000 1 0 892000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_506
timestamp 1670211287
transform 0 -1 776000 1 0 890000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_507
timestamp 1670211287
transform 0 -1 776000 1 0 896000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_508
timestamp 1670211287
transform 0 -1 776000 1 0 894000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_509
timestamp 1670211287
transform 0 -1 776000 1 0 900000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_510
timestamp 1670211287
transform 0 -1 776000 1 0 898000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_511
timestamp 1670211287
transform 0 -1 776000 1 0 904000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_512
timestamp 1670211287
transform 0 -1 776000 1 0 902000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_513
timestamp 1670211287
transform 0 -1 776000 1 0 925000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_514
timestamp 1670211287
transform 0 -1 776000 1 0 921000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_515
timestamp 1670211287
transform 0 -1 776000 1 0 923000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_516
timestamp 1670211287
transform 0 -1 776000 1 0 929000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_517
timestamp 1670211287
transform 0 -1 776000 1 0 927000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_518
timestamp 1670211287
transform 0 -1 776000 1 0 933000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_519
timestamp 1670211287
transform 0 -1 776000 1 0 931000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_520
timestamp 1670211287
transform 0 -1 776000 1 0 937000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_521
timestamp 1670211287
transform 0 -1 776000 1 0 935000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_522
timestamp 1670211287
transform 0 -1 776000 1 0 941000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_523
timestamp 1670211287
transform 0 -1 776000 1 0 939000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_524
timestamp 1670211287
transform -1 0 693000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_525
timestamp 1670211287
transform -1 0 695000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_526
timestamp 1670211287
transform -1 0 705000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_527
timestamp 1670211287
transform -1 0 703000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_528
timestamp 1670211287
transform -1 0 701000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_529
timestamp 1670211287
transform -1 0 699000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_530
timestamp 1670211287
transform -1 0 697000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_531
timestamp 1670211287
transform -1 0 677000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_532
timestamp 1670211287
transform -1 0 679000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_533
timestamp 1670211287
transform -1 0 681000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_534
timestamp 1670211287
transform -1 0 683000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_535
timestamp 1670211287
transform -1 0 685000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_536
timestamp 1670211287
transform -1 0 687000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_537
timestamp 1670211287
transform -1 0 691000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_538
timestamp 1670211287
transform -1 0 689000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_539
timestamp 1670211287
transform -1 0 675000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_540
timestamp 1670211287
transform -1 0 673000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_541
timestamp 1670211287
transform -1 0 671000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_542
timestamp 1670211287
transform -1 0 652000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_543
timestamp 1670211287
transform -1 0 650000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_544
timestamp 1670211287
transform -1 0 648000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_545
timestamp 1670211287
transform -1 0 654000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_546
timestamp 1670211287
transform -1 0 636000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_547
timestamp 1670211287
transform -1 0 634000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_548
timestamp 1670211287
transform -1 0 632000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_549
timestamp 1670211287
transform -1 0 644000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_550
timestamp 1670211287
transform -1 0 642000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_551
timestamp 1670211287
transform -1 0 640000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_552
timestamp 1670211287
transform -1 0 638000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_553
timestamp 1670211287
transform -1 0 646000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_554
timestamp 1670211287
transform -1 0 622000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_555
timestamp 1670211287
transform -1 0 620000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_556
timestamp 1670211287
transform -1 0 618000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_557
timestamp 1670211287
transform -1 0 630000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_558
timestamp 1670211287
transform -1 0 628000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_559
timestamp 1670211287
transform -1 0 626000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_560
timestamp 1670211287
transform -1 0 624000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_561
timestamp 1670211287
transform -1 0 616000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_562
timestamp 1670211287
transform -1 0 587000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_563
timestamp 1670211287
transform -1 0 589000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_564
timestamp 1670211287
transform -1 0 591000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_565
timestamp 1670211287
transform -1 0 593000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_566
timestamp 1670211287
transform -1 0 595000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_567
timestamp 1670211287
transform -1 0 597000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_568
timestamp 1670211287
transform -1 0 599000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_569
timestamp 1670211287
transform -1 0 575000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_570
timestamp 1670211287
transform -1 0 573000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_571
timestamp 1670211287
transform -1 0 581000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_572
timestamp 1670211287
transform -1 0 579000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_573
timestamp 1670211287
transform -1 0 577000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_574
timestamp 1670211287
transform -1 0 583000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_575
timestamp 1670211287
transform -1 0 585000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_576
timestamp 1670211287
transform -1 0 565000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_577
timestamp 1670211287
transform -1 0 563000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_578
timestamp 1670211287
transform -1 0 561000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_579
timestamp 1670211287
transform -1 0 571000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_580
timestamp 1670211287
transform -1 0 569000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_581
timestamp 1670211287
transform -1 0 567000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_582
timestamp 1670211287
transform -1 0 544000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_583
timestamp 1670211287
transform -1 0 542000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_584
timestamp 1670211287
transform -1 0 528000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_585
timestamp 1670211287
transform -1 0 530000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_586
timestamp 1670211287
transform -1 0 526000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_587
timestamp 1670211287
transform -1 0 536000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_588
timestamp 1670211287
transform -1 0 534000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_589
timestamp 1670211287
transform -1 0 532000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_590
timestamp 1670211287
transform -1 0 540000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_591
timestamp 1670211287
transform -1 0 538000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_592
timestamp 1670211287
transform -1 0 512000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_593
timestamp 1670211287
transform -1 0 514000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_594
timestamp 1670211287
transform -1 0 516000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_595
timestamp 1670211287
transform -1 0 518000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_596
timestamp 1670211287
transform -1 0 520000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_597
timestamp 1670211287
transform -1 0 522000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_598
timestamp 1670211287
transform -1 0 524000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_599
timestamp 1670211287
transform -1 0 506000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_600
timestamp 1670211287
transform -1 0 508000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_601
timestamp 1670211287
transform -1 0 510000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_602
timestamp 1670211287
transform -1 0 483000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_603
timestamp 1670211287
transform -1 0 481000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_604
timestamp 1670211287
transform -1 0 485000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_605
timestamp 1670211287
transform -1 0 487000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_606
timestamp 1670211287
transform -1 0 489000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_607
timestamp 1670211287
transform -1 0 467000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_608
timestamp 1670211287
transform -1 0 469000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_609
timestamp 1670211287
transform -1 0 471000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_610
timestamp 1670211287
transform -1 0 473000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_611
timestamp 1670211287
transform -1 0 475000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_612
timestamp 1670211287
transform -1 0 477000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_613
timestamp 1670211287
transform -1 0 479000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_614
timestamp 1670211287
transform -1 0 453000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_615
timestamp 1670211287
transform -1 0 451000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_616
timestamp 1670211287
transform -1 0 461000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_617
timestamp 1670211287
transform -1 0 459000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_618
timestamp 1670211287
transform -1 0 457000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_619
timestamp 1670211287
transform -1 0 455000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_620
timestamp 1670211287
transform -1 0 463000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_621
timestamp 1670211287
transform -1 0 465000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_622
timestamp 1670211287
transform -1 0 422000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_623
timestamp 1670211287
transform -1 0 424000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_624
timestamp 1670211287
transform -1 0 426000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_625
timestamp 1670211287
transform -1 0 428000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_626
timestamp 1670211287
transform -1 0 430000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_627
timestamp 1670211287
transform -1 0 432000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_628
timestamp 1670211287
transform -1 0 434000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_629
timestamp 1670211287
transform -1 0 406000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_630
timestamp 1670211287
transform -1 0 408000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_631
timestamp 1670211287
transform -1 0 410000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_632
timestamp 1670211287
transform -1 0 412000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_633
timestamp 1670211287
transform -1 0 414000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_634
timestamp 1670211287
transform -1 0 416000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_635
timestamp 1670211287
transform -1 0 418000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_636
timestamp 1670211287
transform -1 0 420000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_637
timestamp 1670211287
transform -1 0 400000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_638
timestamp 1670211287
transform -1 0 398000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_639
timestamp 1670211287
transform -1 0 396000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_640
timestamp 1670211287
transform -1 0 402000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_641
timestamp 1670211287
transform -1 0 404000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_642
timestamp 1670211287
transform -1 0 379000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_643
timestamp 1670211287
transform -1 0 377000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_644
timestamp 1670211287
transform -1 0 365000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_645
timestamp 1670211287
transform -1 0 367000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_646
timestamp 1670211287
transform -1 0 363000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_647
timestamp 1670211287
transform -1 0 361000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_648
timestamp 1670211287
transform -1 0 369000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_649
timestamp 1670211287
transform -1 0 375000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_650
timestamp 1670211287
transform -1 0 373000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_651
timestamp 1670211287
transform -1 0 371000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_652
timestamp 1670211287
transform -1 0 353000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_653
timestamp 1670211287
transform -1 0 351000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_654
timestamp 1670211287
transform -1 0 349000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_655
timestamp 1670211287
transform -1 0 347000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_656
timestamp 1670211287
transform -1 0 357000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_657
timestamp 1670211287
transform -1 0 355000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_658
timestamp 1670211287
transform -1 0 359000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_659
timestamp 1670211287
transform -1 0 345000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_660
timestamp 1670211287
transform -1 0 343000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_661
timestamp 1670211287
transform -1 0 341000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_662
timestamp 1670211287
transform -1 0 322000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_663
timestamp 1670211287
transform -1 0 320000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_664
timestamp 1670211287
transform -1 0 318000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_665
timestamp 1670211287
transform -1 0 316000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_666
timestamp 1670211287
transform -1 0 324000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_667
timestamp 1670211287
transform -1 0 302000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_668
timestamp 1670211287
transform -1 0 300000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_669
timestamp 1670211287
transform -1 0 306000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_670
timestamp 1670211287
transform -1 0 304000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_671
timestamp 1670211287
transform -1 0 312000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_672
timestamp 1670211287
transform -1 0 308000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_673
timestamp 1670211287
transform -1 0 310000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_674
timestamp 1670211287
transform -1 0 314000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_675
timestamp 1670211287
transform -1 0 286000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_676
timestamp 1670211287
transform -1 0 290000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_677
timestamp 1670211287
transform -1 0 288000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_678
timestamp 1670211287
transform -1 0 294000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_679
timestamp 1670211287
transform -1 0 292000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_680
timestamp 1670211287
transform -1 0 296000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_681
timestamp 1670211287
transform -1 0 298000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_682
timestamp 1670211287
transform -1 0 255000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_683
timestamp 1670211287
transform -1 0 257000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_684
timestamp 1670211287
transform -1 0 259000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_685
timestamp 1670211287
transform -1 0 261000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_686
timestamp 1670211287
transform -1 0 263000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_687
timestamp 1670211287
transform -1 0 265000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_688
timestamp 1670211287
transform -1 0 267000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_689
timestamp 1670211287
transform -1 0 269000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_690
timestamp 1670211287
transform -1 0 241000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_691
timestamp 1670211287
transform -1 0 243000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_692
timestamp 1670211287
transform -1 0 245000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_693
timestamp 1670211287
transform -1 0 247000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_694
timestamp 1670211287
transform -1 0 251000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_695
timestamp 1670211287
transform -1 0 249000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_696
timestamp 1670211287
transform -1 0 253000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_697
timestamp 1670211287
transform -1 0 237000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_698
timestamp 1670211287
transform -1 0 239000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_699
timestamp 1670211287
transform -1 0 233000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_700
timestamp 1670211287
transform -1 0 235000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_701
timestamp 1670211287
transform -1 0 231000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_702
timestamp 1670211287
transform -1 0 210000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_703
timestamp 1670211287
transform -1 0 212000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_704
timestamp 1670211287
transform -1 0 214000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_705
timestamp 1670211287
transform -1 0 196000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_706
timestamp 1670211287
transform -1 0 208000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_707
timestamp 1670211287
transform -1 0 206000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_708
timestamp 1670211287
transform -1 0 204000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_709
timestamp 1670211287
transform -1 0 202000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_710
timestamp 1670211287
transform -1 0 198000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_711
timestamp 1670211287
transform -1 0 200000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_712
timestamp 1670211287
transform -1 0 180000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_713
timestamp 1670211287
transform -1 0 182000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_714
timestamp 1670211287
transform -1 0 194000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_715
timestamp 1670211287
transform -1 0 190000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_716
timestamp 1670211287
transform -1 0 192000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_717
timestamp 1670211287
transform -1 0 186000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_718
timestamp 1670211287
transform -1 0 188000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_719
timestamp 1670211287
transform -1 0 184000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_720
timestamp 1670211287
transform -1 0 178000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_721
timestamp 1670211287
transform -1 0 176000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_722
timestamp 1670211287
transform -1 0 151000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_723
timestamp 1670211287
transform -1 0 155000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_724
timestamp 1670211287
transform -1 0 153000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_725
timestamp 1670211287
transform -1 0 159000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_726
timestamp 1670211287
transform -1 0 157000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_727
timestamp 1670211287
transform -1 0 139000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_728
timestamp 1670211287
transform -1 0 135000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_729
timestamp 1670211287
transform -1 0 137000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_730
timestamp 1670211287
transform -1 0 141000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_731
timestamp 1670211287
transform -1 0 149000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_732
timestamp 1670211287
transform -1 0 147000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_733
timestamp 1670211287
transform -1 0 143000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_734
timestamp 1670211287
transform -1 0 145000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_735
timestamp 1670211287
transform -1 0 123000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_736
timestamp 1670211287
transform -1 0 125000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_737
timestamp 1670211287
transform -1 0 121000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_738
timestamp 1670211287
transform -1 0 131000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_739
timestamp 1670211287
transform -1 0 133000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_740
timestamp 1670211287
transform -1 0 127000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_741
timestamp 1670211287
transform -1 0 129000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_742
timestamp 1670211287
transform -1 0 90000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_743
timestamp 1670211287
transform -1 0 92000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_744
timestamp 1670211287
transform -1 0 94000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_745
timestamp 1670211287
transform -1 0 96000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_746
timestamp 1670211287
transform -1 0 98000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_747
timestamp 1670211287
transform -1 0 104000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_748
timestamp 1670211287
transform -1 0 102000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_749
timestamp 1670211287
transform -1 0 100000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_750
timestamp 1670211287
transform -1 0 74000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_751
timestamp 1670211287
transform -1 0 76000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_752
timestamp 1670211287
transform -1 0 78000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_753
timestamp 1670211287
transform -1 0 80000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_754
timestamp 1670211287
transform -1 0 82000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_755
timestamp 1670211287
transform -1 0 84000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_756
timestamp 1670211287
transform -1 0 86000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_757
timestamp 1670211287
transform -1 0 88000 0 -1 1014000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_759
timestamp 1670211287
transform 0 1 0 -1 0 940000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_760
timestamp 1670211287
transform 0 1 0 -1 0 942000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_761
timestamp 1670211287
transform 0 1 0 -1 0 102000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_762
timestamp 1670211287
transform 0 1 0 -1 0 934000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_763
timestamp 1670211287
transform 0 1 0 -1 0 936000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_764
timestamp 1670211287
transform 0 1 0 -1 0 938000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_765
timestamp 1670211287
transform 0 1 0 -1 0 932000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_766
timestamp 1670211287
transform 0 1 0 -1 0 928000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_767
timestamp 1670211287
transform 0 1 0 -1 0 930000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_768
timestamp 1670211287
transform 0 1 0 -1 0 922000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_769
timestamp 1670211287
transform 0 1 0 -1 0 926000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_770
timestamp 1670211287
transform 0 1 0 -1 0 924000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_771
timestamp 1670211287
transform 0 1 0 -1 0 903000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_772
timestamp 1670211287
transform 0 1 0 -1 0 905000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_773
timestamp 1670211287
transform 0 1 0 -1 0 104000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_774
timestamp 1670211287
transform 0 1 0 -1 0 895000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_775
timestamp 1670211287
transform 0 1 0 -1 0 893000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_776
timestamp 1670211287
transform 0 1 0 -1 0 899000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_777
timestamp 1670211287
transform 0 1 0 -1 0 901000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_778
timestamp 1670211287
transform 0 1 0 -1 0 897000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_779
timestamp 1670211287
transform 0 1 0 -1 0 889000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_780
timestamp 1670211287
transform 0 1 0 -1 0 891000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_781
timestamp 1670211287
transform 0 1 0 -1 0 881000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_782
timestamp 1670211287
transform 0 1 0 -1 0 887000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_783
timestamp 1670211287
transform 0 1 0 -1 0 883000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_784
timestamp 1670211287
transform 0 1 0 -1 0 885000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_785
timestamp 1670211287
transform 0 1 0 -1 0 106000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_786
timestamp 1670211287
transform 0 1 0 -1 0 860000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_787
timestamp 1670211287
transform 0 1 0 -1 0 862000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_788
timestamp 1670211287
transform 0 1 0 -1 0 864000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_789
timestamp 1670211287
transform 0 1 0 -1 0 854000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_790
timestamp 1670211287
transform 0 1 0 -1 0 858000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_791
timestamp 1670211287
transform 0 1 0 -1 0 856000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_792
timestamp 1670211287
transform 0 1 0 -1 0 846000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_793
timestamp 1670211287
transform 0 1 0 -1 0 850000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_794
timestamp 1670211287
transform 0 1 0 -1 0 848000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_795
timestamp 1670211287
transform 0 1 0 -1 0 852000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_796
timestamp 1670211287
transform 0 1 0 -1 0 842000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_797
timestamp 1670211287
transform 0 1 0 -1 0 840000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_798
timestamp 1670211287
transform 0 1 0 -1 0 844000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_799
timestamp 1670211287
transform 0 1 0 -1 0 817000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_800
timestamp 1670211287
transform 0 1 0 -1 0 108000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_801
timestamp 1670211287
transform 0 1 0 -1 0 823000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_802
timestamp 1670211287
transform 0 1 0 -1 0 821000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_803
timestamp 1670211287
transform 0 1 0 -1 0 819000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_804
timestamp 1670211287
transform 0 1 0 -1 0 815000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_805
timestamp 1670211287
transform 0 1 0 -1 0 811000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_806
timestamp 1670211287
transform 0 1 0 -1 0 813000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_807
timestamp 1670211287
transform 0 1 0 -1 0 809000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_808
timestamp 1670211287
transform 0 1 0 -1 0 805000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_809
timestamp 1670211287
transform 0 1 0 -1 0 803000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_810
timestamp 1670211287
transform 0 1 0 -1 0 807000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_811
timestamp 1670211287
transform 0 1 0 -1 0 801000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_812
timestamp 1670211287
transform 0 1 0 -1 0 799000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_813
timestamp 1670211287
transform 0 1 0 -1 0 776000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_814
timestamp 1670211287
transform 0 1 0 -1 0 774000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_815
timestamp 1670211287
transform 0 1 0 -1 0 778000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_816
timestamp 1670211287
transform 0 1 0 -1 0 780000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_817
timestamp 1670211287
transform 0 1 0 -1 0 782000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_818
timestamp 1670211287
transform 0 1 0 -1 0 110000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_819
timestamp 1670211287
transform 0 1 0 -1 0 772000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_820
timestamp 1670211287
transform 0 1 0 -1 0 760000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_821
timestamp 1670211287
transform 0 1 0 -1 0 764000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_822
timestamp 1670211287
transform 0 1 0 -1 0 762000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_823
timestamp 1670211287
transform 0 1 0 -1 0 768000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_824
timestamp 1670211287
transform 0 1 0 -1 0 766000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_825
timestamp 1670211287
transform 0 1 0 -1 0 770000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_826
timestamp 1670211287
transform 0 1 0 -1 0 758000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_827
timestamp 1670211287
transform 0 1 0 -1 0 112000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_828
timestamp 1670211287
transform 0 1 0 -1 0 741000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_829
timestamp 1670211287
transform 0 1 0 -1 0 739000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_830
timestamp 1670211287
transform 0 1 0 -1 0 737000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_831
timestamp 1670211287
transform 0 1 0 -1 0 733000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_832
timestamp 1670211287
transform 0 1 0 -1 0 735000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_833
timestamp 1670211287
transform 0 1 0 -1 0 731000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_834
timestamp 1670211287
transform 0 1 0 -1 0 729000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_835
timestamp 1670211287
transform 0 1 0 -1 0 725000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_836
timestamp 1670211287
transform 0 1 0 -1 0 727000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_837
timestamp 1670211287
transform 0 1 0 -1 0 721000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_838
timestamp 1670211287
transform 0 1 0 -1 0 723000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_839
timestamp 1670211287
transform 0 1 0 -1 0 719000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_840
timestamp 1670211287
transform 0 1 0 -1 0 717000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_841
timestamp 1670211287
transform 0 1 0 -1 0 700000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_842
timestamp 1670211287
transform 0 1 0 -1 0 698000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_843
timestamp 1670211287
transform 0 1 0 -1 0 696000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_844
timestamp 1670211287
transform 0 1 0 -1 0 692000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_845
timestamp 1670211287
transform 0 1 0 -1 0 694000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_846
timestamp 1670211287
transform 0 1 0 -1 0 690000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_847
timestamp 1670211287
transform 0 1 0 -1 0 114000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_848
timestamp 1670211287
transform 0 1 0 -1 0 688000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_849
timestamp 1670211287
transform 0 1 0 -1 0 684000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_850
timestamp 1670211287
transform 0 1 0 -1 0 680000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_851
timestamp 1670211287
transform 0 1 0 -1 0 682000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_852
timestamp 1670211287
transform 0 1 0 -1 0 676000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_853
timestamp 1670211287
transform 0 1 0 -1 0 678000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_854
timestamp 1670211287
transform 0 1 0 -1 0 686000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_855
timestamp 1670211287
transform 0 1 0 -1 0 659000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_856
timestamp 1670211287
transform 0 1 0 -1 0 116000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_857
timestamp 1670211287
transform 0 1 0 -1 0 653000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_858
timestamp 1670211287
transform 0 1 0 -1 0 651000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_859
timestamp 1670211287
transform 0 1 0 -1 0 655000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_860
timestamp 1670211287
transform 0 1 0 -1 0 657000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_861
timestamp 1670211287
transform 0 1 0 -1 0 645000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_862
timestamp 1670211287
transform 0 1 0 -1 0 649000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_863
timestamp 1670211287
transform 0 1 0 -1 0 647000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_864
timestamp 1670211287
transform 0 1 0 -1 0 637000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_865
timestamp 1670211287
transform 0 1 0 -1 0 641000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_866
timestamp 1670211287
transform 0 1 0 -1 0 639000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_867
timestamp 1670211287
transform 0 1 0 -1 0 643000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_868
timestamp 1670211287
transform 0 1 0 -1 0 635000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_869
timestamp 1670211287
transform 0 1 0 -1 0 616000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_870
timestamp 1670211287
transform 0 1 0 -1 0 618000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_871
timestamp 1670211287
transform 0 1 0 -1 0 118000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_872
timestamp 1670211287
transform 0 1 0 -1 0 612000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_873
timestamp 1670211287
transform 0 1 0 -1 0 610000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_874
timestamp 1670211287
transform 0 1 0 -1 0 614000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_875
timestamp 1670211287
transform 0 1 0 -1 0 608000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_876
timestamp 1670211287
transform 0 1 0 -1 0 604000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_877
timestamp 1670211287
transform 0 1 0 -1 0 602000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_878
timestamp 1670211287
transform 0 1 0 -1 0 606000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_879
timestamp 1670211287
transform 0 1 0 -1 0 596000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_880
timestamp 1670211287
transform 0 1 0 -1 0 594000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_881
timestamp 1670211287
transform 0 1 0 -1 0 600000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_882
timestamp 1670211287
transform 0 1 0 -1 0 598000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_883
timestamp 1670211287
transform 0 1 0 -1 0 573000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_884
timestamp 1670211287
transform 0 1 0 -1 0 575000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_885
timestamp 1670211287
transform 0 1 0 -1 0 577000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_886
timestamp 1670211287
transform 0 1 0 -1 0 120000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_887
timestamp 1670211287
transform 0 1 0 -1 0 571000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_888
timestamp 1670211287
transform 0 1 0 -1 0 569000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_889
timestamp 1670211287
transform 0 1 0 -1 0 559000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_890
timestamp 1670211287
transform 0 1 0 -1 0 563000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_891
timestamp 1670211287
transform 0 1 0 -1 0 561000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_892
timestamp 1670211287
transform 0 1 0 -1 0 565000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_893
timestamp 1670211287
transform 0 1 0 -1 0 567000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_894
timestamp 1670211287
transform 0 1 0 -1 0 555000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_895
timestamp 1670211287
transform 0 1 0 -1 0 557000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_896
timestamp 1670211287
transform 0 1 0 -1 0 553000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_897
timestamp 1670211287
transform 0 1 0 -1 0 530000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_898
timestamp 1670211287
transform 0 1 0 -1 0 532000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_899
timestamp 1670211287
transform 0 1 0 -1 0 534000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_900
timestamp 1670211287
transform 0 1 0 -1 0 536000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_901
timestamp 1670211287
transform 0 1 0 -1 0 122000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_902
timestamp 1670211287
transform 0 1 0 -1 0 526000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_903
timestamp 1670211287
transform 0 1 0 -1 0 528000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_904
timestamp 1670211287
transform 0 1 0 -1 0 518000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_905
timestamp 1670211287
transform 0 1 0 -1 0 516000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_906
timestamp 1670211287
transform 0 1 0 -1 0 522000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_907
timestamp 1670211287
transform 0 1 0 -1 0 520000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_908
timestamp 1670211287
transform 0 1 0 -1 0 524000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_909
timestamp 1670211287
transform 0 1 0 -1 0 512000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_910
timestamp 1670211287
transform 0 1 0 -1 0 514000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_911
timestamp 1670211287
transform 0 1 0 -1 0 489000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_912
timestamp 1670211287
transform 0 1 0 -1 0 487000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_913
timestamp 1670211287
transform 0 1 0 -1 0 491000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_914
timestamp 1670211287
transform 0 1 0 -1 0 493000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_915
timestamp 1670211287
transform 0 1 0 -1 0 495000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_916
timestamp 1670211287
transform 0 1 0 -1 0 124000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_917
timestamp 1670211287
transform 0 1 0 -1 0 473000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_918
timestamp 1670211287
transform 0 1 0 -1 0 477000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_919
timestamp 1670211287
transform 0 1 0 -1 0 475000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_920
timestamp 1670211287
transform 0 1 0 -1 0 481000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_921
timestamp 1670211287
transform 0 1 0 -1 0 479000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_922
timestamp 1670211287
transform 0 1 0 -1 0 483000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_923
timestamp 1670211287
transform 0 1 0 -1 0 485000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_924
timestamp 1670211287
transform 0 1 0 -1 0 471000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_925
timestamp 1670211287
transform 0 1 0 -1 0 126000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_926
timestamp 1670211287
transform 0 1 0 -1 0 454000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_927
timestamp 1670211287
transform 0 1 0 -1 0 452000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_928
timestamp 1670211287
transform 0 1 0 -1 0 450000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_929
timestamp 1670211287
transform 0 1 0 -1 0 448000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_930
timestamp 1670211287
transform 0 1 0 -1 0 444000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_931
timestamp 1670211287
transform 0 1 0 -1 0 446000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_932
timestamp 1670211287
transform 0 1 0 -1 0 442000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_933
timestamp 1670211287
transform 0 1 0 -1 0 438000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_934
timestamp 1670211287
transform 0 1 0 -1 0 440000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_935
timestamp 1670211287
transform 0 1 0 -1 0 436000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_936
timestamp 1670211287
transform 0 1 0 -1 0 434000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_937
timestamp 1670211287
transform 0 1 0 -1 0 430000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_938
timestamp 1670211287
transform 0 1 0 -1 0 432000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_940
timestamp 1670211287
transform 0 1 0 -1 0 405000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_941
timestamp 1670211287
transform 0 1 0 -1 0 407000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_942
timestamp 1670211287
transform 0 1 0 -1 0 413000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_943
timestamp 1670211287
transform 0 1 0 -1 0 411000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_944
timestamp 1670211287
transform 0 1 0 -1 0 409000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_945
timestamp 1670211287
transform 0 1 0 -1 0 401000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_946
timestamp 1670211287
transform 0 1 0 -1 0 403000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_947
timestamp 1670211287
transform 0 1 0 -1 0 399000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_948
timestamp 1670211287
transform 0 1 0 -1 0 397000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_949
timestamp 1670211287
transform 0 1 0 -1 0 393000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_950
timestamp 1670211287
transform 0 1 0 -1 0 395000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_951
timestamp 1670211287
transform 0 1 0 -1 0 391000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_952
timestamp 1670211287
transform 0 1 0 -1 0 389000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_953
timestamp 1670211287
transform 0 1 0 -1 0 372000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_955
timestamp 1670211287
transform 0 1 0 -1 0 366000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_956
timestamp 1670211287
transform 0 1 0 -1 0 368000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_957
timestamp 1670211287
transform 0 1 0 -1 0 370000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_958
timestamp 1670211287
transform 0 1 0 -1 0 362000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_959
timestamp 1670211287
transform 0 1 0 -1 0 360000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_960
timestamp 1670211287
transform 0 1 0 -1 0 364000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_961
timestamp 1670211287
transform 0 1 0 -1 0 358000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_962
timestamp 1670211287
transform 0 1 0 -1 0 354000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_963
timestamp 1670211287
transform 0 1 0 -1 0 352000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_964
timestamp 1670211287
transform 0 1 0 -1 0 356000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_965
timestamp 1670211287
transform 0 1 0 -1 0 350000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_966
timestamp 1670211287
transform 0 1 0 -1 0 348000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_967
timestamp 1670211287
transform 0 1 0 -1 0 329000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_968
timestamp 1670211287
transform 0 1 0 -1 0 331000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_970
timestamp 1670211287
transform 0 1 0 -1 0 325000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_971
timestamp 1670211287
transform 0 1 0 -1 0 323000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_972
timestamp 1670211287
transform 0 1 0 -1 0 327000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_973
timestamp 1670211287
transform 0 1 0 -1 0 321000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_974
timestamp 1670211287
transform 0 1 0 -1 0 317000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_975
timestamp 1670211287
transform 0 1 0 -1 0 315000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_976
timestamp 1670211287
transform 0 1 0 -1 0 319000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_977
timestamp 1670211287
transform 0 1 0 -1 0 313000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_978
timestamp 1670211287
transform 0 1 0 -1 0 309000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_979
timestamp 1670211287
transform 0 1 0 -1 0 307000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_980
timestamp 1670211287
transform 0 1 0 -1 0 311000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_981
timestamp 1670211287
transform 0 1 0 -1 0 286000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_982
timestamp 1670211287
transform 0 1 0 -1 0 288000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_983
timestamp 1670211287
transform 0 1 0 -1 0 290000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_985
timestamp 1670211287
transform 0 1 0 -1 0 284000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_986
timestamp 1670211287
transform 0 1 0 -1 0 272000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_987
timestamp 1670211287
transform 0 1 0 -1 0 276000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_988
timestamp 1670211287
transform 0 1 0 -1 0 274000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_989
timestamp 1670211287
transform 0 1 0 -1 0 280000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_990
timestamp 1670211287
transform 0 1 0 -1 0 278000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_991
timestamp 1670211287
transform 0 1 0 -1 0 282000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_992
timestamp 1670211287
transform 0 1 0 -1 0 270000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_993
timestamp 1670211287
transform 0 1 0 -1 0 266000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_994
timestamp 1670211287
transform 0 1 0 -1 0 268000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_995
timestamp 1670211287
transform 0 1 0 -1 0 245000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_996
timestamp 1670211287
transform 0 1 0 -1 0 247000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_997
timestamp 1670211287
transform 0 1 0 -1 0 249000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_999
timestamp 1670211287
transform 0 1 0 -1 0 243000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1000
timestamp 1670211287
transform 0 1 0 -1 0 231000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1001
timestamp 1670211287
transform 0 1 0 -1 0 235000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1002
timestamp 1670211287
transform 0 1 0 -1 0 233000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1003
timestamp 1670211287
transform 0 1 0 -1 0 239000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1004
timestamp 1670211287
transform 0 1 0 -1 0 237000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1005
timestamp 1670211287
transform 0 1 0 -1 0 241000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1006
timestamp 1670211287
transform 0 1 0 -1 0 227000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1007
timestamp 1670211287
transform 0 1 0 -1 0 229000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1008
timestamp 1670211287
transform 0 1 0 -1 0 225000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1009
timestamp 1670211287
transform 0 1 0 -1 0 206000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1010
timestamp 1670211287
transform 0 1 0 -1 0 204000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1011
timestamp 1670211287
transform 0 1 0 -1 0 202000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1013
timestamp 1670211287
transform 0 1 0 -1 0 208000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1014
timestamp 1670211287
transform 0 1 0 -1 0 200000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1015
timestamp 1670211287
transform 0 1 0 -1 0 188000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1016
timestamp 1670211287
transform 0 1 0 -1 0 190000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1017
timestamp 1670211287
transform 0 1 0 -1 0 196000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1018
timestamp 1670211287
transform 0 1 0 -1 0 198000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1019
timestamp 1670211287
transform 0 1 0 -1 0 192000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1020
timestamp 1670211287
transform 0 1 0 -1 0 194000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1021
timestamp 1670211287
transform 0 1 0 -1 0 184000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1022
timestamp 1670211287
transform 0 1 0 -1 0 186000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1024
timestamp 1670211287
transform 0 1 0 -1 0 167000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1025
timestamp 1670211287
transform 0 1 0 -1 0 165000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1026
timestamp 1670211287
transform 0 1 0 -1 0 163000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1027
timestamp 1670211287
transform 0 1 0 -1 0 159000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1028
timestamp 1670211287
transform 0 1 0 -1 0 161000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1029
timestamp 1670211287
transform 0 1 0 -1 0 157000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1030
timestamp 1670211287
transform 0 1 0 -1 0 155000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1031
timestamp 1670211287
transform 0 1 0 -1 0 151000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1032
timestamp 1670211287
transform 0 1 0 -1 0 153000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1033
timestamp 1670211287
transform 0 1 0 -1 0 149000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1034
timestamp 1670211287
transform 0 1 0 -1 0 147000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1035
timestamp 1670211287
transform 0 1 0 -1 0 143000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1036
timestamp 1670211287
transform 0 1 0 -1 0 145000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1038
timestamp 1670211287
transform 0 1 0 -1 0 85000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1039
timestamp 1670211287
transform 0 1 0 -1 0 83000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1040
timestamp 1670211287
transform 0 1 0 -1 0 81000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1041
timestamp 1670211287
transform 0 1 0 -1 0 79000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1042
timestamp 1670211287
transform 0 1 0 -1 0 77000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1043
timestamp 1670211287
transform 0 1 0 -1 0 73000
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1044
timestamp 1670211287
transform 0 1 0 -1 0 75000
box -32 13097 2032 69968
use gf180mcu_fd_io__in_c  mgmt_clock_input_pad $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 1 0 215000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__cor  mgmt_corner[0] $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 1 0 0 0 1 0
box 0 0 71000 71000
use gf180mcu_fd_io__cor  mgmt_corner[1]
timestamp 1670211287
transform -1 0 776000 0 1 0
box 0 0 71000 71000
use gf180mcu_fd_io__bi_t  mgmt_gpio_pad
timestamp 1670211287
transform 1 0 545000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  mgmt_vccd_pad $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 0 1 0 -1 0 100000
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  mgmt_vdda_pad
timestamp 1670211287
transform 1 0 655000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  mgmt_vddio_pad_0
timestamp 1670211287
transform 0 1 0 -1 0 141000
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  mgmt_vddio_pad_1
timestamp 1670211287
transform 0 1 0 -1 0 838000
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  mgmt_vssa_pad $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 1 0 105000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  mgmt_vssd_pad
timestamp 1670211287
transform 1 0 270000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  mgmt_vssio_pad_0
timestamp 1670211287
transform 1 0 600000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  mgmt_vssio_pad_1
timestamp 1670211287
transform -1 0 394000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[0]
timestamp 1670211287
transform 0 -1 776000 1 0 89000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[1]
timestamp 1670211287
transform 0 -1 776000 1 0 132000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[2]
timestamp 1670211287
transform 0 -1 776000 1 0 175000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[3]
timestamp 1670211287
transform 0 -1 776000 1 0 218000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[4]
timestamp 1670211287
transform 0 -1 776000 1 0 261000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[5]
timestamp 1670211287
transform 0 -1 776000 1 0 304000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[6]
timestamp 1670211287
transform 0 -1 776000 1 0 347000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[7]
timestamp 1670211287
transform 0 -1 776000 1 0 519000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[8]
timestamp 1670211287
transform 0 -1 776000 1 0 562000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[9]
timestamp 1670211287
transform 0 -1 776000 1 0 605000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[10]
timestamp 1670211287
transform 0 -1 776000 1 0 648000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[11]
timestamp 1670211287
transform 0 -1 776000 1 0 691000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[12]
timestamp 1670211287
transform 0 -1 776000 1 0 734000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[13]
timestamp 1670211287
transform 0 -1 776000 1 0 820000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[14]
timestamp 1670211287
transform 0 -1 776000 1 0 906000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[15]
timestamp 1670211287
transform -1 0 669000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[16]
timestamp 1670211287
transform -1 0 559000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[17]
timestamp 1670211287
transform -1 0 504000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[18]
timestamp 1670211287
transform -1 0 449000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[19]
timestamp 1670211287
transform -1 0 339000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[20]
timestamp 1670211287
transform -1 0 284000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[21]
timestamp 1670211287
transform -1 0 229000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[22]
timestamp 1670211287
transform -1 0 174000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[23]
timestamp 1670211287
transform -1 0 119000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[24]
timestamp 1670211287
transform 0 1 0 -1 0 920000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[25]
timestamp 1670211287
transform 0 1 0 -1 0 756000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[26]
timestamp 1670211287
transform 0 1 0 -1 0 715000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[27]
timestamp 1670211287
transform 0 1 0 -1 0 674000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[28]
timestamp 1670211287
transform 0 1 0 -1 0 633000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[29]
timestamp 1670211287
transform 0 1 0 -1 0 592000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[30]
timestamp 1670211287
transform 0 1 0 -1 0 551000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[31]
timestamp 1670211287
transform 0 1 0 -1 0 510000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[32]
timestamp 1670211287
transform 0 1 0 -1 0 387000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[33]
timestamp 1670211287
transform 0 1 0 -1 0 346000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[34]
timestamp 1670211287
transform 0 1 0 -1 0 305000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[35]
timestamp 1670211287
transform 0 1 0 -1 0 264000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[36]
timestamp 1670211287
transform 0 1 0 -1 0 223000
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  mprj_pads[37]
timestamp 1670211287
transform 0 1 0 -1 0 182000
box -32 0 15032 70000
use gf180mcu_fd_io__in_s  resetb_pad $PDKPATH/libs.ref/gf180mcu_fd_io/mag
timestamp 1670211287
transform 1 0 160000 0 1 0
box -32 0 15032 70000
use gf180mcu_fd_io__cor  user1_corner
timestamp 1670211287
transform -1 0 776000 0 -1 1014000
box 0 0 71000 71000
use gf180mcu_fd_io__dvdd  user1_vccd_pad
timestamp 1670211287
transform 0 -1 776000 1 0 863000
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  user1_vdda_pad_0
timestamp 1670211287
transform 0 -1 776000 1 0 777000
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  user1_vdda_pad_1
timestamp 1670211287
transform 0 -1 776000 1 0 476000
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  user1_vssa_pad_0
timestamp 1670211287
transform -1 0 614000 0 -1 1014000
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  user1_vssa_pad_1
timestamp 1670211287
transform 0 -1 776000 1 0 390000
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  user1_vssd_pad
timestamp 1670211287
transform 0 -1 776000 1 0 433000
box -32 0 15032 70000
use gf180mcu_fd_io__cor  user2_corner
timestamp 1670211287
transform 1 0 0 0 -1 1014000
box 0 0 71000 71000
use gf180mcu_fd_io__dvdd  user2_vccd_pad
timestamp 1670211287
transform 0 1 0 -1 0 879000
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  user2_vdda_pad
timestamp 1670211287
transform 0 1 0 -1 0 469000
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  user2_vssa_pad
timestamp 1670211287
transform 0 1 0 -1 0 797000
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  user2_vssd_pad
timestamp 1670211287
transform 0 1 0 -1 0 428000
box -32 0 15032 70000
<< labels >>
flabel metal5 106500 400 118500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 161500 400 173500 12400 0 FreeSans 24000 0 0 0 resetb
port 446 nsew
flabel metal5 271500 400 283500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 326500 400 338500 12400 0 FreeSans 24000 0 0 0 flash_csb
port 5 nsew
flabel metal5 381500 400 393500 12400 0 FreeSans 24000 0 0 0 flash_clk
port 2 nsew
flabel metal5 436500 400 448500 12400 0 FreeSans 24000 0 0 0 flash_io0
port 8 nsew
flabel metal5 491500 400 503500 12400 0 FreeSans 24000 0 0 0 flash_io1
port 13 nsew
flabel metal5 546500 400 558500 12400 0 FreeSans 24000 0 0 0 gpio
port 18 nsew
flabel metal5 601500 400 613500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 656500 400 668500 12400 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 216500 400 228500 12400 0 FreeSans 24000 0 0 0 clock
port 0 nsew
flabel metal2 174172 69924 174248 70200 0 FreeSans 480 90 0 0 resetb_core
port 447 nsew
flabel metal2 229172 69924 229248 70200 0 FreeSans 480 90 0 0 clock_core
port 1 nsew
flabel metal2 393880 69924 393956 70200 0 FreeSans 480 90 0 0 flash_clk_core
port 3 nsew
flabel metal2 394026 69924 394102 70200 0 FreeSans 480 90 0 0 flash_clk_oe_core
port 4 nsew
flabel metal2 338880 69924 338956 70200 0 FreeSans 480 90 0 0 flash_csb_core
port 6 nsew
flabel metal2 339026 69924 339102 70200 0 FreeSans 480 90 0 0 flash_csb_oe_core
port 7 nsew
flabel metal2 437277 69924 437353 70200 0 FreeSans 480 90 0 0 flash_io0_ie_core
port 11 nsew
flabel metal2 448880 69924 448956 70200 0 FreeSans 480 90 0 0 flash_io0_do_core
port 10 nsew
flabel metal2 449026 69924 449102 70200 0 FreeSans 480 90 0 0 flash_io0_oe_core
port 12 nsew
flabel metal2 449171 69924 449247 70200 0 FreeSans 480 90 0 0 flash_io0_di_core
port 9 nsew
flabel metal2 492277 69924 492353 70200 0 FreeSans 480 90 0 0 flash_io1_ie_core
port 16 nsew
flabel metal2 503880 69924 503956 70200 0 FreeSans 480 90 0 0 flash_io1_do_core
port 15 nsew
flabel metal2 504026 69924 504102 70200 0 FreeSans 480 90 0 0 flash_io1_oe_core
port 17 nsew
flabel metal2 504172 69924 504248 70200 0 FreeSans 480 90 0 0 flash_io1_di_core
port 14 nsew
flabel metal2 545672 69924 545748 70200 0 FreeSans 480 90 0 0 gpio_schmitt_select
port 27 nsew
flabel metal2 546193 69924 546269 70200 0 FreeSans 480 90 0 0 gpio_pu_select
port 26 nsew
flabel metal2 546422 69924 546498 70200 0 FreeSans 480 90 0 0 gpio_drive_select_core[0]
port 19 nsew
flabel metal2 546564 69923 546640 70199 0 FreeSans 480 90 0 0 gpio_drive_select_core[1]
port 20 nsew
flabel metal2 547066 69924 547142 70200 0 FreeSans 480 90 0 0 gpio_pd_select
port 25 nsew
flabel metal2 547277 69924 547353 70200 0 FreeSans 480 90 0 0 gpio_inen_core
port 22 nsew
flabel metal2 558734 69924 558810 70200 0 FreeSans 480 90 0 0 gpio_slew_select
port 28 nsew
flabel metal2 558880 69924 558956 70200 0 FreeSans 480 90 0 0 gpio_out_core
port 23 nsew
flabel metal2 559172 69924 559248 70200 0 FreeSans 480 90 0 0 gpio_in_core
port 21 nsew
flabel metal2 559026 69924 559102 70200 0 FreeSans 480 90 0 0 gpio_outen_core
port 24 nsew
flabel metal5 400 906500 12400 918500 0 FreeSans 24000 0 0 0 mprj_io[24]
port 45 nsew
flabel metal5 400 865500 12400 877500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 824500 12400 836500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 783500 12400 795500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 400 742500 12400 754500 0 FreeSans 24000 0 0 0 mprj_io[25]
port 46 nsew
flabel metal5 400 701500 12400 713500 0 FreeSans 24000 0 0 0 mprj_io[26]
port 47 nsew
flabel metal5 400 660500 12400 672500 0 FreeSans 24000 0 0 0 mprj_io[27]
port 48 nsew
flabel metal5 400 619500 12400 631500 0 FreeSans 24000 0 0 0 mprj_io[28]
port 49 nsew
flabel metal5 400 578500 12400 590500 0 FreeSans 24000 0 0 0 mprj_io[29]
port 50 nsew
flabel metal5 400 537500 12400 549500 0 FreeSans 24000 0 0 0 mprj_io[30]
port 52 nsew
flabel metal5 400 496500 12400 508500 0 FreeSans 24000 0 0 0 mprj_io[31]
port 53 nsew
flabel metal5 400 455500 12400 467500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 414500 12400 426500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 400 373500 12400 385500 0 FreeSans 24000 0 0 0 mprj_io[32]
port 54 nsew
flabel metal5 400 332500 12400 344500 0 FreeSans 24000 0 0 0 mprj_io[33]
port 55 nsew
flabel metal5 400 291500 12400 303500 0 FreeSans 24000 0 0 0 mprj_io[34]
port 56 nsew
flabel metal5 400 250500 12400 262500 0 FreeSans 24000 0 0 0 mprj_io[35]
port 57 nsew
flabel metal5 400 209500 12400 221500 0 FreeSans 24000 0 0 0 mprj_io[36]
port 58 nsew
flabel metal5 400 168500 12400 180500 0 FreeSans 24000 0 0 0 mprj_io[37]
port 59 nsew
flabel metal5 400 127500 12400 139500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 86500 12400 98500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal2 69924 167752 70200 167828 0 FreeSans 480 180 0 0 mprj_io_in[37]
port 172 nsew
flabel metal2 69924 167898 70200 167974 0 FreeSans 480 180 0 0 mprj_io_outen[37]
port 286 nsew
flabel metal2 69924 168044 70200 168120 0 FreeSans 480 180 0 0 mprj_io_out[37]
port 248 nsew
flabel metal2 69924 168190 70200 168266 0 FreeSans 480 180 0 0 mprj_io_slew_select[37]
port 438 nsew
flabel metal2 69924 179647 70200 179723 0 FreeSans 480 180 0 0 mprj_io_inen[37]
port 210 nsew
flabel metal2 69924 179858 70200 179934 0 FreeSans 480 180 0 0 mprj_io_pd_select[37]
port 324 nsew
flabel metal2 69924 180360 70200 180436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[75]
port 138 nsew
flabel metal2 69924 180502 70200 180578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[74]
port 137 nsew
flabel metal2 69924 180731 70200 180807 0 FreeSans 480 180 0 0 mprj_io_pu_select[37]
port 362 nsew
flabel metal2 69924 181252 70200 181328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[37]
port 400 nsew
flabel metal2 69924 208752 70200 208828 0 FreeSans 480 180 0 0 mprj_io_in[36]
port 171 nsew
flabel metal2 69924 208898 70200 208974 0 FreeSans 480 180 0 0 mprj_io_outen[36]
port 285 nsew
flabel metal2 69924 209044 70200 209120 0 FreeSans 480 180 0 0 mprj_io_out[36]
port 247 nsew
flabel metal2 69924 209190 70200 209266 0 FreeSans 480 180 0 0 mprj_io_slew_select[36]
port 437 nsew
flabel metal2 69924 220647 70200 220723 0 FreeSans 480 180 0 0 mprj_io_inen[36]
port 209 nsew
flabel metal2 69924 220858 70200 220934 0 FreeSans 480 180 0 0 mprj_io_pd_select[36]
port 323 nsew
flabel metal2 69924 221360 70200 221436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[73]
port 136 nsew
flabel metal2 69924 221502 70200 221578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[72]
port 135 nsew
flabel metal2 69924 221731 70200 221807 0 FreeSans 480 180 0 0 mprj_io_pu_select[36]
port 361 nsew
flabel metal2 69924 222252 70200 222328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[36]
port 399 nsew
flabel metal2 69924 249752 70200 249828 0 FreeSans 480 180 0 0 mprj_io_in[35]
port 170 nsew
flabel metal2 69924 249898 70200 249974 0 FreeSans 480 180 0 0 mprj_io_outen[35]
port 284 nsew
flabel metal2 69924 250044 70200 250120 0 FreeSans 480 180 0 0 mprj_io_out[35]
port 246 nsew
flabel metal2 69924 250190 70200 250266 0 FreeSans 480 180 0 0 mprj_io_slew_select[35]
port 436 nsew
flabel metal2 69924 261647 70200 261723 0 FreeSans 480 180 0 0 mprj_io_inen[35]
port 208 nsew
flabel metal2 69924 261858 70200 261934 0 FreeSans 480 180 0 0 mprj_io_pd_select[35]
port 322 nsew
flabel metal2 69924 262360 70200 262436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[71]
port 134 nsew
flabel metal2 69924 262502 70200 262578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[70]
port 133 nsew
flabel metal2 69924 262731 70200 262807 0 FreeSans 480 180 0 0 mprj_io_pu_select[35]
port 360 nsew
flabel metal2 69924 263252 70200 263328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[35]
port 398 nsew
flabel metal2 69924 290752 70200 290828 0 FreeSans 480 180 0 0 mprj_io_in[34]
port 169 nsew
flabel metal2 69924 290898 70200 290974 0 FreeSans 480 180 0 0 mprj_io_outen[34]
port 283 nsew
flabel metal2 69924 291044 70200 291120 0 FreeSans 480 180 0 0 mprj_io_out[34]
port 245 nsew
flabel metal2 69924 291190 70200 291266 0 FreeSans 480 180 0 0 mprj_io_slew_select[34]
port 435 nsew
flabel metal2 69924 302647 70200 302723 0 FreeSans 480 180 0 0 mprj_io_inen[34]
port 207 nsew
flabel metal2 69924 302858 70200 302934 0 FreeSans 480 180 0 0 mprj_io_pd_select[34]
port 321 nsew
flabel metal2 69924 303360 70200 303436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[69]
port 131 nsew
flabel metal2 69924 303502 70200 303578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[68]
port 130 nsew
flabel metal2 69924 303731 70200 303807 0 FreeSans 480 180 0 0 mprj_io_pu_select[34]
port 359 nsew
flabel metal2 69924 304252 70200 304328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[34]
port 397 nsew
flabel metal2 69924 331752 70200 331828 0 FreeSans 480 180 0 0 mprj_io_in[33]
port 168 nsew
flabel metal2 69924 331898 70200 331974 0 FreeSans 480 180 0 0 mprj_io_outen[33]
port 282 nsew
flabel metal2 69924 332044 70200 332120 0 FreeSans 480 180 0 0 mprj_io_out[33]
port 244 nsew
flabel metal2 69924 332190 70200 332266 0 FreeSans 480 180 0 0 mprj_io_slew_select[33]
port 434 nsew
flabel metal2 69924 343647 70200 343723 0 FreeSans 480 180 0 0 mprj_io_inen[33]
port 206 nsew
flabel metal2 69924 343858 70200 343934 0 FreeSans 480 180 0 0 mprj_io_pd_select[33]
port 320 nsew
flabel metal2 69924 344360 70200 344436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[67]
port 129 nsew
flabel metal2 69924 344502 70200 344578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[66]
port 128 nsew
flabel metal2 69924 344731 70200 344807 0 FreeSans 480 180 0 0 mprj_io_pu_select[33]
port 358 nsew
flabel metal2 69924 345252 70200 345328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[33]
port 396 nsew
flabel metal2 69924 372752 70200 372828 0 FreeSans 480 180 0 0 mprj_io_in[32]
port 167 nsew
flabel metal2 69924 372898 70200 372974 0 FreeSans 480 180 0 0 mprj_io_outen[32]
port 281 nsew
flabel metal2 69924 373044 70200 373120 0 FreeSans 480 180 0 0 mprj_io_out[32]
port 243 nsew
flabel metal2 69924 373190 70200 373266 0 FreeSans 480 180 0 0 mprj_io_slew_select[32]
port 433 nsew
flabel metal2 69924 384647 70200 384723 0 FreeSans 480 180 0 0 mprj_io_inen[32]
port 205 nsew
flabel metal2 69924 384858 70200 384934 0 FreeSans 480 180 0 0 mprj_io_pd_select[32]
port 319 nsew
flabel metal2 69924 385360 70200 385436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[65]
port 127 nsew
flabel metal2 69924 385502 70200 385578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[64]
port 126 nsew
flabel metal2 69924 385731 70200 385807 0 FreeSans 480 180 0 0 mprj_io_pu_select[32]
port 357 nsew
flabel metal2 69924 386252 70200 386328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[32]
port 395 nsew
flabel metal2 69924 495752 70200 495828 0 FreeSans 480 180 0 0 mprj_io_in[31]
port 166 nsew
flabel metal2 69924 495898 70200 495974 0 FreeSans 480 180 0 0 mprj_io_outen[31]
port 280 nsew
flabel metal2 69924 496044 70200 496120 0 FreeSans 480 180 0 0 mprj_io_out[31]
port 242 nsew
flabel metal2 69924 496190 70200 496266 0 FreeSans 480 180 0 0 mprj_io_slew_select[31]
port 432 nsew
flabel metal2 69924 507647 70200 507723 0 FreeSans 480 180 0 0 mprj_io_inen[31]
port 204 nsew
flabel metal2 69924 507858 70200 507934 0 FreeSans 480 180 0 0 mprj_io_pd_select[31]
port 318 nsew
flabel metal2 69924 508360 70200 508436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[63]
port 125 nsew
flabel metal2 69924 508502 70200 508578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[62]
port 124 nsew
flabel metal2 69924 508731 70200 508807 0 FreeSans 480 180 0 0 mprj_io_pu_select[31]
port 356 nsew
flabel metal2 69924 509252 70200 509328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[31]
port 394 nsew
flabel metal2 69924 536752 70200 536828 0 FreeSans 480 180 0 0 mprj_io_in[30]
port 165 nsew
flabel metal2 69924 536898 70200 536974 0 FreeSans 480 180 0 0 mprj_io_outen[30]
port 279 nsew
flabel metal2 69924 537044 70200 537120 0 FreeSans 480 180 0 0 mprj_io_out[30]
port 241 nsew
flabel metal2 69924 537190 70200 537266 0 FreeSans 480 180 0 0 mprj_io_slew_select[30]
port 431 nsew
flabel metal2 69924 548647 70200 548723 0 FreeSans 480 180 0 0 mprj_io_inen[30]
port 203 nsew
flabel metal2 69924 548858 70200 548934 0 FreeSans 480 180 0 0 mprj_io_pd_select[30]
port 317 nsew
flabel metal2 69924 549731 70200 549807 0 FreeSans 480 180 0 0 mprj_io_pu_select[30]
port 355 nsew
flabel metal2 69924 550252 70200 550328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[30]
port 393 nsew
flabel metal2 69924 577752 70200 577828 0 FreeSans 480 180 0 0 mprj_io_in[29]
port 163 nsew
flabel metal2 69924 577898 70200 577974 0 FreeSans 480 180 0 0 mprj_io_outen[29]
port 277 nsew
flabel metal2 69924 578044 70200 578120 0 FreeSans 480 180 0 0 mprj_io_out[29]
port 239 nsew
flabel metal2 69924 578190 70200 578266 0 FreeSans 480 180 0 0 mprj_io_slew_select[29]
port 429 nsew
flabel metal2 69924 589647 70200 589723 0 FreeSans 480 180 0 0 mprj_io_inen[29]
port 201 nsew
flabel metal2 69924 589858 70200 589934 0 FreeSans 480 180 0 0 mprj_io_pd_select[29]
port 315 nsew
flabel metal2 69924 590360 70200 590436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[59]
port 121 nsew
flabel metal2 69924 590502 70200 590578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[58]
port 120 nsew
flabel metal2 69924 590731 70200 590807 0 FreeSans 480 180 0 0 mprj_io_pu_select[29]
port 353 nsew
flabel metal2 69924 591252 70200 591328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[29]
port 391 nsew
flabel metal2 69924 618752 70200 618828 0 FreeSans 480 180 0 0 mprj_io_in[28]
port 162 nsew
flabel metal2 69924 618898 70200 618974 0 FreeSans 480 180 0 0 mprj_io_outen[28]
port 276 nsew
flabel metal2 69924 619044 70200 619120 0 FreeSans 480 180 0 0 mprj_io_out[28]
port 238 nsew
flabel metal2 69924 619190 70200 619266 0 FreeSans 480 180 0 0 mprj_io_slew_select[28]
port 428 nsew
flabel metal2 69924 630647 70200 630723 0 FreeSans 480 180 0 0 mprj_io_inen[28]
port 200 nsew
flabel metal2 69924 630858 70200 630934 0 FreeSans 480 180 0 0 mprj_io_pd_select[28]
port 314 nsew
flabel metal2 69924 631360 70200 631436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[57]
port 119 nsew
flabel metal2 69924 631502 70200 631578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[56]
port 118 nsew
flabel metal2 69924 631731 70200 631807 0 FreeSans 480 180 0 0 mprj_io_pu_select[28]
port 352 nsew
flabel metal2 69924 632252 70200 632328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[28]
port 390 nsew
flabel metal2 69924 659752 70200 659828 0 FreeSans 480 180 0 0 mprj_io_in[27]
port 161 nsew
flabel metal2 69924 659898 70200 659974 0 FreeSans 480 180 0 0 mprj_io_outen[27]
port 275 nsew
flabel metal2 69924 660044 70200 660120 0 FreeSans 480 180 0 0 mprj_io_out[27]
port 237 nsew
flabel metal2 69924 660190 70200 660266 0 FreeSans 480 180 0 0 mprj_io_slew_select[27]
port 427 nsew
flabel metal2 69924 671647 70200 671723 0 FreeSans 480 180 0 0 mprj_io_inen[27]
port 199 nsew
flabel metal2 69924 671858 70200 671934 0 FreeSans 480 180 0 0 mprj_io_pd_select[27]
port 313 nsew
flabel metal2 69924 672360 70200 672436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[55]
port 117 nsew
flabel metal2 69924 672502 70200 672578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[54]
port 116 nsew
flabel metal2 69924 672731 70200 672807 0 FreeSans 480 180 0 0 mprj_io_pu_select[27]
port 351 nsew
flabel metal2 69924 673252 70200 673328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[27]
port 389 nsew
flabel metal2 69924 700752 70200 700828 0 FreeSans 480 180 0 0 mprj_io_in[26]
port 160 nsew
flabel metal2 69924 700898 70200 700974 0 FreeSans 480 180 0 0 mprj_io_outen[26]
port 274 nsew
flabel metal2 69924 701044 70200 701120 0 FreeSans 480 180 0 0 mprj_io_out[26]
port 236 nsew
flabel metal2 69924 701190 70200 701266 0 FreeSans 480 180 0 0 mprj_io_slew_select[26]
port 426 nsew
flabel metal2 69924 712647 70200 712723 0 FreeSans 480 180 0 0 mprj_io_inen[26]
port 198 nsew
flabel metal2 69924 712858 70200 712934 0 FreeSans 480 180 0 0 mprj_io_pd_select[26]
port 312 nsew
flabel metal2 69924 713360 70200 713436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[53]
port 115 nsew
flabel metal2 69924 713502 70200 713578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[52]
port 114 nsew
flabel metal2 69924 713731 70200 713807 0 FreeSans 480 180 0 0 mprj_io_pu_select[26]
port 350 nsew
flabel metal2 69924 714252 70200 714328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[26]
port 388 nsew
flabel metal2 69924 741752 70200 741828 0 FreeSans 480 180 0 0 mprj_io_in[25]
port 159 nsew
flabel metal2 69924 741898 70200 741974 0 FreeSans 480 180 0 0 mprj_io_outen[25]
port 273 nsew
flabel metal2 69924 742044 70200 742120 0 FreeSans 480 180 0 0 mprj_io_out[25]
port 235 nsew
flabel metal2 69924 742190 70200 742266 0 FreeSans 480 180 0 0 mprj_io_slew_select[25]
port 425 nsew
flabel metal2 69924 753647 70200 753723 0 FreeSans 480 180 0 0 mprj_io_inen[25]
port 197 nsew
flabel metal2 69924 753858 70200 753934 0 FreeSans 480 180 0 0 mprj_io_pd_select[25]
port 311 nsew
flabel metal2 69924 754360 70200 754436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[51]
port 112 nsew
flabel metal2 69924 754731 70200 754807 0 FreeSans 480 180 0 0 mprj_io_pu_select[25]
port 349 nsew
flabel metal2 69924 755252 70200 755328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[25]
port 387 nsew
flabel metal2 69924 905752 70200 905828 0 FreeSans 480 180 0 0 mprj_io_in[24]
port 158 nsew
flabel metal2 69924 905898 70200 905974 0 FreeSans 480 180 0 0 mprj_io_outen[24]
port 272 nsew
flabel metal2 69924 906044 70200 906120 0 FreeSans 480 180 0 0 mprj_io_out[24]
port 234 nsew
flabel metal2 69924 906190 70200 906266 0 FreeSans 480 180 0 0 mprj_io_slew_select[24]
port 424 nsew
flabel metal2 69924 917647 70200 917723 0 FreeSans 480 180 0 0 mprj_io_inen[24]
port 196 nsew
flabel metal2 69924 917858 70200 917934 0 FreeSans 480 180 0 0 mprj_io_pd_select[24]
port 310 nsew
flabel metal2 69924 918360 70200 918436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[49]
port 110 nsew
flabel metal2 69924 918502 70200 918578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[48]
port 109 nsew
flabel metal2 69924 918731 70200 918807 0 FreeSans 480 180 0 0 mprj_io_pu_select[24]
port 348 nsew
flabel metal2 69924 919252 70200 919328 0 FreeSans 480 180 0 0 mprj_io_schmitt_select[24]
port 386 nsew
flabel metal5 763600 90500 775600 102500 0 FreeSans 24000 0 0 0 mprj_io[0]
port 29 nsew
flabel metal5 763600 133500 775600 145500 0 FreeSans 24000 0 0 0 mprj_io[1]
port 40 nsew
flabel metal5 763600 176500 775600 188500 0 FreeSans 24000 0 0 0 mprj_io[2]
port 51 nsew
flabel metal5 763600 219500 775600 231500 0 FreeSans 24000 0 0 0 mprj_io[3]
port 60 nsew
flabel metal5 763600 262500 775600 274500 0 FreeSans 24000 0 0 0 mprj_io[4]
port 61 nsew
flabel metal5 763600 305500 775600 317500 0 FreeSans 24000 0 0 0 mprj_io[5]
port 62 nsew
flabel metal5 763600 348500 775600 360500 0 FreeSans 24000 0 0 0 mprj_io[6]
port 63 nsew
flabel metal5 763600 391500 775600 403500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 763600 434500 775600 446500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 763600 477500 775600 489500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 763600 520500 775600 532500 0 FreeSans 24000 0 0 0 mprj_io[7]
port 64 nsew
flabel metal5 763600 563500 775600 575500 0 FreeSans 24000 0 0 0 mprj_io[8]
port 65 nsew
flabel metal5 763600 606500 775600 618500 0 FreeSans 24000 0 0 0 mprj_io[9]
port 66 nsew
flabel metal5 763600 649500 775600 661500 0 FreeSans 24000 0 0 0 mprj_io[10]
port 30 nsew
flabel metal5 763600 692500 775600 704500 0 FreeSans 24000 0 0 0 mprj_io[11]
port 31 nsew
flabel metal5 763600 735500 775600 747500 0 FreeSans 24000 0 0 0 mprj_io[12]
port 32 nsew
flabel metal5 763600 778500 775600 790500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 763600 821500 775600 833500 0 FreeSans 24000 0 0 0 mprj_io[13]
port 33 nsew
flabel metal5 763600 864500 775600 876500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 763600 907500 775600 919500 0 FreeSans 24000 0 0 0 mprj_io[14]
port 34 nsew
flabel metal5 655500 1001600 667500 1013600 0 FreeSans 24000 0 0 0 mprj_io[15]
port 35 nsew
flabel metal5 600500 1001600 612500 1013600 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 545500 1001600 557500 1013600 0 FreeSans 24000 0 0 0 mprj_io[16]
port 36 nsew
flabel metal5 490500 1001600 502500 1013600 0 FreeSans 24000 0 0 0 mprj_io[17]
port 37 nsew
flabel metal5 435500 1001600 447500 1013600 0 FreeSans 24000 0 0 0 mprj_io[18]
port 38 nsew
flabel metal5 380500 1001600 392500 1013600 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 325500 1001600 337500 1013600 0 FreeSans 24000 0 0 0 mprj_io[19]
port 39 nsew
flabel metal5 270500 1001600 282500 1013600 0 FreeSans 24000 0 0 0 mprj_io[20]
port 41 nsew
flabel metal5 215500 1001600 227500 1013600 0 FreeSans 24000 0 0 0 mprj_io[21]
port 42 nsew
flabel metal5 160500 1001600 172500 1013600 0 FreeSans 24000 0 0 0 mprj_io[22]
port 43 nsew
flabel metal5 105500 1001600 117500 1013600 0 FreeSans 24000 0 0 0 mprj_io[23]
port 44 nsew
flabel metal2 705800 89672 706076 89748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[0]
port 370 nsew
flabel metal2 705800 90193 706076 90269 0 FreeSans 480 0 0 0 mprj_io_pu_select[0]
port 332 nsew
flabel metal2 705800 90422 706076 90498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[0]
port 67 nsew
flabel metal2 705800 90564 706076 90640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[1]
port 78 nsew
flabel metal2 705800 91066 706076 91142 0 FreeSans 480 0 0 0 mprj_io_pd_select[0]
port 294 nsew
flabel metal2 705800 91277 706076 91353 0 FreeSans 480 0 0 0 mprj_io_inen[0]
port 180 nsew
flabel metal2 705800 102734 706076 102810 0 FreeSans 480 0 0 0 mprj_io_slew_select[0]
port 408 nsew
flabel metal2 705800 102880 706076 102956 0 FreeSans 480 0 0 0 mprj_io_out[0]
port 218 nsew
flabel metal2 705800 103026 706076 103102 0 FreeSans 480 0 0 0 mprj_io_outen[0]
port 256 nsew
flabel metal2 705800 103172 706076 103248 0 FreeSans 480 0 0 0 mprj_io_in[0]
port 142 nsew
flabel metal2 705621 132672 705897 132748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[1]
port 381 nsew
flabel metal2 705621 133193 705897 133269 0 FreeSans 480 0 0 0 mprj_io_pu_select[1]
port 343 nsew
flabel metal2 705621 133422 705897 133498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[2]
port 89 nsew
flabel metal2 705621 133564 705897 133640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[3]
port 100 nsew
flabel metal2 705621 134066 705897 134142 0 FreeSans 480 0 0 0 mprj_io_pd_select[1]
port 305 nsew
flabel metal2 705621 134277 705897 134353 0 FreeSans 480 0 0 0 mprj_io_inen[1]
port 191 nsew
flabel metal2 705621 145734 705897 145810 0 FreeSans 480 0 0 0 mprj_io_slew_select[1]
port 419 nsew
flabel metal2 705621 145880 705897 145956 0 FreeSans 480 0 0 0 mprj_io_out[1]
port 229 nsew
flabel metal2 705621 146026 705897 146102 0 FreeSans 480 0 0 0 mprj_io_outen[1]
port 267 nsew
flabel metal2 705621 146172 705897 146248 0 FreeSans 480 0 0 0 mprj_io_in[1]
port 153 nsew
flabel metal2 705800 189172 706076 189248 0 FreeSans 480 0 0 0 mprj_io_in[2]
port 164 nsew
flabel metal2 705800 189026 706076 189102 0 FreeSans 480 0 0 0 mprj_io_outen[2]
port 278 nsew
flabel metal2 705800 188880 706076 188956 0 FreeSans 480 0 0 0 mprj_io_out[2]
port 240 nsew
flabel metal2 705800 188734 706076 188810 0 FreeSans 480 0 0 0 mprj_io_slew_select[2]
port 430 nsew
flabel metal2 705800 177277 706076 177353 0 FreeSans 480 0 0 0 mprj_io_inen[2]
port 202 nsew
flabel metal2 705800 177066 706076 177142 0 FreeSans 480 0 0 0 mprj_io_pd_select[2]
port 316 nsew
flabel metal2 705800 176193 706076 176269 0 FreeSans 480 0 0 0 mprj_io_pu_select[2]
port 354 nsew
flabel metal2 705800 175672 706076 175748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[2]
port 392 nsew
flabel metal2 705800 232172 706076 232248 0 FreeSans 480 0 0 0 mprj_io_in[3]
port 173 nsew
flabel metal2 705800 232026 706076 232102 0 FreeSans 480 0 0 0 mprj_io_outen[3]
port 287 nsew
flabel metal2 705800 231880 706076 231956 0 FreeSans 480 0 0 0 mprj_io_out[3]
port 249 nsew
flabel metal2 705800 231734 706076 231810 0 FreeSans 480 0 0 0 mprj_io_slew_select[3]
port 439 nsew
flabel metal2 705800 220277 706076 220353 0 FreeSans 480 0 0 0 mprj_io_inen[3]
port 211 nsew
flabel metal2 705800 220066 706076 220142 0 FreeSans 480 0 0 0 mprj_io_pd_select[3]
port 325 nsew
flabel metal2 705800 219193 706076 219269 0 FreeSans 480 0 0 0 mprj_io_pu_select[3]
port 363 nsew
flabel metal2 705800 218672 706076 218748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[3]
port 401 nsew
flabel metal2 705800 275172 706076 275248 0 FreeSans 480 0 0 0 mprj_io_in[4]
port 174 nsew
flabel metal2 705800 275026 706076 275102 0 FreeSans 480 0 0 0 mprj_io_outen[4]
port 288 nsew
flabel metal2 705800 274880 706076 274956 0 FreeSans 480 0 0 0 mprj_io_out[4]
port 250 nsew
flabel metal2 705800 274734 706076 274810 0 FreeSans 480 0 0 0 mprj_io_slew_select[4]
port 440 nsew
flabel metal2 705800 263277 706076 263353 0 FreeSans 480 0 0 0 mprj_io_inen[4]
port 212 nsew
flabel metal2 705800 263066 706076 263142 0 FreeSans 480 0 0 0 mprj_io_pd_select[4]
port 326 nsew
flabel metal2 705800 262193 706076 262269 0 FreeSans 480 0 0 0 mprj_io_pu_select[4]
port 364 nsew
flabel metal2 705800 261672 706076 261748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[4]
port 402 nsew
flabel metal2 705800 318172 706076 318248 0 FreeSans 480 0 0 0 mprj_io_in[5]
port 175 nsew
flabel metal2 705800 318026 706076 318102 0 FreeSans 480 0 0 0 mprj_io_outen[5]
port 289 nsew
flabel metal2 705800 317880 706076 317956 0 FreeSans 480 0 0 0 mprj_io_out[5]
port 251 nsew
flabel metal2 705800 317734 706076 317810 0 FreeSans 480 0 0 0 mprj_io_slew_select[5]
port 441 nsew
flabel metal2 705800 306277 706076 306353 0 FreeSans 480 0 0 0 mprj_io_inen[5]
port 213 nsew
flabel metal2 705800 306066 706076 306142 0 FreeSans 480 0 0 0 mprj_io_pd_select[5]
port 327 nsew
flabel metal2 705800 305193 706076 305269 0 FreeSans 480 0 0 0 mprj_io_pu_select[5]
port 365 nsew
flabel metal2 705800 304672 706076 304748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[5]
port 403 nsew
flabel metal2 705800 361172 706076 361248 0 FreeSans 480 0 0 0 mprj_io_in[6]
port 176 nsew
flabel metal2 705800 361026 706076 361102 0 FreeSans 480 0 0 0 mprj_io_outen[6]
port 290 nsew
flabel metal2 705800 360880 706076 360956 0 FreeSans 480 0 0 0 mprj_io_out[6]
port 252 nsew
flabel metal2 705800 360734 706076 360810 0 FreeSans 480 0 0 0 mprj_io_slew_select[6]
port 442 nsew
flabel metal2 705800 349277 706076 349353 0 FreeSans 480 0 0 0 mprj_io_inen[6]
port 214 nsew
flabel metal2 705800 349066 706076 349142 0 FreeSans 480 0 0 0 mprj_io_pd_select[6]
port 328 nsew
flabel metal2 705800 348193 706076 348269 0 FreeSans 480 0 0 0 mprj_io_pu_select[6]
port 366 nsew
flabel metal2 705800 347672 706076 347748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[6]
port 404 nsew
flabel metal2 705800 533172 706076 533248 0 FreeSans 480 0 0 0 mprj_io_in[7]
port 177 nsew
flabel metal2 705800 533026 706076 533102 0 FreeSans 480 0 0 0 mprj_io_outen[7]
port 291 nsew
flabel metal2 705800 532880 706076 532956 0 FreeSans 480 0 0 0 mprj_io_out[7]
port 253 nsew
flabel metal2 705800 532734 706076 532810 0 FreeSans 480 0 0 0 mprj_io_slew_select[7]
port 443 nsew
flabel metal2 705800 521277 706076 521353 0 FreeSans 480 0 0 0 mprj_io_inen[7]
port 215 nsew
flabel metal2 705800 521066 706076 521142 0 FreeSans 480 0 0 0 mprj_io_pd_select[7]
port 329 nsew
flabel metal2 705800 520193 706076 520269 0 FreeSans 480 0 0 0 mprj_io_pu_select[7]
port 367 nsew
flabel metal2 705800 519672 706076 519748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[7]
port 405 nsew
flabel metal2 705800 576172 706076 576248 0 FreeSans 480 0 0 0 mprj_io_in[8]
port 178 nsew
flabel metal2 705800 576026 706076 576102 0 FreeSans 480 0 0 0 mprj_io_outen[8]
port 292 nsew
flabel metal2 705800 575880 706076 575956 0 FreeSans 480 0 0 0 mprj_io_out[8]
port 254 nsew
flabel metal2 705800 575734 706076 575810 0 FreeSans 480 0 0 0 mprj_io_slew_select[8]
port 444 nsew
flabel metal2 705800 564277 706076 564353 0 FreeSans 480 0 0 0 mprj_io_inen[8]
port 216 nsew
flabel metal2 705800 564066 706076 564142 0 FreeSans 480 0 0 0 mprj_io_pd_select[8]
port 330 nsew
flabel metal2 705800 563193 706076 563269 0 FreeSans 480 0 0 0 mprj_io_pu_select[8]
port 368 nsew
flabel metal2 705800 562672 706076 562748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[8]
port 406 nsew
flabel metal2 705800 619172 706076 619248 0 FreeSans 480 0 0 0 mprj_io_in[9]
port 179 nsew
flabel metal2 705800 619026 706076 619102 0 FreeSans 480 0 0 0 mprj_io_outen[9]
port 293 nsew
flabel metal2 705800 618880 706076 618956 0 FreeSans 480 0 0 0 mprj_io_out[9]
port 255 nsew
flabel metal2 705800 618734 706076 618810 0 FreeSans 480 0 0 0 mprj_io_slew_select[9]
port 445 nsew
flabel metal2 705800 607277 706076 607353 0 FreeSans 480 0 0 0 mprj_io_inen[9]
port 217 nsew
flabel metal2 705800 607066 706076 607142 0 FreeSans 480 0 0 0 mprj_io_pd_select[9]
port 331 nsew
flabel metal2 705800 606193 706076 606269 0 FreeSans 480 0 0 0 mprj_io_pu_select[9]
port 369 nsew
flabel metal2 705800 605672 706076 605748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[9]
port 407 nsew
flabel metal2 705800 662172 706076 662248 0 FreeSans 480 0 0 0 mprj_io_in[10]
port 143 nsew
flabel metal2 705800 662026 706076 662102 0 FreeSans 480 0 0 0 mprj_io_outen[10]
port 257 nsew
flabel metal2 705800 661880 706076 661956 0 FreeSans 480 0 0 0 mprj_io_out[10]
port 219 nsew
flabel metal2 705800 661734 706076 661810 0 FreeSans 480 0 0 0 mprj_io_slew_select[10]
port 409 nsew
flabel metal2 705800 650277 706076 650353 0 FreeSans 480 0 0 0 mprj_io_inen[10]
port 181 nsew
flabel metal2 705800 650066 706076 650142 0 FreeSans 480 0 0 0 mprj_io_pd_select[10]
port 295 nsew
flabel metal2 705800 649193 706076 649269 0 FreeSans 480 0 0 0 mprj_io_pu_select[10]
port 333 nsew
flabel metal2 705800 648672 706076 648748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[10]
port 371 nsew
flabel metal2 705800 705172 706076 705248 0 FreeSans 480 0 0 0 mprj_io_in[11]
port 144 nsew
flabel metal2 705800 705026 706076 705102 0 FreeSans 480 0 0 0 mprj_io_outen[11]
port 258 nsew
flabel metal2 705800 704880 706076 704956 0 FreeSans 480 0 0 0 mprj_io_out[11]
port 220 nsew
flabel metal2 705800 704734 706076 704810 0 FreeSans 480 0 0 0 mprj_io_slew_select[11]
port 410 nsew
flabel metal2 705800 693277 706076 693353 0 FreeSans 480 0 0 0 mprj_io_inen[11]
port 182 nsew
flabel metal2 705800 693066 706076 693142 0 FreeSans 480 0 0 0 mprj_io_pd_select[11]
port 296 nsew
flabel metal2 705800 692193 706076 692269 0 FreeSans 480 0 0 0 mprj_io_pu_select[11]
port 334 nsew
flabel metal2 705800 691672 706076 691748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[11]
port 372 nsew
flabel metal2 705800 906672 706076 906748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[14]
port 375 nsew
flabel metal2 705800 907193 706076 907269 0 FreeSans 480 0 0 0 mprj_io_pu_select[14]
port 337 nsew
flabel metal2 705800 907422 706076 907498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[28]
port 87 nsew
flabel metal2 705800 907564 706076 907640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[29]
port 88 nsew
flabel metal2 705800 908066 706076 908142 0 FreeSans 480 0 0 0 mprj_io_pd_select[14]
port 299 nsew
flabel metal2 705800 908277 706076 908353 0 FreeSans 480 0 0 0 mprj_io_inen[14]
port 185 nsew
flabel metal2 705800 919734 706076 919810 0 FreeSans 480 0 0 0 mprj_io_slew_select[14]
port 413 nsew
flabel metal2 705800 919880 706076 919956 0 FreeSans 480 0 0 0 mprj_io_out[14]
port 223 nsew
flabel metal2 705800 920026 706076 920102 0 FreeSans 480 0 0 0 mprj_io_outen[14]
port 261 nsew
flabel metal2 705800 920172 706076 920248 0 FreeSans 480 0 0 0 mprj_io_in[14]
port 147 nsew
flabel metal2 668252 943800 668328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[15]
port 376 nsew
flabel metal2 667731 943800 667807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[15]
port 338 nsew
flabel metal2 667502 943800 667578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[30]
port 90 nsew
flabel metal2 667360 943800 667436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[31]
port 91 nsew
flabel metal2 666858 943800 666934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[15]
port 300 nsew
flabel metal2 666647 943800 666723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[15]
port 186 nsew
flabel metal2 655190 943800 655266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[15]
port 414 nsew
flabel metal2 655044 943800 655120 944076 0 FreeSans 480 270 0 0 mprj_io_out[15]
port 224 nsew
flabel metal2 654898 943800 654974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[15]
port 262 nsew
flabel metal2 654752 943800 654828 944076 0 FreeSans 480 270 0 0 mprj_io_in[15]
port 148 nsew
flabel metal2 558252 943800 558328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[16]
port 377 nsew
flabel metal2 557731 943800 557807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[16]
port 339 nsew
flabel metal2 557502 943800 557578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[32]
port 92 nsew
flabel metal2 557360 943800 557436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[33]
port 93 nsew
flabel metal2 556858 943800 556934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[16]
port 301 nsew
flabel metal2 556647 943800 556723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[16]
port 187 nsew
flabel metal2 545190 943800 545266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[16]
port 415 nsew
flabel metal2 545044 943800 545120 944076 0 FreeSans 480 270 0 0 mprj_io_out[16]
port 225 nsew
flabel metal2 544898 943800 544974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[16]
port 263 nsew
flabel metal2 544752 943800 544828 944076 0 FreeSans 480 270 0 0 mprj_io_in[16]
port 149 nsew
flabel metal2 503252 943800 503328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[17]
port 378 nsew
flabel metal2 502731 943800 502807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[17]
port 340 nsew
flabel metal2 502502 943800 502578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[34]
port 94 nsew
flabel metal2 502360 943800 502436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[35]
port 95 nsew
flabel metal2 501858 943800 501934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[17]
port 302 nsew
flabel metal2 501647 943800 501723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[17]
port 188 nsew
flabel metal2 490190 943800 490266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[17]
port 416 nsew
flabel metal2 490044 943800 490120 944076 0 FreeSans 480 270 0 0 mprj_io_out[17]
port 226 nsew
flabel metal2 489898 943800 489974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[17]
port 264 nsew
flabel metal2 489752 943800 489828 944076 0 FreeSans 480 270 0 0 mprj_io_in[17]
port 150 nsew
flabel metal2 448252 943800 448328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[18]
port 379 nsew
flabel metal2 447731 943800 447807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[18]
port 341 nsew
flabel metal2 447502 943800 447578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[36]
port 96 nsew
flabel metal2 447360 943800 447436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[37]
port 97 nsew
flabel metal2 446858 943800 446934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[18]
port 303 nsew
flabel metal2 446647 943800 446723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[18]
port 189 nsew
flabel metal2 435190 943800 435266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[18]
port 417 nsew
flabel metal2 435044 943800 435120 944076 0 FreeSans 480 270 0 0 mprj_io_out[18]
port 227 nsew
flabel metal2 434898 943800 434974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[18]
port 265 nsew
flabel metal2 434752 943800 434828 944076 0 FreeSans 480 270 0 0 mprj_io_in[18]
port 151 nsew
flabel metal2 338252 943800 338328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[19]
port 380 nsew
flabel metal2 337731 943800 337807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[19]
port 342 nsew
flabel metal2 337502 943800 337578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[38]
port 98 nsew
flabel metal2 337360 943800 337436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[39]
port 99 nsew
flabel metal2 336858 943800 336934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[19]
port 304 nsew
flabel metal2 336647 943800 336723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[19]
port 190 nsew
flabel metal2 325190 943800 325266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[19]
port 418 nsew
flabel metal2 325044 943800 325120 944076 0 FreeSans 480 270 0 0 mprj_io_out[19]
port 228 nsew
flabel metal2 324898 943800 324974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[19]
port 266 nsew
flabel metal2 324752 943800 324828 944076 0 FreeSans 480 270 0 0 mprj_io_in[19]
port 152 nsew
flabel metal2 283252 943800 283328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[20]
port 382 nsew
flabel metal2 282731 943800 282807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[20]
port 344 nsew
flabel metal2 282502 943800 282578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[40]
port 101 nsew
flabel metal2 282360 943800 282436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[41]
port 102 nsew
flabel metal2 281858 943800 281934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[20]
port 306 nsew
flabel metal2 281647 943800 281723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[20]
port 192 nsew
flabel metal2 270190 943800 270266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[20]
port 420 nsew
flabel metal2 270044 943800 270120 944076 0 FreeSans 480 270 0 0 mprj_io_out[20]
port 230 nsew
flabel metal2 269898 943800 269974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[20]
port 268 nsew
flabel metal2 269752 943800 269828 944076 0 FreeSans 480 270 0 0 mprj_io_in[20]
port 154 nsew
flabel metal2 228252 943800 228328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[21]
port 383 nsew
flabel metal2 227731 943800 227807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[21]
port 345 nsew
flabel metal2 227502 943800 227578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[42]
port 103 nsew
flabel metal2 227360 943800 227436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[43]
port 104 nsew
flabel metal2 226858 943800 226934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[21]
port 307 nsew
flabel metal2 226647 943800 226723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[21]
port 193 nsew
flabel metal2 215190 943800 215266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[21]
port 421 nsew
flabel metal2 215044 943800 215120 944076 0 FreeSans 480 270 0 0 mprj_io_out[21]
port 231 nsew
flabel metal2 214898 943800 214974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[21]
port 269 nsew
flabel metal2 214752 943800 214828 944076 0 FreeSans 480 270 0 0 mprj_io_in[21]
port 155 nsew
flabel metal2 173252 943800 173328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[22]
port 384 nsew
flabel metal2 172731 943800 172807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[22]
port 346 nsew
flabel metal2 172502 943800 172578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[44]
port 105 nsew
flabel metal2 172360 943800 172436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[45]
port 106 nsew
flabel metal2 171858 943800 171934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[22]
port 308 nsew
flabel metal2 171647 943800 171723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[22]
port 194 nsew
flabel metal2 160190 943800 160266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[22]
port 422 nsew
flabel metal2 160044 943800 160120 944076 0 FreeSans 480 270 0 0 mprj_io_out[22]
port 232 nsew
flabel metal2 159898 943800 159974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[22]
port 270 nsew
flabel metal2 159752 943800 159828 944076 0 FreeSans 480 270 0 0 mprj_io_in[22]
port 156 nsew
flabel metal2 118252 943800 118328 944076 0 FreeSans 480 270 0 0 mprj_io_schmitt_select[23]
port 385 nsew
flabel metal2 117731 943800 117807 944076 0 FreeSans 480 270 0 0 mprj_io_pu_select[23]
port 347 nsew
flabel metal2 117502 943800 117578 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[46]
port 107 nsew
flabel metal2 117360 943800 117436 944076 0 FreeSans 480 270 0 0 mprj_io_drive_sel[47]
port 108 nsew
flabel metal2 116858 943800 116934 944076 0 FreeSans 480 270 0 0 mprj_io_pd_select[23]
port 309 nsew
flabel metal2 116647 943800 116723 944076 0 FreeSans 480 270 0 0 mprj_io_inen[23]
port 195 nsew
flabel metal2 105190 943800 105266 944076 0 FreeSans 480 270 0 0 mprj_io_slew_select[23]
port 423 nsew
flabel metal2 105044 943800 105120 944076 0 FreeSans 480 270 0 0 mprj_io_out[23]
port 233 nsew
flabel metal2 104898 943800 104974 944076 0 FreeSans 480 270 0 0 mprj_io_outen[23]
port 271 nsew
flabel metal2 104752 943800 104828 944076 0 FreeSans 480 270 0 0 mprj_io_in[23]
port 157 nsew
flabel metal2 162066 70000 162142 70225 0 FreeSans 480 90 0 0 const_zero[5]
port 451 nsew
flabel metal2 216193 70000 216269 70199 0 FreeSans 480 90 0 0 const_zero[4]
port 452 nsew
flabel metal2 338733 69924 338810 70202 0 FreeSans 480 90 0 0 const_zero[3]
port 453 nsew
flabel metal2 393734 69924 393810 70198 0 FreeSans 480 90 0 0 const_zero[2]
port 454 nsew
flabel metal2 448734 69924 448810 70198 0 FreeSans 480 90 0 0 const_zero[1]
port 455 nsew
flabel metal2 503734 69924 503810 70198 0 FreeSans 480 90 0 0 const_zero[0]
port 456 nsew
flabel metal2 326193 69924 326269 70156 0 FreeSans 480 90 0 0 const_one[1]
port 457 nsew
flabel metal2 161193 70000 161269 70225 0 FreeSans 480 90 0 0 const_one[0]
port 450 nsew
flabel metal2 705800 748172 706076 748248 0 FreeSans 480 0 0 0 mprj_io_in[12]
port 145 nsew
flabel metal2 705800 748026 706076 748102 0 FreeSans 480 0 0 0 mprj_io_outen[12]
port 259 nsew
flabel metal2 705800 747880 706076 747956 0 FreeSans 480 0 0 0 mprj_io_out[12]
port 221 nsew
flabel metal2 705800 747734 706076 747810 0 FreeSans 480 0 0 0 mprj_io_slew_select[12]
port 411 nsew
flabel metal2 705800 736277 706076 736353 0 FreeSans 480 0 0 0 mprj_io_inen[12]
port 183 nsew
flabel metal2 705800 736066 706076 736142 0 FreeSans 480 0 0 0 mprj_io_pd_select[12]
port 297 nsew
flabel metal2 705800 735193 706076 735269 0 FreeSans 480 0 0 0 mprj_io_pu_select[12]
port 335 nsew
flabel metal2 705800 734672 706076 734748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[12]
port 373 nsew
flabel metal2 705800 834172 706076 834248 0 FreeSans 480 0 0 0 mprj_io_in[13]
port 146 nsew
flabel metal2 705800 834026 706076 834102 0 FreeSans 480 0 0 0 mprj_io_outen[13]
port 260 nsew
flabel metal2 705800 833880 706076 833956 0 FreeSans 480 0 0 0 mprj_io_out[13]
port 222 nsew
flabel metal2 705800 833734 706076 833810 0 FreeSans 480 0 0 0 mprj_io_slew_select[13]
port 412 nsew
flabel metal2 705800 822277 706076 822353 0 FreeSans 480 0 0 0 mprj_io_inen[13]
port 184 nsew
flabel metal2 705800 822066 706076 822142 0 FreeSans 480 0 0 0 mprj_io_pd_select[13]
port 298 nsew
flabel metal2 705800 821564 706076 821640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[27]
port 86 nsew
flabel metal2 705800 821422 706076 821498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[26]
port 85 nsew
flabel metal2 705800 821193 706076 821269 0 FreeSans 480 0 0 0 mprj_io_pu_select[13]
port 336 nsew
flabel metal2 705800 820672 706076 820748 0 FreeSans 480 0 0 0 mprj_io_schmitt_select[13]
port 374 nsew
flabel metal2 705800 176422 706076 176498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[4]
port 111 nsew
flabel metal2 705800 176564 706076 176640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[5]
port 122 nsew
flabel metal2 705800 219422 706076 219498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[6]
port 132 nsew
flabel metal2 705800 219564 706076 219640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[7]
port 139 nsew
flabel metal2 705800 262422 706076 262498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[8]
port 140 nsew
flabel metal2 705800 262564 706076 262640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[9]
port 141 nsew
flabel metal2 705800 305422 706076 305498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[10]
port 68 nsew
flabel metal2 705800 305564 706076 305640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[11]
port 69 nsew
flabel metal2 705800 348422 706076 348498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[12]
port 70 nsew
flabel metal2 705800 348564 706076 348640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[13]
port 71 nsew
flabel metal2 705800 520422 706076 520498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[14]
port 72 nsew
flabel metal2 705800 520564 706076 520640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[15]
port 73 nsew
flabel metal2 705800 563422 706076 563498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[16]
port 74 nsew
flabel metal2 705800 563564 706076 563640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[17]
port 75 nsew
flabel metal2 705800 606422 706076 606498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[18]
port 76 nsew
flabel metal2 705800 606564 706076 606640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[19]
port 77 nsew
flabel metal2 705800 649422 706076 649498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[20]
port 79 nsew
flabel metal2 705800 649564 706076 649640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[21]
port 80 nsew
flabel metal2 705800 692422 706076 692498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[22]
port 81 nsew
flabel metal2 705800 692564 706076 692640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[23]
port 82 nsew
flabel metal2 705800 735422 706076 735498 0 FreeSans 480 0 0 0 mprj_io_drive_sel[24]
port 83 nsew
flabel metal2 705800 735564 706076 735640 0 FreeSans 480 0 0 0 mprj_io_drive_sel[25]
port 84 nsew
flabel metal2 69924 754502 70200 754578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[50]
port 113 nsew
flabel metal2 69924 549360 70200 549436 0 FreeSans 480 180 0 0 mprj_io_drive_sel[61]
port 123 nsew
flabel metal2 69924 549502 70200 549578 0 FreeSans 480 180 0 0 mprj_io_drive_sel[60]
port 458 nsew
<< end >>
