magic
tech gf180mcuC
magscale 6 5
timestamp 1654634570
<< metal5 >>
rect 0 648 324 756
rect 216 0 324 648
<< properties >>
string FIXED_BBOX 0 0 432 756
<< end >>
