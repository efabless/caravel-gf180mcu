magic
tech gf180mcuD
magscale 1 10
timestamp 1670447154
<< metal4 >>
rect 94 93 10733 373
<< metal5 >>
rect 6066 10173 6300 10266
tri 5460 10080 5553 10173 se
rect 5553 10080 6300 10173
tri 5366 9893 5460 9986 se
rect 5460 9893 6300 10080
tri 4593 9800 4686 9893 se
rect 4686 9800 5693 9893
rect 4593 9753 5693 9800
tri 4500 9613 4593 9706 se
rect 4593 9660 5600 9753
tri 5600 9660 5693 9753 nw
rect 4593 9613 4806 9660
tri 4806 9613 4853 9660 nw
rect 4200 9473 4806 9613
rect 6066 9566 6300 9893
rect 6066 9520 7280 9566
rect 4200 9380 4713 9473
tri 4713 9380 4806 9473 nw
tri 5693 9426 5786 9520 se
rect 5786 9426 7280 9520
tri 5180 9380 5226 9426 se
rect 5226 9380 7280 9426
tri 4760 8960 5180 9380 se
rect 5180 9333 7280 9380
rect 5180 9053 7093 9333
tri 7093 9240 7186 9333 nw
rect 5180 8960 7000 9053
tri 7000 8960 7093 9053 nw
tri 4666 8586 4760 8680 se
rect 4760 8586 7000 8960
rect 4666 8400 7000 8586
tri 7000 8400 7093 8493 sw
rect 2706 7746 2940 8213
rect 4666 8026 7093 8400
tri 4666 7933 4760 8026 ne
rect 4760 7933 7093 8026
tri 7093 7933 7280 8120 sw
rect 4760 7840 5693 7933
tri 5693 7840 5786 7933 nw
rect 6066 7840 7280 7933
rect 4760 7746 5315 7840
rect 2426 7466 3173 7746
tri 2426 7373 2520 7466 ne
rect 2520 7186 3080 7466
tri 3080 7373 3173 7466 nw
tri 4760 7404 5102 7746 ne
rect 5102 7404 5315 7746
tri 5315 7695 5460 7840 nw
rect 6066 7326 6346 7840
tri 6813 7653 7000 7840 ne
rect 7000 7653 7280 7840
tri 9893 7746 10173 8026 se
rect 10173 7746 10386 8026
tri 9800 7653 9893 7746 se
tri 9613 7466 9800 7653 se
rect 9800 7466 9893 7653
tri 9473 7326 9613 7466 se
rect 9613 7326 9893 7466
tri 9893 7373 10266 7746 nw
rect 6066 7280 7933 7326
tri 5693 7186 5786 7280 se
rect 5786 7186 7933 7280
rect 2706 6953 2940 7186
rect 4946 7093 7933 7186
tri 9240 7093 9473 7326 se
rect 9473 7280 9893 7326
rect 9473 7093 9800 7280
tri 9800 7186 9893 7280 nw
tri 4900 6954 4946 7000 se
rect 4946 6954 7466 7093
rect 2706 6906 3733 6953
tri 4853 6906 4900 6953 se
rect 4900 6906 7466 6954
tri 7466 6906 7653 7093 nw
tri 9147 7000 9240 7093 se
rect 9240 7000 9800 7093
tri 1960 6813 2053 6906 se
rect 2053 6813 3733 6906
rect 1400 6720 3733 6813
tri 4574 6720 4760 6906 se
rect 4760 6720 7466 6906
tri 933 6160 1400 6626 se
rect 1400 6253 3360 6720
tri 3360 6626 3453 6720 nw
tri 4480 6626 4574 6720 se
rect 4574 6626 7186 6720
rect 1400 6160 3266 6253
tri 3266 6160 3360 6253 nw
tri 4013 6160 4480 6626 se
rect 4480 6160 7186 6626
tri 7186 6440 7466 6720 nw
rect 8446 6673 8680 7000
tri 8960 6813 9147 7000 se
rect 9147 6813 9706 7000
tri 9706 6906 9800 7000 nw
tri 8913 6673 8960 6720 se
rect 8960 6673 9706 6813
rect 8446 6533 9706 6673
tri 840 5786 933 5880 se
rect 933 5786 3266 6160
rect 840 5413 3266 5786
tri 3640 5693 4013 6066 se
rect 4013 5693 7093 6160
tri 7093 6066 7186 6160 nw
tri 8353 6160 8446 6253 se
rect 8446 6160 9613 6533
tri 9613 6440 9706 6533 nw
tri 8306 6066 8353 6113 se
rect 8353 6066 9613 6160
tri 3266 5413 3360 5506 sw
rect 840 4946 3360 5413
tri 840 4853 933 4946 ne
rect 933 4573 3360 4946
tri 933 4433 1073 4573 ne
rect 1073 4480 3360 4573
tri 3593 5273 3640 5320 se
rect 3640 5273 7093 5693
rect 3593 4573 7093 5273
tri 7746 5413 8306 5973 se
rect 8306 5413 9520 6066
tri 9520 5973 9613 6066 nw
tri 7560 5040 7746 5226 se
rect 7746 5040 9520 5413
tri 7420 4853 7560 4993 se
rect 7560 4853 9520 5040
tri 7326 4573 7420 4666 se
rect 7420 4573 9520 4853
rect 3593 4480 9520 4573
tri 9520 4480 9613 4573 sw
rect 1073 4433 2053 4480
rect 187 4386 467 4433
tri 467 4386 514 4433 sw
tri 1073 4386 1120 4433 ne
rect 1120 4386 2053 4433
tri 2053 4386 2146 4480 nw
tri 2426 4386 2520 4480 ne
rect 2520 4386 9613 4480
rect 187 4293 560 4386
tri 560 4293 654 4386 sw
tri 1120 4293 1213 4386 ne
rect 1213 4293 1773 4386
rect 187 4200 747 4293
tri 374 4080 494 4200 ne
rect 494 4106 747 4200
tri 747 4106 933 4293 sw
rect 1306 4106 1773 4293
tri 1773 4200 1960 4386 nw
rect 2706 4293 9613 4386
rect 494 4080 1026 4106
tri 587 3893 774 4080 ne
rect 774 4060 1026 4080
tri 1026 4060 1073 4106 sw
rect 1306 4060 1726 4106
tri 1726 4060 1773 4106 nw
rect 774 3893 1726 4060
tri 866 3826 933 3893 ne
rect 933 3826 1726 3893
tri 1026 3733 1120 3826 ne
rect 1120 3733 2280 3826
tri 1213 3640 1306 3733 ne
rect 1306 3640 2280 3733
tri 2280 3640 2466 3826 sw
rect 2706 3640 2986 4293
tri 3226 4200 3320 4293 ne
rect 3320 4200 9613 4293
tri 3360 4013 3546 4200 ne
rect 3546 4013 9613 4200
rect 1306 3453 2986 3640
rect 3546 3920 7840 4013
tri 7840 3920 7933 4013 nw
rect 3546 3826 7560 3920
tri 7560 3826 7653 3920 nw
tri 3546 3453 3920 3826 ne
rect 3920 3480 7560 3826
tri 7560 3480 7746 3666 sw
rect 3920 3453 7746 3480
rect 1493 3360 2986 3453
tri 2986 3360 3080 3453 sw
rect 3920 3360 5600 3453
tri 5600 3360 5693 3453 nw
tri 5973 3360 6066 3453 ne
rect 6066 3360 7746 3453
tri 1493 3266 1586 3360 ne
rect 1586 3266 3266 3360
tri 3266 3266 3360 3360 sw
tri 1773 2706 2333 3266 ne
rect 2333 2520 3640 3266
rect 3920 3173 4853 3360
tri 4853 3266 4946 3360 nw
tri 3920 2893 4200 3173 ne
rect 4200 2893 4573 3173
tri 4573 2893 4853 3173 nw
rect 6160 3173 7746 3360
tri 3640 2520 4013 2893 sw
tri 4200 2800 4293 2893 ne
rect 4293 2520 4573 2893
tri 2240 2333 2333 2426 se
rect 2333 2333 4573 2520
rect 2240 2240 4573 2333
tri 4573 2240 4853 2520 sw
rect 2240 2146 5040 2240
tri 5040 2146 5133 2240 sw
rect 2240 2053 5413 2146
tri 5413 2053 5506 2146 sw
rect 6160 2053 6533 3173
tri 6813 3080 6906 3173 ne
rect 6906 3080 7746 3173
tri 7746 3080 8026 3360 sw
tri 7280 2893 7466 3080 ne
rect 7466 2986 8026 3080
rect 8400 2986 8680 4013
tri 8960 3920 9053 4013 ne
rect 9053 3920 9613 4013
tri 9613 3920 9800 4106 sw
tri 9213 3546 9586 3920 ne
rect 9586 3546 9800 3920
tri 9146 3080 9333 3266 se
rect 9333 3173 10173 3266
tri 10173 3173 10266 3266 sw
rect 9333 3080 10266 3173
tri 8960 2986 9053 3080 se
rect 9053 2986 10266 3080
rect 7466 2940 10266 2986
rect 7466 2893 10173 2940
tri 7746 2706 7933 2893 ne
rect 7933 2706 10173 2893
rect 7933 2473 10733 2706
rect 7933 2426 10266 2473
tri 7280 2053 7653 2426 se
rect 7653 2333 10266 2426
rect 7653 2053 10173 2333
tri 10173 2240 10266 2333 nw
rect 2240 1866 10173 2053
rect 2240 1773 4806 1866
tri 2240 1680 2333 1773 ne
rect 2333 1586 4806 1773
rect 5040 1773 10173 1866
rect 5040 1586 5366 1773
rect 2333 1493 5366 1586
rect 5600 1680 9986 1773
tri 9986 1680 10080 1773 nw
rect 5600 1493 5973 1680
rect 2333 1400 5973 1493
rect 6206 1400 6533 1680
rect 6766 1400 7093 1680
rect 7326 1400 9986 1680
rect 2333 1306 9986 1400
tri 2333 1213 2426 1306 ne
rect 2426 1026 9893 1306
tri 9893 1213 9986 1306 nw
tri 2426 933 2520 1026 ne
rect 2520 840 9613 1026
tri 2520 560 2800 840 ne
rect 2800 466 9613 840
tri 9613 746 9893 1026 nw
tri 2800 373 2893 466 ne
rect 2893 373 9613 466
<< fillblock >>
rect 0 0 10840 10373
<< end >>
