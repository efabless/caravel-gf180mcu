magic
tech gf180mcuD
magscale 1 10
timestamp 1655309791
<< nwell >>
rect 7000 607 7056 1270
<< metal1 >>
rect 374 2361 25324 2408
rect 374 2152 24613 2361
rect 24853 2152 25324 2361
rect 374 2108 25324 2152
rect 374 1478 17790 2108
rect 409 680 556 1478
rect 1397 1313 1443 1478
rect 1825 1309 1871 1478
rect 2258 1311 2304 1478
rect 2686 1311 2732 1478
rect 3064 923 3218 1478
rect 4908 1310 4954 1478
rect 5336 1311 5382 1478
rect 5764 1310 5810 1478
rect 6192 1310 6238 1478
rect 6358 933 6509 1478
rect 7361 704 7508 1478
rect 15845 888 17277 948
rect 7186 460 7580 473
rect 393 -357 505 381
rect 871 -357 1008 221
rect 1018 -357 1248 381
rect 3238 217 3468 381
rect 1607 -357 1653 -173
rect 2095 -357 2141 -176
rect 2583 -357 2629 -171
rect 3071 -357 3117 -171
rect 3238 -357 3601 217
rect 3977 -357 6761 381
rect 7186 287 7201 460
rect 7363 287 7580 460
rect 7186 273 7580 287
rect 15845 -357 15911 888
rect 351 -431 15911 -357
rect 17191 -357 17277 888
rect 17191 -431 25373 -357
rect 351 -657 25373 -431
rect 562 -825 758 -657
rect 837 -836 1320 -773
rect 1397 -836 1880 -773
rect 1957 -836 2440 -773
rect 2517 -779 3000 -773
rect 2517 -831 2643 -779
rect 2882 -831 3000 -779
rect 2517 -836 3000 -831
rect 3077 -836 3560 -773
rect 3637 -836 4120 -773
rect 4197 -836 4680 -773
rect 4757 -836 5240 -773
rect 5317 -836 5800 -773
rect 5877 -836 6360 -773
rect 6437 -836 6920 -773
rect 6997 -836 7480 -773
rect 7557 -836 8040 -773
rect 8117 -836 8600 -773
rect 8677 -836 9160 -773
rect 9237 -836 9720 -773
rect 9797 -836 10280 -773
rect 10357 -836 10840 -773
rect 10917 -836 11400 -773
rect 11477 -836 11960 -773
rect 12037 -836 12520 -773
rect 12597 -836 13080 -773
rect 13157 -836 13640 -773
rect 13717 -836 14200 -773
rect 14277 -836 14760 -773
rect 14837 -836 15320 -773
rect 15397 -836 15880 -773
rect 15957 -836 16440 -773
rect 16517 -836 17000 -773
rect 17077 -836 17560 -773
rect 17637 -836 18120 -773
rect 18197 -836 18680 -773
rect 18757 -836 19240 -773
rect 19317 -836 19800 -773
rect 19877 -836 20360 -773
rect 20437 -836 20920 -773
rect 20997 -836 21480 -773
rect 21557 -836 22040 -773
rect 22117 -836 22600 -773
rect 22677 -836 23160 -773
rect 23237 -836 23720 -773
rect 23797 -836 24280 -773
rect 24357 -836 24840 -773
rect 24917 -778 25124 -772
rect 24917 -830 24935 -778
rect 25100 -830 25124 -778
rect 24917 -833 25124 -830
rect 555 -6001 1038 -5938
rect 1115 -6001 1598 -5938
rect 1675 -6001 2158 -5938
rect 2235 -6001 2718 -5938
rect 2795 -6001 3278 -5938
rect 3355 -6001 3838 -5938
rect 3915 -6001 4398 -5938
rect 4475 -6001 4958 -5938
rect 5035 -6001 5518 -5938
rect 5595 -6001 6078 -5938
rect 6155 -6001 6638 -5938
rect 6715 -6001 7198 -5938
rect 7275 -6001 7758 -5938
rect 7835 -6001 8318 -5938
rect 8395 -6001 8878 -5938
rect 8955 -6001 9438 -5938
rect 9515 -6001 9998 -5938
rect 10075 -6001 10558 -5938
rect 10635 -6001 11118 -5938
rect 11195 -6001 11678 -5938
rect 11755 -6001 12238 -5938
rect 12315 -6001 12798 -5938
rect 12875 -6001 13358 -5938
rect 13435 -6001 13918 -5938
rect 13995 -6001 14478 -5938
rect 14555 -6001 15038 -5938
rect 15115 -6001 15598 -5938
rect 15675 -6001 16158 -5938
rect 16235 -6001 16718 -5938
rect 16795 -6001 17278 -5938
rect 17355 -6001 17838 -5938
rect 17915 -6001 18398 -5938
rect 18475 -6001 18958 -5938
rect 19035 -6001 19518 -5938
rect 19595 -6001 20078 -5938
rect 20155 -6001 20638 -5938
rect 20715 -6001 21198 -5938
rect 21275 -6001 21758 -5938
rect 21835 -6001 22318 -5938
rect 22395 -6001 22878 -5938
rect 22955 -6001 23438 -5938
rect 23515 -6001 23998 -5938
rect 24075 -6001 24558 -5938
rect 24635 -6001 25118 -5938
<< via1 >>
rect 24613 2152 24853 2361
rect 7201 287 7363 460
rect 15911 -431 17191 888
rect 2643 -831 2882 -779
rect 24935 -830 25100 -778
<< metal2 >>
rect 24594 2361 24869 2392
rect 24594 2152 24613 2361
rect 24853 2152 24869 2361
rect 24594 2127 24869 2152
rect 654 749 711 1267
rect 921 1004 2919 1206
rect 3432 1017 3716 1217
rect 1037 869 1093 1004
rect 804 749 860 849
rect 1037 813 3380 869
rect 3785 749 3841 825
rect 654 693 3841 749
rect 654 562 711 693
rect 3926 622 3982 1275
rect 607 505 711 562
rect 3296 566 3982 622
rect 4145 862 4203 1264
rect 4433 1027 5997 1208
rect 4145 806 4270 862
rect 4541 861 4602 1027
rect 6726 1023 7022 1218
rect 4145 739 4203 806
rect 4541 803 6672 861
rect 7091 739 7149 853
rect 4145 681 7149 739
rect 607 119 664 505
rect 3296 290 3352 566
rect 4145 507 4203 681
rect 3858 449 4203 507
rect 7220 473 7278 1272
rect 15845 888 17277 948
rect 7186 460 7633 473
rect 1437 222 3796 290
rect 3296 107 3352 222
rect 1393 -83 3352 107
rect 1393 -86 3341 -83
rect 3858 -195 3916 449
rect 7186 287 7201 460
rect 7363 287 7633 460
rect 7186 273 7633 287
rect 724 -510 787 -234
rect 15845 -431 15911 888
rect 17191 -431 17277 888
rect 24641 -202 24800 2127
rect 24641 -361 25100 -202
rect 15845 -500 17277 -431
rect 724 -573 2781 -510
rect 2718 -773 2781 -573
rect 24941 -772 25100 -361
rect 2624 -779 2903 -773
rect 2624 -831 2643 -779
rect 2882 -831 2903 -779
rect 2624 -835 2903 -831
rect 24916 -778 25123 -772
rect 24916 -830 24935 -778
rect 25100 -830 25123 -778
rect 24916 -834 25123 -830
<< via2 >>
rect 15911 -431 17191 888
<< metal3 >>
rect 15845 888 17277 948
rect 15845 -431 15911 888
rect 17191 -431 17277 888
rect 15845 -500 17277 -431
<< via3 >>
rect 15996 -431 17191 888
<< metal4 >>
rect 15955 888 17277 948
rect 15955 -431 15996 888
rect 17191 -431 17277 888
rect 15955 -500 17277 -431
use nmos_6p0_B4TB5U  XM0 primitives
timestamp 1655304105
transform 1 0 754 0 1 -4
box -334 -432 334 432
use pmos_6p0_CYEQN4  XM1 primitives
timestamp 1655304105
transform 1 0 3815 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM3
timestamp 1655304105
transform 1 0 806 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM4
timestamp 1655304105
transform 1 0 3313 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM7
timestamp 1655304105
transform 1 0 6605 0 1 1093
box -368 -486 378 486
use pmos_6p0_CYEQN4  XM9
timestamp 1655304105
transform 1 0 4317 0 1 1093
box -368 -486 378 486
use nmos_6p0_BJPB5U  nmos_6p0_BJPB5U_0 primitives
timestamp 1655307388
transform 1 0 3722 0 1 -4
box -334 -432 334 432
use nmos_6p0_BJXXPT  nmos_6p0_BJXXPT_0 primitives
timestamp 1655304105
transform 1 0 2242 0 1 8
box -1066 -432 1066 432
use pmos_6p0_CYEQN4  pmos_6p0_CYEQN4_0
timestamp 1655304105
transform 1 0 7107 0 1 1093
box -368 -486 378 486
use pmos_6p0_EYEQQM  pmos_6p0_EYEQQM_0 primitives
timestamp 1655304105
transform 1 0 5501 0 1 1093
box -1050 -486 980 486
use pmos_6p0_HUEQQM  pmos_6p0_HUEQQM_0 primitives
timestamp 1655304105
transform 1 0 2068 0 1 1093
box -1128 -486 1121 486
use ppolyf_u_1k_6p0_TRTT7C  ppolyf_u_1k_6p0_TRTT7C_0 primitives
timestamp 1655304105
transform 1 0 12839 0 1 -3388
box -12578 -2920 12578 2920
use via_cont_0p6um  via_cont_0p6um_0 primitives
timestamp 1655304105
transform 1 0 724 0 1 -55
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_1
timestamp 1655304105
transform 1 0 1483 0 1 432
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_2
timestamp 1655304105
transform 1 0 1730 0 1 434
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_3
timestamp 1655304105
transform 1 0 1974 0 1 436
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_4
timestamp 1655304105
transform 1 0 2221 0 1 439
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_5
timestamp 1655304105
transform 1 0 2455 0 1 438
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_6
timestamp 1655304105
transform 1 0 2717 0 1 439
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_7
timestamp 1655304105
transform 1 0 2952 0 1 437
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_8
timestamp 1655304105
transform 1 0 3698 0 1 423
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_9
timestamp 1655304105
transform 1 0 814 0 1 1030
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_10
timestamp 1655304105
transform 1 0 1270 0 1 1026
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_11
timestamp 1655304105
transform 1 0 1486 0 1 1025
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_12
timestamp 1655304105
transform 1 0 1696 0 1 1025
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_13
timestamp 1655304105
transform 1 0 1910 0 1 1028
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_14
timestamp 1655304105
transform 1 0 2136 0 1 1027
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_15
timestamp 1655304105
transform 1 0 2348 0 1 1028
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_16
timestamp 1655304105
transform 1 0 2561 0 1 1031
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_17
timestamp 1655304105
transform 1 0 2778 0 1 1030
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_18
timestamp 1655304105
transform 1 0 3283 0 1 1029
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_19
timestamp 1655304105
transform 1 0 3768 0 1 1025
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_20
timestamp 1655304105
transform 1 0 4799 0 1 1022
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_21
timestamp 1655304105
transform 1 0 5016 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_22
timestamp 1655304105
transform 1 0 5229 0 1 1017
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_23
timestamp 1655304105
transform 1 0 5437 0 1 1022
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_24
timestamp 1655304105
transform 1 0 5654 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_25
timestamp 1655304105
transform 1 0 5865 0 1 1022
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_26
timestamp 1655304105
transform 1 0 6083 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_27
timestamp 1655304105
transform 1 0 6572 0 1 1019
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_28
timestamp 1655304105
transform 1 0 4291 0 1 1020
box -43 -214 99 -158
use via_cont_0p6um  via_cont_0p6um_29
timestamp 1655304105
transform 1 0 7063 0 1 1032
box -43 -214 99 -158
use via_cont_2um  via_cont_2um_0 primitives
timestamp 1655304105
transform 1 0 696 0 1 -46
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_1
timestamp 1655304105
transform 1 0 1450 0 1 -78
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_2
timestamp 1655304105
transform 1 0 1938 0 1 -82
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_3
timestamp 1655304105
transform 1 0 2423 0 1 -75
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_4
timestamp 1655304105
transform 1 0 2916 0 1 -77
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_5
timestamp 1655304105
transform 1 0 766 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_6
timestamp 1655304105
transform 1 0 972 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_7
timestamp 1655304105
transform 1 0 1263 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_8
timestamp 1655304105
transform 1 0 1698 0 1 1034
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_9
timestamp 1655304105
transform 1 0 2127 0 1 1036
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_10
timestamp 1655304105
transform 1 0 2563 0 1 1041
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_11
timestamp 1655304105
transform 1 0 2987 0 1 1033
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_12
timestamp 1655304105
transform 1 0 3904 0 1 -110
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_13
timestamp 1655304105
transform 1 0 4273 0 1 1029
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_14
timestamp 1655304105
transform 1 0 3493 0 1 1041
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_15
timestamp 1655304105
transform 1 0 3774 0 1 1038
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_16
timestamp 1655304105
transform 1 0 4016 0 1 1044
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_17
timestamp 1655304105
transform 1 0 4780 0 1 1032
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_18
timestamp 1655304105
transform 1 0 5211 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_19
timestamp 1655304105
transform 1 0 5637 0 1 1035
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_20
timestamp 1655304105
transform 1 0 6064 0 1 1040
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_21
timestamp 1655304105
transform 1 0 7070 0 1 1038
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_22
timestamp 1655304105
transform 1 0 6784 0 1 1058
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_23
timestamp 1655304105
transform 1 0 4499 0 1 1030
box -92 -99 -36 240
use via_cont_2um  via_cont_2um_24
timestamp 1655304105
transform 1 0 7288 0 1 1038
box -92 -99 -36 240
<< labels >>
flabel metal1 404 -608 604 -408 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 412 1527 612 1727 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 7380 273 7580 473 0 FreeSans 1280 0 0 0 Vout
port 2 nsew
<< end >>
