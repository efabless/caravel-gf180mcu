magic
tech gf180mcuC
magscale 1 5
timestamp 1655473187
<< obsm1 >>
rect 93 1538 29979 74941
<< metal2 >>
rect 84 74600 140 75000
rect 308 74600 364 75000
rect 532 74600 588 75000
rect 756 74600 812 75000
rect 1036 74600 1092 75000
rect 1260 74600 1316 75000
rect 1484 74600 1540 75000
rect 1764 74600 1820 75000
rect 1988 74600 2044 75000
rect 2212 74600 2268 75000
rect 2436 74600 2492 75000
rect 2716 74600 2772 75000
rect 2940 74600 2996 75000
rect 3164 74600 3220 75000
rect 3444 74600 3500 75000
rect 3668 74600 3724 75000
rect 3892 74600 3948 75000
rect 4116 74600 4172 75000
rect 4396 74600 4452 75000
rect 4620 74600 4676 75000
rect 4844 74600 4900 75000
rect 5124 74600 5180 75000
rect 5348 74600 5404 75000
rect 5572 74600 5628 75000
rect 5796 74600 5852 75000
rect 6076 74600 6132 75000
rect 6300 74600 6356 75000
rect 6524 74600 6580 75000
rect 6804 74600 6860 75000
rect 7028 74600 7084 75000
rect 7252 74600 7308 75000
rect 7476 74600 7532 75000
rect 7756 74600 7812 75000
rect 7980 74600 8036 75000
rect 8204 74600 8260 75000
rect 8484 74600 8540 75000
rect 8708 74600 8764 75000
rect 8932 74600 8988 75000
rect 9156 74600 9212 75000
rect 9436 74600 9492 75000
rect 9660 74600 9716 75000
rect 9884 74600 9940 75000
rect 10164 74600 10220 75000
rect 10388 74600 10444 75000
rect 10612 74600 10668 75000
rect 10836 74600 10892 75000
rect 11116 74600 11172 75000
rect 11340 74600 11396 75000
rect 11564 74600 11620 75000
rect 11844 74600 11900 75000
rect 12068 74600 12124 75000
rect 12292 74600 12348 75000
rect 12516 74600 12572 75000
rect 12796 74600 12852 75000
rect 13020 74600 13076 75000
rect 13244 74600 13300 75000
rect 13524 74600 13580 75000
rect 13748 74600 13804 75000
rect 13972 74600 14028 75000
rect 14196 74600 14252 75000
rect 14476 74600 14532 75000
rect 14700 74600 14756 75000
rect 14924 74600 14980 75000
rect 15204 74600 15260 75000
rect 15428 74600 15484 75000
rect 15652 74600 15708 75000
rect 15932 74600 15988 75000
rect 16156 74600 16212 75000
rect 16380 74600 16436 75000
rect 16604 74600 16660 75000
rect 16884 74600 16940 75000
rect 17108 74600 17164 75000
rect 17332 74600 17388 75000
rect 17612 74600 17668 75000
rect 17836 74600 17892 75000
rect 18060 74600 18116 75000
rect 18284 74600 18340 75000
rect 18564 74600 18620 75000
rect 18788 74600 18844 75000
rect 19012 74600 19068 75000
rect 19292 74600 19348 75000
rect 19516 74600 19572 75000
rect 19740 74600 19796 75000
rect 19964 74600 20020 75000
rect 20244 74600 20300 75000
rect 20468 74600 20524 75000
rect 20692 74600 20748 75000
rect 20972 74600 21028 75000
rect 21196 74600 21252 75000
rect 21420 74600 21476 75000
rect 21644 74600 21700 75000
rect 21924 74600 21980 75000
rect 22148 74600 22204 75000
rect 22372 74600 22428 75000
rect 22652 74600 22708 75000
rect 22876 74600 22932 75000
rect 23100 74600 23156 75000
rect 23324 74600 23380 75000
rect 23604 74600 23660 75000
rect 23828 74600 23884 75000
rect 24052 74600 24108 75000
rect 24332 74600 24388 75000
rect 24556 74600 24612 75000
rect 24780 74600 24836 75000
rect 25004 74600 25060 75000
rect 25284 74600 25340 75000
rect 25508 74600 25564 75000
rect 25732 74600 25788 75000
rect 26012 74600 26068 75000
rect 26236 74600 26292 75000
rect 26460 74600 26516 75000
rect 26684 74600 26740 75000
rect 26964 74600 27020 75000
rect 27188 74600 27244 75000
rect 27412 74600 27468 75000
rect 27692 74600 27748 75000
rect 27916 74600 27972 75000
rect 28140 74600 28196 75000
rect 28364 74600 28420 75000
rect 28644 74600 28700 75000
rect 28868 74600 28924 75000
rect 29092 74600 29148 75000
rect 29372 74600 29428 75000
rect 29596 74600 29652 75000
rect 29820 74600 29876 75000
rect 140 0 196 400
rect 476 0 532 400
rect 812 0 868 400
rect 1148 0 1204 400
rect 1484 0 1540 400
rect 1820 0 1876 400
rect 2156 0 2212 400
rect 2492 0 2548 400
rect 2828 0 2884 400
rect 3164 0 3220 400
rect 3500 0 3556 400
rect 3836 0 3892 400
rect 4172 0 4228 400
rect 4508 0 4564 400
rect 4844 0 4900 400
rect 5180 0 5236 400
rect 5516 0 5572 400
rect 5852 0 5908 400
rect 6188 0 6244 400
rect 6524 0 6580 400
rect 6860 0 6916 400
rect 7196 0 7252 400
rect 7532 0 7588 400
rect 7868 0 7924 400
rect 8204 0 8260 400
rect 8540 0 8596 400
rect 8876 0 8932 400
rect 9212 0 9268 400
rect 9548 0 9604 400
rect 9884 0 9940 400
rect 10220 0 10276 400
rect 10556 0 10612 400
rect 10892 0 10948 400
rect 11228 0 11284 400
rect 11564 0 11620 400
rect 11900 0 11956 400
rect 12236 0 12292 400
rect 12572 0 12628 400
rect 12908 0 12964 400
rect 13244 0 13300 400
rect 13580 0 13636 400
rect 13916 0 13972 400
rect 14252 0 14308 400
rect 14588 0 14644 400
rect 14924 0 14980 400
rect 15316 0 15372 400
rect 15652 0 15708 400
rect 15988 0 16044 400
rect 16324 0 16380 400
rect 16660 0 16716 400
rect 16996 0 17052 400
rect 17332 0 17388 400
rect 17668 0 17724 400
rect 18004 0 18060 400
rect 18340 0 18396 400
rect 18676 0 18732 400
rect 19012 0 19068 400
rect 19348 0 19404 400
rect 19684 0 19740 400
rect 20020 0 20076 400
rect 20356 0 20412 400
rect 20692 0 20748 400
rect 21028 0 21084 400
rect 21364 0 21420 400
rect 21700 0 21756 400
rect 22036 0 22092 400
rect 22372 0 22428 400
rect 22708 0 22764 400
rect 23044 0 23100 400
rect 23380 0 23436 400
rect 23716 0 23772 400
rect 24052 0 24108 400
rect 24388 0 24444 400
rect 24724 0 24780 400
rect 25060 0 25116 400
rect 25396 0 25452 400
rect 25732 0 25788 400
rect 26068 0 26124 400
rect 26404 0 26460 400
rect 26740 0 26796 400
rect 27076 0 27132 400
rect 27412 0 27468 400
rect 27748 0 27804 400
rect 28084 0 28140 400
rect 28420 0 28476 400
rect 28756 0 28812 400
rect 29092 0 29148 400
rect 29428 0 29484 400
rect 29764 0 29820 400
<< obsm2 >>
rect 42 74570 54 74947
rect 170 74570 278 74947
rect 394 74570 502 74947
rect 618 74570 726 74947
rect 842 74570 1006 74947
rect 1122 74570 1230 74947
rect 1346 74570 1454 74947
rect 1570 74570 1734 74947
rect 1850 74570 1958 74947
rect 2074 74570 2182 74947
rect 2298 74570 2406 74947
rect 2522 74570 2686 74947
rect 2802 74570 2910 74947
rect 3026 74570 3134 74947
rect 3250 74570 3414 74947
rect 3530 74570 3638 74947
rect 3754 74570 3862 74947
rect 3978 74570 4086 74947
rect 4202 74570 4366 74947
rect 4482 74570 4590 74947
rect 4706 74570 4814 74947
rect 4930 74570 5094 74947
rect 5210 74570 5318 74947
rect 5434 74570 5542 74947
rect 5658 74570 5766 74947
rect 5882 74570 6046 74947
rect 6162 74570 6270 74947
rect 6386 74570 6494 74947
rect 6610 74570 6774 74947
rect 6890 74570 6998 74947
rect 7114 74570 7222 74947
rect 7338 74570 7446 74947
rect 7562 74570 7726 74947
rect 7842 74570 7950 74947
rect 8066 74570 8174 74947
rect 8290 74570 8454 74947
rect 8570 74570 8678 74947
rect 8794 74570 8902 74947
rect 9018 74570 9126 74947
rect 9242 74570 9406 74947
rect 9522 74570 9630 74947
rect 9746 74570 9854 74947
rect 9970 74570 10134 74947
rect 10250 74570 10358 74947
rect 10474 74570 10582 74947
rect 10698 74570 10806 74947
rect 10922 74570 11086 74947
rect 11202 74570 11310 74947
rect 11426 74570 11534 74947
rect 11650 74570 11814 74947
rect 11930 74570 12038 74947
rect 12154 74570 12262 74947
rect 12378 74570 12486 74947
rect 12602 74570 12766 74947
rect 12882 74570 12990 74947
rect 13106 74570 13214 74947
rect 13330 74570 13494 74947
rect 13610 74570 13718 74947
rect 13834 74570 13942 74947
rect 14058 74570 14166 74947
rect 14282 74570 14446 74947
rect 14562 74570 14670 74947
rect 14786 74570 14894 74947
rect 15010 74570 15174 74947
rect 15290 74570 15398 74947
rect 15514 74570 15622 74947
rect 15738 74570 15902 74947
rect 16018 74570 16126 74947
rect 16242 74570 16350 74947
rect 16466 74570 16574 74947
rect 16690 74570 16854 74947
rect 16970 74570 17078 74947
rect 17194 74570 17302 74947
rect 17418 74570 17582 74947
rect 17698 74570 17806 74947
rect 17922 74570 18030 74947
rect 18146 74570 18254 74947
rect 18370 74570 18534 74947
rect 18650 74570 18758 74947
rect 18874 74570 18982 74947
rect 19098 74570 19262 74947
rect 19378 74570 19486 74947
rect 19602 74570 19710 74947
rect 19826 74570 19934 74947
rect 20050 74570 20214 74947
rect 20330 74570 20438 74947
rect 20554 74570 20662 74947
rect 20778 74570 20942 74947
rect 21058 74570 21166 74947
rect 21282 74570 21390 74947
rect 21506 74570 21614 74947
rect 21730 74570 21894 74947
rect 22010 74570 22118 74947
rect 22234 74570 22342 74947
rect 22458 74570 22622 74947
rect 22738 74570 22846 74947
rect 22962 74570 23070 74947
rect 23186 74570 23294 74947
rect 23410 74570 23574 74947
rect 23690 74570 23798 74947
rect 23914 74570 24022 74947
rect 24138 74570 24302 74947
rect 24418 74570 24526 74947
rect 24642 74570 24750 74947
rect 24866 74570 24974 74947
rect 25090 74570 25254 74947
rect 25370 74570 25478 74947
rect 25594 74570 25702 74947
rect 25818 74570 25982 74947
rect 26098 74570 26206 74947
rect 26322 74570 26430 74947
rect 26546 74570 26654 74947
rect 26770 74570 26934 74947
rect 27050 74570 27158 74947
rect 27274 74570 27382 74947
rect 27498 74570 27662 74947
rect 27778 74570 27886 74947
rect 28002 74570 28110 74947
rect 28226 74570 28334 74947
rect 28450 74570 28614 74947
rect 28730 74570 28838 74947
rect 28954 74570 29062 74947
rect 29178 74570 29342 74947
rect 29458 74570 29566 74947
rect 29682 74570 29790 74947
rect 29906 74570 29974 74947
rect 42 430 29974 74570
rect 42 373 110 430
rect 226 373 446 430
rect 562 373 782 430
rect 898 373 1118 430
rect 1234 373 1454 430
rect 1570 373 1790 430
rect 1906 373 2126 430
rect 2242 373 2462 430
rect 2578 373 2798 430
rect 2914 373 3134 430
rect 3250 373 3470 430
rect 3586 373 3806 430
rect 3922 373 4142 430
rect 4258 373 4478 430
rect 4594 373 4814 430
rect 4930 373 5150 430
rect 5266 373 5486 430
rect 5602 373 5822 430
rect 5938 373 6158 430
rect 6274 373 6494 430
rect 6610 373 6830 430
rect 6946 373 7166 430
rect 7282 373 7502 430
rect 7618 373 7838 430
rect 7954 373 8174 430
rect 8290 373 8510 430
rect 8626 373 8846 430
rect 8962 373 9182 430
rect 9298 373 9518 430
rect 9634 373 9854 430
rect 9970 373 10190 430
rect 10306 373 10526 430
rect 10642 373 10862 430
rect 10978 373 11198 430
rect 11314 373 11534 430
rect 11650 373 11870 430
rect 11986 373 12206 430
rect 12322 373 12542 430
rect 12658 373 12878 430
rect 12994 373 13214 430
rect 13330 373 13550 430
rect 13666 373 13886 430
rect 14002 373 14222 430
rect 14338 373 14558 430
rect 14674 373 14894 430
rect 15010 373 15286 430
rect 15402 373 15622 430
rect 15738 373 15958 430
rect 16074 373 16294 430
rect 16410 373 16630 430
rect 16746 373 16966 430
rect 17082 373 17302 430
rect 17418 373 17638 430
rect 17754 373 17974 430
rect 18090 373 18310 430
rect 18426 373 18646 430
rect 18762 373 18982 430
rect 19098 373 19318 430
rect 19434 373 19654 430
rect 19770 373 19990 430
rect 20106 373 20326 430
rect 20442 373 20662 430
rect 20778 373 20998 430
rect 21114 373 21334 430
rect 21450 373 21670 430
rect 21786 373 22006 430
rect 22122 373 22342 430
rect 22458 373 22678 430
rect 22794 373 23014 430
rect 23130 373 23350 430
rect 23466 373 23686 430
rect 23802 373 24022 430
rect 24138 373 24358 430
rect 24474 373 24694 430
rect 24810 373 25030 430
rect 25146 373 25366 430
rect 25482 373 25702 430
rect 25818 373 26038 430
rect 26154 373 26374 430
rect 26490 373 26710 430
rect 26826 373 27046 430
rect 27162 373 27382 430
rect 27498 373 27718 430
rect 27834 373 28054 430
rect 28170 373 28390 430
rect 28506 373 28726 430
rect 28842 373 29062 430
rect 29178 373 29398 430
rect 29514 373 29734 430
rect 29850 373 29974 430
<< metal3 >>
rect 0 74396 400 74452
rect 29600 74396 30000 74452
rect 0 73276 400 73332
rect 29600 73220 30000 73276
rect 0 72156 400 72212
rect 29600 72100 30000 72156
rect 0 70980 400 71036
rect 29600 70924 30000 70980
rect 0 69860 400 69916
rect 29600 69804 30000 69860
rect 0 68740 400 68796
rect 29600 68628 30000 68684
rect 0 67564 400 67620
rect 29600 67452 30000 67508
rect 0 66444 400 66500
rect 29600 66332 30000 66388
rect 0 65324 400 65380
rect 29600 65156 30000 65212
rect 0 64204 400 64260
rect 29600 64036 30000 64092
rect 0 63028 400 63084
rect 29600 62860 30000 62916
rect 0 61908 400 61964
rect 29600 61684 30000 61740
rect 0 60788 400 60844
rect 29600 60564 30000 60620
rect 0 59612 400 59668
rect 29600 59388 30000 59444
rect 0 58492 400 58548
rect 29600 58268 30000 58324
rect 0 57372 400 57428
rect 29600 57092 30000 57148
rect 0 56252 400 56308
rect 29600 55916 30000 55972
rect 0 55076 400 55132
rect 29600 54796 30000 54852
rect 0 53956 400 54012
rect 29600 53620 30000 53676
rect 0 52836 400 52892
rect 29600 52500 30000 52556
rect 0 51660 400 51716
rect 29600 51324 30000 51380
rect 0 50540 400 50596
rect 29600 50148 30000 50204
rect 0 49420 400 49476
rect 29600 49028 30000 49084
rect 0 48300 400 48356
rect 29600 47852 30000 47908
rect 0 47124 400 47180
rect 29600 46732 30000 46788
rect 0 46004 400 46060
rect 29600 45556 30000 45612
rect 0 44884 400 44940
rect 29600 44380 30000 44436
rect 0 43708 400 43764
rect 29600 43260 30000 43316
rect 0 42588 400 42644
rect 29600 42084 30000 42140
rect 0 41468 400 41524
rect 29600 40964 30000 41020
rect 0 40348 400 40404
rect 29600 39788 30000 39844
rect 0 39172 400 39228
rect 29600 38612 30000 38668
rect 0 38052 400 38108
rect 29600 37492 30000 37548
rect 0 36932 400 36988
rect 29600 36316 30000 36372
rect 0 35756 400 35812
rect 29600 35196 30000 35252
rect 0 34636 400 34692
rect 29600 34020 30000 34076
rect 0 33516 400 33572
rect 29600 32844 30000 32900
rect 0 32396 400 32452
rect 29600 31724 30000 31780
rect 0 31220 400 31276
rect 29600 30548 30000 30604
rect 0 30100 400 30156
rect 29600 29428 30000 29484
rect 0 28980 400 29036
rect 29600 28252 30000 28308
rect 0 27804 400 27860
rect 29600 27076 30000 27132
rect 0 26684 400 26740
rect 29600 25956 30000 26012
rect 0 25564 400 25620
rect 29600 24780 30000 24836
rect 0 24444 400 24500
rect 29600 23660 30000 23716
rect 0 23268 400 23324
rect 29600 22484 30000 22540
rect 0 22148 400 22204
rect 29600 21308 30000 21364
rect 0 21028 400 21084
rect 29600 20188 30000 20244
rect 0 19852 400 19908
rect 29600 19012 30000 19068
rect 0 18732 400 18788
rect 29600 17892 30000 17948
rect 0 17612 400 17668
rect 29600 16716 30000 16772
rect 0 16492 400 16548
rect 29600 15540 30000 15596
rect 0 15316 400 15372
rect 29600 14420 30000 14476
rect 0 14196 400 14252
rect 29600 13244 30000 13300
rect 0 13076 400 13132
rect 29600 12124 30000 12180
rect 0 11900 400 11956
rect 29600 10948 30000 11004
rect 0 10780 400 10836
rect 29600 9772 30000 9828
rect 0 9660 400 9716
rect 29600 8652 30000 8708
rect 0 8540 400 8596
rect 29600 7476 30000 7532
rect 0 7364 400 7420
rect 29600 6356 30000 6412
rect 0 6244 400 6300
rect 0 5124 400 5180
rect 29600 5180 30000 5236
rect 0 3948 400 4004
rect 29600 4004 30000 4060
rect 0 2828 400 2884
rect 29600 2884 30000 2940
rect 0 1708 400 1764
rect 29600 1708 30000 1764
rect 0 588 400 644
rect 29600 588 30000 644
<< obsm3 >>
rect 0 74482 29979 74998
rect 430 74366 29570 74482
rect 0 73362 29979 74366
rect 430 73306 29979 73362
rect 430 73246 29570 73306
rect 0 73190 29570 73246
rect 0 72242 29979 73190
rect 430 72186 29979 72242
rect 430 72126 29570 72186
rect 0 72070 29570 72126
rect 0 71066 29979 72070
rect 430 71010 29979 71066
rect 430 70950 29570 71010
rect 0 70894 29570 70950
rect 0 69946 29979 70894
rect 430 69890 29979 69946
rect 430 69830 29570 69890
rect 0 69774 29570 69830
rect 0 68826 29979 69774
rect 430 68714 29979 68826
rect 430 68710 29570 68714
rect 0 68598 29570 68710
rect 0 67650 29979 68598
rect 430 67538 29979 67650
rect 430 67534 29570 67538
rect 0 67422 29570 67534
rect 0 66530 29979 67422
rect 430 66418 29979 66530
rect 430 66414 29570 66418
rect 0 66302 29570 66414
rect 0 65410 29979 66302
rect 430 65294 29979 65410
rect 0 65242 29979 65294
rect 0 65126 29570 65242
rect 0 64290 29979 65126
rect 430 64174 29979 64290
rect 0 64122 29979 64174
rect 0 64006 29570 64122
rect 0 63114 29979 64006
rect 430 62998 29979 63114
rect 0 62946 29979 62998
rect 0 62830 29570 62946
rect 0 61994 29979 62830
rect 430 61878 29979 61994
rect 0 61770 29979 61878
rect 0 61654 29570 61770
rect 0 60874 29979 61654
rect 430 60758 29979 60874
rect 0 60650 29979 60758
rect 0 60534 29570 60650
rect 0 59698 29979 60534
rect 430 59582 29979 59698
rect 0 59474 29979 59582
rect 0 59358 29570 59474
rect 0 58578 29979 59358
rect 430 58462 29979 58578
rect 0 58354 29979 58462
rect 0 58238 29570 58354
rect 0 57458 29979 58238
rect 430 57342 29979 57458
rect 0 57178 29979 57342
rect 0 57062 29570 57178
rect 0 56338 29979 57062
rect 430 56222 29979 56338
rect 0 56070 29979 56222
rect -14 56002 29979 56070
rect -14 55886 29570 56002
rect -14 55818 29979 55886
rect 0 55162 29979 55818
rect 430 55046 29979 55162
rect 0 54882 29979 55046
rect 0 54766 29570 54882
rect 0 54042 29979 54766
rect 430 53926 29979 54042
rect 0 53706 29979 53926
rect 0 53590 29570 53706
rect 0 52922 29979 53590
rect 430 52806 29979 52922
rect 0 52586 29979 52806
rect 0 52470 29570 52586
rect 0 51746 29979 52470
rect 430 51630 29979 51746
rect 0 51410 29979 51630
rect 0 51294 29570 51410
rect 0 50626 29979 51294
rect 430 50510 29979 50626
rect 0 50234 29979 50510
rect 0 50118 29570 50234
rect 0 49506 29979 50118
rect 430 49390 29979 49506
rect 0 49114 29979 49390
rect 0 48998 29570 49114
rect 0 48386 29979 48998
rect 430 48270 29979 48386
rect 0 47938 29979 48270
rect 0 47822 29570 47938
rect 0 47210 29979 47822
rect 430 47094 29979 47210
rect 0 46818 29979 47094
rect 0 46702 29570 46818
rect 0 46090 29979 46702
rect 430 45974 29979 46090
rect 0 45642 29979 45974
rect 0 45526 29570 45642
rect 0 44970 29979 45526
rect 430 44854 29979 44970
rect 0 44466 29979 44854
rect 0 44350 29570 44466
rect 0 43794 29979 44350
rect 430 43678 29979 43794
rect 0 43346 29979 43678
rect 0 43230 29570 43346
rect 0 42674 29979 43230
rect 430 42558 29979 42674
rect 0 42170 29979 42558
rect 0 42054 29570 42170
rect 0 41554 29979 42054
rect 430 41438 29979 41554
rect 0 41050 29979 41438
rect 0 40934 29570 41050
rect 0 40434 29979 40934
rect 430 40318 29979 40434
rect 0 39874 29979 40318
rect 0 39758 29570 39874
rect 0 39258 29979 39758
rect 430 39142 29979 39258
rect 0 38698 29979 39142
rect 0 38582 29570 38698
rect 0 38138 29979 38582
rect 430 38022 29979 38138
rect 0 37578 29979 38022
rect 0 37462 29570 37578
rect 0 37018 29979 37462
rect 430 36902 29979 37018
rect 0 36402 29979 36902
rect 0 36286 29570 36402
rect 0 35842 29979 36286
rect 430 35726 29979 35842
rect 0 35282 29979 35726
rect 0 35166 29570 35282
rect 0 34722 29979 35166
rect 430 34606 29979 34722
rect 0 34106 29979 34606
rect 0 33990 29570 34106
rect 0 33602 29979 33990
rect 430 33486 29979 33602
rect 0 32930 29979 33486
rect 0 32814 29570 32930
rect 0 32482 29979 32814
rect 430 32366 29979 32482
rect 0 31810 29979 32366
rect 0 31694 29570 31810
rect 0 31306 29979 31694
rect 430 31190 29979 31306
rect 0 30634 29979 31190
rect 0 30518 29570 30634
rect 0 30186 29979 30518
rect 430 30070 29979 30186
rect 0 29514 29979 30070
rect 0 29398 29570 29514
rect 0 29066 29979 29398
rect 430 28950 29979 29066
rect 0 28338 29979 28950
rect 0 28222 29570 28338
rect 0 27890 29979 28222
rect 430 27774 29979 27890
rect 0 27162 29979 27774
rect 0 27046 29570 27162
rect 0 26770 29979 27046
rect 430 26654 29979 26770
rect 0 26042 29979 26654
rect 0 25926 29570 26042
rect 0 25650 29979 25926
rect 430 25534 29979 25650
rect 0 24866 29979 25534
rect 0 24750 29570 24866
rect 0 24530 29979 24750
rect 430 24414 29979 24530
rect 0 23746 29979 24414
rect 0 23630 29570 23746
rect 0 23354 29979 23630
rect 430 23238 29979 23354
rect 0 22570 29979 23238
rect 0 22454 29570 22570
rect 0 22234 29979 22454
rect 430 22118 29979 22234
rect 0 21394 29979 22118
rect 0 21278 29570 21394
rect 0 21114 29979 21278
rect 430 20998 29979 21114
rect 0 20274 29979 20998
rect 0 20158 29570 20274
rect 0 19938 29979 20158
rect 430 19822 29979 19938
rect 0 19098 29979 19822
rect 0 18982 29570 19098
rect 0 18818 29979 18982
rect 430 18702 29979 18818
rect 0 17978 29979 18702
rect 0 17862 29570 17978
rect 0 17698 29979 17862
rect 430 17582 29979 17698
rect 0 16802 29979 17582
rect 0 16686 29570 16802
rect 0 16578 29979 16686
rect 430 16462 29979 16578
rect 0 15626 29979 16462
rect 0 15510 29570 15626
rect 0 15402 29979 15510
rect 430 15286 29979 15402
rect 0 14506 29979 15286
rect 0 14390 29570 14506
rect 0 14282 29979 14390
rect 430 14166 29979 14282
rect 0 13330 29979 14166
rect 0 13214 29570 13330
rect 0 13162 29979 13214
rect 430 13046 29979 13162
rect 0 12210 29979 13046
rect 0 12094 29570 12210
rect 0 11986 29979 12094
rect 430 11870 29979 11986
rect 0 11034 29979 11870
rect 0 10918 29570 11034
rect 0 10866 29979 10918
rect 430 10750 29979 10866
rect 0 9858 29979 10750
rect 0 9746 29570 9858
rect 430 9742 29570 9746
rect 430 9630 29979 9742
rect 0 8738 29979 9630
rect 0 8626 29570 8738
rect 430 8622 29570 8626
rect 430 8510 29979 8622
rect 0 7562 29979 8510
rect 0 7450 29570 7562
rect 430 7446 29570 7450
rect 430 7334 29979 7446
rect 0 6442 29979 7334
rect 0 6330 29570 6442
rect 430 6326 29570 6330
rect 430 6214 29979 6326
rect 0 5266 29979 6214
rect 0 5210 29570 5266
rect 430 5150 29570 5210
rect 430 5094 29979 5150
rect 0 4090 29979 5094
rect 0 4034 29570 4090
rect 430 3974 29570 4034
rect 430 3918 29979 3974
rect 0 2970 29979 3918
rect 0 2914 29570 2970
rect 430 2854 29570 2914
rect 430 2798 29979 2854
rect 0 1794 29979 2798
rect 430 1678 29570 1794
rect 0 674 29979 1678
rect 430 558 29570 674
rect 0 322 29979 558
<< metal4 >>
rect 2224 1538 2384 73334
rect 9904 1538 10064 73334
rect 17584 1538 17744 73334
rect 25264 1538 25424 73334
<< obsm4 >>
rect 42 73364 29974 74989
rect 42 1508 2194 73364
rect 2414 1508 9874 73364
rect 10094 1508 17554 73364
rect 17774 1508 25234 73364
rect 25454 1508 29974 73364
rect 42 317 29974 1508
<< metal5 >>
rect 642 72084 29318 72244
rect 642 64425 29318 64585
rect 642 56766 29318 56926
rect 642 49107 29318 49267
rect 642 41448 29318 41608
rect 642 33789 29318 33949
rect 642 26130 29318 26290
rect 642 18471 29318 18631
rect 642 10812 29318 10972
rect 642 3153 29318 3313
<< obsm5 >>
rect 34 72294 29982 74992
rect 34 72034 592 72294
rect 29368 72034 29982 72294
rect 34 64635 29982 72034
rect 34 64375 592 64635
rect 29368 64375 29982 64635
rect 34 56976 29982 64375
rect 34 56716 592 56976
rect 29368 56716 29982 56976
rect 34 49317 29982 56716
rect 34 49057 592 49317
rect 29368 49057 29982 49317
rect 34 41658 29982 49057
rect 34 41398 592 41658
rect 29368 41398 29982 41658
rect 34 33999 29982 41398
rect 34 33739 592 33999
rect 29368 33739 29982 33999
rect 34 26340 29982 33739
rect 34 26080 592 26340
rect 29368 26080 29982 26340
rect 34 18681 29982 26080
rect 34 18421 592 18681
rect 29368 18421 29982 18681
rect 34 11022 29982 18421
rect 34 10762 592 11022
rect 29368 10762 29982 11022
rect 34 3363 29982 10762
rect 34 3103 592 3363
rect 29368 3103 29982 3363
rect 34 1688 29982 3103
<< labels >>
rlabel metal4 s 2224 1538 2384 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 73334 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 3153 29318 3313 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 18471 29318 18631 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 33789 29318 33949 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 49107 29318 49267 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 642 64425 29318 64585 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 73334 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 10812 29318 10972 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 26130 29318 26290 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 41448 29318 41608 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 56766 29318 56926 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 642 72084 29318 72244 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 588 400 644 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 1708 400 1764 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 2828 400 2884 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 3948 400 4004 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 6244 400 6300 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 7364 400 7420 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 8540 400 8596 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 19012 0 19068 400 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 22372 0 22428 400 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 22708 0 22764 400 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 23044 0 23100 400 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 23380 0 23436 400 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 23716 0 23772 400 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 24052 0 24108 400 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 24388 0 24444 400 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 24724 0 24780 400 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 25060 0 25116 400 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 25396 0 25452 400 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 19348 0 19404 400 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 25732 0 25788 400 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 26068 0 26124 400 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 26404 0 26460 400 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 26740 0 26796 400 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 27076 0 27132 400 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 27412 0 27468 400 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 27748 0 27804 400 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 28084 0 28140 400 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 28420 0 28476 400 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 28756 0 28812 400 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 19684 0 19740 400 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 29092 0 29148 400 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 29428 0 29484 400 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 20020 0 20076 400 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 20356 0 20412 400 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 20692 0 20748 400 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 21028 0 21084 400 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 21364 0 21420 400 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 21700 0 21756 400 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 22036 0 22092 400 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 29600 6356 30000 6412 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 29600 40964 30000 41020 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 29600 44380 30000 44436 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 29600 47852 30000 47908 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 29600 51324 30000 51380 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 29600 54796 30000 54852 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 29600 58268 30000 58324 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 29600 61684 30000 61740 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 29600 65156 30000 65212 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 29600 68628 30000 68684 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 29600 72100 30000 72156 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 29600 9772 30000 9828 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal2 s 17108 74600 17164 75000 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal2 s 17836 74600 17892 75000 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal2 s 18564 74600 18620 75000 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal2 s 19292 74600 19348 75000 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal2 s 19964 74600 20020 75000 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal2 s 20692 74600 20748 75000 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal2 s 21420 74600 21476 75000 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal2 s 22148 74600 22204 75000 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal2 s 22876 74600 22932 75000 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal2 s 23604 74600 23660 75000 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 29600 13244 30000 13300 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal2 s 24332 74600 24388 75000 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal2 s 25004 74600 25060 75000 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal2 s 25732 74600 25788 75000 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal2 s 26460 74600 26516 75000 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal2 s 27188 74600 27244 75000 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal2 s 27916 74600 27972 75000 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal2 s 28644 74600 28700 75000 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal2 s 29372 74600 29428 75000 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 29600 16716 30000 16772 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 29600 20188 30000 20244 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 29600 23660 30000 23716 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 29600 27076 30000 27132 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 29600 30548 30000 30604 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 29600 34020 30000 34076 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 29600 37492 30000 37548 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 29600 7476 30000 7532 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 29600 42084 30000 42140 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 29600 45556 30000 45612 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 29600 49028 30000 49084 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 29600 52500 30000 52556 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 29600 55916 30000 55972 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 29600 59388 30000 59444 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 29600 62860 30000 62916 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 29600 66332 30000 66388 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 29600 69804 30000 69860 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 29600 73220 30000 73276 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 29600 10948 30000 11004 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal2 s 17332 74600 17388 75000 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal2 s 18060 74600 18116 75000 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal2 s 18788 74600 18844 75000 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal2 s 19516 74600 19572 75000 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal2 s 20244 74600 20300 75000 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal2 s 20972 74600 21028 75000 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal2 s 21644 74600 21700 75000 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal2 s 22372 74600 22428 75000 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal2 s 23100 74600 23156 75000 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal2 s 23828 74600 23884 75000 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 29600 14420 30000 14476 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal2 s 24556 74600 24612 75000 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal2 s 25284 74600 25340 75000 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal2 s 26012 74600 26068 75000 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal2 s 26684 74600 26740 75000 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal2 s 27412 74600 27468 75000 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal2 s 28140 74600 28196 75000 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal2 s 28868 74600 28924 75000 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal2 s 29596 74600 29652 75000 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 29600 17892 30000 17948 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 29600 21308 30000 21364 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 29600 24780 30000 24836 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 29600 28252 30000 28308 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 29600 31724 30000 31780 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 29600 35196 30000 35252 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 29600 38612 30000 38668 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 29600 8652 30000 8708 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 29600 43260 30000 43316 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 29600 46732 30000 46788 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 29600 50148 30000 50204 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 29600 53620 30000 53676 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 29600 57092 30000 57148 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 29600 60564 30000 60620 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 29600 64036 30000 64092 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 29600 67452 30000 67508 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 29600 70924 30000 70980 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 29600 74396 30000 74452 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 29600 12124 30000 12180 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal2 s 17612 74600 17668 75000 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal2 s 18284 74600 18340 75000 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal2 s 19012 74600 19068 75000 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal2 s 19740 74600 19796 75000 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal2 s 20468 74600 20524 75000 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal2 s 21196 74600 21252 75000 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal2 s 21924 74600 21980 75000 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal2 s 22652 74600 22708 75000 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal2 s 23324 74600 23380 75000 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal2 s 24052 74600 24108 75000 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 29600 15540 30000 15596 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal2 s 24780 74600 24836 75000 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal2 s 25508 74600 25564 75000 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal2 s 26236 74600 26292 75000 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal2 s 26964 74600 27020 75000 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal2 s 27692 74600 27748 75000 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal2 s 28364 74600 28420 75000 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal2 s 29092 74600 29148 75000 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal2 s 29820 74600 29876 75000 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 29600 19012 30000 19068 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 29600 22484 30000 22540 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 29600 25956 30000 26012 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 29600 29428 30000 29484 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 29600 32844 30000 32900 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 29600 36316 30000 36372 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 29600 39788 30000 39844 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 140 0 196 400 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 476 0 532 400 6 pad_flash_clk_oe
port 157 nsew signal output
rlabel metal2 s 812 0 868 400 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 1148 0 1204 400 6 pad_flash_csb_oe
port 159 nsew signal output
rlabel metal2 s 1484 0 1540 400 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 1820 0 1876 400 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 2156 0 2212 400 6 pad_flash_io0_ie
port 162 nsew signal output
rlabel metal2 s 2492 0 2548 400 6 pad_flash_io0_oe
port 163 nsew signal output
rlabel metal2 s 2828 0 2884 400 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 3164 0 3220 400 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 3500 0 3556 400 6 pad_flash_io1_ie
port 166 nsew signal output
rlabel metal2 s 3836 0 3892 400 6 pad_flash_io1_oe
port 167 nsew signal output
rlabel metal2 s 8204 0 8260 400 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 8540 0 8596 400 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 8876 0 8932 400 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 18004 0 18060 400 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 5180 0 5236 400 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 5516 0 5572 400 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 5852 0 5908 400 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 6188 0 6244 400 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 6524 0 6580 400 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 6860 0 6916 400 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 4844 0 4900 400 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 7196 0 7252 400 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 7532 0 7588 400 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 7868 0 7924 400 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 9212 0 9268 400 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 12572 0 12628 400 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 12908 0 12964 400 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 13244 0 13300 400 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 13580 0 13636 400 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 13916 0 13972 400 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 14252 0 14308 400 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 14588 0 14644 400 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 14924 0 14980 400 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 15316 0 15372 400 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 15652 0 15708 400 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 9548 0 9604 400 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 15988 0 16044 400 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 16324 0 16380 400 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 16660 0 16716 400 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 16996 0 17052 400 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 17332 0 17388 400 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 17668 0 17724 400 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 9884 0 9940 400 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 10220 0 10276 400 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 10556 0 10612 400 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 10892 0 10948 400 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 11228 0 11284 400 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 11564 0 11620 400 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 11900 0 11956 400 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 12236 0 12292 400 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 4172 0 4228 400 6 porb
port 208 nsew signal input
rlabel metal2 s 29764 0 29820 400 6 pwr_ctrl_out
port 209 nsew signal output
rlabel metal3 s 0 17612 400 17668 6 qspi_enabled
port 210 nsew signal input
rlabel metal2 s 4508 0 4564 400 6 reset
port 211 nsew signal output
rlabel metal3 s 0 16492 400 16548 6 ser_rx
port 212 nsew signal output
rlabel metal3 s 0 15316 400 15372 6 ser_tx
port 213 nsew signal input
rlabel metal3 s 29600 588 30000 644 6 serial_clock
port 214 nsew signal output
rlabel metal3 s 29600 4004 30000 4060 6 serial_data_1
port 215 nsew signal output
rlabel metal3 s 29600 5180 30000 5236 6 serial_data_2
port 216 nsew signal output
rlabel metal3 s 29600 2884 30000 2940 6 serial_load
port 217 nsew signal output
rlabel metal3 s 29600 1708 30000 1764 6 serial_resetn
port 218 nsew signal output
rlabel metal3 s 0 13076 400 13132 6 spi_csb
port 219 nsew signal input
rlabel metal3 s 0 19852 400 19908 6 spi_enabled
port 220 nsew signal input
rlabel metal3 s 0 11900 400 11956 6 spi_sck
port 221 nsew signal input
rlabel metal3 s 0 14196 400 14252 6 spi_sdi
port 222 nsew signal output
rlabel metal3 s 0 10780 400 10836 6 spi_sdo
port 223 nsew signal input
rlabel metal3 s 0 9660 400 9716 6 spi_sdoenb
port 224 nsew signal input
rlabel metal3 s 0 59612 400 59668 6 spimemio_flash_clk
port 225 nsew signal input
rlabel metal3 s 0 60788 400 60844 6 spimemio_flash_csb
port 226 nsew signal input
rlabel metal3 s 0 61908 400 61964 6 spimemio_flash_io0_di
port 227 nsew signal output
rlabel metal3 s 0 63028 400 63084 6 spimemio_flash_io0_do
port 228 nsew signal input
rlabel metal3 s 0 64204 400 64260 6 spimemio_flash_io0_oeb
port 229 nsew signal input
rlabel metal3 s 0 65324 400 65380 6 spimemio_flash_io1_di
port 230 nsew signal output
rlabel metal3 s 0 66444 400 66500 6 spimemio_flash_io1_do
port 231 nsew signal input
rlabel metal3 s 0 67564 400 67620 6 spimemio_flash_io1_oeb
port 232 nsew signal input
rlabel metal3 s 0 68740 400 68796 6 spimemio_flash_io2_di
port 233 nsew signal output
rlabel metal3 s 0 69860 400 69916 6 spimemio_flash_io2_do
port 234 nsew signal input
rlabel metal3 s 0 70980 400 71036 6 spimemio_flash_io2_oeb
port 235 nsew signal input
rlabel metal3 s 0 72156 400 72212 6 spimemio_flash_io3_di
port 236 nsew signal output
rlabel metal3 s 0 73276 400 73332 6 spimemio_flash_io3_do
port 237 nsew signal input
rlabel metal3 s 0 74396 400 74452 6 spimemio_flash_io3_oeb
port 238 nsew signal input
rlabel metal3 s 0 5124 400 5180 6 trap
port 239 nsew signal input
rlabel metal3 s 0 18732 400 18788 6 uart_enabled
port 240 nsew signal input
rlabel metal2 s 16884 74600 16940 75000 6 user_clock
port 241 nsew signal input
rlabel metal3 s 0 21028 400 21084 6 wb_ack_o
port 242 nsew signal output
rlabel metal2 s 84 74600 140 75000 6 wb_adr_i[0]
port 243 nsew signal input
rlabel metal2 s 2436 74600 2492 75000 6 wb_adr_i[10]
port 244 nsew signal input
rlabel metal2 s 2716 74600 2772 75000 6 wb_adr_i[11]
port 245 nsew signal input
rlabel metal2 s 2940 74600 2996 75000 6 wb_adr_i[12]
port 246 nsew signal input
rlabel metal2 s 3164 74600 3220 75000 6 wb_adr_i[13]
port 247 nsew signal input
rlabel metal2 s 3444 74600 3500 75000 6 wb_adr_i[14]
port 248 nsew signal input
rlabel metal2 s 3668 74600 3724 75000 6 wb_adr_i[15]
port 249 nsew signal input
rlabel metal2 s 3892 74600 3948 75000 6 wb_adr_i[16]
port 250 nsew signal input
rlabel metal2 s 4116 74600 4172 75000 6 wb_adr_i[17]
port 251 nsew signal input
rlabel metal2 s 4396 74600 4452 75000 6 wb_adr_i[18]
port 252 nsew signal input
rlabel metal2 s 4620 74600 4676 75000 6 wb_adr_i[19]
port 253 nsew signal input
rlabel metal2 s 308 74600 364 75000 6 wb_adr_i[1]
port 254 nsew signal input
rlabel metal2 s 4844 74600 4900 75000 6 wb_adr_i[20]
port 255 nsew signal input
rlabel metal2 s 5124 74600 5180 75000 6 wb_adr_i[21]
port 256 nsew signal input
rlabel metal2 s 5348 74600 5404 75000 6 wb_adr_i[22]
port 257 nsew signal input
rlabel metal2 s 5572 74600 5628 75000 6 wb_adr_i[23]
port 258 nsew signal input
rlabel metal2 s 5796 74600 5852 75000 6 wb_adr_i[24]
port 259 nsew signal input
rlabel metal2 s 6076 74600 6132 75000 6 wb_adr_i[25]
port 260 nsew signal input
rlabel metal2 s 6300 74600 6356 75000 6 wb_adr_i[26]
port 261 nsew signal input
rlabel metal2 s 6524 74600 6580 75000 6 wb_adr_i[27]
port 262 nsew signal input
rlabel metal2 s 6804 74600 6860 75000 6 wb_adr_i[28]
port 263 nsew signal input
rlabel metal2 s 7028 74600 7084 75000 6 wb_adr_i[29]
port 264 nsew signal input
rlabel metal2 s 532 74600 588 75000 6 wb_adr_i[2]
port 265 nsew signal input
rlabel metal2 s 7252 74600 7308 75000 6 wb_adr_i[30]
port 266 nsew signal input
rlabel metal2 s 7476 74600 7532 75000 6 wb_adr_i[31]
port 267 nsew signal input
rlabel metal2 s 756 74600 812 75000 6 wb_adr_i[3]
port 268 nsew signal input
rlabel metal2 s 1036 74600 1092 75000 6 wb_adr_i[4]
port 269 nsew signal input
rlabel metal2 s 1260 74600 1316 75000 6 wb_adr_i[5]
port 270 nsew signal input
rlabel metal2 s 1484 74600 1540 75000 6 wb_adr_i[6]
port 271 nsew signal input
rlabel metal2 s 1764 74600 1820 75000 6 wb_adr_i[7]
port 272 nsew signal input
rlabel metal2 s 1988 74600 2044 75000 6 wb_adr_i[8]
port 273 nsew signal input
rlabel metal2 s 2212 74600 2268 75000 6 wb_adr_i[9]
port 274 nsew signal input
rlabel metal2 s 18340 0 18396 400 6 wb_clk_i
port 275 nsew signal input
rlabel metal2 s 16604 74600 16660 75000 6 wb_cyc_i
port 276 nsew signal input
rlabel metal2 s 7756 74600 7812 75000 6 wb_dat_i[0]
port 277 nsew signal input
rlabel metal2 s 10164 74600 10220 75000 6 wb_dat_i[10]
port 278 nsew signal input
rlabel metal2 s 10388 74600 10444 75000 6 wb_dat_i[11]
port 279 nsew signal input
rlabel metal2 s 10612 74600 10668 75000 6 wb_dat_i[12]
port 280 nsew signal input
rlabel metal2 s 10836 74600 10892 75000 6 wb_dat_i[13]
port 281 nsew signal input
rlabel metal2 s 11116 74600 11172 75000 6 wb_dat_i[14]
port 282 nsew signal input
rlabel metal2 s 11340 74600 11396 75000 6 wb_dat_i[15]
port 283 nsew signal input
rlabel metal2 s 11564 74600 11620 75000 6 wb_dat_i[16]
port 284 nsew signal input
rlabel metal2 s 11844 74600 11900 75000 6 wb_dat_i[17]
port 285 nsew signal input
rlabel metal2 s 12068 74600 12124 75000 6 wb_dat_i[18]
port 286 nsew signal input
rlabel metal2 s 12292 74600 12348 75000 6 wb_dat_i[19]
port 287 nsew signal input
rlabel metal2 s 7980 74600 8036 75000 6 wb_dat_i[1]
port 288 nsew signal input
rlabel metal2 s 12516 74600 12572 75000 6 wb_dat_i[20]
port 289 nsew signal input
rlabel metal2 s 12796 74600 12852 75000 6 wb_dat_i[21]
port 290 nsew signal input
rlabel metal2 s 13020 74600 13076 75000 6 wb_dat_i[22]
port 291 nsew signal input
rlabel metal2 s 13244 74600 13300 75000 6 wb_dat_i[23]
port 292 nsew signal input
rlabel metal2 s 13524 74600 13580 75000 6 wb_dat_i[24]
port 293 nsew signal input
rlabel metal2 s 13748 74600 13804 75000 6 wb_dat_i[25]
port 294 nsew signal input
rlabel metal2 s 13972 74600 14028 75000 6 wb_dat_i[26]
port 295 nsew signal input
rlabel metal2 s 14196 74600 14252 75000 6 wb_dat_i[27]
port 296 nsew signal input
rlabel metal2 s 14476 74600 14532 75000 6 wb_dat_i[28]
port 297 nsew signal input
rlabel metal2 s 14700 74600 14756 75000 6 wb_dat_i[29]
port 298 nsew signal input
rlabel metal2 s 8204 74600 8260 75000 6 wb_dat_i[2]
port 299 nsew signal input
rlabel metal2 s 14924 74600 14980 75000 6 wb_dat_i[30]
port 300 nsew signal input
rlabel metal2 s 15204 74600 15260 75000 6 wb_dat_i[31]
port 301 nsew signal input
rlabel metal2 s 8484 74600 8540 75000 6 wb_dat_i[3]
port 302 nsew signal input
rlabel metal2 s 8708 74600 8764 75000 6 wb_dat_i[4]
port 303 nsew signal input
rlabel metal2 s 8932 74600 8988 75000 6 wb_dat_i[5]
port 304 nsew signal input
rlabel metal2 s 9156 74600 9212 75000 6 wb_dat_i[6]
port 305 nsew signal input
rlabel metal2 s 9436 74600 9492 75000 6 wb_dat_i[7]
port 306 nsew signal input
rlabel metal2 s 9660 74600 9716 75000 6 wb_dat_i[8]
port 307 nsew signal input
rlabel metal2 s 9884 74600 9940 75000 6 wb_dat_i[9]
port 308 nsew signal input
rlabel metal3 s 0 23268 400 23324 6 wb_dat_o[0]
port 309 nsew signal output
rlabel metal3 s 0 34636 400 34692 6 wb_dat_o[10]
port 310 nsew signal output
rlabel metal3 s 0 35756 400 35812 6 wb_dat_o[11]
port 311 nsew signal output
rlabel metal3 s 0 36932 400 36988 6 wb_dat_o[12]
port 312 nsew signal output
rlabel metal3 s 0 38052 400 38108 6 wb_dat_o[13]
port 313 nsew signal output
rlabel metal3 s 0 39172 400 39228 6 wb_dat_o[14]
port 314 nsew signal output
rlabel metal3 s 0 40348 400 40404 6 wb_dat_o[15]
port 315 nsew signal output
rlabel metal3 s 0 41468 400 41524 6 wb_dat_o[16]
port 316 nsew signal output
rlabel metal3 s 0 42588 400 42644 6 wb_dat_o[17]
port 317 nsew signal output
rlabel metal3 s 0 43708 400 43764 6 wb_dat_o[18]
port 318 nsew signal output
rlabel metal3 s 0 44884 400 44940 6 wb_dat_o[19]
port 319 nsew signal output
rlabel metal3 s 0 24444 400 24500 6 wb_dat_o[1]
port 320 nsew signal output
rlabel metal3 s 0 46004 400 46060 6 wb_dat_o[20]
port 321 nsew signal output
rlabel metal3 s 0 47124 400 47180 6 wb_dat_o[21]
port 322 nsew signal output
rlabel metal3 s 0 48300 400 48356 6 wb_dat_o[22]
port 323 nsew signal output
rlabel metal3 s 0 49420 400 49476 6 wb_dat_o[23]
port 324 nsew signal output
rlabel metal3 s 0 50540 400 50596 6 wb_dat_o[24]
port 325 nsew signal output
rlabel metal3 s 0 51660 400 51716 6 wb_dat_o[25]
port 326 nsew signal output
rlabel metal3 s 0 52836 400 52892 6 wb_dat_o[26]
port 327 nsew signal output
rlabel metal3 s 0 53956 400 54012 6 wb_dat_o[27]
port 328 nsew signal output
rlabel metal3 s 0 55076 400 55132 6 wb_dat_o[28]
port 329 nsew signal output
rlabel metal3 s 0 56252 400 56308 6 wb_dat_o[29]
port 330 nsew signal output
rlabel metal3 s 0 25564 400 25620 6 wb_dat_o[2]
port 331 nsew signal output
rlabel metal3 s 0 57372 400 57428 6 wb_dat_o[30]
port 332 nsew signal output
rlabel metal3 s 0 58492 400 58548 6 wb_dat_o[31]
port 333 nsew signal output
rlabel metal3 s 0 26684 400 26740 6 wb_dat_o[3]
port 334 nsew signal output
rlabel metal3 s 0 27804 400 27860 6 wb_dat_o[4]
port 335 nsew signal output
rlabel metal3 s 0 28980 400 29036 6 wb_dat_o[5]
port 336 nsew signal output
rlabel metal3 s 0 30100 400 30156 6 wb_dat_o[6]
port 337 nsew signal output
rlabel metal3 s 0 31220 400 31276 6 wb_dat_o[7]
port 338 nsew signal output
rlabel metal3 s 0 32396 400 32452 6 wb_dat_o[8]
port 339 nsew signal output
rlabel metal3 s 0 33516 400 33572 6 wb_dat_o[9]
port 340 nsew signal output
rlabel metal2 s 18676 0 18732 400 6 wb_rstn_i
port 341 nsew signal input
rlabel metal2 s 15428 74600 15484 75000 6 wb_sel_i[0]
port 342 nsew signal input
rlabel metal2 s 15652 74600 15708 75000 6 wb_sel_i[1]
port 343 nsew signal input
rlabel metal2 s 15932 74600 15988 75000 6 wb_sel_i[2]
port 344 nsew signal input
rlabel metal2 s 16156 74600 16212 75000 6 wb_sel_i[3]
port 345 nsew signal input
rlabel metal3 s 0 22148 400 22204 6 wb_stb_i
port 346 nsew signal input
rlabel metal2 s 16380 74600 16436 75000 6 wb_we_i
port 347 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 75000
string GDS_END 15847012
string GDS_FILE ../gds/housekeeping.gds.gz
string GDS_START 400576
string LEFclass BLOCK
string LEFview TRUE
<< end >>
