magic
tech gf180mcuC
magscale 1 5
timestamp 1669509657
use caravel_core  chip_core
timestamp 0
transform 1 0 35500 0 1 35500
box -400 -422 317400 436400
use chip_io  padframe
timestamp 0
transform 1 0 0 0 1 0
box 0 0 388000 507000
<< properties >>
string FIXED_BBOX 0 0 389000 510000
<< end >>
