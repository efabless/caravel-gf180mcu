magic
tech gf180mcuD
magscale 6 5
timestamp 1654634570
<< metal5 >>
rect 72 720 324 756
rect 36 684 324 720
rect 0 612 324 684
rect 0 144 108 612
rect 0 72 324 144
rect 36 36 324 72
rect 72 0 324 36
<< properties >>
string FIXED_BBOX 0 0 432 756
<< end >>
