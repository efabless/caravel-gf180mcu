VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_logo
  CLASS BLOCK ;
  FOREIGN caravel_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 58.400 BY 51.865 ;
  OBS
      LAYER Metal4 ;
        RECT -3.730 0.465 49.465 1.865 ;
      LAYER Metal5 ;
        RECT 26.130 50.865 27.300 51.330 ;
        POLYGON 23.565 50.865 23.565 50.400 23.100 50.400 ;
        RECT 23.565 50.400 27.300 50.865 ;
        POLYGON 23.100 49.930 23.100 49.465 22.630 49.465 ;
        RECT 23.100 49.465 27.300 50.400 ;
        POLYGON 19.230 49.465 19.230 49.000 18.765 49.000 ;
        RECT 19.230 49.000 24.265 49.465 ;
        RECT 18.765 48.765 24.265 49.000 ;
        POLYGON 18.765 48.530 18.765 48.065 18.300 48.065 ;
        RECT 18.765 48.300 23.800 48.765 ;
        POLYGON 23.800 48.765 24.265 48.765 23.800 48.300 ;
        RECT 18.765 48.065 19.830 48.300 ;
        POLYGON 19.830 48.300 20.065 48.300 19.830 48.065 ;
        RECT 16.800 47.365 19.830 48.065 ;
        RECT 26.130 47.830 27.300 49.465 ;
        RECT 26.130 47.600 32.200 47.830 ;
        RECT 16.800 46.900 19.365 47.365 ;
        POLYGON 19.365 47.365 19.830 47.365 19.365 46.900 ;
        POLYGON 24.730 47.600 24.730 47.130 24.265 47.130 ;
        RECT 24.730 47.130 32.200 47.600 ;
        POLYGON 21.930 47.130 21.930 46.900 21.700 46.900 ;
        RECT 21.930 46.900 32.200 47.130 ;
        POLYGON 21.700 46.900 21.700 44.800 19.600 44.800 ;
        RECT 21.700 46.665 32.200 46.900 ;
        RECT 21.700 45.265 31.265 46.665 ;
        POLYGON 31.265 46.665 31.730 46.665 31.265 46.200 ;
        RECT 21.700 44.800 30.800 45.265 ;
        POLYGON 30.800 45.265 31.265 45.265 30.800 44.800 ;
        POLYGON 19.600 43.400 19.600 42.930 19.130 42.930 ;
        RECT 19.600 42.930 30.800 44.800 ;
        RECT 19.130 42.000 30.800 42.930 ;
        POLYGON 30.800 42.465 31.265 42.000 30.800 42.000 ;
        RECT 9.330 38.730 10.500 41.065 ;
        RECT 19.130 40.130 31.265 42.000 ;
        POLYGON 19.130 40.130 19.600 40.130 19.600 39.665 ;
        RECT 19.600 39.665 31.265 40.130 ;
        POLYGON 31.265 40.600 32.200 39.665 31.265 39.665 ;
        RECT 19.600 39.200 24.265 39.665 ;
        POLYGON 24.265 39.665 24.730 39.665 24.265 39.200 ;
        RECT 26.130 39.200 32.200 39.665 ;
        RECT 19.600 38.730 22.375 39.200 ;
        RECT 7.930 37.330 11.665 38.730 ;
        POLYGON 7.930 37.330 8.400 37.330 8.400 36.865 ;
        RECT 8.400 35.930 11.200 37.330 ;
        POLYGON 11.200 37.330 11.665 37.330 11.200 36.865 ;
        POLYGON 19.600 38.730 21.310 38.730 21.310 37.020 ;
        RECT 21.310 37.020 22.375 38.730 ;
        POLYGON 22.375 39.200 23.100 39.200 22.375 38.475 ;
        RECT 26.130 36.630 27.530 39.200 ;
        POLYGON 29.865 39.200 30.800 39.200 30.800 38.265 ;
        RECT 30.800 38.265 32.200 39.200 ;
        POLYGON 46.665 40.130 46.665 38.730 45.265 38.730 ;
        RECT 46.665 38.730 47.730 40.130 ;
        POLYGON 45.265 38.730 45.265 38.265 44.800 38.265 ;
        POLYGON 44.800 38.265 44.800 37.330 43.865 37.330 ;
        RECT 44.800 37.330 45.265 38.265 ;
        POLYGON 43.865 37.330 43.865 36.630 43.165 36.630 ;
        RECT 43.865 36.630 45.265 37.330 ;
        POLYGON 45.265 38.730 47.130 38.730 45.265 36.865 ;
        RECT 26.130 36.400 35.465 36.630 ;
        POLYGON 24.730 36.400 24.730 35.930 24.265 35.930 ;
        RECT 24.730 35.930 35.465 36.400 ;
        RECT 9.330 34.765 10.500 35.930 ;
        RECT 20.530 35.465 35.465 35.930 ;
        POLYGON 43.165 36.630 43.165 35.465 42.000 35.465 ;
        RECT 43.165 36.400 45.265 36.630 ;
        RECT 43.165 35.465 44.800 36.400 ;
        POLYGON 44.800 36.400 45.265 36.400 44.800 35.930 ;
        POLYGON 20.530 35.000 20.530 34.770 20.300 34.770 ;
        RECT 20.530 34.770 33.130 35.465 ;
        RECT 9.330 34.530 14.465 34.765 ;
        POLYGON 20.300 34.765 20.300 34.530 20.065 34.530 ;
        RECT 20.300 34.530 33.130 34.770 ;
        POLYGON 33.130 35.465 34.065 35.465 33.130 34.530 ;
        POLYGON 42.000 35.465 42.000 35.000 41.535 35.000 ;
        RECT 42.000 35.000 44.800 35.465 ;
        POLYGON 6.065 34.530 6.065 34.065 5.600 34.065 ;
        RECT 6.065 34.065 14.465 34.530 ;
        RECT 2.800 33.600 14.465 34.065 ;
        POLYGON 19.600 34.530 19.600 33.600 18.670 33.600 ;
        RECT 19.600 33.600 33.130 34.530 ;
        POLYGON 2.800 33.130 2.800 30.800 0.465 30.800 ;
        RECT 2.800 31.265 12.600 33.600 ;
        POLYGON 12.600 33.600 13.065 33.600 12.600 33.130 ;
        POLYGON 18.670 33.600 18.670 33.130 18.200 33.130 ;
        RECT 18.670 33.130 31.730 33.600 ;
        RECT 2.800 30.800 12.130 31.265 ;
        POLYGON 12.130 31.265 12.600 31.265 12.130 30.800 ;
        POLYGON 18.200 33.130 18.200 30.800 15.865 30.800 ;
        RECT 18.200 30.800 31.730 33.130 ;
        POLYGON 31.730 33.600 33.130 33.600 31.730 32.200 ;
        RECT 38.030 33.365 39.200 35.000 ;
        POLYGON 41.535 35.000 41.535 34.065 40.600 34.065 ;
        RECT 41.535 34.065 44.330 35.000 ;
        POLYGON 44.330 35.000 44.800 35.000 44.330 34.530 ;
        POLYGON 40.600 33.600 40.600 33.365 40.365 33.365 ;
        RECT 40.600 33.365 44.330 34.065 ;
        RECT 38.030 32.665 44.330 33.365 ;
        POLYGON 0.465 29.400 0.465 28.930 0.000 28.930 ;
        RECT 0.465 28.930 12.130 30.800 ;
        RECT 0.000 27.065 12.130 28.930 ;
        POLYGON 15.865 30.330 15.865 28.465 14.000 28.465 ;
        RECT 15.865 28.465 31.265 30.800 ;
        POLYGON 31.265 30.800 31.730 30.800 31.265 30.330 ;
        POLYGON 38.030 31.265 38.030 30.800 37.565 30.800 ;
        RECT 38.030 30.800 43.865 32.665 ;
        POLYGON 43.865 32.665 44.330 32.665 43.865 32.200 ;
        POLYGON 37.565 30.565 37.565 30.330 37.330 30.330 ;
        RECT 37.565 30.330 43.865 30.800 ;
        POLYGON 12.130 27.530 12.600 27.065 12.130 27.065 ;
        RECT 0.000 24.730 12.600 27.065 ;
        POLYGON 0.000 24.730 0.465 24.730 0.465 24.265 ;
        RECT 0.465 22.865 12.600 24.730 ;
        POLYGON 0.465 22.865 1.165 22.865 1.165 22.165 ;
        RECT 1.165 22.400 12.600 22.865 ;
        POLYGON 14.000 26.600 14.000 26.365 13.765 26.365 ;
        RECT 14.000 26.365 31.265 28.465 ;
        RECT 13.765 22.865 31.265 26.365 ;
        POLYGON 37.330 29.865 37.330 27.065 34.530 27.065 ;
        RECT 37.330 27.065 43.400 30.330 ;
        POLYGON 43.400 30.330 43.865 30.330 43.400 29.865 ;
        POLYGON 34.530 26.130 34.530 25.200 33.600 25.200 ;
        RECT 34.530 25.200 43.400 27.065 ;
        POLYGON 33.600 24.965 33.600 24.265 32.900 24.265 ;
        RECT 33.600 24.265 43.400 25.200 ;
        POLYGON 32.900 23.330 32.900 22.865 32.430 22.865 ;
        RECT 32.900 22.865 43.400 24.265 ;
        RECT 13.765 22.400 43.400 22.865 ;
        POLYGON 43.400 22.865 43.865 22.400 43.400 22.400 ;
        RECT 1.165 22.165 6.065 22.400 ;
        RECT -3.265 21.930 -1.865 22.165 ;
        POLYGON -1.865 22.165 -1.630 21.930 -1.865 21.930 ;
        POLYGON 1.165 22.165 1.400 22.165 1.400 21.930 ;
        RECT 1.400 21.930 6.065 22.165 ;
        POLYGON 6.065 22.400 6.530 22.400 6.065 21.930 ;
        POLYGON 7.930 22.400 8.400 22.400 8.400 21.930 ;
        RECT 8.400 21.930 43.865 22.400 ;
        RECT -3.265 21.465 -1.400 21.930 ;
        POLYGON -1.400 21.930 -0.930 21.465 -1.400 21.465 ;
        POLYGON 1.400 21.930 1.865 21.930 1.865 21.465 ;
        RECT 1.865 21.465 4.665 21.930 ;
        RECT -3.265 21.000 -0.465 21.465 ;
        POLYGON -2.330 21.000 -1.730 21.000 -1.730 20.400 ;
        RECT -1.730 20.530 -0.465 21.000 ;
        POLYGON -0.465 21.465 0.465 20.530 -0.465 20.530 ;
        RECT 2.330 20.530 4.665 21.465 ;
        POLYGON 4.665 21.930 5.600 21.930 4.665 21.000 ;
        RECT 9.330 21.465 43.865 21.930 ;
        RECT -1.730 20.400 0.930 20.530 ;
        POLYGON -1.265 20.400 -0.330 20.400 -0.330 19.465 ;
        RECT -0.330 20.300 0.930 20.400 ;
        POLYGON 0.930 20.530 1.165 20.300 0.930 20.300 ;
        RECT 2.330 20.300 4.430 20.530 ;
        POLYGON 4.430 20.530 4.665 20.530 4.430 20.300 ;
        RECT -0.330 19.465 4.430 20.300 ;
        POLYGON 0.130 19.465 0.465 19.465 0.465 19.130 ;
        RECT 0.465 19.130 4.430 19.465 ;
        POLYGON 0.930 19.130 1.400 19.130 1.400 18.665 ;
        RECT 1.400 18.665 7.200 19.130 ;
        POLYGON 1.865 18.665 2.330 18.665 2.330 18.200 ;
        RECT 2.330 18.200 7.200 18.665 ;
        POLYGON 7.200 19.130 8.130 18.200 7.200 18.200 ;
        RECT 9.330 18.200 10.730 21.465 ;
        POLYGON 11.930 21.465 12.400 21.465 12.400 21.000 ;
        RECT 12.400 21.000 43.865 21.465 ;
        POLYGON 12.600 21.000 13.530 21.000 13.530 20.065 ;
        RECT 13.530 20.065 43.865 21.000 ;
        RECT 2.330 17.265 10.730 18.200 ;
        RECT 13.530 19.600 35.000 20.065 ;
        POLYGON 35.000 20.065 35.465 20.065 35.000 19.600 ;
        RECT 13.530 19.130 33.600 19.600 ;
        POLYGON 33.600 19.600 34.065 19.600 33.600 19.130 ;
        POLYGON 13.530 19.130 15.400 19.130 15.400 17.265 ;
        RECT 15.400 17.400 33.600 19.130 ;
        POLYGON 33.600 18.330 34.530 17.400 33.600 17.400 ;
        RECT 15.400 17.265 34.530 17.400 ;
        RECT 3.265 16.800 10.730 17.265 ;
        POLYGON 10.730 17.265 11.200 16.800 10.730 16.800 ;
        RECT 15.400 16.800 23.800 17.265 ;
        POLYGON 23.800 17.265 24.265 17.265 23.800 16.800 ;
        POLYGON 25.665 17.265 26.130 17.265 26.130 16.800 ;
        RECT 26.130 16.800 34.530 17.265 ;
        POLYGON 3.265 16.800 3.730 16.800 3.730 16.330 ;
        RECT 3.730 16.330 12.130 16.800 ;
        POLYGON 12.130 16.800 12.600 16.330 12.130 16.330 ;
        POLYGON 4.665 16.330 7.465 16.330 7.465 13.530 ;
        RECT 7.465 12.600 14.000 16.330 ;
        RECT 15.400 15.865 20.065 16.800 ;
        POLYGON 20.065 16.800 20.530 16.800 20.065 16.330 ;
        POLYGON 15.400 15.865 16.800 15.865 16.800 14.465 ;
        RECT 16.800 14.465 18.665 15.865 ;
        POLYGON 18.665 15.865 20.065 15.865 18.665 14.465 ;
        RECT 26.600 15.865 34.530 16.800 ;
        POLYGON 14.000 14.465 15.865 12.600 14.000 12.600 ;
        POLYGON 16.800 14.465 17.265 14.465 17.265 14.000 ;
        RECT 17.265 12.600 18.665 14.465 ;
        POLYGON 7.465 12.130 7.465 11.665 7.000 11.665 ;
        RECT 7.465 11.665 18.665 12.600 ;
        RECT 7.000 11.200 18.665 11.665 ;
        POLYGON 18.665 12.600 20.065 11.200 18.665 11.200 ;
        RECT 7.000 10.730 21.000 11.200 ;
        POLYGON 21.000 11.200 21.465 10.730 21.000 10.730 ;
        RECT 7.000 10.265 22.865 10.730 ;
        POLYGON 22.865 10.730 23.330 10.265 22.865 10.265 ;
        RECT 26.600 10.265 28.465 15.865 ;
        POLYGON 29.865 15.865 30.330 15.865 30.330 15.400 ;
        RECT 30.330 15.400 34.530 15.865 ;
        POLYGON 34.530 16.800 35.930 15.400 34.530 15.400 ;
        POLYGON 32.200 15.400 33.130 15.400 33.130 14.465 ;
        RECT 33.130 14.930 35.930 15.400 ;
        RECT 37.800 14.930 39.200 20.065 ;
        POLYGON 40.600 20.065 41.065 20.065 41.065 19.600 ;
        RECT 41.065 19.600 43.865 20.065 ;
        POLYGON 43.865 20.530 44.800 19.600 43.865 19.600 ;
        POLYGON 41.865 19.600 43.730 19.600 43.730 17.730 ;
        RECT 43.730 17.730 44.800 19.600 ;
        POLYGON 42.465 16.330 42.465 15.400 41.530 15.400 ;
        RECT 42.465 15.865 46.665 16.330 ;
        POLYGON 46.665 16.330 47.130 15.865 46.665 15.865 ;
        RECT 42.465 15.400 47.130 15.865 ;
        POLYGON 41.065 15.400 41.065 14.930 40.600 14.930 ;
        RECT 41.065 14.930 47.130 15.400 ;
        RECT 33.130 14.700 47.130 14.930 ;
        RECT 33.130 14.465 46.665 14.700 ;
        POLYGON 34.530 14.465 35.465 14.465 35.465 13.530 ;
        RECT 35.465 13.530 46.665 14.465 ;
        RECT 35.465 12.365 49.465 13.530 ;
        RECT 35.465 12.130 47.130 12.365 ;
        POLYGON 34.065 12.130 34.065 10.265 32.200 10.265 ;
        RECT 34.065 11.665 47.130 12.130 ;
        RECT 34.065 10.265 46.665 11.665 ;
        POLYGON 46.665 11.665 47.130 11.665 46.665 11.200 ;
        RECT 7.000 9.330 46.665 10.265 ;
        RECT 7.000 8.865 19.830 9.330 ;
        POLYGON 7.000 8.865 7.465 8.865 7.465 8.400 ;
        RECT 7.465 7.930 19.830 8.865 ;
        RECT 21.000 8.865 46.665 9.330 ;
        RECT 21.000 7.930 22.630 8.865 ;
        RECT 7.465 7.465 22.630 7.930 ;
        RECT 23.800 8.400 45.730 8.865 ;
        POLYGON 45.730 8.865 46.200 8.865 45.730 8.400 ;
        RECT 23.800 7.465 25.665 8.400 ;
        RECT 7.465 7.000 25.665 7.465 ;
        RECT 26.830 7.000 28.465 8.400 ;
        RECT 29.630 7.000 31.265 8.400 ;
        RECT 32.430 7.000 45.730 8.400 ;
        RECT 7.465 6.530 45.730 7.000 ;
        POLYGON 7.465 6.530 7.930 6.530 7.930 6.065 ;
        RECT 7.930 5.130 45.265 6.530 ;
        POLYGON 45.265 6.530 45.730 6.530 45.265 6.065 ;
        POLYGON 7.930 5.130 8.400 5.130 8.400 4.665 ;
        RECT 8.400 4.200 43.865 5.130 ;
        POLYGON 8.400 4.200 9.800 4.200 9.800 2.800 ;
        RECT 9.800 2.330 43.865 4.200 ;
        POLYGON 43.865 5.130 45.265 5.130 43.865 3.730 ;
        POLYGON 9.800 2.330 10.265 2.330 10.265 1.865 ;
        RECT 10.265 1.865 43.865 2.330 ;
  END
END caravel_logo
END LIBRARY

