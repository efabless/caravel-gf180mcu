// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none
module chip_io(
`ifdef USE_POWER_PINS
	// Power buses
	inout  vss,	// Common padframe/ESD 5.0V ground
	inout  vdd,	// Management padframe/ESD 5.0V supply
`endif

	inout  gpio,
	input  clock,
	input  resetb,
	output flash_csb,
	output flash_clk,
	inout  flash_io0,
	inout  flash_io1,

	// Chip Core Interface
	output resetb_core,
	output clock_core,
	output gpio_in_core,
	input  gpio_out_core,
	input  gpio_outen_core,
	input  gpio_inen_core,
	input  gpio_pu_select,
	input  gpio_pd_select,
	input  gpio_schmitt_select,
	input  gpio_slew_select,
	input  [1:0] gpio_drive_select_core,
	input  flash_csb_core,
	input  flash_clk_core,
	input  flash_csb_oe_core,
	input  flash_clk_oe_core,
	input  flash_io0_oe_core,
	input  flash_io1_oe_core,
	input  flash_io0_ie_core,
	input  flash_io1_ie_core,
	input  flash_io0_do_core,
	input  flash_io1_do_core,
	output flash_io0_di_core,
	output flash_io1_di_core,

	// Constant value inputs for fixed GPIO configuration
	input [5:0] const_zero,
	input [1:0] const_one,

	// User project IOs
	inout [`MPRJ_IO_PADS-1:0] mprj_io,
	input [`MPRJ_IO_PADS-1:0] mprj_io_out,
	input [`MPRJ_IO_PADS-1:0] mprj_io_outen,
	input [`MPRJ_IO_PADS-1:0] mprj_io_inen,
	input [`MPRJ_IO_PADS-1:0] mprj_io_schmitt_select,
	input [`MPRJ_IO_PADS-1:0] mprj_io_slew_select,
	input [`MPRJ_IO_PADS-1:0] mprj_io_pu_select,
	input [`MPRJ_IO_PADS-1:0] mprj_io_pd_select,
	input [`MPRJ_IO_PADS*2-1:0] mprj_io_drive_sel,
	output [`MPRJ_IO_PADS-1:0] mprj_io_in
);

	// Instantiate power and ground pads for management domain
	// 12 pads:  vddio, vssio, vdda, vssa, vccd, vssd correspond
	// to names used with sky130, with multiple voltages for each
	// domain.  The instance names reflect where these pads
	// match the position of corresponding pads on the sky130
	// caravel, but note that there is actually only one
	// 5V supply, VDD and one common ground, VSS.

	// NOTE:  Global Foundries only supplies two pads, DVDD and
	// DVSS for 5V.  Only 5V digital cells are available for this
	// process.  Therefore, all power supplies are on the 5V
	// domain.  The VDD breaker cell divides VDD domains;
	// however, all VSS domains are tied together.

    	gf180mcu_fd_io__dvdd mgmt_vddio_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

	// lies in user area---Does not belong to management domain
	// like it does on the Sky130 version.
    	gf180mcu_fd_io__dvdd mgmt_vddio_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd mgmt_vdda_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd mgmt_vccd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssio_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssio_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssa_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

	// Instantiate power and ground pads for user 1 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	gf180mcu_fd_io__dvdd user1_vdda_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

		gf180mcu_fd_io__dvdd user1_vdda_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd user1_vccd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvss user1_vssa_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);


    	gf180mcu_fd_io__dvss user1_vssa_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss user1_vssd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

	// Instantiate power and ground pads for user 2 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	gf180mcu_fd_io__dvdd user2_vdda_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd user2_vccd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvss user2_vssa_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss user2_vssd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

	// Management clock input pad
	gf180mcu_fd_io__in_c mgmt_clock_input_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PU(const_zero[4]),
		.PD(const_zero[4]),
		.PAD(clock),
		.Y(clock_core)
	);

	// Management GPIO pad
	gf180mcu_fd_io__bi_t mgmt_gpio_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(gpio),
		.CS(gpio_schmitt_select),
		.SL(gpio_slew_select),
		.IE(gpio_inen_core),
		.OE(gpio_outen_core),
		.PU(gpio_pu_select),
		.PD(gpio_pd_select),
		.PDRV0(gpio_drive_select_core[0]),
		.PDRV1(gpio_drive_select_core[1]),
		.A(gpio_out_core),
		.Y(gpio_in_core)
	);

	// Management Flash SPI pads
	gf180mcu_fd_io__bi_t flash_io0_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_io0),
		.CS(const_zero[1]),
		.SL(const_zero[1]),
		.IE(flash_io0_ie_core),
		.OE(flash_io0_oe_core),
		.PU(const_zero[1]),
		.PD(const_zero[1]),
		.PDRV0(const_zero[1]),
		.PDRV1(const_zero[1]),
		.A(flash_io0_do_core),
		.Y(flash_io0_di_core)
	);
	
	gf180mcu_fd_io__bi_t flash_io1_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_io1),
		.CS(const_zero[0]),
		.SL(const_zero[0]),
		.IE(flash_io1_ie_core),
		.OE(flash_io1_oe_core),
		.PU(const_zero[0]),
		.PD(const_zero[0]),
		.PDRV0(const_zero[0]),
		.PDRV1(const_zero[0]),
		.A(flash_io1_do_core),
		.Y(flash_io1_di_core)
	);

	gf180mcu_fd_io__bi_t flash_csb_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_csb),
		.CS(const_zero[3]),
		.SL(const_zero[3]),
		.IE(const_zero[3]),
		.OE(flash_csb_oe_core),
		.PU(const_one[1]),
		.PD(const_zero[3]),
		.PDRV0(const_zero[3]),
		.PDRV1(const_zero[3]),
		.A(flash_csb_core),
		.Y()
	);

	gf180mcu_fd_io__bi_t flash_clk_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_clk),
		.CS(const_zero[2]),
		.SL(const_zero[2]),
		.IE(const_zero[2]),
		.OE(flash_clk_oe_core),
		.PU(const_zero[2]),
		.PD(const_zero[2]),
		.PDRV0(const_zero[2]),
		.PDRV1(const_zero[2]),
		.A(flash_clk_core),
		.Y()
	);

	// NOTE:  Resetb is active low and is configured as a pull-up

	gf180mcu_fd_io__in_s resetb_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PU(const_one[0]),
		.PD(const_zero[5]),
		.PAD(resetb),
		.Y(resetb_core)
	);

	// Corner cells (These are overlay cells;  it is not clear what is normally
    	// supposed to go under them.)

	gf180mcu_fd_io__cor mgmt_corner [1:0] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	);

	gf180mcu_fd_io__cor user1_corner (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
    	);

	gf180mcu_fd_io__cor user2_corner (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
    	);

	// generated by running ./scripts/update_chip_io_rtl.py then copying ./scripts/chip_io.txt and pasting here
	gf180mcu_fd_io__bi_t mprj_pads[0] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[0]),
		.CS(mprj_io_schmitt_select[0]),
		.SL(mprj_io_slew_select[0]),
		.IE(mprj_io_inen[0]),
		.OE(mprj_io_outen[0]),
		.PU(mprj_io_pu_select[0]),
		.PD(mprj_io_pd_select[0]),
		.PDRV0(mprj_io_drive_sel[0]),
		.PDRV1(mprj_io_drive_sel[1]),
		.A(mprj_io_out[0]),
		.Y(mprj_io_in[0]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[1] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[1]),
		.CS(mprj_io_schmitt_select[1]),
		.SL(mprj_io_slew_select[1]),
		.IE(mprj_io_inen[1]),
		.OE(mprj_io_outen[1]),
		.PU(mprj_io_pu_select[1]),
		.PD(mprj_io_pd_select[1]),
		.PDRV0(mprj_io_drive_sel[2]),
		.PDRV1(mprj_io_drive_sel[3]),
		.A(mprj_io_out[1]),
		.Y(mprj_io_in[1]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[2] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[2]),
		.CS(mprj_io_schmitt_select[2]),
		.SL(mprj_io_slew_select[2]),
		.IE(mprj_io_inen[2]),
		.OE(mprj_io_outen[2]),
		.PU(mprj_io_pu_select[2]),
		.PD(mprj_io_pd_select[2]),
		.PDRV0(mprj_io_drive_sel[4]),
		.PDRV1(mprj_io_drive_sel[5]),
		.A(mprj_io_out[2]),
		.Y(mprj_io_in[2]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[3] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[3]),
		.CS(mprj_io_schmitt_select[3]),
		.SL(mprj_io_slew_select[3]),
		.IE(mprj_io_inen[3]),
		.OE(mprj_io_outen[3]),
		.PU(mprj_io_pu_select[3]),
		.PD(mprj_io_pd_select[3]),
		.PDRV0(mprj_io_drive_sel[6]),
		.PDRV1(mprj_io_drive_sel[7]),
		.A(mprj_io_out[3]),
		.Y(mprj_io_in[3]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[4] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[4]),
		.CS(mprj_io_schmitt_select[4]),
		.SL(mprj_io_slew_select[4]),
		.IE(mprj_io_inen[4]),
		.OE(mprj_io_outen[4]),
		.PU(mprj_io_pu_select[4]),
		.PD(mprj_io_pd_select[4]),
		.PDRV0(mprj_io_drive_sel[8]),
		.PDRV1(mprj_io_drive_sel[9]),
		.A(mprj_io_out[4]),
		.Y(mprj_io_in[4]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[5] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[5]),
		.CS(mprj_io_schmitt_select[5]),
		.SL(mprj_io_slew_select[5]),
		.IE(mprj_io_inen[5]),
		.OE(mprj_io_outen[5]),
		.PU(mprj_io_pu_select[5]),
		.PD(mprj_io_pd_select[5]),
		.PDRV0(mprj_io_drive_sel[10]),
		.PDRV1(mprj_io_drive_sel[11]),
		.A(mprj_io_out[5]),
		.Y(mprj_io_in[5]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[6] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[6]),
		.CS(mprj_io_schmitt_select[6]),
		.SL(mprj_io_slew_select[6]),
		.IE(mprj_io_inen[6]),
		.OE(mprj_io_outen[6]),
		.PU(mprj_io_pu_select[6]),
		.PD(mprj_io_pd_select[6]),
		.PDRV0(mprj_io_drive_sel[12]),
		.PDRV1(mprj_io_drive_sel[13]),
		.A(mprj_io_out[6]),
		.Y(mprj_io_in[6]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[7] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[7]),
		.CS(mprj_io_schmitt_select[7]),
		.SL(mprj_io_slew_select[7]),
		.IE(mprj_io_inen[7]),
		.OE(mprj_io_outen[7]),
		.PU(mprj_io_pu_select[7]),
		.PD(mprj_io_pd_select[7]),
		.PDRV0(mprj_io_drive_sel[14]),
		.PDRV1(mprj_io_drive_sel[15]),
		.A(mprj_io_out[7]),
		.Y(mprj_io_in[7]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[8] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[8]),
		.CS(mprj_io_schmitt_select[8]),
		.SL(mprj_io_slew_select[8]),
		.IE(mprj_io_inen[8]),
		.OE(mprj_io_outen[8]),
		.PU(mprj_io_pu_select[8]),
		.PD(mprj_io_pd_select[8]),
		.PDRV0(mprj_io_drive_sel[16]),
		.PDRV1(mprj_io_drive_sel[17]),
		.A(mprj_io_out[8]),
		.Y(mprj_io_in[8]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[9] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[9]),
		.CS(mprj_io_schmitt_select[9]),
		.SL(mprj_io_slew_select[9]),
		.IE(mprj_io_inen[9]),
		.OE(mprj_io_outen[9]),
		.PU(mprj_io_pu_select[9]),
		.PD(mprj_io_pd_select[9]),
		.PDRV0(mprj_io_drive_sel[18]),
		.PDRV1(mprj_io_drive_sel[19]),
		.A(mprj_io_out[9]),
		.Y(mprj_io_in[9]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[10] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[10]),
		.CS(mprj_io_schmitt_select[10]),
		.SL(mprj_io_slew_select[10]),
		.IE(mprj_io_inen[10]),
		.OE(mprj_io_outen[10]),
		.PU(mprj_io_pu_select[10]),
		.PD(mprj_io_pd_select[10]),
		.PDRV0(mprj_io_drive_sel[20]),
		.PDRV1(mprj_io_drive_sel[21]),
		.A(mprj_io_out[10]),
		.Y(mprj_io_in[10]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[11] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[11]),
		.CS(mprj_io_schmitt_select[11]),
		.SL(mprj_io_slew_select[11]),
		.IE(mprj_io_inen[11]),
		.OE(mprj_io_outen[11]),
		.PU(mprj_io_pu_select[11]),
		.PD(mprj_io_pd_select[11]),
		.PDRV0(mprj_io_drive_sel[22]),
		.PDRV1(mprj_io_drive_sel[23]),
		.A(mprj_io_out[11]),
		.Y(mprj_io_in[11]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[12] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[12]),
		.CS(mprj_io_schmitt_select[12]),
		.SL(mprj_io_slew_select[12]),
		.IE(mprj_io_inen[12]),
		.OE(mprj_io_outen[12]),
		.PU(mprj_io_pu_select[12]),
		.PD(mprj_io_pd_select[12]),
		.PDRV0(mprj_io_drive_sel[24]),
		.PDRV1(mprj_io_drive_sel[25]),
		.A(mprj_io_out[12]),
		.Y(mprj_io_in[12]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[13] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[13]),
		.CS(mprj_io_schmitt_select[13]),
		.SL(mprj_io_slew_select[13]),
		.IE(mprj_io_inen[13]),
		.OE(mprj_io_outen[13]),
		.PU(mprj_io_pu_select[13]),
		.PD(mprj_io_pd_select[13]),
		.PDRV0(mprj_io_drive_sel[26]),
		.PDRV1(mprj_io_drive_sel[27]),
		.A(mprj_io_out[13]),
		.Y(mprj_io_in[13]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[14] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[14]),
		.CS(mprj_io_schmitt_select[14]),
		.SL(mprj_io_slew_select[14]),
		.IE(mprj_io_inen[14]),
		.OE(mprj_io_outen[14]),
		.PU(mprj_io_pu_select[14]),
		.PD(mprj_io_pd_select[14]),
		.PDRV0(mprj_io_drive_sel[28]),
		.PDRV1(mprj_io_drive_sel[29]),
		.A(mprj_io_out[14]),
		.Y(mprj_io_in[14]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[15] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[15]),
		.CS(mprj_io_schmitt_select[15]),
		.SL(mprj_io_slew_select[15]),
		.IE(mprj_io_inen[15]),
		.OE(mprj_io_outen[15]),
		.PU(mprj_io_pu_select[15]),
		.PD(mprj_io_pd_select[15]),
		.PDRV0(mprj_io_drive_sel[30]),
		.PDRV1(mprj_io_drive_sel[31]),
		.A(mprj_io_out[15]),
		.Y(mprj_io_in[15]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[16] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[16]),
		.CS(mprj_io_schmitt_select[16]),
		.SL(mprj_io_slew_select[16]),
		.IE(mprj_io_inen[16]),
		.OE(mprj_io_outen[16]),
		.PU(mprj_io_pu_select[16]),
		.PD(mprj_io_pd_select[16]),
		.PDRV0(mprj_io_drive_sel[32]),
		.PDRV1(mprj_io_drive_sel[33]),
		.A(mprj_io_out[16]),
		.Y(mprj_io_in[16]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[17] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[17]),
		.CS(mprj_io_schmitt_select[17]),
		.SL(mprj_io_slew_select[17]),
		.IE(mprj_io_inen[17]),
		.OE(mprj_io_outen[17]),
		.PU(mprj_io_pu_select[17]),
		.PD(mprj_io_pd_select[17]),
		.PDRV0(mprj_io_drive_sel[34]),
		.PDRV1(mprj_io_drive_sel[35]),
		.A(mprj_io_out[17]),
		.Y(mprj_io_in[17]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[18] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[18]),
		.CS(mprj_io_schmitt_select[18]),
		.SL(mprj_io_slew_select[18]),
		.IE(mprj_io_inen[18]),
		.OE(mprj_io_outen[18]),
		.PU(mprj_io_pu_select[18]),
		.PD(mprj_io_pd_select[18]),
		.PDRV0(mprj_io_drive_sel[36]),
		.PDRV1(mprj_io_drive_sel[37]),
		.A(mprj_io_out[18]),
		.Y(mprj_io_in[18]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[19] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[19]),
		.CS(mprj_io_schmitt_select[19]),
		.SL(mprj_io_slew_select[19]),
		.IE(mprj_io_inen[19]),
		.OE(mprj_io_outen[19]),
		.PU(mprj_io_pu_select[19]),
		.PD(mprj_io_pd_select[19]),
		.PDRV0(mprj_io_drive_sel[38]),
		.PDRV1(mprj_io_drive_sel[39]),
		.A(mprj_io_out[19]),
		.Y(mprj_io_in[19]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[20] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[20]),
		.CS(mprj_io_schmitt_select[20]),
		.SL(mprj_io_slew_select[20]),
		.IE(mprj_io_inen[20]),
		.OE(mprj_io_outen[20]),
		.PU(mprj_io_pu_select[20]),
		.PD(mprj_io_pd_select[20]),
		.PDRV0(mprj_io_drive_sel[40]),
		.PDRV1(mprj_io_drive_sel[41]),
		.A(mprj_io_out[20]),
		.Y(mprj_io_in[20]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[21] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[21]),
		.CS(mprj_io_schmitt_select[21]),
		.SL(mprj_io_slew_select[21]),
		.IE(mprj_io_inen[21]),
		.OE(mprj_io_outen[21]),
		.PU(mprj_io_pu_select[21]),
		.PD(mprj_io_pd_select[21]),
		.PDRV0(mprj_io_drive_sel[42]),
		.PDRV1(mprj_io_drive_sel[43]),
		.A(mprj_io_out[21]),
		.Y(mprj_io_in[21]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[22] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[22]),
		.CS(mprj_io_schmitt_select[22]),
		.SL(mprj_io_slew_select[22]),
		.IE(mprj_io_inen[22]),
		.OE(mprj_io_outen[22]),
		.PU(mprj_io_pu_select[22]),
		.PD(mprj_io_pd_select[22]),
		.PDRV0(mprj_io_drive_sel[44]),
		.PDRV1(mprj_io_drive_sel[45]),
		.A(mprj_io_out[22]),
		.Y(mprj_io_in[22]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[23] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[23]),
		.CS(mprj_io_schmitt_select[23]),
		.SL(mprj_io_slew_select[23]),
		.IE(mprj_io_inen[23]),
		.OE(mprj_io_outen[23]),
		.PU(mprj_io_pu_select[23]),
		.PD(mprj_io_pd_select[23]),
		.PDRV0(mprj_io_drive_sel[46]),
		.PDRV1(mprj_io_drive_sel[47]),
		.A(mprj_io_out[23]),
		.Y(mprj_io_in[23]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[24] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[24]),
		.CS(mprj_io_schmitt_select[24]),
		.SL(mprj_io_slew_select[24]),
		.IE(mprj_io_inen[24]),
		.OE(mprj_io_outen[24]),
		.PU(mprj_io_pu_select[24]),
		.PD(mprj_io_pd_select[24]),
		.PDRV0(mprj_io_drive_sel[48]),
		.PDRV1(mprj_io_drive_sel[49]),
		.A(mprj_io_out[24]),
		.Y(mprj_io_in[24]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[25] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[25]),
		.CS(mprj_io_schmitt_select[25]),
		.SL(mprj_io_slew_select[25]),
		.IE(mprj_io_inen[25]),
		.OE(mprj_io_outen[25]),
		.PU(mprj_io_pu_select[25]),
		.PD(mprj_io_pd_select[25]),
		.PDRV0(mprj_io_drive_sel[50]),
		.PDRV1(mprj_io_drive_sel[51]),
		.A(mprj_io_out[25]),
		.Y(mprj_io_in[25]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[26] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[26]),
		.CS(mprj_io_schmitt_select[26]),
		.SL(mprj_io_slew_select[26]),
		.IE(mprj_io_inen[26]),
		.OE(mprj_io_outen[26]),
		.PU(mprj_io_pu_select[26]),
		.PD(mprj_io_pd_select[26]),
		.PDRV0(mprj_io_drive_sel[52]),
		.PDRV1(mprj_io_drive_sel[53]),
		.A(mprj_io_out[26]),
		.Y(mprj_io_in[26]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[27] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[27]),
		.CS(mprj_io_schmitt_select[27]),
		.SL(mprj_io_slew_select[27]),
		.IE(mprj_io_inen[27]),
		.OE(mprj_io_outen[27]),
		.PU(mprj_io_pu_select[27]),
		.PD(mprj_io_pd_select[27]),
		.PDRV0(mprj_io_drive_sel[54]),
		.PDRV1(mprj_io_drive_sel[55]),
		.A(mprj_io_out[27]),
		.Y(mprj_io_in[27]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[28] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[28]),
		.CS(mprj_io_schmitt_select[28]),
		.SL(mprj_io_slew_select[28]),
		.IE(mprj_io_inen[28]),
		.OE(mprj_io_outen[28]),
		.PU(mprj_io_pu_select[28]),
		.PD(mprj_io_pd_select[28]),
		.PDRV0(mprj_io_drive_sel[56]),
		.PDRV1(mprj_io_drive_sel[57]),
		.A(mprj_io_out[28]),
		.Y(mprj_io_in[28]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[29] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[29]),
		.CS(mprj_io_schmitt_select[29]),
		.SL(mprj_io_slew_select[29]),
		.IE(mprj_io_inen[29]),
		.OE(mprj_io_outen[29]),
		.PU(mprj_io_pu_select[29]),
		.PD(mprj_io_pd_select[29]),
		.PDRV0(mprj_io_drive_sel[58]),
		.PDRV1(mprj_io_drive_sel[59]),
		.A(mprj_io_out[29]),
		.Y(mprj_io_in[29]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[30] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[30]),
		.CS(mprj_io_schmitt_select[30]),
		.SL(mprj_io_slew_select[30]),
		.IE(mprj_io_inen[30]),
		.OE(mprj_io_outen[30]),
		.PU(mprj_io_pu_select[30]),
		.PD(mprj_io_pd_select[30]),
		.PDRV0(mprj_io_drive_sel[60]),
		.PDRV1(mprj_io_drive_sel[61]),
		.A(mprj_io_out[30]),
		.Y(mprj_io_in[30]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[31] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[31]),
		.CS(mprj_io_schmitt_select[31]),
		.SL(mprj_io_slew_select[31]),
		.IE(mprj_io_inen[31]),
		.OE(mprj_io_outen[31]),
		.PU(mprj_io_pu_select[31]),
		.PD(mprj_io_pd_select[31]),
		.PDRV0(mprj_io_drive_sel[62]),
		.PDRV1(mprj_io_drive_sel[63]),
		.A(mprj_io_out[31]),
		.Y(mprj_io_in[31]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[32] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[32]),
		.CS(mprj_io_schmitt_select[32]),
		.SL(mprj_io_slew_select[32]),
		.IE(mprj_io_inen[32]),
		.OE(mprj_io_outen[32]),
		.PU(mprj_io_pu_select[32]),
		.PD(mprj_io_pd_select[32]),
		.PDRV0(mprj_io_drive_sel[64]),
		.PDRV1(mprj_io_drive_sel[65]),
		.A(mprj_io_out[32]),
		.Y(mprj_io_in[32]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[33] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[33]),
		.CS(mprj_io_schmitt_select[33]),
		.SL(mprj_io_slew_select[33]),
		.IE(mprj_io_inen[33]),
		.OE(mprj_io_outen[33]),
		.PU(mprj_io_pu_select[33]),
		.PD(mprj_io_pd_select[33]),
		.PDRV0(mprj_io_drive_sel[66]),
		.PDRV1(mprj_io_drive_sel[67]),
		.A(mprj_io_out[33]),
		.Y(mprj_io_in[33]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[34] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[34]),
		.CS(mprj_io_schmitt_select[34]),
		.SL(mprj_io_slew_select[34]),
		.IE(mprj_io_inen[34]),
		.OE(mprj_io_outen[34]),
		.PU(mprj_io_pu_select[34]),
		.PD(mprj_io_pd_select[34]),
		.PDRV0(mprj_io_drive_sel[68]),
		.PDRV1(mprj_io_drive_sel[69]),
		.A(mprj_io_out[34]),
		.Y(mprj_io_in[34]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[35] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[35]),
		.CS(mprj_io_schmitt_select[35]),
		.SL(mprj_io_slew_select[35]),
		.IE(mprj_io_inen[35]),
		.OE(mprj_io_outen[35]),
		.PU(mprj_io_pu_select[35]),
		.PD(mprj_io_pd_select[35]),
		.PDRV0(mprj_io_drive_sel[70]),
		.PDRV1(mprj_io_drive_sel[71]),
		.A(mprj_io_out[35]),
		.Y(mprj_io_in[35]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[36] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[36]),
		.CS(mprj_io_schmitt_select[36]),
		.SL(mprj_io_slew_select[36]),
		.IE(mprj_io_inen[36]),
		.OE(mprj_io_outen[36]),
		.PU(mprj_io_pu_select[36]),
		.PD(mprj_io_pd_select[36]),
		.PDRV0(mprj_io_drive_sel[72]),
		.PDRV1(mprj_io_drive_sel[73]),
		.A(mprj_io_out[36]),
		.Y(mprj_io_in[36]),
	);
	gf180mcu_fd_io__bi_t mprj_pads[37] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(mprj_io[37]),
		.CS(mprj_io_schmitt_select[37]),
		.SL(mprj_io_slew_select[37]),
		.IE(mprj_io_inen[37]),
		.OE(mprj_io_outen[37]),
		.PU(mprj_io_pu_select[37]),
		.PD(mprj_io_pd_select[37]),
		.PDRV0(mprj_io_drive_sel[74]),
		.PDRV1(mprj_io_drive_sel[75]),
		.A(mprj_io_out[37]),
		.Y(mprj_io_in[37]),
	);
	gf180mcu_fd_io__fill5 gf180mcu_fd_io__fill5_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill5 gf180mcu_fd_io__fill5_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill5 gf180mcu_fd_io__fill5_2 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_2 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_3 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_4 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_5 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_6 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_7 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_8 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_9 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_10 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_11 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_12 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_13 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_14 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_15 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_16 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_17 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_18 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_19 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_20 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_21 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_22 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_23 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_24 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_25 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_26 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_27 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_28 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_29 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_30 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_31 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_32 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_33 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_34 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_35 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_36 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_37 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_38 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_39 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_40 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_41 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_42 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_43 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_44 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_45 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_46 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_47 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_48 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_49 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_50 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_51 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_52 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_53 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_54 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_55 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_56 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_57 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_58 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_59 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_60 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_61 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_62 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_63 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_64 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_65 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_66 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_67 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_68 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_69 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_70 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_71 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_72 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_73 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_74 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_75 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_76 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_77 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_78 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_79 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_80 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_81 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_82 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_83 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_84 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_85 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_86 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_87 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_88 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_89 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_90 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_91 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_92 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_93 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_94 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_95 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_96 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_97 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_98 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_99 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_100 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_101 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_102 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_103 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_104 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_105 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_106 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_107 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_108 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_109 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_110 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_111 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_112 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_113 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_114 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_115 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_116 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_117 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_118 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_119 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_120 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_121 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_122 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_123 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_124 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_125 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_126 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_127 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_128 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_129 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_130 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_131 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_132 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_133 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_134 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_135 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_136 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_137 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_138 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_139 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_140 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_141 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_142 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_143 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_144 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_145 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_146 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_147 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_148 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_149 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_150 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_151 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_152 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_153 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_154 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_155 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_156 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_157 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_158 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_159 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_160 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_161 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_162 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_163 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_164 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_165 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_166 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_167 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_168 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_169 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_170 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_171 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_172 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_173 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_174 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_175 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_176 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_177 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_178 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_179 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_180 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_181 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_182 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_183 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_184 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_185 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_186 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_187 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_188 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_189 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_190 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_191 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_192 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_193 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_194 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_195 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_196 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_197 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_198 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_199 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_200 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_201 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_202 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_203 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_204 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_205 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_206 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_207 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_208 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_209 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_210 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_211 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_212 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_213 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_214 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_215 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_216 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_217 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_218 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_219 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_220 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_221 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_222 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_223 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_224 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_225 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_226 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_227 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_228 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_229 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_230 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_231 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_232 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_233 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_234 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_238 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_239 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_240 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_241 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_242 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_243 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_244 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_245 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_246 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_247 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_248 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_249 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_250 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_251 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_252 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_253 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_254 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_255 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_256 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_257 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_258 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_259 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_260 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_261 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_262 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_263 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_264 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_265 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_266 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_267 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_268 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_269 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_270 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_271 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_272 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_273 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_274 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_275 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_276 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_277 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_278 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_279 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_280 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_281 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_282 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_283 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_284 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_285 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_286 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_287 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_288 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_289 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_290 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_291 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_292 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_293 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_294 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_295 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_296 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_297 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_298 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_299 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_300 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_301 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_302 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_303 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_304 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_305 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_306 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_307 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_308 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_309 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_310 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_311 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_312 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_313 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_314 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_315 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_316 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_317 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_318 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_319 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_320 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_321 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_322 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_323 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_324 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_325 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_326 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_327 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_328 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_329 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_330 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_331 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_332 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_333 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_334 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_335 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_336 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_337 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_338 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_339 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_340 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_341 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_342 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_343 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_344 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_345 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_346 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_347 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_348 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_349 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_350 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_351 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_352 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_353 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_354 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_355 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_356 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_357 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_358 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_359 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_360 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_361 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_362 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_363 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_364 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_365 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_366 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_367 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_368 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_369 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_370 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_371 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_372 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_373 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_374 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_375 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_376 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_377 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_378 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_379 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_380 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_381 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_382 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_383 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_384 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_385 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_386 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_387 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_388 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_389 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_390 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_391 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_392 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_393 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_394 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_395 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_396 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_397 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_398 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_399 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_400 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_401 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_402 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_403 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_404 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_405 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_406 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_407 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_408 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_409 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_410 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_411 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_412 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_413 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_414 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_415 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_416 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_417 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_418 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_419 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_420 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_421 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_422 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_423 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_424 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_425 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_426 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_427 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_428 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_429 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_430 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_431 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_432 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_433 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_434 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_435 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_436 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_437 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_438 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_439 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_440 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_441 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_442 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_443 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_444 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_445 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_446 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_447 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_448 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_449 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_450 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_451 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_452 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_453 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_454 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_455 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_456 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_457 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_458 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_459 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_460 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_461 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_462 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_463 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_464 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_465 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_466 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_467 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_468 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_469 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_470 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_471 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_472 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_473 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_474 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_475 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_476 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_477 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_478 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_479 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_480 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_481 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_482 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_483 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_484 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_485 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_486 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_487 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_488 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_489 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_490 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_491 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_492 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_493 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_494 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_495 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_496 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_497 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_498 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_499 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_500 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_501 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_502 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_503 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_504 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_505 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_506 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_507 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_508 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_509 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_510 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_511 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_512 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_513 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_514 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_515 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_516 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_517 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_518 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_519 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_520 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_521 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_522 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_523 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_524 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_525 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_526 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_527 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_528 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_529 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_530 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_531 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_532 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_533 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_534 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_535 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_536 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_537 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_538 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_539 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_540 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_541 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_542 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_543 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_544 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_545 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_546 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_547 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_548 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_549 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_550 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_551 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_552 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_553 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_554 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_555 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_556 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_557 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_558 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_559 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_560 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_561 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_562 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_563 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_564 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_565 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_566 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_567 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_568 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_569 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_570 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_571 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_572 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_573 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_574 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_575 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_576 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_577 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_578 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_579 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_580 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_581 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_582 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_583 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_584 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_585 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_586 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_587 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_588 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_589 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_590 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_591 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_592 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_593 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_594 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_595 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_596 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_597 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_598 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_599 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_600 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_601 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_602 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_603 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_604 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_605 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_606 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_607 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_608 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_609 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_610 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_611 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_612 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_613 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_614 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_615 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_616 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_617 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_618 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_619 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_620 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_621 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_622 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_623 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_624 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_625 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_626 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_627 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_628 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_629 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_630 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_631 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_632 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_633 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_634 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_635 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_636 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_637 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_638 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_639 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_640 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_641 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_642 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_643 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_644 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_645 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_646 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_647 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_648 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_649 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_650 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_651 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_652 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_653 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_654 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_655 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_656 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_657 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_658 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_659 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_660 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_661 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_662 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_663 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_664 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_665 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_666 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_667 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_668 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_669 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_670 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_671 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_672 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_673 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_674 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_675 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_676 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_677 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_678 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_679 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_680 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_681 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_682 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_683 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_684 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_685 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_686 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_687 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_688 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_689 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_690 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_691 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_692 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_693 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_694 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_695 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_696 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_697 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_698 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_699 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_700 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_701 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_702 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_703 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_704 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_705 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_706 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_707 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_708 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_709 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_710 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_711 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_712 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_713 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_714 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_715 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_716 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_717 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_718 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_719 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_720 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_721 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_722 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_723 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_724 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_725 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_726 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_727 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_728 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_729 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_730 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_731 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_732 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_733 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_734 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_735 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_736 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_737 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_738 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_739 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_740 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_741 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_742 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_743 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_744 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_745 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_746 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_747 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_748 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_749 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_750 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_751 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_752 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_753 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_754 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_755 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_756 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_757 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_759 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_760 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_761 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_762 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_763 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_764 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_765 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_766 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_767 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_768 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_769 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_770 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_771 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_772 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_773 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_774 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_775 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_776 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_777 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_778 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_779 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_780 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_781 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_782 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_783 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_784 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_785 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_786 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_787 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_788 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_789 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_790 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_791 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_792 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_793 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_794 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_795 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_796 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_797 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_798 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_799 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_800 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_801 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_802 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_803 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_804 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_805 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_806 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_807 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_808 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_809 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_810 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_811 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_812 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_813 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_814 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_815 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_816 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_817 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_818 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_819 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_820 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_821 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_822 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_823 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_824 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_825 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_826 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_827 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_828 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_829 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_830 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_831 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_832 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_833 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_834 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_835 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_836 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_837 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_838 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_839 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_840 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_841 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_842 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_843 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_844 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_845 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_846 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_847 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_848 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_849 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_850 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_851 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_852 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_853 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_854 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_855 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_856 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_857 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_858 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_859 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_860 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_861 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_862 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_863 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_864 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_865 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_866 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_867 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_868 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_869 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_870 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_871 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_872 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_873 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_874 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_875 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_876 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_877 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_878 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_879 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_880 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_881 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_882 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_883 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_884 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_885 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_886 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_887 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_888 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_889 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_890 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_891 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_892 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_893 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_894 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_895 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_896 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_897 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_898 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_899 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_900 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_901 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_902 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_903 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_904 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_905 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_906 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_907 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_908 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_909 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_910 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_911 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_912 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_913 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_914 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_915 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_916 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_917 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_918 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_919 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_920 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_921 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_922 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_923 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_924 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_925 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_926 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_927 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_928 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_929 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_930 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_931 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_932 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_933 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_934 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_935 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_936 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_937 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_938 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_940 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_941 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_942 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_943 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_944 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_945 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_946 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_947 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_948 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_949 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_950 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_951 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_952 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_953 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_955 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_956 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_957 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_958 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_959 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_960 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_961 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_962 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_963 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_964 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_965 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_966 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_967 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_968 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_970 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_971 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_972 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_973 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_974 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_975 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_976 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_977 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_978 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_979 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_980 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_981 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_982 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_983 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_985 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_986 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_987 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_988 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_989 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_990 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_991 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_992 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_993 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_994 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_995 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_996 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_997 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_999 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1000 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1001 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1002 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1003 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1004 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1005 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1006 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1007 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1008 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1009 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1010 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1011 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1013 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1014 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1015 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1016 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1017 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1018 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1019 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1020 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1021 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1022 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1024 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1025 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1026 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1027 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1028 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1029 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1030 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1031 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1032 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1033 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1034 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1035 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1036 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1038 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1039 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1040 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1041 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1042 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1043 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1044 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	);

endmodule
// `default_nettype wire
