magic
tech gf180mcuC
magscale 1 10
timestamp 1669743582
<< obsm1 >>
rect 578 5428 633790 870770
<< metal2 >>
rect 33752 871200 33828 872800
rect 33898 871200 33974 872800
rect 34044 871200 34120 872800
rect 34190 871200 34266 872800
rect 45647 871200 45723 872800
rect 45858 871200 45934 872800
rect 46360 871200 46436 872800
rect 46502 871200 46578 872800
rect 46731 871200 46807 872800
rect 47252 871200 47328 872800
rect 88752 871200 88828 872800
rect 88898 871200 88974 872800
rect 89044 871200 89120 872800
rect 89190 871200 89266 872800
rect 100647 871200 100723 872800
rect 100858 871200 100934 872800
rect 101360 871200 101436 872800
rect 101502 871200 101578 872800
rect 101731 871200 101807 872800
rect 102252 871200 102328 872800
rect 143752 871200 143828 872800
rect 143898 871200 143974 872800
rect 144044 871200 144120 872800
rect 144190 871200 144266 872800
rect 155647 871200 155723 872800
rect 155858 871200 155934 872800
rect 156360 871200 156436 872800
rect 156502 871200 156578 872800
rect 156731 871200 156807 872800
rect 157252 871200 157328 872800
rect 198752 871200 198828 872800
rect 198898 871200 198974 872800
rect 199044 871200 199120 872800
rect 199190 871200 199266 872800
rect 210647 871200 210723 872800
rect 210858 871200 210934 872800
rect 211360 871200 211436 872800
rect 211502 871200 211578 872800
rect 211731 871200 211807 872800
rect 212252 871200 212328 872800
rect 253752 871200 253828 872800
rect 253898 871200 253974 872800
rect 254044 871200 254120 872800
rect 254190 871200 254266 872800
rect 265647 871200 265723 872800
rect 265858 871200 265934 872800
rect 266360 871200 266436 872800
rect 266502 871200 266578 872800
rect 266731 871200 266807 872800
rect 267252 871200 267328 872800
rect 363752 871200 363828 872800
rect 363898 871200 363974 872800
rect 364044 871200 364120 872800
rect 364190 871200 364266 872800
rect 375647 871200 375723 872800
rect 375858 871200 375934 872800
rect 376360 871200 376436 872800
rect 376502 871200 376578 872800
rect 376731 871200 376807 872800
rect 377252 871200 377328 872800
rect 418752 871200 418828 872800
rect 418898 871200 418974 872800
rect 419044 871200 419120 872800
rect 419190 871200 419266 872800
rect 430647 871200 430723 872800
rect 430858 871200 430934 872800
rect 431360 871200 431436 872800
rect 431502 871200 431578 872800
rect 431731 871200 431807 872800
rect 432252 871200 432328 872800
rect 473752 871200 473828 872800
rect 473898 871200 473974 872800
rect 474044 871200 474120 872800
rect 474190 871200 474266 872800
rect 485647 871200 485723 872800
rect 485858 871200 485934 872800
rect 486360 871200 486436 872800
rect 486502 871200 486578 872800
rect 486731 871200 486807 872800
rect 487252 871200 487328 872800
rect 583752 871200 583828 872800
rect 583898 871200 583974 872800
rect 584044 871200 584120 872800
rect 584190 871200 584266 872800
rect 595647 871200 595723 872800
rect 595858 871200 595934 872800
rect 596360 871200 596436 872800
rect 596502 871200 596578 872800
rect 596731 871200 596807 872800
rect 597252 871200 597328 872800
rect 632200 849172 634800 849248
rect 632700 849026 634800 849102
rect 633200 848880 634800 848956
rect 633700 848734 634800 848810
rect -800 848252 300 848328
rect -800 847731 800 847807
rect -800 847502 1300 847578
rect -800 847360 1800 847436
rect -800 846858 2300 846934
rect -800 846647 2800 846723
rect 631200 837277 634800 837353
rect 631700 837066 634800 837142
rect 632200 836564 634800 836640
rect 632700 836422 634800 836498
rect 633200 836193 634800 836269
rect 633700 835672 634800 835748
rect -800 835190 300 835266
rect -800 835044 800 835120
rect -800 834898 1300 834974
rect -800 834752 1800 834828
rect 632200 763172 634800 763248
rect 632700 763026 634800 763102
rect 633200 762880 634800 762956
rect 633700 762734 634800 762810
rect 631200 751277 634800 751353
rect 631700 751066 634800 751142
rect 632200 750564 634800 750640
rect 632700 750422 634800 750498
rect 633200 750193 634800 750269
rect 633700 749672 634800 749748
rect -800 684252 300 684328
rect -800 683731 800 683807
rect -800 683502 1300 683578
rect -800 683360 1800 683436
rect -800 682858 2300 682934
rect -800 682647 2800 682723
rect 632200 677172 634800 677248
rect 632700 677026 634800 677102
rect 633200 676880 634800 676956
rect 633700 676734 634800 676810
rect -800 671190 300 671266
rect -800 671044 800 671120
rect -800 670898 1300 670974
rect -800 670752 1800 670828
rect 631200 665277 634800 665353
rect 631700 665066 634800 665142
rect 632200 664564 634800 664640
rect 632700 664422 634800 664498
rect 633200 664193 634800 664269
rect 633700 663672 634800 663748
rect -800 643252 300 643328
rect -800 642731 800 642807
rect -800 642502 1300 642578
rect -800 642360 1800 642436
rect -800 641858 2300 641934
rect -800 641647 2800 641723
rect 632200 634172 634800 634248
rect 632700 634026 634800 634102
rect 633200 633880 634800 633956
rect 633700 633734 634800 633810
rect -800 630190 300 630266
rect -800 630044 800 630120
rect -800 629898 1300 629974
rect -800 629752 1800 629828
rect 631200 622277 634800 622353
rect 631700 622066 634800 622142
rect 632200 621564 634800 621640
rect 632700 621422 634800 621498
rect 633200 621193 634800 621269
rect 633700 620672 634800 620748
rect -800 602252 300 602328
rect -800 601731 800 601807
rect -800 601502 1300 601578
rect -800 601360 1800 601436
rect -800 600858 2300 600934
rect -800 600647 2800 600723
rect 632200 591172 634800 591248
rect 632700 591026 634800 591102
rect 633200 590880 634800 590956
rect 633700 590734 634800 590810
rect -800 589190 300 589266
rect -800 589044 800 589120
rect -800 588898 1300 588974
rect -800 588752 1800 588828
rect 631200 579277 634800 579353
rect 631700 579066 634800 579142
rect 632200 578564 634800 578640
rect 632700 578422 634800 578498
rect 633200 578193 634800 578269
rect 633700 577672 634800 577748
rect -800 561252 300 561328
rect -800 560731 800 560807
rect -800 560502 1300 560578
rect -800 560360 1800 560436
rect -800 559858 2300 559934
rect -800 559647 2800 559723
rect -800 548190 300 548266
rect -800 548044 800 548120
rect 632200 548172 634800 548248
rect -800 547898 1300 547974
rect 632700 548026 634800 548102
rect -800 547752 1800 547828
rect 633200 547880 634800 547956
rect 633700 547734 634800 547810
rect 631200 536277 634800 536353
rect 631700 536066 634800 536142
rect 632200 535564 634800 535640
rect 632700 535422 634800 535498
rect 633200 535193 634800 535269
rect 633700 534672 634800 534748
rect -800 520252 300 520328
rect -800 519731 800 519807
rect -800 519502 1300 519578
rect -800 519360 1800 519436
rect -800 518858 2300 518934
rect -800 518647 2800 518723
rect -800 507190 300 507266
rect -800 507044 800 507120
rect -800 506898 1300 506974
rect -800 506752 1800 506828
rect 632200 505172 634800 505248
rect 632700 505026 634800 505102
rect 633200 504880 634800 504956
rect 633700 504734 634800 504810
rect 631200 493277 634800 493353
rect 631700 493066 634800 493142
rect 632200 492564 634800 492640
rect 632700 492422 634800 492498
rect 633200 492193 634800 492269
rect 633700 491672 634800 491748
rect -800 479252 300 479328
rect -800 478731 800 478807
rect -800 478502 1300 478578
rect -800 478360 1800 478436
rect -800 477858 2300 477934
rect -800 477647 2800 477723
rect -800 466190 300 466266
rect -800 466044 800 466120
rect -800 465898 1300 465974
rect -800 465752 1800 465828
rect 632200 462172 634800 462248
rect 632700 462026 634800 462102
rect 633200 461880 634800 461956
rect 633700 461734 634800 461810
rect 631200 450277 634800 450353
rect 631700 450066 634800 450142
rect 632200 449564 634800 449640
rect 632700 449422 634800 449498
rect 633200 449193 634800 449269
rect 633700 448672 634800 448748
rect -800 438252 300 438328
rect -800 437731 800 437807
rect -800 437502 1300 437578
rect -800 437360 1800 437436
rect -800 436858 2300 436934
rect -800 436647 2800 436723
rect -800 425190 300 425266
rect -800 425044 800 425120
rect -800 424898 1300 424974
rect -800 424752 1800 424828
rect -800 315252 300 315328
rect -800 314731 800 314807
rect -800 314502 1300 314578
rect -800 314360 1800 314436
rect -800 313858 2300 313934
rect -800 313647 2800 313723
rect -800 302190 300 302266
rect -800 302044 800 302120
rect -800 301898 1300 301974
rect -800 301752 1800 301828
rect 632200 290172 634800 290248
rect 632700 290026 634800 290102
rect 633200 289880 634800 289956
rect 633700 289734 634800 289810
rect 631200 278277 634800 278353
rect 631700 278066 634800 278142
rect 632200 277564 634800 277640
rect 632700 277422 634800 277498
rect 633200 277193 634800 277269
rect 633700 276672 634800 276748
rect -800 274252 300 274328
rect -800 273731 800 273807
rect -800 273502 1300 273578
rect -800 273360 1800 273436
rect -800 272858 2300 272934
rect -800 272647 2800 272723
rect -800 261190 300 261266
rect -800 261044 800 261120
rect -800 260898 1300 260974
rect -800 260752 1800 260828
rect 632200 247172 634800 247248
rect 632700 247026 634800 247102
rect 633200 246880 634800 246956
rect 633700 246734 634800 246810
rect 631200 235277 634800 235353
rect 631700 235066 634800 235142
rect 632200 234564 634800 234640
rect 632700 234422 634800 234498
rect 633200 234193 634800 234269
rect 633700 233672 634800 233748
rect -800 233252 300 233328
rect -800 232731 800 232807
rect -800 232502 1300 232578
rect -800 232360 1800 232436
rect -800 231858 2300 231934
rect -800 231647 2800 231723
rect -800 220190 300 220266
rect -800 220044 800 220120
rect -800 219898 1300 219974
rect -800 219752 1800 219828
rect 632200 204172 634800 204248
rect 632700 204026 634800 204102
rect 633200 203880 634800 203956
rect 633700 203734 634800 203810
rect -800 192252 300 192328
rect 631200 192277 634800 192353
rect 631700 192066 634800 192142
rect -800 191731 800 191807
rect -800 191502 1300 191578
rect 632200 191564 634800 191640
rect -800 191360 1800 191436
rect 632700 191422 634800 191498
rect 633200 191193 634800 191269
rect -800 190858 2300 190934
rect -800 190647 2800 190723
rect 633700 190672 634800 190748
rect -800 179190 300 179266
rect -800 179044 800 179120
rect -800 178898 1300 178974
rect -800 178752 1800 178828
rect 632200 161172 634800 161248
rect 632700 161026 634800 161102
rect 633200 160880 634800 160956
rect 633700 160734 634800 160810
rect -800 151252 300 151328
rect -800 150731 800 150807
rect -800 150502 1300 150578
rect -800 150360 1800 150436
rect -800 149858 2300 149934
rect -800 149647 2800 149723
rect 631200 149277 634800 149353
rect 631700 149066 634800 149142
rect 632200 148564 634800 148640
rect 632700 148422 634800 148498
rect 633200 148193 634800 148269
rect 633700 147672 634800 147748
rect -800 138190 300 138266
rect -800 138044 800 138120
rect -800 137898 1300 137974
rect -800 137752 1800 137828
rect 632200 118172 634800 118248
rect 632700 118026 634800 118102
rect 633200 117880 634800 117956
rect 633700 117734 634800 117810
rect -800 110252 300 110328
rect -800 109731 800 109807
rect -800 109502 1300 109578
rect -800 109360 1800 109436
rect -800 108858 2300 108934
rect -800 108647 2800 108723
rect 631200 106277 634800 106353
rect 631700 106066 634800 106142
rect 632200 105564 634800 105640
rect 632700 105422 634800 105498
rect 633200 105193 634800 105269
rect 633700 104672 634800 104748
rect -800 97190 300 97266
rect -800 97044 800 97120
rect -800 96898 1300 96974
rect -800 96752 1800 96828
rect 632200 75172 634800 75248
rect 632700 75026 634800 75102
rect 633200 74880 634800 74956
rect 633700 74734 634800 74810
rect 631200 63277 634800 63353
rect 631700 63066 634800 63142
rect 632200 62564 634800 62640
rect 632700 62422 634800 62498
rect 633200 62193 634800 62269
rect 633700 61672 634800 61748
rect 632200 32172 634800 32248
rect 632700 32026 634800 32102
rect 633200 31880 634800 31956
rect 633700 31734 634800 31810
rect 631200 20277 634800 20353
rect 631700 20066 634800 20142
rect 632200 19564 634800 19640
rect 632700 19422 634800 19498
rect 633200 19193 634800 19269
rect 633700 18672 634800 18748
rect 90193 -800 90269 800
rect 91066 -800 91142 800
rect 103172 -800 103248 800
rect 145193 -810 145269 800
rect 158172 -800 158248 800
rect 255193 -844 255269 800
rect 267733 -800 267811 800
rect 267880 -800 267956 800
rect 268026 -800 268102 800
rect 322734 -802 322810 800
rect 322880 -800 322956 800
rect 323026 -800 323102 800
rect 366277 -800 366353 800
rect 377734 -802 377810 800
rect 377880 -800 377956 800
rect 378026 -800 378102 800
rect 378171 -800 378247 800
rect 421277 -800 421353 800
rect 432734 -802 432810 800
rect 432880 -800 432956 800
rect 433026 -800 433102 800
rect 433172 -800 433248 800
rect 474672 -802 474748 800
rect 475193 -802 475269 800
rect 475422 -800 475498 800
rect 475564 -800 475640 800
rect 476066 -802 476142 800
rect 476277 -800 476353 800
rect 487734 -802 487810 800
rect 487880 -800 487956 800
rect 488026 -800 488102 800
rect 488172 -800 488248 800
<< obsm2 >>
rect 140 871140 33692 871332
rect 34326 871140 45587 871332
rect 45783 871140 45798 871332
rect 45994 871140 46300 871332
rect 46638 871140 46671 871332
rect 46867 871140 47192 871332
rect 47388 871140 88692 871332
rect 89326 871140 100587 871332
rect 100783 871140 100798 871332
rect 100994 871140 101300 871332
rect 101638 871140 101671 871332
rect 101867 871140 102192 871332
rect 102388 871140 143692 871332
rect 144326 871140 155587 871332
rect 155783 871140 155798 871332
rect 155994 871140 156300 871332
rect 156638 871140 156671 871332
rect 156867 871140 157192 871332
rect 157388 871140 198692 871332
rect 199326 871140 210587 871332
rect 210783 871140 210798 871332
rect 210994 871140 211300 871332
rect 211638 871140 211671 871332
rect 211867 871140 212192 871332
rect 212388 871140 253692 871332
rect 254326 871140 265587 871332
rect 265783 871140 265798 871332
rect 265994 871140 266300 871332
rect 266638 871140 266671 871332
rect 266867 871140 267192 871332
rect 267388 871140 363692 871332
rect 364326 871140 375587 871332
rect 375783 871140 375798 871332
rect 375994 871140 376300 871332
rect 376638 871140 376671 871332
rect 376867 871140 377192 871332
rect 377388 871140 418692 871332
rect 419326 871140 430587 871332
rect 430783 871140 430798 871332
rect 430994 871140 431300 871332
rect 431638 871140 431671 871332
rect 431867 871140 432192 871332
rect 432388 871140 473692 871332
rect 474326 871140 485587 871332
rect 485783 871140 485798 871332
rect 485994 871140 486300 871332
rect 486638 871140 486671 871332
rect 486867 871140 487192 871332
rect 487388 871140 583692 871332
rect 584326 871140 595587 871332
rect 595783 871140 595798 871332
rect 595994 871140 596300 871332
rect 596638 871140 596671 871332
rect 596867 871140 597192 871332
rect 597388 871140 633892 871332
rect 140 849308 633892 871140
rect 140 849112 632140 849308
rect 140 848966 632640 849112
rect 140 848820 633140 848966
rect 140 848674 633640 848820
rect 140 848388 633892 848674
rect 360 848192 633892 848388
rect 140 847867 633892 848192
rect 860 847671 633892 847867
rect 140 847638 633892 847671
rect 1360 847496 633892 847638
rect 1860 847300 633892 847496
rect 140 846994 633892 847300
rect 2360 846798 633892 846994
rect 140 846783 633892 846798
rect 2860 846587 633892 846783
rect 140 837413 633892 846587
rect 140 837217 631140 837413
rect 140 837202 633892 837217
rect 140 837006 631640 837202
rect 140 836700 633892 837006
rect 140 836504 632140 836700
rect 140 836362 632640 836504
rect 140 836329 633892 836362
rect 140 836133 633140 836329
rect 140 835808 633892 836133
rect 140 835612 633640 835808
rect 140 835326 633892 835612
rect 360 835180 633892 835326
rect 860 835034 633892 835180
rect 1360 834888 633892 835034
rect 1860 834692 633892 834888
rect 140 763308 633892 834692
rect 140 763112 632140 763308
rect 140 762966 632640 763112
rect 140 762820 633140 762966
rect 140 762674 633640 762820
rect 140 751413 633892 762674
rect 140 751217 631140 751413
rect 140 751202 633892 751217
rect 140 751006 631640 751202
rect 140 750700 633892 751006
rect 140 750504 632140 750700
rect 140 750362 632640 750504
rect 140 750329 633892 750362
rect 140 750133 633140 750329
rect 140 749808 633892 750133
rect 140 749612 633640 749808
rect 140 684388 633892 749612
rect 360 684192 633892 684388
rect 140 683867 633892 684192
rect 860 683671 633892 683867
rect 140 683638 633892 683671
rect 1360 683496 633892 683638
rect 1860 683300 633892 683496
rect 140 682994 633892 683300
rect 2360 682798 633892 682994
rect 140 682783 633892 682798
rect 2860 682587 633892 682783
rect 140 677308 633892 682587
rect 140 677112 632140 677308
rect 140 676966 632640 677112
rect 140 676820 633140 676966
rect 140 676674 633640 676820
rect 140 671326 633892 676674
rect 360 671180 633892 671326
rect 860 671034 633892 671180
rect 1360 670888 633892 671034
rect 1860 670692 633892 670888
rect 140 665413 633892 670692
rect 140 665217 631140 665413
rect 140 665202 633892 665217
rect 140 665006 631640 665202
rect 140 664700 633892 665006
rect 140 664504 632140 664700
rect 140 664362 632640 664504
rect 140 664329 633892 664362
rect 140 664133 633140 664329
rect 140 663808 633892 664133
rect 140 663612 633640 663808
rect 140 643388 633892 663612
rect 360 643192 633892 643388
rect 140 642867 633892 643192
rect 860 642671 633892 642867
rect 140 642638 633892 642671
rect 1360 642496 633892 642638
rect 1860 642300 633892 642496
rect 140 641994 633892 642300
rect 2360 641798 633892 641994
rect 140 641783 633892 641798
rect 2860 641587 633892 641783
rect 140 634308 633892 641587
rect 140 634112 632140 634308
rect 140 633966 632640 634112
rect 140 633820 633140 633966
rect 140 633674 633640 633820
rect 140 630326 633892 633674
rect 360 630180 633892 630326
rect 860 630034 633892 630180
rect 1360 629888 633892 630034
rect 1860 629692 633892 629888
rect 140 622413 633892 629692
rect 140 622217 631140 622413
rect 140 622202 633892 622217
rect 140 622006 631640 622202
rect 140 621700 633892 622006
rect 140 621504 632140 621700
rect 140 621362 632640 621504
rect 140 621329 633892 621362
rect 140 621133 633140 621329
rect 140 620808 633892 621133
rect 140 620612 633640 620808
rect 140 602388 633892 620612
rect 360 602192 633892 602388
rect 140 601867 633892 602192
rect 860 601671 633892 601867
rect 140 601638 633892 601671
rect 1360 601496 633892 601638
rect 1860 601300 633892 601496
rect 140 600994 633892 601300
rect 2360 600798 633892 600994
rect 140 600783 633892 600798
rect 2860 600587 633892 600783
rect 140 591308 633892 600587
rect 140 591112 632140 591308
rect 140 590966 632640 591112
rect 140 590820 633140 590966
rect 140 590674 633640 590820
rect 140 589326 633892 590674
rect 360 589180 633892 589326
rect 860 589034 633892 589180
rect 1360 588888 633892 589034
rect 1860 588692 633892 588888
rect 140 579413 633892 588692
rect 140 579217 631140 579413
rect 140 579202 633892 579217
rect 140 579006 631640 579202
rect 140 578700 633892 579006
rect 140 578504 632140 578700
rect 140 578362 632640 578504
rect 140 578329 633892 578362
rect 140 578133 633140 578329
rect 140 577808 633892 578133
rect 140 577612 633640 577808
rect 140 561388 633892 577612
rect 360 561192 633892 561388
rect 140 560867 633892 561192
rect 860 560671 633892 560867
rect 140 560638 633892 560671
rect 1360 560496 633892 560638
rect 1860 560300 633892 560496
rect 140 559994 633892 560300
rect 2360 559798 633892 559994
rect 140 559783 633892 559798
rect 2860 559587 633892 559783
rect 140 548326 633892 559587
rect 360 548308 633892 548326
rect 360 548180 632140 548308
rect 860 548112 632140 548180
rect 860 548034 632640 548112
rect 1360 547966 632640 548034
rect 1360 547888 633140 547966
rect 1860 547820 633140 547888
rect 1860 547692 633640 547820
rect 140 547674 633640 547692
rect 140 536413 633892 547674
rect 140 536217 631140 536413
rect 140 536202 633892 536217
rect 140 536006 631640 536202
rect 140 535700 633892 536006
rect 140 535504 632140 535700
rect 140 535362 632640 535504
rect 140 535329 633892 535362
rect 140 535133 633140 535329
rect 140 534808 633892 535133
rect 140 534612 633640 534808
rect 140 520388 633892 534612
rect 360 520192 633892 520388
rect 140 519867 633892 520192
rect 860 519671 633892 519867
rect 140 519638 633892 519671
rect 1360 519496 633892 519638
rect 1860 519300 633892 519496
rect 140 518994 633892 519300
rect 2360 518798 633892 518994
rect 140 518783 633892 518798
rect 2860 518587 633892 518783
rect 140 507326 633892 518587
rect 360 507180 633892 507326
rect 860 507034 633892 507180
rect 1360 506888 633892 507034
rect 1860 506692 633892 506888
rect 140 505308 633892 506692
rect 140 505112 632140 505308
rect 140 504966 632640 505112
rect 140 504820 633140 504966
rect 140 504674 633640 504820
rect 140 493413 633892 504674
rect 140 493217 631140 493413
rect 140 493202 633892 493217
rect 140 493006 631640 493202
rect 140 492700 633892 493006
rect 140 492504 632140 492700
rect 140 492362 632640 492504
rect 140 492329 633892 492362
rect 140 492133 633140 492329
rect 140 491808 633892 492133
rect 140 491612 633640 491808
rect 140 479388 633892 491612
rect 360 479192 633892 479388
rect 140 478867 633892 479192
rect 860 478671 633892 478867
rect 140 478638 633892 478671
rect 1360 478496 633892 478638
rect 1860 478300 633892 478496
rect 140 477994 633892 478300
rect 2360 477798 633892 477994
rect 140 477783 633892 477798
rect 2860 477587 633892 477783
rect 140 466326 633892 477587
rect 360 466180 633892 466326
rect 860 466034 633892 466180
rect 1360 465888 633892 466034
rect 1860 465692 633892 465888
rect 140 462308 633892 465692
rect 140 462112 632140 462308
rect 140 461966 632640 462112
rect 140 461820 633140 461966
rect 140 461674 633640 461820
rect 140 450413 633892 461674
rect 140 450217 631140 450413
rect 140 450202 633892 450217
rect 140 450006 631640 450202
rect 140 449700 633892 450006
rect 140 449504 632140 449700
rect 140 449362 632640 449504
rect 140 449329 633892 449362
rect 140 449133 633140 449329
rect 140 448808 633892 449133
rect 140 448612 633640 448808
rect 140 438388 633892 448612
rect 360 438192 633892 438388
rect 140 437867 633892 438192
rect 860 437671 633892 437867
rect 140 437638 633892 437671
rect 1360 437496 633892 437638
rect 1860 437300 633892 437496
rect 140 436994 633892 437300
rect 2360 436798 633892 436994
rect 140 436783 633892 436798
rect 2860 436587 633892 436783
rect 140 425326 633892 436587
rect 360 425180 633892 425326
rect 860 425034 633892 425180
rect 1360 424888 633892 425034
rect 1860 424692 633892 424888
rect 140 315388 633892 424692
rect 360 315192 633892 315388
rect 140 314867 633892 315192
rect 860 314671 633892 314867
rect 140 314638 633892 314671
rect 1360 314496 633892 314638
rect 1860 314300 633892 314496
rect 140 313994 633892 314300
rect 2360 313798 633892 313994
rect 140 313783 633892 313798
rect 2860 313587 633892 313783
rect 140 302326 633892 313587
rect 360 302180 633892 302326
rect 860 302034 633892 302180
rect 1360 301888 633892 302034
rect 1860 301692 633892 301888
rect 140 290308 633892 301692
rect 140 290112 632140 290308
rect 140 289966 632640 290112
rect 140 289820 633140 289966
rect 140 289674 633640 289820
rect 140 278413 633892 289674
rect 140 278217 631140 278413
rect 140 278202 633892 278217
rect 140 278006 631640 278202
rect 140 277700 633892 278006
rect 140 277504 632140 277700
rect 140 277362 632640 277504
rect 140 277329 633892 277362
rect 140 277133 633140 277329
rect 140 276808 633892 277133
rect 140 276612 633640 276808
rect 140 274388 633892 276612
rect 360 274192 633892 274388
rect 140 273867 633892 274192
rect 860 273671 633892 273867
rect 140 273638 633892 273671
rect 1360 273496 633892 273638
rect 1860 273300 633892 273496
rect 140 272994 633892 273300
rect 2360 272798 633892 272994
rect 140 272783 633892 272798
rect 2860 272587 633892 272783
rect 140 261326 633892 272587
rect 360 261180 633892 261326
rect 860 261034 633892 261180
rect 1360 260888 633892 261034
rect 1860 260692 633892 260888
rect 140 247308 633892 260692
rect 140 247112 632140 247308
rect 140 246966 632640 247112
rect 140 246820 633140 246966
rect 140 246674 633640 246820
rect 140 235413 633892 246674
rect 140 235217 631140 235413
rect 140 235202 633892 235217
rect 140 235006 631640 235202
rect 140 234700 633892 235006
rect 140 234504 632140 234700
rect 140 234362 632640 234504
rect 140 234329 633892 234362
rect 140 234133 633140 234329
rect 140 233808 633892 234133
rect 140 233612 633640 233808
rect 140 233388 633892 233612
rect 360 233192 633892 233388
rect 140 232867 633892 233192
rect 860 232671 633892 232867
rect 140 232638 633892 232671
rect 1360 232496 633892 232638
rect 1860 232300 633892 232496
rect 140 231994 633892 232300
rect 2360 231798 633892 231994
rect 140 231783 633892 231798
rect 2860 231587 633892 231783
rect 140 220326 633892 231587
rect 360 220180 633892 220326
rect 860 220034 633892 220180
rect 1360 219888 633892 220034
rect 1860 219692 633892 219888
rect 140 204308 633892 219692
rect 140 204112 632140 204308
rect 140 203966 632640 204112
rect 140 203820 633140 203966
rect 140 203674 633640 203820
rect 140 192413 633892 203674
rect 140 192388 631140 192413
rect 360 192217 631140 192388
rect 360 192202 633892 192217
rect 360 192192 631640 192202
rect 140 192006 631640 192192
rect 140 191867 633892 192006
rect 860 191700 633892 191867
rect 860 191671 632140 191700
rect 140 191638 632140 191671
rect 1360 191504 632140 191638
rect 1360 191496 632640 191504
rect 1860 191362 632640 191496
rect 1860 191329 633892 191362
rect 1860 191300 633140 191329
rect 140 191133 633140 191300
rect 140 190994 633892 191133
rect 2360 190808 633892 190994
rect 2360 190798 633640 190808
rect 140 190783 633640 190798
rect 2860 190612 633640 190783
rect 2860 190587 633892 190612
rect 140 179326 633892 190587
rect 360 179180 633892 179326
rect 860 179034 633892 179180
rect 1360 178888 633892 179034
rect 1860 178692 633892 178888
rect 140 161308 633892 178692
rect 140 161112 632140 161308
rect 140 160966 632640 161112
rect 140 160820 633140 160966
rect 140 160674 633640 160820
rect 140 151388 633892 160674
rect 360 151192 633892 151388
rect 140 150867 633892 151192
rect 860 150671 633892 150867
rect 140 150638 633892 150671
rect 1360 150496 633892 150638
rect 1860 150300 633892 150496
rect 140 149994 633892 150300
rect 2360 149798 633892 149994
rect 140 149783 633892 149798
rect 2860 149587 633892 149783
rect 140 149413 633892 149587
rect 140 149217 631140 149413
rect 140 149202 633892 149217
rect 140 149006 631640 149202
rect 140 148700 633892 149006
rect 140 148504 632140 148700
rect 140 148362 632640 148504
rect 140 148329 633892 148362
rect 140 148133 633140 148329
rect 140 147808 633892 148133
rect 140 147612 633640 147808
rect 140 138326 633892 147612
rect 360 138180 633892 138326
rect 860 138034 633892 138180
rect 1360 137888 633892 138034
rect 1860 137692 633892 137888
rect 140 118308 633892 137692
rect 140 118112 632140 118308
rect 140 117966 632640 118112
rect 140 117820 633140 117966
rect 140 117674 633640 117820
rect 140 110388 633892 117674
rect 360 110192 633892 110388
rect 140 109867 633892 110192
rect 860 109671 633892 109867
rect 140 109638 633892 109671
rect 1360 109496 633892 109638
rect 1860 109300 633892 109496
rect 140 108994 633892 109300
rect 2360 108798 633892 108994
rect 140 108783 633892 108798
rect 2860 108587 633892 108783
rect 140 106413 633892 108587
rect 140 106217 631140 106413
rect 140 106202 633892 106217
rect 140 106006 631640 106202
rect 140 105700 633892 106006
rect 140 105504 632140 105700
rect 140 105362 632640 105504
rect 140 105329 633892 105362
rect 140 105133 633140 105329
rect 140 104808 633892 105133
rect 140 104612 633640 104808
rect 140 97326 633892 104612
rect 360 97180 633892 97326
rect 860 97034 633892 97180
rect 1360 96888 633892 97034
rect 1860 96692 633892 96888
rect 140 75308 633892 96692
rect 140 75112 632140 75308
rect 140 74966 632640 75112
rect 140 74820 633140 74966
rect 140 74674 633640 74820
rect 140 63413 633892 74674
rect 140 63217 631140 63413
rect 140 63202 633892 63217
rect 140 63006 631640 63202
rect 140 62700 633892 63006
rect 140 62504 632140 62700
rect 140 62362 632640 62504
rect 140 62329 633892 62362
rect 140 62133 633140 62329
rect 140 61808 633892 62133
rect 140 61612 633640 61808
rect 140 32308 633892 61612
rect 140 32112 632140 32308
rect 140 31966 632640 32112
rect 140 31820 633140 31966
rect 140 31674 633640 31820
rect 140 20413 633892 31674
rect 140 20217 631140 20413
rect 140 20202 633892 20217
rect 140 20006 631640 20202
rect 140 19700 633892 20006
rect 140 19504 632140 19700
rect 140 19362 632640 19504
rect 140 19329 633892 19362
rect 140 19133 633140 19329
rect 140 18808 633892 19133
rect 140 18612 633640 18808
rect 140 860 633892 18612
rect 140 700 90133 860
rect 90329 700 91006 860
rect 91202 700 103112 860
rect 103308 700 145133 860
rect 145329 700 158112 860
rect 158308 700 255133 860
rect 255329 700 267673 860
rect 268162 700 322674 860
rect 323162 700 366217 860
rect 366413 700 377674 860
rect 378307 700 421217 860
rect 421413 700 432674 860
rect 433308 700 474612 860
rect 474808 700 475133 860
rect 475329 700 475362 860
rect 475700 700 476006 860
rect 476202 700 476217 860
rect 476413 700 487674 860
rect 488308 700 633892 860
<< obsm3 >>
rect 130 5068 633902 871108
<< metal4 >>
rect 416 1088 2416 870720
rect 2816 3488 4816 868320
rect 7216 1088 7816 870720
rect 9016 1088 9616 870720
rect 12188 1088 12788 870720
rect 13988 1088 14588 870720
rect 21216 856576 21816 870720
rect 25616 856576 26216 870720
rect 37216 856576 37816 870720
rect 41616 856576 42216 870720
rect 53216 856576 53816 870720
rect 57616 856576 58216 870720
rect 61316 856576 61916 870720
rect 62716 856576 63316 870720
rect 69216 856576 69816 870720
rect 73616 856576 74216 870720
rect 85216 856576 85816 870720
rect 89616 856576 90216 870720
rect 101216 856576 101816 870720
rect 105616 856576 106216 870720
rect 111256 856576 111856 870720
rect 112656 856576 113256 870720
rect 117216 856576 117816 870720
rect 121616 856576 122216 870720
rect 133216 856576 133816 870720
rect 137616 856576 138216 870720
rect 149216 856576 149816 870720
rect 153616 856576 154216 870720
rect 165216 856576 165816 870720
rect 169616 856576 170216 870720
rect 172956 856576 173556 870720
rect 174356 856576 174956 870720
rect 181216 856576 181816 870720
rect 185616 856576 186216 870720
rect 197216 856576 197816 870720
rect 201616 856576 202216 870720
rect 213216 856576 213816 870720
rect 217616 856576 218216 870720
rect 223296 856576 223896 870720
rect 224696 856576 225296 870720
rect 229216 856576 229816 870720
rect 233616 856576 234216 870720
rect 245216 856576 245816 870720
rect 249616 856576 250216 870720
rect 261216 856576 261816 870720
rect 265616 856576 266216 870720
rect 271876 856576 272476 870720
rect 273276 856576 273876 870720
rect 277216 856576 277816 870720
rect 281616 856576 282216 870720
rect 293216 856576 293816 870720
rect 297616 856576 298216 870720
rect 309216 856576 309816 870720
rect 313616 856576 314216 870720
rect 325216 856576 325816 870720
rect 329616 856576 330216 870720
rect 341216 856576 341816 870720
rect 345616 856576 346216 870720
rect 357216 856576 357816 870720
rect 361616 856576 362216 870720
rect 373216 856576 373816 870720
rect 377616 856576 378216 870720
rect 383276 856576 383876 870720
rect 384676 856576 385276 870720
rect 389216 856576 389816 870720
rect 393616 856576 394216 870720
rect 405216 856576 405816 870720
rect 409616 856576 410216 870720
rect 421216 856576 421816 870720
rect 425616 856576 426216 870720
rect 432616 856576 433216 870720
rect 434016 856576 434616 870720
rect 437216 856576 437816 870720
rect 441616 856576 442216 870720
rect 453216 856576 453816 870720
rect 457616 856576 458216 870720
rect 466216 856576 466816 870720
rect 469216 856576 469816 870720
rect 470616 856576 471216 870720
rect 473616 856576 474216 870720
rect 485216 856576 485816 870720
rect 489616 856576 490216 870720
rect 501216 856576 501816 870720
rect 505616 856576 506216 870720
rect 517216 856576 517816 870720
rect 521616 856576 522216 870720
rect 533216 856576 533816 870720
rect 537616 856576 538216 870720
rect 549216 856576 549816 870720
rect 553616 856576 554216 870720
rect 565216 856576 565816 870720
rect 569616 856576 570216 870720
rect 576116 856576 576716 870720
rect 578516 856576 579116 870720
rect 581216 856576 581816 870720
rect 585616 856576 586216 870720
rect 597216 856576 597816 870720
rect 601616 856576 602216 870720
rect 21216 1088 21816 253264
rect 25616 1088 26216 253264
rect 37216 1088 37816 253264
rect 41616 1088 42216 253264
rect 53216 1088 53816 253264
rect 57616 1088 58216 253264
rect 61316 1088 61916 253264
rect 62716 1088 63316 253264
rect 69216 1088 69816 253264
rect 73616 1088 74216 253264
rect 85216 1088 85816 253264
rect 89616 1088 90216 253264
rect 101216 1088 101816 253264
rect 105616 1088 106216 253264
rect 111256 1088 111856 253264
rect 112656 1088 113256 253264
rect 117216 1088 117816 253264
rect 121616 1088 122216 253264
rect 133216 1088 133816 253264
rect 137616 1088 138216 253264
rect 149216 1088 149816 253264
rect 153616 1088 154216 253264
rect 165216 1088 165816 253264
rect 169616 1088 170216 253264
rect 172956 1088 173556 253264
rect 174356 1088 174956 253264
rect 181216 1088 181816 253264
rect 185616 1088 186216 253264
rect 197216 1088 197816 253264
rect 201616 1088 202216 253264
rect 213216 1088 213816 253264
rect 217616 1088 218216 253264
rect 223296 196656 223896 253264
rect 224696 196656 225296 253264
rect 223296 1088 223896 178344
rect 224696 1088 225296 178344
rect 229216 1088 229816 253264
rect 233616 1088 234216 253264
rect 245216 1088 245816 253264
rect 249616 1088 250216 253264
rect 261216 1088 261816 253264
rect 265616 1088 266216 253264
rect 271876 1088 272476 253264
rect 273276 1088 273876 253264
rect 277216 1088 277816 253264
rect 281616 1088 282216 253264
rect 293216 1088 293816 253264
rect 297616 1088 298216 253264
rect 309216 1088 309816 253264
rect 313616 1088 314216 253264
rect 325216 1088 325816 253264
rect 329616 1088 330216 253264
rect 341216 1088 341816 253264
rect 345616 1088 346216 253264
rect 357216 1088 357816 253264
rect 361616 1088 362216 253264
rect 373216 1088 373816 253264
rect 377616 1088 378216 253264
rect 383276 1088 383876 253264
rect 384676 1088 385276 253264
rect 389216 1088 389816 253264
rect 393616 1088 394216 253264
rect 405216 1088 405816 253264
rect 409616 1088 410216 253264
rect 421216 1088 421816 253264
rect 425616 1088 426216 253264
rect 432616 224656 433216 253264
rect 434016 224656 434616 253264
rect 432616 1088 433216 206344
rect 434016 1088 434616 206344
rect 437216 1088 437816 253264
rect 441616 1088 442216 253264
rect 453216 1088 453816 253264
rect 457616 1088 458216 253264
rect 466216 1088 466816 253264
rect 469216 1088 469816 253264
rect 470616 1088 471216 253264
rect 473616 1088 474216 253264
rect 485216 1088 485816 253264
rect 489616 199856 490216 253264
rect 501216 199856 501816 253264
rect 505616 199856 506216 253264
rect 517216 199856 517816 253264
rect 521616 199856 522216 253264
rect 533216 199856 533816 253264
rect 537616 199856 538216 253264
rect 549216 199856 549816 253264
rect 553616 199856 554216 253264
rect 565216 199856 565816 253264
rect 569616 199856 570216 253264
rect 576116 199856 576716 253264
rect 578516 199856 579116 253264
rect 581216 199856 581816 253264
rect 585616 199856 586216 253264
rect 597216 199856 597816 253264
rect 601616 199856 602216 253264
rect 489616 1088 490216 40544
rect 501216 1088 501816 40544
rect 505616 1088 506216 40544
rect 517216 1088 517816 40544
rect 521616 1088 522216 40544
rect 533216 1088 533816 40544
rect 537616 1088 538216 40544
rect 549216 1088 549816 40544
rect 553616 1088 554216 40544
rect 565216 1088 565816 40544
rect 569616 1088 570216 40544
rect 576116 1088 576716 40544
rect 578516 1088 579116 40544
rect 581216 28945 581816 40544
rect 585616 28945 586216 40544
rect 581216 1088 581816 17346
rect 585616 1088 586216 17346
rect 597216 1088 597816 40544
rect 601616 1088 602216 40544
rect 619816 1088 620416 870720
rect 621616 1088 622216 870720
rect 625324 1088 625924 870720
rect 627124 1088 627724 870720
rect 629104 3488 631104 868320
rect 631504 1088 633504 870720
<< obsm4 >>
rect 2604 12114 2756 865966
rect 4876 12114 7156 865966
rect 7876 12114 8956 865966
rect 9676 12114 12128 865966
rect 12848 12114 13928 865966
rect 14648 856516 21156 865966
rect 21876 856516 25556 865966
rect 26276 856516 37156 865966
rect 37876 856516 41556 865966
rect 42276 856516 53156 865966
rect 53876 856516 57556 865966
rect 58276 856516 61256 865966
rect 61976 856516 62656 865966
rect 63376 856516 69156 865966
rect 69876 856516 73556 865966
rect 74276 856516 85156 865966
rect 85876 856516 89556 865966
rect 90276 856516 101156 865966
rect 101876 856516 105556 865966
rect 106276 856516 111196 865966
rect 111916 856516 112596 865966
rect 113316 856516 117156 865966
rect 117876 856516 121556 865966
rect 122276 856516 133156 865966
rect 133876 856516 137556 865966
rect 138276 856516 149156 865966
rect 149876 856516 153556 865966
rect 154276 856516 165156 865966
rect 165876 856516 169556 865966
rect 170276 856516 172896 865966
rect 173616 856516 174296 865966
rect 175016 856516 181156 865966
rect 181876 856516 185556 865966
rect 186276 856516 197156 865966
rect 197876 856516 201556 865966
rect 202276 856516 213156 865966
rect 213876 856516 217556 865966
rect 218276 856516 223236 865966
rect 223956 856516 224636 865966
rect 225356 856516 229156 865966
rect 229876 856516 233556 865966
rect 234276 856516 245156 865966
rect 245876 856516 249556 865966
rect 250276 856516 261156 865966
rect 261876 856516 265556 865966
rect 266276 856516 271816 865966
rect 272536 856516 273216 865966
rect 273936 856516 277156 865966
rect 277876 856516 281556 865966
rect 282276 856516 293156 865966
rect 293876 856516 297556 865966
rect 298276 856516 309156 865966
rect 309876 856516 313556 865966
rect 314276 856516 325156 865966
rect 325876 856516 329556 865966
rect 330276 856516 341156 865966
rect 341876 856516 345556 865966
rect 346276 856516 357156 865966
rect 357876 856516 361556 865966
rect 362276 856516 373156 865966
rect 373876 856516 377556 865966
rect 378276 856516 383216 865966
rect 383936 856516 384616 865966
rect 385336 856516 389156 865966
rect 389876 856516 393556 865966
rect 394276 856516 405156 865966
rect 405876 856516 409556 865966
rect 410276 856516 421156 865966
rect 421876 856516 425556 865966
rect 426276 856516 432556 865966
rect 433276 856516 433956 865966
rect 434676 856516 437156 865966
rect 437876 856516 441556 865966
rect 442276 856516 453156 865966
rect 453876 856516 457556 865966
rect 458276 856516 466156 865966
rect 466876 856516 469156 865966
rect 469876 856516 470556 865966
rect 471276 856516 473556 865966
rect 474276 856516 485156 865966
rect 485876 856516 489556 865966
rect 490276 856516 501156 865966
rect 501876 856516 505556 865966
rect 506276 856516 517156 865966
rect 517876 856516 521556 865966
rect 522276 856516 533156 865966
rect 533876 856516 537556 865966
rect 538276 856516 549156 865966
rect 549876 856516 553556 865966
rect 554276 856516 565156 865966
rect 565876 856516 569556 865966
rect 570276 856516 576056 865966
rect 576776 856516 578456 865966
rect 579176 856516 581156 865966
rect 581876 856516 585556 865966
rect 586276 856516 597156 865966
rect 597876 856516 601556 865966
rect 602276 856516 619756 865966
rect 14648 253324 619756 856516
rect 14648 12114 21156 253324
rect 21876 12114 25556 253324
rect 26276 12114 37156 253324
rect 37876 12114 41556 253324
rect 42276 12114 53156 253324
rect 53876 12114 57556 253324
rect 58276 12114 61256 253324
rect 61976 12114 62656 253324
rect 63376 12114 69156 253324
rect 69876 12114 73556 253324
rect 74276 12114 85156 253324
rect 85876 12114 89556 253324
rect 90276 12114 101156 253324
rect 101876 12114 105556 253324
rect 106276 12114 111196 253324
rect 111916 12114 112596 253324
rect 113316 12114 117156 253324
rect 117876 12114 121556 253324
rect 122276 12114 133156 253324
rect 133876 12114 137556 253324
rect 138276 12114 149156 253324
rect 149876 12114 153556 253324
rect 154276 12114 165156 253324
rect 165876 12114 169556 253324
rect 170276 12114 172896 253324
rect 173616 12114 174296 253324
rect 175016 12114 181156 253324
rect 181876 12114 185556 253324
rect 186276 12114 197156 253324
rect 197876 12114 201556 253324
rect 202276 12114 213156 253324
rect 213876 12114 217556 253324
rect 218276 196596 223236 253324
rect 223956 196596 224636 253324
rect 225356 196596 229156 253324
rect 218276 178404 229156 196596
rect 218276 12114 223236 178404
rect 223956 12114 224636 178404
rect 225356 12114 229156 178404
rect 229876 12114 233556 253324
rect 234276 12114 245156 253324
rect 245876 12114 249556 253324
rect 250276 12114 261156 253324
rect 261876 12114 265556 253324
rect 266276 12114 271816 253324
rect 272536 12114 273216 253324
rect 273936 12114 277156 253324
rect 277876 12114 281556 253324
rect 282276 12114 293156 253324
rect 293876 12114 297556 253324
rect 298276 12114 309156 253324
rect 309876 12114 313556 253324
rect 314276 12114 325156 253324
rect 325876 12114 329556 253324
rect 330276 12114 341156 253324
rect 341876 12114 345556 253324
rect 346276 12114 357156 253324
rect 357876 12114 361556 253324
rect 362276 12114 373156 253324
rect 373876 12114 377556 253324
rect 378276 12114 383216 253324
rect 383936 12114 384616 253324
rect 385336 12114 389156 253324
rect 389876 12114 393556 253324
rect 394276 12114 405156 253324
rect 405876 12114 409556 253324
rect 410276 12114 421156 253324
rect 421876 12114 425556 253324
rect 426276 224596 432556 253324
rect 433276 224596 433956 253324
rect 434676 224596 437156 253324
rect 426276 206404 437156 224596
rect 426276 12114 432556 206404
rect 433276 12114 433956 206404
rect 434676 12114 437156 206404
rect 437876 12114 441556 253324
rect 442276 12114 453156 253324
rect 453876 12114 457556 253324
rect 458276 12114 466156 253324
rect 466876 12114 469156 253324
rect 469876 12114 470556 253324
rect 471276 12114 473556 253324
rect 474276 12114 485156 253324
rect 485876 199796 489556 253324
rect 490276 199796 501156 253324
rect 501876 199796 505556 253324
rect 506276 199796 517156 253324
rect 517876 199796 521556 253324
rect 522276 199796 533156 253324
rect 533876 199796 537556 253324
rect 538276 199796 549156 253324
rect 549876 199796 553556 253324
rect 554276 199796 565156 253324
rect 565876 199796 569556 253324
rect 570276 199796 576056 253324
rect 576776 199796 578456 253324
rect 579176 199796 581156 253324
rect 581876 199796 585556 253324
rect 586276 199796 597156 253324
rect 597876 199796 601556 253324
rect 602276 199796 619756 253324
rect 485876 40604 619756 199796
rect 485876 12114 489556 40604
rect 490276 12114 501156 40604
rect 501876 12114 505556 40604
rect 506276 12114 517156 40604
rect 517876 12114 521556 40604
rect 522276 12114 533156 40604
rect 533876 12114 537556 40604
rect 538276 12114 549156 40604
rect 549876 12114 553556 40604
rect 554276 12114 565156 40604
rect 565876 12114 569556 40604
rect 570276 12114 576056 40604
rect 576776 12114 578456 40604
rect 579176 28885 581156 40604
rect 581876 28885 585556 40604
rect 586276 28885 597156 40604
rect 579176 17406 597156 28885
rect 579176 12114 581156 17406
rect 581876 12114 585556 17406
rect 586276 12114 597156 17406
rect 597876 12114 601556 40604
rect 602276 12114 619756 40604
rect 620476 12114 621556 865966
rect 622276 12114 625264 865966
rect 625984 12114 627064 865966
rect 627784 12114 629044 865966
rect 631164 12114 631428 865966
<< metal5 >>
rect 416 868720 633504 870720
rect 2816 866320 631104 868320
rect 416 863318 633504 863918
rect 416 857318 633504 857918
rect 416 851318 18628 851918
rect 615372 851318 633504 851918
rect 416 845318 18628 845918
rect 615372 845318 633504 845918
rect 416 839318 18628 839918
rect 615372 839318 633504 839918
rect 416 833318 18628 833918
rect 615372 833318 633504 833918
rect 416 827318 18628 827918
rect 615372 827318 633504 827918
rect 416 821318 18628 821918
rect 615372 821318 633504 821918
rect 416 815318 18628 815918
rect 615372 815318 633504 815918
rect 416 809318 18628 809918
rect 615372 809318 633504 809918
rect 416 803318 18628 803918
rect 615372 803318 633504 803918
rect 416 797318 18628 797918
rect 615372 797318 633504 797918
rect 416 791318 18628 791918
rect 615372 791318 633504 791918
rect 416 785318 18628 785918
rect 615372 785318 633504 785918
rect 416 779318 18628 779918
rect 615372 779318 633504 779918
rect 416 773318 18628 773918
rect 615372 773318 633504 773918
rect 416 767318 18628 767918
rect 615372 767318 633504 767918
rect 416 761318 18628 761918
rect 615372 761318 633504 761918
rect 416 755318 18628 755918
rect 615372 755318 633504 755918
rect 416 749318 18628 749918
rect 615372 749318 633504 749918
rect 416 743318 18628 743918
rect 615372 743318 633504 743918
rect 416 737318 18628 737918
rect 615372 737318 633504 737918
rect 416 731318 18628 731918
rect 615372 731318 633504 731918
rect 416 725318 18628 725918
rect 615372 725318 633504 725918
rect 416 719318 18628 719918
rect 615372 719318 633504 719918
rect 416 713318 18628 713918
rect 615372 713318 633504 713918
rect 416 707318 18628 707918
rect 615372 707318 633504 707918
rect 416 701318 18628 701918
rect 615372 701318 633504 701918
rect 416 695318 18628 695918
rect 615372 695318 633504 695918
rect 416 689318 18628 689918
rect 615372 689318 633504 689918
rect 416 683318 18628 683918
rect 615372 683318 633504 683918
rect 416 677318 18628 677918
rect 615372 677318 633504 677918
rect 416 671318 18628 671918
rect 615372 671318 633504 671918
rect 416 665318 18628 665918
rect 615372 665318 633504 665918
rect 416 659318 18628 659918
rect 615372 659318 633504 659918
rect 416 653318 18628 653918
rect 615372 653318 633504 653918
rect 416 647318 18628 647918
rect 615372 647318 633504 647918
rect 416 641318 18628 641918
rect 615372 641318 633504 641918
rect 416 635318 18628 635918
rect 615372 635318 633504 635918
rect 416 629318 18628 629918
rect 615372 629318 633504 629918
rect 416 623318 18628 623918
rect 615372 623318 633504 623918
rect 416 617318 18628 617918
rect 615372 617318 633504 617918
rect 416 611318 18628 611918
rect 615372 611318 633504 611918
rect 416 605318 18628 605918
rect 615372 605318 633504 605918
rect 416 599318 18628 599918
rect 615372 599318 633504 599918
rect 416 593318 18628 593918
rect 615372 593318 633504 593918
rect 416 587318 18628 587918
rect 615372 587318 633504 587918
rect 416 581318 18628 581918
rect 615372 581318 633504 581918
rect 416 575318 18628 575918
rect 615372 575318 633504 575918
rect 416 569318 18628 569918
rect 615372 569318 633504 569918
rect 416 563318 18628 563918
rect 615372 563318 633504 563918
rect 416 557318 18628 557918
rect 615372 557318 633504 557918
rect 416 551318 18628 551918
rect 615372 551318 633504 551918
rect 416 545318 18628 545918
rect 615372 545318 633504 545918
rect 416 539318 18628 539918
rect 615372 539318 633504 539918
rect 416 533318 18628 533918
rect 615372 533318 633504 533918
rect 416 527318 18628 527918
rect 615372 527318 633504 527918
rect 416 521318 18628 521918
rect 615372 521318 633504 521918
rect 416 515318 18628 515918
rect 615372 515318 633504 515918
rect 416 509318 18628 509918
rect 615372 509318 633504 509918
rect 416 503318 18628 503918
rect 615372 503318 633504 503918
rect 416 497318 18628 497918
rect 615372 497318 633504 497918
rect 416 491318 18628 491918
rect 615372 491318 633504 491918
rect 416 485318 18628 485918
rect 615372 485318 633504 485918
rect 416 479318 18628 479918
rect 615372 479318 633504 479918
rect 416 473318 18628 473918
rect 615372 473318 633504 473918
rect 416 467318 18628 467918
rect 615372 467318 633504 467918
rect 416 461318 18628 461918
rect 615372 461318 633504 461918
rect 416 455318 18628 455918
rect 615372 455318 633504 455918
rect 416 449318 18628 449918
rect 615372 449318 633504 449918
rect 416 443318 18628 443918
rect 615372 443318 633504 443918
rect 416 437318 18628 437918
rect 615372 437318 633504 437918
rect 416 431318 18628 431918
rect 615372 431318 633504 431918
rect 416 425318 18628 425918
rect 615372 425318 633504 425918
rect 416 419318 18628 419918
rect 615372 419318 633504 419918
rect 416 413318 18628 413918
rect 615372 413318 633504 413918
rect 416 407318 18628 407918
rect 615372 407318 633504 407918
rect 416 401318 18628 401918
rect 615372 401318 633504 401918
rect 416 395318 18628 395918
rect 615372 395318 633504 395918
rect 416 389318 18628 389918
rect 615372 389318 633504 389918
rect 416 383318 18628 383918
rect 615372 383318 633504 383918
rect 416 377318 18628 377918
rect 615372 377318 633504 377918
rect 416 371318 18628 371918
rect 615372 371318 633504 371918
rect 416 365318 18628 365918
rect 615372 365318 633504 365918
rect 416 359318 18628 359918
rect 615372 359318 633504 359918
rect 416 353318 18628 353918
rect 615372 353318 633504 353918
rect 416 347318 18628 347918
rect 615372 347318 633504 347918
rect 416 341318 18628 341918
rect 615372 341318 633504 341918
rect 416 335318 18628 335918
rect 615372 335318 633504 335918
rect 416 329318 18628 329918
rect 615372 329318 633504 329918
rect 416 323318 18628 323918
rect 615372 323318 633504 323918
rect 416 317318 18628 317918
rect 615372 317318 633504 317918
rect 416 311318 18628 311918
rect 615372 311318 633504 311918
rect 416 305318 18628 305918
rect 615372 305318 633504 305918
rect 416 299318 18628 299918
rect 615372 299318 633504 299918
rect 416 293318 18628 293918
rect 615372 293318 633504 293918
rect 416 287318 18628 287918
rect 615372 287318 633504 287918
rect 416 281318 18628 281918
rect 615372 281318 633504 281918
rect 416 275318 18628 275918
rect 615372 275318 633504 275918
rect 416 269318 18628 269918
rect 615372 269318 633504 269918
rect 416 263318 18628 263918
rect 615372 263318 633504 263918
rect 416 257318 18628 257918
rect 615372 257318 633504 257918
rect 416 251318 633504 251918
rect 416 245318 633504 245918
rect 416 239318 633504 239918
rect 416 233318 633504 233918
rect 416 227318 633504 227918
rect 416 221318 312308 221918
rect 326492 221318 424208 221918
rect 438392 221318 633504 221918
rect 416 215318 312308 215918
rect 326492 215318 424208 215918
rect 438392 215318 633504 215918
rect 416 209318 312308 209918
rect 326492 209318 424208 209918
rect 438392 209318 633504 209918
rect 416 203318 633504 203918
rect 416 197318 488944 197918
rect 612656 197318 633504 197918
rect 416 191318 120308 191918
rect 134492 191318 216308 191918
rect 230492 191318 488944 191918
rect 612656 191318 633504 191918
rect 416 185318 120308 185918
rect 134492 185318 216308 185918
rect 230492 185318 488944 185918
rect 612656 185318 633504 185918
rect 416 179318 120308 179918
rect 134492 179318 216308 179918
rect 230492 179318 488944 179918
rect 612656 179318 633504 179918
rect 416 173318 488944 173918
rect 612656 173318 633504 173918
rect 416 167318 488944 167918
rect 612656 167318 633504 167918
rect 416 161318 488944 161918
rect 612656 161318 633504 161918
rect 416 155318 488944 155918
rect 612656 155318 633504 155918
rect 416 149318 488944 149918
rect 612656 149318 633504 149918
rect 416 143318 488944 143918
rect 612656 143318 633504 143918
rect 416 137318 488944 137918
rect 612656 137318 633504 137918
rect 416 131318 488944 131918
rect 612656 131318 633504 131918
rect 416 125318 488944 125918
rect 612656 125318 633504 125918
rect 416 119318 488944 119918
rect 612656 119318 633504 119918
rect 416 113318 488944 113918
rect 612656 113318 633504 113918
rect 416 107318 488944 107918
rect 612656 107318 633504 107918
rect 416 101318 488944 101918
rect 612656 101318 633504 101918
rect 416 95318 488944 95918
rect 612656 95318 633504 95918
rect 416 89318 488944 89918
rect 612656 89318 633504 89918
rect 416 83318 488944 83918
rect 612656 83318 633504 83918
rect 416 77318 488944 77918
rect 612656 77318 633504 77918
rect 416 71318 488944 71918
rect 612656 71318 633504 71918
rect 416 65318 488944 65918
rect 612656 65318 633504 65918
rect 416 59318 488944 59918
rect 612656 59318 633504 59918
rect 416 53318 488944 53918
rect 612656 53318 633504 53918
rect 416 47318 488944 47918
rect 612656 47318 633504 47918
rect 416 41318 488944 41918
rect 612656 41318 633504 41918
rect 416 35318 633504 35918
rect 416 29318 579271 29918
rect 593399 29318 633504 29918
rect 416 23318 579271 23918
rect 593399 23318 633504 23918
rect 416 17318 579371 17918
rect 593399 17318 633504 17918
rect 416 11318 633504 11918
rect 2816 3488 631104 5488
rect 416 1088 633504 3088
<< obsm5 >>
rect 2588 864018 631332 864404
rect 2588 858018 631332 863218
rect 2588 852018 631332 857218
rect 18728 851218 615272 852018
rect 2588 846018 631332 851218
rect 18728 845218 615272 846018
rect 2588 840018 631332 845218
rect 18728 839218 615272 840018
rect 2588 834018 631332 839218
rect 18728 833218 615272 834018
rect 2588 828018 631332 833218
rect 18728 827218 615272 828018
rect 2588 822018 631332 827218
rect 18728 821218 615272 822018
rect 2588 816018 631332 821218
rect 18728 815218 615272 816018
rect 2588 810018 631332 815218
rect 18728 809218 615272 810018
rect 2588 804018 631332 809218
rect 18728 803218 615272 804018
rect 2588 798018 631332 803218
rect 18728 797218 615272 798018
rect 2588 792018 631332 797218
rect 18728 791218 615272 792018
rect 2588 786018 631332 791218
rect 18728 785218 615272 786018
rect 2588 780018 631332 785218
rect 18728 779218 615272 780018
rect 2588 774018 631332 779218
rect 18728 773218 615272 774018
rect 2588 768018 631332 773218
rect 18728 767218 615272 768018
rect 2588 762018 631332 767218
rect 18728 761218 615272 762018
rect 2588 756018 631332 761218
rect 18728 755218 615272 756018
rect 2588 750018 631332 755218
rect 18728 749218 615272 750018
rect 2588 744018 631332 749218
rect 18728 743218 615272 744018
rect 2588 738018 631332 743218
rect 18728 737218 615272 738018
rect 2588 732018 631332 737218
rect 18728 731218 615272 732018
rect 2588 726018 631332 731218
rect 18728 725218 615272 726018
rect 2588 720018 631332 725218
rect 18728 719218 615272 720018
rect 2588 714018 631332 719218
rect 18728 713218 615272 714018
rect 2588 708018 631332 713218
rect 18728 707218 615272 708018
rect 2588 702018 631332 707218
rect 18728 701218 615272 702018
rect 2588 696018 631332 701218
rect 18728 695218 615272 696018
rect 2588 690018 631332 695218
rect 18728 689218 615272 690018
rect 2588 684018 631332 689218
rect 18728 683218 615272 684018
rect 2588 678018 631332 683218
rect 18728 677218 615272 678018
rect 2588 672018 631332 677218
rect 18728 671218 615272 672018
rect 2588 666018 631332 671218
rect 18728 665218 615272 666018
rect 2588 660018 631332 665218
rect 18728 659218 615272 660018
rect 2588 654018 631332 659218
rect 18728 653218 615272 654018
rect 2588 648018 631332 653218
rect 18728 647218 615272 648018
rect 2588 642018 631332 647218
rect 18728 641218 615272 642018
rect 2588 636018 631332 641218
rect 18728 635218 615272 636018
rect 2588 630018 631332 635218
rect 18728 629218 615272 630018
rect 2588 624018 631332 629218
rect 18728 623218 615272 624018
rect 2588 618018 631332 623218
rect 18728 617218 615272 618018
rect 2588 612018 631332 617218
rect 18728 611218 615272 612018
rect 2588 606018 631332 611218
rect 18728 605218 615272 606018
rect 2588 600018 631332 605218
rect 18728 599218 615272 600018
rect 2588 594018 631332 599218
rect 18728 593218 615272 594018
rect 2588 588018 631332 593218
rect 18728 587218 615272 588018
rect 2588 582018 631332 587218
rect 18728 581218 615272 582018
rect 2588 576018 631332 581218
rect 18728 575218 615272 576018
rect 2588 570018 631332 575218
rect 18728 569218 615272 570018
rect 2588 564018 631332 569218
rect 18728 563218 615272 564018
rect 2588 558018 631332 563218
rect 18728 557218 615272 558018
rect 2588 552018 631332 557218
rect 18728 551218 615272 552018
rect 2588 546018 631332 551218
rect 18728 545218 615272 546018
rect 2588 540018 631332 545218
rect 18728 539218 615272 540018
rect 2588 534018 631332 539218
rect 18728 533218 615272 534018
rect 2588 528018 631332 533218
rect 18728 527218 615272 528018
rect 2588 522018 631332 527218
rect 18728 521218 615272 522018
rect 2588 516018 631332 521218
rect 18728 515218 615272 516018
rect 2588 510018 631332 515218
rect 18728 509218 615272 510018
rect 2588 504018 631332 509218
rect 18728 503218 615272 504018
rect 2588 498018 631332 503218
rect 18728 497218 615272 498018
rect 2588 492018 631332 497218
rect 18728 491218 615272 492018
rect 2588 486018 631332 491218
rect 18728 485218 615272 486018
rect 2588 480018 631332 485218
rect 18728 479218 615272 480018
rect 2588 474018 631332 479218
rect 18728 473218 615272 474018
rect 2588 468018 631332 473218
rect 18728 467218 615272 468018
rect 2588 462018 631332 467218
rect 18728 461218 615272 462018
rect 2588 456018 631332 461218
rect 18728 455218 615272 456018
rect 2588 450018 631332 455218
rect 18728 449218 615272 450018
rect 2588 444018 631332 449218
rect 18728 443218 615272 444018
rect 2588 438018 631332 443218
rect 18728 437218 615272 438018
rect 2588 432018 631332 437218
rect 18728 431218 615272 432018
rect 2588 426018 631332 431218
rect 18728 425218 615272 426018
rect 2588 420018 631332 425218
rect 18728 419218 615272 420018
rect 2588 414018 631332 419218
rect 18728 413218 615272 414018
rect 2588 408018 631332 413218
rect 18728 407218 615272 408018
rect 2588 402018 631332 407218
rect 18728 401218 615272 402018
rect 2588 396018 631332 401218
rect 18728 395218 615272 396018
rect 2588 390018 631332 395218
rect 18728 389218 615272 390018
rect 2588 384018 631332 389218
rect 18728 383218 615272 384018
rect 2588 378018 631332 383218
rect 18728 377218 615272 378018
rect 2588 372018 631332 377218
rect 18728 371218 615272 372018
rect 2588 366018 631332 371218
rect 18728 365218 615272 366018
rect 2588 360018 631332 365218
rect 18728 359218 615272 360018
rect 2588 354018 631332 359218
rect 18728 353218 615272 354018
rect 2588 348018 631332 353218
rect 18728 347218 615272 348018
rect 2588 342018 631332 347218
rect 18728 341218 615272 342018
rect 2588 336018 631332 341218
rect 18728 335218 615272 336018
rect 2588 330018 631332 335218
rect 18728 329218 615272 330018
rect 2588 324018 631332 329218
rect 18728 323218 615272 324018
rect 2588 318018 631332 323218
rect 18728 317218 615272 318018
rect 2588 312018 631332 317218
rect 18728 311218 615272 312018
rect 2588 306018 631332 311218
rect 18728 305218 615272 306018
rect 2588 300018 631332 305218
rect 18728 299218 615272 300018
rect 2588 294018 631332 299218
rect 18728 293218 615272 294018
rect 2588 288018 631332 293218
rect 18728 287218 615272 288018
rect 2588 282018 631332 287218
rect 18728 281218 615272 282018
rect 2588 276018 631332 281218
rect 18728 275218 615272 276018
rect 2588 270018 631332 275218
rect 18728 269218 615272 270018
rect 2588 264018 631332 269218
rect 18728 263218 615272 264018
rect 2588 258018 631332 263218
rect 18728 257218 615272 258018
rect 2588 252018 631332 257218
rect 2588 246018 631332 251218
rect 2588 240018 631332 245218
rect 2588 234018 631332 239218
rect 2588 228018 631332 233218
rect 2588 222018 631332 227218
rect 312408 221218 326392 222018
rect 424308 221218 438292 222018
rect 2588 216018 631332 221218
rect 312408 215218 326392 216018
rect 424308 215218 438292 216018
rect 2588 210018 631332 215218
rect 312408 209218 326392 210018
rect 424308 209218 438292 210018
rect 2588 204018 631332 209218
rect 2588 198018 631332 203218
rect 489044 197218 612556 198018
rect 2588 192018 631332 197218
rect 120408 191218 134392 192018
rect 216408 191218 230392 192018
rect 489044 191218 612556 192018
rect 2588 186018 631332 191218
rect 120408 185218 134392 186018
rect 216408 185218 230392 186018
rect 489044 185218 612556 186018
rect 2588 180018 631332 185218
rect 120408 179218 134392 180018
rect 216408 179218 230392 180018
rect 489044 179218 612556 180018
rect 2588 174018 631332 179218
rect 489044 173218 612556 174018
rect 2588 168018 631332 173218
rect 489044 167218 612556 168018
rect 2588 162018 631332 167218
rect 489044 161218 612556 162018
rect 2588 156018 631332 161218
rect 489044 155218 612556 156018
rect 2588 150018 631332 155218
rect 489044 149218 612556 150018
rect 2588 144018 631332 149218
rect 489044 143218 612556 144018
rect 2588 138018 631332 143218
rect 489044 137218 612556 138018
rect 2588 132018 631332 137218
rect 489044 131218 612556 132018
rect 2588 126018 631332 131218
rect 489044 125218 612556 126018
rect 2588 120018 631332 125218
rect 489044 119218 612556 120018
rect 2588 114018 631332 119218
rect 489044 113218 612556 114018
rect 2588 108018 631332 113218
rect 489044 107218 612556 108018
rect 2588 102018 631332 107218
rect 489044 101218 612556 102018
rect 2588 96018 631332 101218
rect 489044 95218 612556 96018
rect 2588 90018 631332 95218
rect 489044 89218 612556 90018
rect 2588 84018 631332 89218
rect 489044 83218 612556 84018
rect 2588 78018 631332 83218
rect 489044 77218 612556 78018
rect 2588 72018 631332 77218
rect 489044 71218 612556 72018
rect 2588 66018 631332 71218
rect 489044 65218 612556 66018
rect 2588 60018 631332 65218
rect 489044 59218 612556 60018
rect 2588 54018 631332 59218
rect 489044 53218 612556 54018
rect 2588 48018 631332 53218
rect 489044 47218 612556 48018
rect 2588 42018 631332 47218
rect 489044 41218 612556 42018
rect 2588 36018 631332 41218
rect 2588 30018 631332 35218
rect 579371 29218 593299 30018
rect 2588 24018 631332 29218
rect 579371 23218 593299 24018
rect 2588 19002 631332 23218
<< labels >>
rlabel metal4 s 2816 3488 4816 868320 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 2816 3488 631104 5488 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 2816 866320 631104 868320 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 629104 3488 631104 868320 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 21216 1088 21816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 21216 856576 21816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 37216 1088 37816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 37216 856576 37816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 53216 1088 53816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 53216 856576 53816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 69216 1088 69816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 69216 856576 69816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 85216 1088 85816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 85216 856576 85816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 101216 1088 101816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 101216 856576 101816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 117216 1088 117816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 117216 856576 117816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 133216 1088 133816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 133216 856576 133816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 149216 1088 149816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 149216 856576 149816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 165216 1088 165816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 165216 856576 165816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 181216 1088 181816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 181216 856576 181816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 197216 1088 197816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 197216 856576 197816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 213216 1088 213816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 213216 856576 213816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 229216 1088 229816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 229216 856576 229816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 245216 1088 245816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 245216 856576 245816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 261216 1088 261816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 261216 856576 261816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 277216 1088 277816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 277216 856576 277816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 293216 1088 293816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 293216 856576 293816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 309216 1088 309816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 309216 856576 309816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 325216 1088 325816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 325216 856576 325816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 341216 1088 341816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 341216 856576 341816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 357216 1088 357816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 357216 856576 357816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 373216 1088 373816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 373216 856576 373816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 389216 1088 389816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 389216 856576 389816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 405216 1088 405816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 405216 856576 405816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 421216 1088 421816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 421216 856576 421816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 437216 1088 437816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 437216 856576 437816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 453216 1088 453816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 453216 856576 453816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 469216 1088 469816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 469216 856576 469816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 485216 1088 485816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 485216 856576 485816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 501216 1088 501816 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 501216 199856 501816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 501216 856576 501816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 517216 1088 517816 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 517216 199856 517816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 517216 856576 517816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 533216 1088 533816 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 533216 199856 533816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 533216 856576 533816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 549216 1088 549816 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 549216 199856 549816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 549216 856576 549816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 565216 1088 565816 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 565216 199856 565816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 565216 856576 565816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 581216 1088 581816 17346 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 581216 28945 581816 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 581216 199856 581816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 581216 856576 581816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 597216 1088 597816 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 597216 199856 597816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 597216 856576 597816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 619816 1088 620416 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 625324 1088 625924 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 7216 1088 7816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 12188 1088 12788 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 11318 633504 11918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 23318 579271 23918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 35318 633504 35918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 47318 488944 47918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 59318 488944 59918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 71318 488944 71918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 83318 488944 83918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 95318 488944 95918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 107318 488944 107918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 119318 488944 119918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 131318 488944 131918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 143318 488944 143918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 155318 488944 155918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 167318 488944 167918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 179318 120308 179918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 191318 120308 191918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 203318 633504 203918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 215318 312308 215918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 227318 633504 227918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 239318 633504 239918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 251318 633504 251918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 263318 18628 263918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 275318 18628 275918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 287318 18628 287918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 299318 18628 299918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 311318 18628 311918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 323318 18628 323918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 335318 18628 335918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 347318 18628 347918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 359318 18628 359918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 371318 18628 371918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 383318 18628 383918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 395318 18628 395918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 407318 18628 407918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 419318 18628 419918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 431318 18628 431918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 443318 18628 443918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 455318 18628 455918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 467318 18628 467918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 479318 18628 479918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 491318 18628 491918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 503318 18628 503918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 515318 18628 515918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 527318 18628 527918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 539318 18628 539918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 551318 18628 551918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 563318 18628 563918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 575318 18628 575918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 587318 18628 587918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 599318 18628 599918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 611318 18628 611918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 623318 18628 623918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 635318 18628 635918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 647318 18628 647918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 659318 18628 659918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 671318 18628 671918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 683318 18628 683918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 695318 18628 695918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 707318 18628 707918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 719318 18628 719918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 731318 18628 731918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 743318 18628 743918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 755318 18628 755918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 767318 18628 767918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 779318 18628 779918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 791318 18628 791918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 803318 18628 803918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 815318 18628 815918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 827318 18628 827918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 839318 18628 839918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 851318 18628 851918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 416 863318 633504 863918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 134492 179318 216308 179918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 134492 191318 216308 191918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 230492 179318 488944 179918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 230492 191318 488944 191918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 326492 215318 424208 215918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 438392 215318 633504 215918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 593399 23318 633504 23918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 47318 633504 47918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 59318 633504 59918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 71318 633504 71918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 83318 633504 83918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 95318 633504 95918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 107318 633504 107918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 119318 633504 119918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 131318 633504 131918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 143318 633504 143918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 155318 633504 155918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 167318 633504 167918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 179318 633504 179918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 612656 191318 633504 191918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 263318 633504 263918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 275318 633504 275918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 287318 633504 287918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 299318 633504 299918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 311318 633504 311918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 323318 633504 323918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 335318 633504 335918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 347318 633504 347918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 359318 633504 359918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 371318 633504 371918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 383318 633504 383918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 395318 633504 395918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 407318 633504 407918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 419318 633504 419918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 431318 633504 431918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 443318 633504 443918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 455318 633504 455918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 467318 633504 467918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 479318 633504 479918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 491318 633504 491918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 503318 633504 503918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 515318 633504 515918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 527318 633504 527918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 539318 633504 539918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 551318 633504 551918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 563318 633504 563918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 575318 633504 575918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 587318 633504 587918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 599318 633504 599918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 611318 633504 611918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 623318 633504 623918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 635318 633504 635918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 647318 633504 647918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 659318 633504 659918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 671318 633504 671918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 683318 633504 683918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 695318 633504 695918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 707318 633504 707918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 719318 633504 719918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 731318 633504 731918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 743318 633504 743918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 755318 633504 755918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 767318 633504 767918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 779318 633504 779918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 791318 633504 791918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 803318 633504 803918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 815318 633504 815918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 827318 633504 827918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 839318 633504 839918 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 615372 851318 633504 851918 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 466216 1088 466816 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 466216 856576 466816 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 576116 1088 576716 40544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 576116 199856 576716 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 576116 856576 576716 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 432616 1088 433216 206344 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 432616 224656 433216 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 432616 856576 433216 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 383276 1088 383876 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 383276 856576 383876 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 271876 1088 272476 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 271876 856576 272476 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 223296 1088 223896 178344 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 223296 196656 223896 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 223296 856576 223896 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 172956 1088 173556 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 172956 856576 173556 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 111256 1088 111856 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 111256 856576 111856 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 61316 1088 61916 253264 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 61316 856576 61916 870720 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 416 1088 2416 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 1088 633504 3088 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 868720 633504 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 631504 1088 633504 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25616 1088 26216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25616 856576 26216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 41616 1088 42216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 41616 856576 42216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 57616 1088 58216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 57616 856576 58216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 73616 1088 74216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 73616 856576 74216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 89616 1088 90216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 89616 856576 90216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 105616 1088 106216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 105616 856576 106216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 121616 1088 122216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 121616 856576 122216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 137616 1088 138216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 137616 856576 138216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 153616 1088 154216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 153616 856576 154216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 169616 1088 170216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 169616 856576 170216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 185616 1088 186216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 185616 856576 186216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 201616 1088 202216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 201616 856576 202216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 217616 1088 218216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 217616 856576 218216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 233616 1088 234216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 233616 856576 234216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 249616 1088 250216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 249616 856576 250216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 265616 1088 266216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 265616 856576 266216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 281616 1088 282216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 281616 856576 282216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 297616 1088 298216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 297616 856576 298216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 313616 1088 314216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 313616 856576 314216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 329616 1088 330216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 329616 856576 330216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 345616 1088 346216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 345616 856576 346216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 361616 1088 362216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 361616 856576 362216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 377616 1088 378216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 377616 856576 378216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 393616 1088 394216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 393616 856576 394216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 409616 1088 410216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 409616 856576 410216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 425616 1088 426216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 425616 856576 426216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 441616 1088 442216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 441616 856576 442216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 457616 1088 458216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 457616 856576 458216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 473616 1088 474216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 473616 856576 474216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 489616 1088 490216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 489616 199856 490216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 489616 856576 490216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 505616 1088 506216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 505616 199856 506216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 505616 856576 506216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 521616 1088 522216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 521616 199856 522216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 521616 856576 522216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 537616 1088 538216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 537616 199856 538216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 537616 856576 538216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 553616 1088 554216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 553616 199856 554216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 553616 856576 554216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 569616 1088 570216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 569616 199856 570216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 569616 856576 570216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 585616 1088 586216 17346 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 585616 28945 586216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 585616 199856 586216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 585616 856576 586216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 601616 1088 602216 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 601616 199856 602216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 601616 856576 602216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 621616 1088 622216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 627124 1088 627724 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 9016 1088 9616 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 13988 1088 14588 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 17318 579371 17918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 29318 579271 29918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 41318 488944 41918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 53318 488944 53918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 65318 488944 65918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 77318 488944 77918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 89318 488944 89918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 101318 488944 101918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 113318 488944 113918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 125318 488944 125918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 137318 488944 137918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 149318 488944 149918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 161318 488944 161918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 173318 488944 173918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 185318 120308 185918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 197318 488944 197918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 209318 312308 209918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 221318 312308 221918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 233318 633504 233918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 245318 633504 245918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 257318 18628 257918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 269318 18628 269918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 281318 18628 281918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 293318 18628 293918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 305318 18628 305918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 317318 18628 317918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 329318 18628 329918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 341318 18628 341918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 353318 18628 353918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 365318 18628 365918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 377318 18628 377918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 389318 18628 389918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 401318 18628 401918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 413318 18628 413918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 425318 18628 425918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 437318 18628 437918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 449318 18628 449918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 461318 18628 461918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 473318 18628 473918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 485318 18628 485918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 497318 18628 497918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 509318 18628 509918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 521318 18628 521918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 533318 18628 533918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 545318 18628 545918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 557318 18628 557918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 569318 18628 569918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 581318 18628 581918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 593318 18628 593918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 605318 18628 605918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 617318 18628 617918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 629318 18628 629918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 641318 18628 641918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 653318 18628 653918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 665318 18628 665918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 677318 18628 677918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 689318 18628 689918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 701318 18628 701918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 713318 18628 713918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 725318 18628 725918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 737318 18628 737918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 749318 18628 749918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 761318 18628 761918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 773318 18628 773918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 785318 18628 785918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 797318 18628 797918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 809318 18628 809918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 821318 18628 821918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 833318 18628 833918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 845318 18628 845918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 416 857318 633504 857918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 134492 185318 216308 185918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 230492 185318 488944 185918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 326492 209318 424208 209918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 326492 221318 424208 221918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 438392 209318 633504 209918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 438392 221318 633504 221918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 593399 17318 633504 17918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 593399 29318 633504 29918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 41318 633504 41918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 53318 633504 53918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 65318 633504 65918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 77318 633504 77918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 89318 633504 89918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 101318 633504 101918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 113318 633504 113918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 125318 633504 125918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 137318 633504 137918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 149318 633504 149918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 161318 633504 161918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 173318 633504 173918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 185318 633504 185918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 612656 197318 633504 197918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 257318 633504 257918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 269318 633504 269918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 281318 633504 281918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 293318 633504 293918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 305318 633504 305918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 317318 633504 317918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 329318 633504 329918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 341318 633504 341918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 353318 633504 353918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 365318 633504 365918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 377318 633504 377918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 389318 633504 389918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 401318 633504 401918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 413318 633504 413918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 425318 633504 425918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 437318 633504 437918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 449318 633504 449918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 461318 633504 461918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 473318 633504 473918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 485318 633504 485918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 497318 633504 497918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 509318 633504 509918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 521318 633504 521918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 533318 633504 533918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 545318 633504 545918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 557318 633504 557918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 569318 633504 569918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 581318 633504 581918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 593318 633504 593918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 605318 633504 605918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 617318 633504 617918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 629318 633504 629918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 641318 633504 641918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 653318 633504 653918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 665318 633504 665918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 677318 633504 677918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 689318 633504 689918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 701318 633504 701918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 713318 633504 713918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 725318 633504 725918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 737318 633504 737918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 749318 633504 749918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 761318 633504 761918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 773318 633504 773918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 785318 633504 785918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 797318 633504 797918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 809318 633504 809918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 821318 633504 821918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 833318 633504 833918 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 615372 845318 633504 845918 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 470616 1088 471216 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 470616 856576 471216 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 578516 1088 579116 40544 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 578516 199856 579116 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 578516 856576 579116 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 434016 1088 434616 206344 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 434016 224656 434616 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 434016 856576 434616 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 384676 1088 385276 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 384676 856576 385276 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 273276 1088 273876 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 273276 856576 273876 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 224696 1088 225296 178344 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 224696 196656 225296 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 224696 856576 225296 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 174356 1088 174956 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 174356 856576 174956 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 112656 1088 113256 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 112656 856576 113256 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 62716 1088 63316 253264 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 62716 856576 63316 870720 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 158172 -800 158248 800 8 clock_core
port 3 nsew signal input
rlabel metal2 s 90193 -800 90269 800 8 const_one[0]
port 4 nsew signal output
rlabel metal2 s 255193 -844 255269 800 8 const_one[1]
port 5 nsew signal output
rlabel metal2 s 432734 -802 432810 800 8 const_zero[0]
port 6 nsew signal output
rlabel metal2 s 377734 -802 377810 800 8 const_zero[1]
port 7 nsew signal output
rlabel metal2 s 322734 -802 322810 800 8 const_zero[2]
port 8 nsew signal output
rlabel metal2 s 267733 -800 267811 800 8 const_zero[3]
port 9 nsew signal output
rlabel metal2 s 145193 -810 145269 800 8 const_zero[4]
port 10 nsew signal output
rlabel metal2 s 91066 -800 91142 800 8 const_zero[5]
port 11 nsew signal output
rlabel metal2 s 474672 -802 474748 800 8 const_zero[6]
port 12 nsew signal output
rlabel metal2 s 475193 -802 475269 800 8 const_zero[7]
port 13 nsew signal output
rlabel metal2 s 476066 -802 476142 800 8 const_zero[8]
port 14 nsew signal output
rlabel metal2 s 487734 -802 487810 800 8 const_zero[9]
port 15 nsew signal output
rlabel metal2 s 322880 -800 322956 800 8 flash_clk_frame
port 16 nsew signal output
rlabel metal2 s 323026 -800 323102 800 8 flash_clk_oe
port 17 nsew signal output
rlabel metal2 s 267880 -800 267956 800 8 flash_csb_frame
port 18 nsew signal output
rlabel metal2 s 268026 -800 268102 800 8 flash_csb_oe
port 19 nsew signal output
rlabel metal2 s 378171 -800 378247 800 8 flash_io0_di
port 20 nsew signal input
rlabel metal2 s 377880 -800 377956 800 8 flash_io0_do
port 21 nsew signal output
rlabel metal2 s 366277 -800 366353 800 8 flash_io0_ie
port 22 nsew signal output
rlabel metal2 s 378026 -800 378102 800 8 flash_io0_oe
port 23 nsew signal output
rlabel metal2 s 433172 -800 433248 800 8 flash_io1_di
port 24 nsew signal input
rlabel metal2 s 432880 -800 432956 800 8 flash_io1_do
port 25 nsew signal output
rlabel metal2 s 421277 -800 421353 800 8 flash_io1_ie
port 26 nsew signal output
rlabel metal2 s 433026 -800 433102 800 8 flash_io1_oe
port 27 nsew signal output
rlabel metal2 s 475422 -800 475498 800 8 gpio_drive_select_core[0]
port 28 nsew signal output
rlabel metal2 s 475564 -800 475640 800 8 gpio_drive_select_core[1]
port 29 nsew signal output
rlabel metal2 s 488172 -800 488248 800 8 gpio_in_core
port 30 nsew signal input
rlabel metal2 s 476277 -800 476353 800 8 gpio_inenb_core
port 31 nsew signal output
rlabel metal2 s 487880 -800 487956 800 8 gpio_out_core
port 32 nsew signal output
rlabel metal2 s 488026 -800 488102 800 8 gpio_outenb_core
port 33 nsew signal output
rlabel metal2 s 632700 19422 634800 19498 6 mprj_io_drive_sel[0]
port 34 nsew signal output
rlabel metal2 s 632700 234422 634800 234498 6 mprj_io_drive_sel[10]
port 35 nsew signal output
rlabel metal2 s 632200 234564 634800 234640 6 mprj_io_drive_sel[11]
port 36 nsew signal output
rlabel metal2 s 632700 277422 634800 277498 6 mprj_io_drive_sel[12]
port 37 nsew signal output
rlabel metal2 s 632200 277564 634800 277640 6 mprj_io_drive_sel[13]
port 38 nsew signal output
rlabel metal2 s 632700 449422 634800 449498 6 mprj_io_drive_sel[14]
port 39 nsew signal output
rlabel metal2 s 632200 449564 634800 449640 6 mprj_io_drive_sel[15]
port 40 nsew signal output
rlabel metal2 s 632700 492422 634800 492498 6 mprj_io_drive_sel[16]
port 41 nsew signal output
rlabel metal2 s 632200 492564 634800 492640 6 mprj_io_drive_sel[17]
port 42 nsew signal output
rlabel metal2 s 632700 535422 634800 535498 6 mprj_io_drive_sel[18]
port 43 nsew signal output
rlabel metal2 s 632200 535564 634800 535640 6 mprj_io_drive_sel[19]
port 44 nsew signal output
rlabel metal2 s 632200 19564 634800 19640 6 mprj_io_drive_sel[1]
port 45 nsew signal output
rlabel metal2 s 632700 578422 634800 578498 6 mprj_io_drive_sel[20]
port 46 nsew signal output
rlabel metal2 s 632200 578564 634800 578640 6 mprj_io_drive_sel[21]
port 47 nsew signal output
rlabel metal2 s 632700 621422 634800 621498 6 mprj_io_drive_sel[22]
port 48 nsew signal output
rlabel metal2 s 632200 621564 634800 621640 6 mprj_io_drive_sel[23]
port 49 nsew signal output
rlabel metal2 s 632700 664422 634800 664498 6 mprj_io_drive_sel[24]
port 50 nsew signal output
rlabel metal2 s 632200 664564 634800 664640 6 mprj_io_drive_sel[25]
port 51 nsew signal output
rlabel metal2 s 632700 750422 634800 750498 6 mprj_io_drive_sel[26]
port 52 nsew signal output
rlabel metal2 s 632200 750564 634800 750640 6 mprj_io_drive_sel[27]
port 53 nsew signal output
rlabel metal2 s 632700 836422 634800 836498 6 mprj_io_drive_sel[28]
port 54 nsew signal output
rlabel metal2 s 632200 836564 634800 836640 6 mprj_io_drive_sel[29]
port 55 nsew signal output
rlabel metal2 s 632700 62422 634800 62498 6 mprj_io_drive_sel[2]
port 56 nsew signal output
rlabel metal2 s 596502 871200 596578 872800 6 mprj_io_drive_sel[30]
port 57 nsew signal output
rlabel metal2 s 596360 871200 596436 872800 6 mprj_io_drive_sel[31]
port 58 nsew signal output
rlabel metal2 s 486502 871200 486578 872800 6 mprj_io_drive_sel[32]
port 59 nsew signal output
rlabel metal2 s 486360 871200 486436 872800 6 mprj_io_drive_sel[33]
port 60 nsew signal output
rlabel metal2 s 431502 871200 431578 872800 6 mprj_io_drive_sel[34]
port 61 nsew signal output
rlabel metal2 s 431360 871200 431436 872800 6 mprj_io_drive_sel[35]
port 62 nsew signal output
rlabel metal2 s 376502 871200 376578 872800 6 mprj_io_drive_sel[36]
port 63 nsew signal output
rlabel metal2 s 376360 871200 376436 872800 6 mprj_io_drive_sel[37]
port 64 nsew signal output
rlabel metal2 s 266502 871200 266578 872800 6 mprj_io_drive_sel[38]
port 65 nsew signal output
rlabel metal2 s 266360 871200 266436 872800 6 mprj_io_drive_sel[39]
port 66 nsew signal output
rlabel metal2 s 632200 62564 634800 62640 6 mprj_io_drive_sel[3]
port 67 nsew signal output
rlabel metal2 s 211502 871200 211578 872800 6 mprj_io_drive_sel[40]
port 68 nsew signal output
rlabel metal2 s 211360 871200 211436 872800 6 mprj_io_drive_sel[41]
port 69 nsew signal output
rlabel metal2 s 156502 871200 156578 872800 6 mprj_io_drive_sel[42]
port 70 nsew signal output
rlabel metal2 s 156360 871200 156436 872800 6 mprj_io_drive_sel[43]
port 71 nsew signal output
rlabel metal2 s 101502 871200 101578 872800 6 mprj_io_drive_sel[44]
port 72 nsew signal output
rlabel metal2 s 101360 871200 101436 872800 6 mprj_io_drive_sel[45]
port 73 nsew signal output
rlabel metal2 s 46502 871200 46578 872800 6 mprj_io_drive_sel[46]
port 74 nsew signal output
rlabel metal2 s 46360 871200 46436 872800 6 mprj_io_drive_sel[47]
port 75 nsew signal output
rlabel metal2 s -800 847502 1300 847578 6 mprj_io_drive_sel[48]
port 76 nsew signal output
rlabel metal2 s -800 847360 1800 847436 6 mprj_io_drive_sel[49]
port 77 nsew signal output
rlabel metal2 s 632700 105422 634800 105498 6 mprj_io_drive_sel[4]
port 78 nsew signal output
rlabel metal2 s -800 683502 1300 683578 6 mprj_io_drive_sel[50]
port 79 nsew signal output
rlabel metal2 s -800 683360 1800 683436 6 mprj_io_drive_sel[51]
port 80 nsew signal output
rlabel metal2 s -800 642502 1300 642578 6 mprj_io_drive_sel[52]
port 81 nsew signal output
rlabel metal2 s -800 642360 1800 642436 6 mprj_io_drive_sel[53]
port 82 nsew signal output
rlabel metal2 s -800 601502 1300 601578 6 mprj_io_drive_sel[54]
port 83 nsew signal output
rlabel metal2 s -800 601360 1800 601436 6 mprj_io_drive_sel[55]
port 84 nsew signal output
rlabel metal2 s -800 560502 1300 560578 6 mprj_io_drive_sel[56]
port 85 nsew signal output
rlabel metal2 s -800 560360 1800 560436 6 mprj_io_drive_sel[57]
port 86 nsew signal output
rlabel metal2 s -800 519502 1300 519578 6 mprj_io_drive_sel[58]
port 87 nsew signal output
rlabel metal2 s -800 519360 1800 519436 6 mprj_io_drive_sel[59]
port 88 nsew signal output
rlabel metal2 s 632200 105564 634800 105640 6 mprj_io_drive_sel[5]
port 89 nsew signal output
rlabel metal2 s -800 478502 1300 478578 6 mprj_io_drive_sel[60]
port 90 nsew signal output
rlabel metal2 s -800 478360 1800 478436 6 mprj_io_drive_sel[61]
port 91 nsew signal output
rlabel metal2 s -800 437502 1300 437578 6 mprj_io_drive_sel[62]
port 92 nsew signal output
rlabel metal2 s -800 437360 1800 437436 6 mprj_io_drive_sel[63]
port 93 nsew signal output
rlabel metal2 s -800 314502 1300 314578 6 mprj_io_drive_sel[64]
port 94 nsew signal output
rlabel metal2 s -800 314360 1800 314436 6 mprj_io_drive_sel[65]
port 95 nsew signal output
rlabel metal2 s -800 273502 1300 273578 6 mprj_io_drive_sel[66]
port 96 nsew signal output
rlabel metal2 s -800 273360 1800 273436 6 mprj_io_drive_sel[67]
port 97 nsew signal output
rlabel metal2 s -800 232502 1300 232578 6 mprj_io_drive_sel[68]
port 98 nsew signal output
rlabel metal2 s -800 232360 1800 232436 6 mprj_io_drive_sel[69]
port 99 nsew signal output
rlabel metal2 s 632700 148422 634800 148498 6 mprj_io_drive_sel[6]
port 100 nsew signal output
rlabel metal2 s -800 191502 1300 191578 6 mprj_io_drive_sel[70]
port 101 nsew signal output
rlabel metal2 s -800 191360 1800 191436 6 mprj_io_drive_sel[71]
port 102 nsew signal output
rlabel metal2 s -800 150502 1300 150578 6 mprj_io_drive_sel[72]
port 103 nsew signal output
rlabel metal2 s -800 150360 1800 150436 6 mprj_io_drive_sel[73]
port 104 nsew signal output
rlabel metal2 s -800 109502 1300 109578 6 mprj_io_drive_sel[74]
port 105 nsew signal output
rlabel metal2 s -800 109360 1800 109436 6 mprj_io_drive_sel[75]
port 106 nsew signal output
rlabel metal2 s 632200 148564 634800 148640 6 mprj_io_drive_sel[7]
port 107 nsew signal output
rlabel metal2 s 632700 191422 634800 191498 6 mprj_io_drive_sel[8]
port 108 nsew signal output
rlabel metal2 s 632200 191564 634800 191640 6 mprj_io_drive_sel[9]
port 109 nsew signal output
rlabel metal2 s 631200 20277 634800 20353 6 mprj_io_ie[0]
port 110 nsew signal output
rlabel metal2 s 631200 579277 634800 579353 6 mprj_io_ie[10]
port 111 nsew signal output
rlabel metal2 s 631200 622277 634800 622353 6 mprj_io_ie[11]
port 112 nsew signal output
rlabel metal2 s 631200 665277 634800 665353 6 mprj_io_ie[12]
port 113 nsew signal output
rlabel metal2 s 631200 751277 634800 751353 6 mprj_io_ie[13]
port 114 nsew signal output
rlabel metal2 s 631200 837277 634800 837353 6 mprj_io_ie[14]
port 115 nsew signal output
rlabel metal2 s 595647 871200 595723 872800 6 mprj_io_ie[15]
port 116 nsew signal output
rlabel metal2 s 485647 871200 485723 872800 6 mprj_io_ie[16]
port 117 nsew signal output
rlabel metal2 s 430647 871200 430723 872800 6 mprj_io_ie[17]
port 118 nsew signal output
rlabel metal2 s 375647 871200 375723 872800 6 mprj_io_ie[18]
port 119 nsew signal output
rlabel metal2 s 265647 871200 265723 872800 6 mprj_io_ie[19]
port 120 nsew signal output
rlabel metal2 s 631200 63277 634800 63353 6 mprj_io_ie[1]
port 121 nsew signal output
rlabel metal2 s 210647 871200 210723 872800 6 mprj_io_ie[20]
port 122 nsew signal output
rlabel metal2 s 155647 871200 155723 872800 6 mprj_io_ie[21]
port 123 nsew signal output
rlabel metal2 s 100647 871200 100723 872800 6 mprj_io_ie[22]
port 124 nsew signal output
rlabel metal2 s 45647 871200 45723 872800 6 mprj_io_ie[23]
port 125 nsew signal output
rlabel metal2 s -800 846647 2800 846723 6 mprj_io_ie[24]
port 126 nsew signal output
rlabel metal2 s -800 682647 2800 682723 6 mprj_io_ie[25]
port 127 nsew signal output
rlabel metal2 s -800 641647 2800 641723 6 mprj_io_ie[26]
port 128 nsew signal output
rlabel metal2 s -800 600647 2800 600723 6 mprj_io_ie[27]
port 129 nsew signal output
rlabel metal2 s -800 559647 2800 559723 6 mprj_io_ie[28]
port 130 nsew signal output
rlabel metal2 s -800 518647 2800 518723 6 mprj_io_ie[29]
port 131 nsew signal output
rlabel metal2 s 631200 106277 634800 106353 6 mprj_io_ie[2]
port 132 nsew signal output
rlabel metal2 s -800 477647 2800 477723 6 mprj_io_ie[30]
port 133 nsew signal output
rlabel metal2 s -800 436647 2800 436723 6 mprj_io_ie[31]
port 134 nsew signal output
rlabel metal2 s -800 313647 2800 313723 6 mprj_io_ie[32]
port 135 nsew signal output
rlabel metal2 s -800 272647 2800 272723 6 mprj_io_ie[33]
port 136 nsew signal output
rlabel metal2 s -800 231647 2800 231723 6 mprj_io_ie[34]
port 137 nsew signal output
rlabel metal2 s -800 190647 2800 190723 6 mprj_io_ie[35]
port 138 nsew signal output
rlabel metal2 s -800 149647 2800 149723 6 mprj_io_ie[36]
port 139 nsew signal output
rlabel metal2 s -800 108647 2800 108723 6 mprj_io_ie[37]
port 140 nsew signal output
rlabel metal2 s 631200 149277 634800 149353 6 mprj_io_ie[3]
port 141 nsew signal output
rlabel metal2 s 631200 192277 634800 192353 6 mprj_io_ie[4]
port 142 nsew signal output
rlabel metal2 s 631200 235277 634800 235353 6 mprj_io_ie[5]
port 143 nsew signal output
rlabel metal2 s 631200 278277 634800 278353 6 mprj_io_ie[6]
port 144 nsew signal output
rlabel metal2 s 631200 450277 634800 450353 6 mprj_io_ie[7]
port 145 nsew signal output
rlabel metal2 s 631200 493277 634800 493353 6 mprj_io_ie[8]
port 146 nsew signal output
rlabel metal2 s 631200 536277 634800 536353 6 mprj_io_ie[9]
port 147 nsew signal output
rlabel metal2 s 632200 32172 634800 32248 6 mprj_io_in[0]
port 148 nsew signal input
rlabel metal2 s 632200 591172 634800 591248 6 mprj_io_in[10]
port 149 nsew signal input
rlabel metal2 s 632200 634172 634800 634248 6 mprj_io_in[11]
port 150 nsew signal input
rlabel metal2 s 632200 677172 634800 677248 6 mprj_io_in[12]
port 151 nsew signal input
rlabel metal2 s 632200 763172 634800 763248 6 mprj_io_in[13]
port 152 nsew signal input
rlabel metal2 s 632200 849172 634800 849248 6 mprj_io_in[14]
port 153 nsew signal input
rlabel metal2 s 583752 871200 583828 872800 6 mprj_io_in[15]
port 154 nsew signal input
rlabel metal2 s 473752 871200 473828 872800 6 mprj_io_in[16]
port 155 nsew signal input
rlabel metal2 s 418752 871200 418828 872800 6 mprj_io_in[17]
port 156 nsew signal input
rlabel metal2 s 363752 871200 363828 872800 6 mprj_io_in[18]
port 157 nsew signal input
rlabel metal2 s 253752 871200 253828 872800 6 mprj_io_in[19]
port 158 nsew signal input
rlabel metal2 s 632200 75172 634800 75248 6 mprj_io_in[1]
port 159 nsew signal input
rlabel metal2 s 198752 871200 198828 872800 6 mprj_io_in[20]
port 160 nsew signal input
rlabel metal2 s 143752 871200 143828 872800 6 mprj_io_in[21]
port 161 nsew signal input
rlabel metal2 s 88752 871200 88828 872800 6 mprj_io_in[22]
port 162 nsew signal input
rlabel metal2 s 33752 871200 33828 872800 6 mprj_io_in[23]
port 163 nsew signal input
rlabel metal2 s -800 834752 1800 834828 6 mprj_io_in[24]
port 164 nsew signal input
rlabel metal2 s -800 670752 1800 670828 6 mprj_io_in[25]
port 165 nsew signal input
rlabel metal2 s -800 629752 1800 629828 6 mprj_io_in[26]
port 166 nsew signal input
rlabel metal2 s -800 588752 1800 588828 6 mprj_io_in[27]
port 167 nsew signal input
rlabel metal2 s -800 547752 1800 547828 6 mprj_io_in[28]
port 168 nsew signal input
rlabel metal2 s -800 506752 1800 506828 6 mprj_io_in[29]
port 169 nsew signal input
rlabel metal2 s 632200 118172 634800 118248 6 mprj_io_in[2]
port 170 nsew signal input
rlabel metal2 s -800 465752 1800 465828 6 mprj_io_in[30]
port 171 nsew signal input
rlabel metal2 s -800 424752 1800 424828 6 mprj_io_in[31]
port 172 nsew signal input
rlabel metal2 s -800 301752 1800 301828 6 mprj_io_in[32]
port 173 nsew signal input
rlabel metal2 s -800 260752 1800 260828 6 mprj_io_in[33]
port 174 nsew signal input
rlabel metal2 s -800 219752 1800 219828 6 mprj_io_in[34]
port 175 nsew signal input
rlabel metal2 s -800 178752 1800 178828 6 mprj_io_in[35]
port 176 nsew signal input
rlabel metal2 s -800 137752 1800 137828 6 mprj_io_in[36]
port 177 nsew signal input
rlabel metal2 s -800 96752 1800 96828 6 mprj_io_in[37]
port 178 nsew signal input
rlabel metal2 s 632200 161172 634800 161248 6 mprj_io_in[3]
port 179 nsew signal input
rlabel metal2 s 632200 204172 634800 204248 6 mprj_io_in[4]
port 180 nsew signal input
rlabel metal2 s 632200 247172 634800 247248 6 mprj_io_in[5]
port 181 nsew signal input
rlabel metal2 s 632200 290172 634800 290248 6 mprj_io_in[6]
port 182 nsew signal input
rlabel metal2 s 632200 462172 634800 462248 6 mprj_io_in[7]
port 183 nsew signal input
rlabel metal2 s 632200 505172 634800 505248 6 mprj_io_in[8]
port 184 nsew signal input
rlabel metal2 s 632200 548172 634800 548248 6 mprj_io_in[9]
port 185 nsew signal input
rlabel metal2 s 632700 32026 634800 32102 6 mprj_io_oe[0]
port 186 nsew signal output
rlabel metal2 s 632700 591026 634800 591102 6 mprj_io_oe[10]
port 187 nsew signal output
rlabel metal2 s 632700 634026 634800 634102 6 mprj_io_oe[11]
port 188 nsew signal output
rlabel metal2 s 632700 677026 634800 677102 6 mprj_io_oe[12]
port 189 nsew signal output
rlabel metal2 s 632700 763026 634800 763102 6 mprj_io_oe[13]
port 190 nsew signal output
rlabel metal2 s 632700 849026 634800 849102 6 mprj_io_oe[14]
port 191 nsew signal output
rlabel metal2 s 583898 871200 583974 872800 6 mprj_io_oe[15]
port 192 nsew signal output
rlabel metal2 s 473898 871200 473974 872800 6 mprj_io_oe[16]
port 193 nsew signal output
rlabel metal2 s 418898 871200 418974 872800 6 mprj_io_oe[17]
port 194 nsew signal output
rlabel metal2 s 363898 871200 363974 872800 6 mprj_io_oe[18]
port 195 nsew signal output
rlabel metal2 s 253898 871200 253974 872800 6 mprj_io_oe[19]
port 196 nsew signal output
rlabel metal2 s 632700 75026 634800 75102 6 mprj_io_oe[1]
port 197 nsew signal output
rlabel metal2 s 198898 871200 198974 872800 6 mprj_io_oe[20]
port 198 nsew signal output
rlabel metal2 s 143898 871200 143974 872800 6 mprj_io_oe[21]
port 199 nsew signal output
rlabel metal2 s 88898 871200 88974 872800 6 mprj_io_oe[22]
port 200 nsew signal output
rlabel metal2 s 33898 871200 33974 872800 6 mprj_io_oe[23]
port 201 nsew signal output
rlabel metal2 s -800 834898 1300 834974 6 mprj_io_oe[24]
port 202 nsew signal output
rlabel metal2 s -800 670898 1300 670974 6 mprj_io_oe[25]
port 203 nsew signal output
rlabel metal2 s -800 629898 1300 629974 6 mprj_io_oe[26]
port 204 nsew signal output
rlabel metal2 s -800 588898 1300 588974 6 mprj_io_oe[27]
port 205 nsew signal output
rlabel metal2 s -800 547898 1300 547974 6 mprj_io_oe[28]
port 206 nsew signal output
rlabel metal2 s -800 506898 1300 506974 6 mprj_io_oe[29]
port 207 nsew signal output
rlabel metal2 s 632700 118026 634800 118102 6 mprj_io_oe[2]
port 208 nsew signal output
rlabel metal2 s -800 465898 1300 465974 6 mprj_io_oe[30]
port 209 nsew signal output
rlabel metal2 s -800 424898 1300 424974 6 mprj_io_oe[31]
port 210 nsew signal output
rlabel metal2 s -800 301898 1300 301974 6 mprj_io_oe[32]
port 211 nsew signal output
rlabel metal2 s -800 260898 1300 260974 6 mprj_io_oe[33]
port 212 nsew signal output
rlabel metal2 s -800 219898 1300 219974 6 mprj_io_oe[34]
port 213 nsew signal output
rlabel metal2 s -800 178898 1300 178974 6 mprj_io_oe[35]
port 214 nsew signal output
rlabel metal2 s -800 137898 1300 137974 6 mprj_io_oe[36]
port 215 nsew signal output
rlabel metal2 s -800 96898 1300 96974 6 mprj_io_oe[37]
port 216 nsew signal output
rlabel metal2 s 632700 161026 634800 161102 6 mprj_io_oe[3]
port 217 nsew signal output
rlabel metal2 s 632700 204026 634800 204102 6 mprj_io_oe[4]
port 218 nsew signal output
rlabel metal2 s 632700 247026 634800 247102 6 mprj_io_oe[5]
port 219 nsew signal output
rlabel metal2 s 632700 290026 634800 290102 6 mprj_io_oe[6]
port 220 nsew signal output
rlabel metal2 s 632700 462026 634800 462102 6 mprj_io_oe[7]
port 221 nsew signal output
rlabel metal2 s 632700 505026 634800 505102 6 mprj_io_oe[8]
port 222 nsew signal output
rlabel metal2 s 632700 548026 634800 548102 6 mprj_io_oe[9]
port 223 nsew signal output
rlabel metal2 s 633200 31880 634800 31956 6 mprj_io_out[0]
port 224 nsew signal output
rlabel metal2 s 633200 590880 634800 590956 6 mprj_io_out[10]
port 225 nsew signal output
rlabel metal2 s 633200 633880 634800 633956 6 mprj_io_out[11]
port 226 nsew signal output
rlabel metal2 s 633200 676880 634800 676956 6 mprj_io_out[12]
port 227 nsew signal output
rlabel metal2 s 633200 762880 634800 762956 6 mprj_io_out[13]
port 228 nsew signal output
rlabel metal2 s 633200 848880 634800 848956 6 mprj_io_out[14]
port 229 nsew signal output
rlabel metal2 s 584044 871200 584120 872800 6 mprj_io_out[15]
port 230 nsew signal output
rlabel metal2 s 474044 871200 474120 872800 6 mprj_io_out[16]
port 231 nsew signal output
rlabel metal2 s 419044 871200 419120 872800 6 mprj_io_out[17]
port 232 nsew signal output
rlabel metal2 s 364044 871200 364120 872800 6 mprj_io_out[18]
port 233 nsew signal output
rlabel metal2 s 254044 871200 254120 872800 6 mprj_io_out[19]
port 234 nsew signal output
rlabel metal2 s 633200 74880 634800 74956 6 mprj_io_out[1]
port 235 nsew signal output
rlabel metal2 s 199044 871200 199120 872800 6 mprj_io_out[20]
port 236 nsew signal output
rlabel metal2 s 144044 871200 144120 872800 6 mprj_io_out[21]
port 237 nsew signal output
rlabel metal2 s 89044 871200 89120 872800 6 mprj_io_out[22]
port 238 nsew signal output
rlabel metal2 s 34044 871200 34120 872800 6 mprj_io_out[23]
port 239 nsew signal output
rlabel metal2 s -800 835044 800 835120 4 mprj_io_out[24]
port 240 nsew signal output
rlabel metal2 s -800 671044 800 671120 4 mprj_io_out[25]
port 241 nsew signal output
rlabel metal2 s -800 630044 800 630120 4 mprj_io_out[26]
port 242 nsew signal output
rlabel metal2 s -800 589044 800 589120 4 mprj_io_out[27]
port 243 nsew signal output
rlabel metal2 s -800 548044 800 548120 4 mprj_io_out[28]
port 244 nsew signal output
rlabel metal2 s -800 507044 800 507120 4 mprj_io_out[29]
port 245 nsew signal output
rlabel metal2 s 633200 117880 634800 117956 6 mprj_io_out[2]
port 246 nsew signal output
rlabel metal2 s -800 466044 800 466120 4 mprj_io_out[30]
port 247 nsew signal output
rlabel metal2 s -800 425044 800 425120 4 mprj_io_out[31]
port 248 nsew signal output
rlabel metal2 s -800 302044 800 302120 4 mprj_io_out[32]
port 249 nsew signal output
rlabel metal2 s -800 261044 800 261120 4 mprj_io_out[33]
port 250 nsew signal output
rlabel metal2 s -800 220044 800 220120 4 mprj_io_out[34]
port 251 nsew signal output
rlabel metal2 s -800 179044 800 179120 4 mprj_io_out[35]
port 252 nsew signal output
rlabel metal2 s -800 138044 800 138120 4 mprj_io_out[36]
port 253 nsew signal output
rlabel metal2 s -800 97044 800 97120 4 mprj_io_out[37]
port 254 nsew signal output
rlabel metal2 s 633200 160880 634800 160956 6 mprj_io_out[3]
port 255 nsew signal output
rlabel metal2 s 633200 203880 634800 203956 6 mprj_io_out[4]
port 256 nsew signal output
rlabel metal2 s 633200 246880 634800 246956 6 mprj_io_out[5]
port 257 nsew signal output
rlabel metal2 s 633200 289880 634800 289956 6 mprj_io_out[6]
port 258 nsew signal output
rlabel metal2 s 633200 461880 634800 461956 6 mprj_io_out[7]
port 259 nsew signal output
rlabel metal2 s 633200 504880 634800 504956 6 mprj_io_out[8]
port 260 nsew signal output
rlabel metal2 s 633200 547880 634800 547956 6 mprj_io_out[9]
port 261 nsew signal output
rlabel metal2 s 631700 20066 634800 20142 6 mprj_io_pulldown_sel[0]
port 262 nsew signal output
rlabel metal2 s 631700 579066 634800 579142 6 mprj_io_pulldown_sel[10]
port 263 nsew signal output
rlabel metal2 s 631700 622066 634800 622142 6 mprj_io_pulldown_sel[11]
port 264 nsew signal output
rlabel metal2 s 631700 665066 634800 665142 6 mprj_io_pulldown_sel[12]
port 265 nsew signal output
rlabel metal2 s 631700 751066 634800 751142 6 mprj_io_pulldown_sel[13]
port 266 nsew signal output
rlabel metal2 s 631700 837066 634800 837142 6 mprj_io_pulldown_sel[14]
port 267 nsew signal output
rlabel metal2 s 595858 871200 595934 872800 6 mprj_io_pulldown_sel[15]
port 268 nsew signal output
rlabel metal2 s 485858 871200 485934 872800 6 mprj_io_pulldown_sel[16]
port 269 nsew signal output
rlabel metal2 s 430858 871200 430934 872800 6 mprj_io_pulldown_sel[17]
port 270 nsew signal output
rlabel metal2 s 375858 871200 375934 872800 6 mprj_io_pulldown_sel[18]
port 271 nsew signal output
rlabel metal2 s 265858 871200 265934 872800 6 mprj_io_pulldown_sel[19]
port 272 nsew signal output
rlabel metal2 s 631700 63066 634800 63142 6 mprj_io_pulldown_sel[1]
port 273 nsew signal output
rlabel metal2 s 210858 871200 210934 872800 6 mprj_io_pulldown_sel[20]
port 274 nsew signal output
rlabel metal2 s 155858 871200 155934 872800 6 mprj_io_pulldown_sel[21]
port 275 nsew signal output
rlabel metal2 s 100858 871200 100934 872800 6 mprj_io_pulldown_sel[22]
port 276 nsew signal output
rlabel metal2 s 45858 871200 45934 872800 6 mprj_io_pulldown_sel[23]
port 277 nsew signal output
rlabel metal2 s -800 846858 2300 846934 6 mprj_io_pulldown_sel[24]
port 278 nsew signal output
rlabel metal2 s -800 682858 2300 682934 6 mprj_io_pulldown_sel[25]
port 279 nsew signal output
rlabel metal2 s -800 641858 2300 641934 6 mprj_io_pulldown_sel[26]
port 280 nsew signal output
rlabel metal2 s -800 600858 2300 600934 6 mprj_io_pulldown_sel[27]
port 281 nsew signal output
rlabel metal2 s -800 559858 2300 559934 6 mprj_io_pulldown_sel[28]
port 282 nsew signal output
rlabel metal2 s -800 518858 2300 518934 6 mprj_io_pulldown_sel[29]
port 283 nsew signal output
rlabel metal2 s 631700 106066 634800 106142 6 mprj_io_pulldown_sel[2]
port 284 nsew signal output
rlabel metal2 s -800 477858 2300 477934 6 mprj_io_pulldown_sel[30]
port 285 nsew signal output
rlabel metal2 s -800 436858 2300 436934 6 mprj_io_pulldown_sel[31]
port 286 nsew signal output
rlabel metal2 s -800 313858 2300 313934 6 mprj_io_pulldown_sel[32]
port 287 nsew signal output
rlabel metal2 s -800 272858 2300 272934 6 mprj_io_pulldown_sel[33]
port 288 nsew signal output
rlabel metal2 s -800 231858 2300 231934 6 mprj_io_pulldown_sel[34]
port 289 nsew signal output
rlabel metal2 s -800 190858 2300 190934 6 mprj_io_pulldown_sel[35]
port 290 nsew signal output
rlabel metal2 s -800 149858 2300 149934 6 mprj_io_pulldown_sel[36]
port 291 nsew signal output
rlabel metal2 s -800 108858 2300 108934 6 mprj_io_pulldown_sel[37]
port 292 nsew signal output
rlabel metal2 s 631700 149066 634800 149142 6 mprj_io_pulldown_sel[3]
port 293 nsew signal output
rlabel metal2 s 631700 192066 634800 192142 6 mprj_io_pulldown_sel[4]
port 294 nsew signal output
rlabel metal2 s 631700 235066 634800 235142 6 mprj_io_pulldown_sel[5]
port 295 nsew signal output
rlabel metal2 s 631700 278066 634800 278142 6 mprj_io_pulldown_sel[6]
port 296 nsew signal output
rlabel metal2 s 631700 450066 634800 450142 6 mprj_io_pulldown_sel[7]
port 297 nsew signal output
rlabel metal2 s 631700 493066 634800 493142 6 mprj_io_pulldown_sel[8]
port 298 nsew signal output
rlabel metal2 s 631700 536066 634800 536142 6 mprj_io_pulldown_sel[9]
port 299 nsew signal output
rlabel metal2 s 633200 19193 634800 19269 6 mprj_io_pullup_sel[0]
port 300 nsew signal output
rlabel metal2 s 633200 578193 634800 578269 6 mprj_io_pullup_sel[10]
port 301 nsew signal output
rlabel metal2 s 633200 621193 634800 621269 6 mprj_io_pullup_sel[11]
port 302 nsew signal output
rlabel metal2 s 633200 664193 634800 664269 6 mprj_io_pullup_sel[12]
port 303 nsew signal output
rlabel metal2 s 633200 750193 634800 750269 6 mprj_io_pullup_sel[13]
port 304 nsew signal output
rlabel metal2 s 633200 836193 634800 836269 6 mprj_io_pullup_sel[14]
port 305 nsew signal output
rlabel metal2 s 596731 871200 596807 872800 6 mprj_io_pullup_sel[15]
port 306 nsew signal output
rlabel metal2 s 486731 871200 486807 872800 6 mprj_io_pullup_sel[16]
port 307 nsew signal output
rlabel metal2 s 431731 871200 431807 872800 6 mprj_io_pullup_sel[17]
port 308 nsew signal output
rlabel metal2 s 376731 871200 376807 872800 6 mprj_io_pullup_sel[18]
port 309 nsew signal output
rlabel metal2 s 266731 871200 266807 872800 6 mprj_io_pullup_sel[19]
port 310 nsew signal output
rlabel metal2 s 633200 62193 634800 62269 6 mprj_io_pullup_sel[1]
port 311 nsew signal output
rlabel metal2 s 211731 871200 211807 872800 6 mprj_io_pullup_sel[20]
port 312 nsew signal output
rlabel metal2 s 156731 871200 156807 872800 6 mprj_io_pullup_sel[21]
port 313 nsew signal output
rlabel metal2 s 101731 871200 101807 872800 6 mprj_io_pullup_sel[22]
port 314 nsew signal output
rlabel metal2 s 46731 871200 46807 872800 6 mprj_io_pullup_sel[23]
port 315 nsew signal output
rlabel metal2 s -800 847731 800 847807 4 mprj_io_pullup_sel[24]
port 316 nsew signal output
rlabel metal2 s -800 683731 800 683807 4 mprj_io_pullup_sel[25]
port 317 nsew signal output
rlabel metal2 s -800 642731 800 642807 4 mprj_io_pullup_sel[26]
port 318 nsew signal output
rlabel metal2 s -800 601731 800 601807 4 mprj_io_pullup_sel[27]
port 319 nsew signal output
rlabel metal2 s -800 560731 800 560807 4 mprj_io_pullup_sel[28]
port 320 nsew signal output
rlabel metal2 s -800 519731 800 519807 4 mprj_io_pullup_sel[29]
port 321 nsew signal output
rlabel metal2 s 633200 105193 634800 105269 6 mprj_io_pullup_sel[2]
port 322 nsew signal output
rlabel metal2 s -800 478731 800 478807 4 mprj_io_pullup_sel[30]
port 323 nsew signal output
rlabel metal2 s -800 437731 800 437807 4 mprj_io_pullup_sel[31]
port 324 nsew signal output
rlabel metal2 s -800 314731 800 314807 4 mprj_io_pullup_sel[32]
port 325 nsew signal output
rlabel metal2 s -800 273731 800 273807 4 mprj_io_pullup_sel[33]
port 326 nsew signal output
rlabel metal2 s -800 232731 800 232807 4 mprj_io_pullup_sel[34]
port 327 nsew signal output
rlabel metal2 s -800 191731 800 191807 4 mprj_io_pullup_sel[35]
port 328 nsew signal output
rlabel metal2 s -800 150731 800 150807 4 mprj_io_pullup_sel[36]
port 329 nsew signal output
rlabel metal2 s -800 109731 800 109807 4 mprj_io_pullup_sel[37]
port 330 nsew signal output
rlabel metal2 s 633200 148193 634800 148269 6 mprj_io_pullup_sel[3]
port 331 nsew signal output
rlabel metal2 s 633200 191193 634800 191269 6 mprj_io_pullup_sel[4]
port 332 nsew signal output
rlabel metal2 s 633200 234193 634800 234269 6 mprj_io_pullup_sel[5]
port 333 nsew signal output
rlabel metal2 s 633200 277193 634800 277269 6 mprj_io_pullup_sel[6]
port 334 nsew signal output
rlabel metal2 s 633200 449193 634800 449269 6 mprj_io_pullup_sel[7]
port 335 nsew signal output
rlabel metal2 s 633200 492193 634800 492269 6 mprj_io_pullup_sel[8]
port 336 nsew signal output
rlabel metal2 s 633200 535193 634800 535269 6 mprj_io_pullup_sel[9]
port 337 nsew signal output
rlabel metal2 s 633700 18672 634800 18748 6 mprj_io_schmitt_sel[0]
port 338 nsew signal output
rlabel metal2 s 633700 577672 634800 577748 6 mprj_io_schmitt_sel[10]
port 339 nsew signal output
rlabel metal2 s 633700 620672 634800 620748 6 mprj_io_schmitt_sel[11]
port 340 nsew signal output
rlabel metal2 s 633700 663672 634800 663748 6 mprj_io_schmitt_sel[12]
port 341 nsew signal output
rlabel metal2 s 633700 749672 634800 749748 6 mprj_io_schmitt_sel[13]
port 342 nsew signal output
rlabel metal2 s 633700 835672 634800 835748 6 mprj_io_schmitt_sel[14]
port 343 nsew signal output
rlabel metal2 s 597252 871200 597328 872800 6 mprj_io_schmitt_sel[15]
port 344 nsew signal output
rlabel metal2 s 487252 871200 487328 872800 6 mprj_io_schmitt_sel[16]
port 345 nsew signal output
rlabel metal2 s 432252 871200 432328 872800 6 mprj_io_schmitt_sel[17]
port 346 nsew signal output
rlabel metal2 s 377252 871200 377328 872800 6 mprj_io_schmitt_sel[18]
port 347 nsew signal output
rlabel metal2 s 267252 871200 267328 872800 6 mprj_io_schmitt_sel[19]
port 348 nsew signal output
rlabel metal2 s 633700 61672 634800 61748 6 mprj_io_schmitt_sel[1]
port 349 nsew signal output
rlabel metal2 s 212252 871200 212328 872800 6 mprj_io_schmitt_sel[20]
port 350 nsew signal output
rlabel metal2 s 157252 871200 157328 872800 6 mprj_io_schmitt_sel[21]
port 351 nsew signal output
rlabel metal2 s 102252 871200 102328 872800 6 mprj_io_schmitt_sel[22]
port 352 nsew signal output
rlabel metal2 s 47252 871200 47328 872800 6 mprj_io_schmitt_sel[23]
port 353 nsew signal output
rlabel metal2 s -800 848252 300 848328 4 mprj_io_schmitt_sel[24]
port 354 nsew signal output
rlabel metal2 s -800 684252 300 684328 4 mprj_io_schmitt_sel[25]
port 355 nsew signal output
rlabel metal2 s -800 643252 300 643328 4 mprj_io_schmitt_sel[26]
port 356 nsew signal output
rlabel metal2 s -800 602252 300 602328 4 mprj_io_schmitt_sel[27]
port 357 nsew signal output
rlabel metal2 s -800 561252 300 561328 4 mprj_io_schmitt_sel[28]
port 358 nsew signal output
rlabel metal2 s -800 520252 300 520328 4 mprj_io_schmitt_sel[29]
port 359 nsew signal output
rlabel metal2 s 633700 104672 634800 104748 6 mprj_io_schmitt_sel[2]
port 360 nsew signal output
rlabel metal2 s -800 479252 300 479328 4 mprj_io_schmitt_sel[30]
port 361 nsew signal output
rlabel metal2 s -800 438252 300 438328 4 mprj_io_schmitt_sel[31]
port 362 nsew signal output
rlabel metal2 s -800 315252 300 315328 4 mprj_io_schmitt_sel[32]
port 363 nsew signal output
rlabel metal2 s -800 274252 300 274328 4 mprj_io_schmitt_sel[33]
port 364 nsew signal output
rlabel metal2 s -800 233252 300 233328 4 mprj_io_schmitt_sel[34]
port 365 nsew signal output
rlabel metal2 s -800 192252 300 192328 4 mprj_io_schmitt_sel[35]
port 366 nsew signal output
rlabel metal2 s -800 151252 300 151328 4 mprj_io_schmitt_sel[36]
port 367 nsew signal output
rlabel metal2 s -800 110252 300 110328 4 mprj_io_schmitt_sel[37]
port 368 nsew signal output
rlabel metal2 s 633700 147672 634800 147748 6 mprj_io_schmitt_sel[3]
port 369 nsew signal output
rlabel metal2 s 633700 190672 634800 190748 6 mprj_io_schmitt_sel[4]
port 370 nsew signal output
rlabel metal2 s 633700 233672 634800 233748 6 mprj_io_schmitt_sel[5]
port 371 nsew signal output
rlabel metal2 s 633700 276672 634800 276748 6 mprj_io_schmitt_sel[6]
port 372 nsew signal output
rlabel metal2 s 633700 448672 634800 448748 6 mprj_io_schmitt_sel[7]
port 373 nsew signal output
rlabel metal2 s 633700 491672 634800 491748 6 mprj_io_schmitt_sel[8]
port 374 nsew signal output
rlabel metal2 s 633700 534672 634800 534748 6 mprj_io_schmitt_sel[9]
port 375 nsew signal output
rlabel metal2 s 633700 31734 634800 31810 6 mprj_io_slew_sel[0]
port 376 nsew signal output
rlabel metal2 s 633700 590734 634800 590810 6 mprj_io_slew_sel[10]
port 377 nsew signal output
rlabel metal2 s 633700 633734 634800 633810 6 mprj_io_slew_sel[11]
port 378 nsew signal output
rlabel metal2 s 633700 676734 634800 676810 6 mprj_io_slew_sel[12]
port 379 nsew signal output
rlabel metal2 s 633700 762734 634800 762810 6 mprj_io_slew_sel[13]
port 380 nsew signal output
rlabel metal2 s 633700 848734 634800 848810 6 mprj_io_slew_sel[14]
port 381 nsew signal output
rlabel metal2 s 584190 871200 584266 872800 6 mprj_io_slew_sel[15]
port 382 nsew signal output
rlabel metal2 s 474190 871200 474266 872800 6 mprj_io_slew_sel[16]
port 383 nsew signal output
rlabel metal2 s 419190 871200 419266 872800 6 mprj_io_slew_sel[17]
port 384 nsew signal output
rlabel metal2 s 364190 871200 364266 872800 6 mprj_io_slew_sel[18]
port 385 nsew signal output
rlabel metal2 s 254190 871200 254266 872800 6 mprj_io_slew_sel[19]
port 386 nsew signal output
rlabel metal2 s 633700 74734 634800 74810 6 mprj_io_slew_sel[1]
port 387 nsew signal output
rlabel metal2 s 199190 871200 199266 872800 6 mprj_io_slew_sel[20]
port 388 nsew signal output
rlabel metal2 s 144190 871200 144266 872800 6 mprj_io_slew_sel[21]
port 389 nsew signal output
rlabel metal2 s 89190 871200 89266 872800 6 mprj_io_slew_sel[22]
port 390 nsew signal output
rlabel metal2 s 34190 871200 34266 872800 6 mprj_io_slew_sel[23]
port 391 nsew signal output
rlabel metal2 s -800 835190 300 835266 4 mprj_io_slew_sel[24]
port 392 nsew signal output
rlabel metal2 s -800 671190 300 671266 4 mprj_io_slew_sel[25]
port 393 nsew signal output
rlabel metal2 s -800 630190 300 630266 4 mprj_io_slew_sel[26]
port 394 nsew signal output
rlabel metal2 s -800 589190 300 589266 4 mprj_io_slew_sel[27]
port 395 nsew signal output
rlabel metal2 s -800 548190 300 548266 4 mprj_io_slew_sel[28]
port 396 nsew signal output
rlabel metal2 s -800 507190 300 507266 4 mprj_io_slew_sel[29]
port 397 nsew signal output
rlabel metal2 s 633700 117734 634800 117810 6 mprj_io_slew_sel[2]
port 398 nsew signal output
rlabel metal2 s -800 466190 300 466266 4 mprj_io_slew_sel[30]
port 399 nsew signal output
rlabel metal2 s -800 425190 300 425266 4 mprj_io_slew_sel[31]
port 400 nsew signal output
rlabel metal2 s -800 302190 300 302266 4 mprj_io_slew_sel[32]
port 401 nsew signal output
rlabel metal2 s -800 261190 300 261266 4 mprj_io_slew_sel[33]
port 402 nsew signal output
rlabel metal2 s -800 220190 300 220266 4 mprj_io_slew_sel[34]
port 403 nsew signal output
rlabel metal2 s -800 179190 300 179266 4 mprj_io_slew_sel[35]
port 404 nsew signal output
rlabel metal2 s -800 138190 300 138266 4 mprj_io_slew_sel[36]
port 405 nsew signal output
rlabel metal2 s -800 97190 300 97266 4 mprj_io_slew_sel[37]
port 406 nsew signal output
rlabel metal2 s 633700 160734 634800 160810 6 mprj_io_slew_sel[3]
port 407 nsew signal output
rlabel metal2 s 633700 203734 634800 203810 6 mprj_io_slew_sel[4]
port 408 nsew signal output
rlabel metal2 s 633700 246734 634800 246810 6 mprj_io_slew_sel[5]
port 409 nsew signal output
rlabel metal2 s 633700 289734 634800 289810 6 mprj_io_slew_sel[6]
port 410 nsew signal output
rlabel metal2 s 633700 461734 634800 461810 6 mprj_io_slew_sel[7]
port 411 nsew signal output
rlabel metal2 s 633700 504734 634800 504810 6 mprj_io_slew_sel[8]
port 412 nsew signal output
rlabel metal2 s 633700 547734 634800 547810 6 mprj_io_slew_sel[9]
port 413 nsew signal output
rlabel metal2 s 103172 -800 103248 800 8 rstb
port 414 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 634000 872000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 106434896
string GDS_FILE /home/hosni/GF180/PnR_2/caravel-gf180mcu/openlane/caravel_core/runs/RUN_2022.11.29_17.28.14/results/signoff/caravel_core.magic.gds
string GDS_START 41779966
<< end >>

