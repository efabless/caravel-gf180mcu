magic
tech gf180mcuC
magscale 1 10
timestamp 1668623937
<< checkpaint >>
rect -8119 -2000 786119 1022000
<< metal1 >>
rect 73210 946038 73222 946090
rect 73274 946038 73286 946090
rect 73225 945751 73271 946038
rect 77578 945751 77590 945754
rect 73225 945705 77590 945751
rect 77578 945702 77590 945705
rect 77642 945702 77654 945754
rect 105802 942342 105814 942394
rect 105866 942391 105878 942394
rect 196522 942391 196534 942394
rect 105866 942345 196534 942391
rect 105866 942342 105878 942345
rect 196522 942342 196534 942345
rect 196586 942342 196598 942394
rect 216346 942342 216358 942394
rect 216410 942391 216422 942394
rect 306506 942391 306518 942394
rect 216410 942345 306518 942391
rect 216410 942342 216422 942345
rect 306506 942342 306518 942345
rect 306570 942342 306582 942394
rect 161130 942230 161142 942282
rect 161194 942279 161206 942282
rect 251290 942279 251302 942282
rect 161194 942233 251302 942279
rect 161194 942230 161206 942233
rect 251290 942230 251302 942233
rect 251354 942230 251366 942282
rect 270442 942230 270454 942282
rect 270506 942279 270518 942282
rect 361162 942279 361174 942282
rect 270506 942233 361174 942279
rect 270506 942230 270518 942233
rect 361162 942230 361174 942233
rect 361226 942230 361238 942282
rect 160346 942118 160358 942170
rect 160410 942167 160422 942170
rect 251066 942167 251078 942170
rect 160410 942121 251078 942167
rect 160410 942118 160422 942121
rect 251066 942118 251078 942121
rect 251130 942118 251142 942170
rect 271338 942118 271350 942170
rect 271402 942167 271414 942170
rect 335850 942167 335862 942170
rect 271402 942121 335862 942167
rect 271402 942118 271414 942121
rect 335850 942118 335862 942121
rect 335914 942118 335926 942170
rect 106362 942006 106374 942058
rect 106426 942055 106438 942058
rect 196298 942055 196310 942058
rect 106426 942009 196310 942055
rect 106426 942006 106438 942009
rect 196298 942006 196310 942009
rect 196362 942006 196374 942058
rect 215562 942006 215574 942058
rect 215626 942055 215638 942058
rect 306058 942055 306070 942058
rect 215626 942009 306070 942055
rect 215626 942006 215638 942009
rect 306058 942006 306070 942009
rect 306122 942006 306134 942058
rect 177034 938198 177046 938250
rect 177098 938247 177110 938250
rect 687754 938247 687766 938250
rect 177098 938201 687766 938247
rect 177098 938198 177110 938201
rect 687754 938198 687766 938201
rect 687818 938198 687830 938250
rect 341002 937414 341014 937466
rect 341066 937463 341078 937466
rect 344586 937463 344598 937466
rect 341066 937417 344598 937463
rect 341066 937414 341078 937417
rect 344586 937414 344598 937417
rect 344650 937414 344662 937466
rect 120922 937302 120934 937354
rect 120986 937351 120998 937354
rect 688202 937351 688214 937354
rect 120986 937305 688214 937351
rect 120986 937302 120998 937305
rect 688202 937302 688214 937305
rect 688266 937302 688278 937354
rect 505642 936966 505654 937018
rect 505706 937015 505718 937018
rect 689210 937015 689222 937018
rect 505706 936969 689222 937015
rect 505706 936966 505718 936969
rect 689210 936966 689222 936969
rect 689274 936966 689286 937018
rect 453562 936854 453574 936906
rect 453626 936903 453638 936906
rect 687306 936903 687318 936906
rect 453626 936857 687318 936903
rect 453626 936854 453638 936857
rect 687306 936854 687318 936857
rect 687370 936854 687382 936906
rect 450202 936742 450214 936794
rect 450266 936791 450278 936794
rect 687642 936791 687654 936794
rect 450266 936745 687654 936791
rect 450266 936742 450278 936745
rect 687642 936742 687654 936745
rect 687706 936742 687718 936794
rect 344698 936630 344710 936682
rect 344762 936679 344774 936682
rect 687530 936679 687542 936682
rect 344762 936633 687542 936679
rect 344762 936630 344774 936633
rect 687530 936630 687542 936633
rect 687594 936630 687606 936682
rect 84746 936518 84758 936570
rect 84810 936567 84822 936570
rect 141530 936567 141542 936570
rect 84810 936521 141542 936567
rect 84810 936518 84822 936521
rect 141530 936518 141542 936521
rect 141594 936518 141606 936570
rect 233818 936518 233830 936570
rect 233882 936567 233894 936570
rect 688090 936567 688102 936570
rect 233882 936521 688102 936567
rect 233882 936518 233894 936521
rect 688090 936518 688102 936521
rect 688154 936518 688166 936570
rect 176698 935622 176710 935674
rect 176762 935671 176774 935674
rect 185770 935671 185782 935674
rect 176762 935625 185782 935671
rect 176762 935622 176774 935625
rect 185770 935622 185782 935625
rect 185834 935622 185846 935674
rect 176474 935398 176486 935450
rect 176538 935447 176550 935450
rect 208058 935447 208070 935450
rect 176538 935401 208070 935447
rect 176538 935398 176550 935401
rect 208058 935398 208070 935401
rect 208122 935398 208134 935450
rect 630410 935398 630422 935450
rect 630474 935447 630486 935450
rect 674090 935447 674102 935450
rect 630474 935401 674102 935447
rect 630474 935398 630486 935401
rect 674090 935398 674102 935401
rect 674154 935398 674166 935450
rect 341002 935286 341014 935338
rect 341066 935286 341078 935338
rect 289146 935174 289158 935226
rect 289210 935223 289222 935226
rect 296314 935223 296326 935226
rect 289210 935177 296326 935223
rect 289210 935174 289222 935177
rect 296314 935174 296326 935177
rect 296378 935174 296390 935226
rect 282426 935062 282438 935114
rect 282490 935111 282502 935114
rect 318938 935111 318950 935114
rect 282490 935065 318950 935111
rect 282490 935062 282502 935065
rect 318938 935062 318950 935065
rect 319002 935062 319014 935114
rect 341017 934999 341063 935286
rect 385242 934999 385254 935002
rect 341017 934953 385254 934999
rect 385242 934950 385254 934953
rect 385306 934950 385318 935002
rect 497354 934950 497366 935002
rect 497418 934999 497430 935002
rect 507434 934999 507446 935002
rect 497418 934953 507446 934999
rect 497418 934950 497430 934953
rect 507434 934950 507446 934953
rect 507498 934950 507510 935002
rect 342570 934838 342582 934890
rect 342634 934887 342646 934890
rect 407418 934887 407430 934890
rect 342634 934841 407430 934887
rect 342634 934838 342646 934841
rect 407418 934838 407430 934841
rect 407482 934838 407494 934890
rect 453338 934838 453350 934890
rect 453402 934887 453414 934890
rect 458490 934887 458502 934890
rect 453402 934841 458502 934887
rect 453402 934838 453414 934841
rect 458490 934838 458502 934841
rect 458554 934838 458566 934890
rect 700410 739062 700422 739114
rect 700474 739111 700486 739114
rect 701306 739111 701318 739114
rect 700474 739065 701318 739111
rect 700474 739062 700486 739065
rect 701306 739062 701318 739065
rect 701370 739062 701382 739114
rect 700410 712070 700422 712122
rect 700474 712119 700486 712122
rect 704554 712119 704566 712122
rect 700474 712073 704566 712119
rect 700474 712070 700486 712073
rect 704554 712070 704566 712073
rect 704618 712070 704630 712122
rect 72986 618102 72998 618154
rect 73050 618102 73062 618154
rect 73434 618102 73446 618154
rect 73498 618151 73510 618154
rect 77690 618151 77702 618154
rect 73498 618105 77702 618151
rect 73498 618102 73510 618105
rect 77690 618102 77702 618105
rect 77754 618102 77766 618154
rect 73001 618039 73047 618102
rect 78362 618039 78374 618042
rect 73001 617993 78374 618039
rect 78362 617990 78374 617993
rect 78426 617990 78438 618042
rect 73210 536118 73222 536170
rect 73274 536118 73286 536170
rect 73225 535831 73271 536118
rect 77466 535831 77478 535834
rect 73225 535785 77478 535831
rect 77466 535782 77478 535785
rect 77530 535782 77542 535834
rect 72986 413142 72998 413194
rect 73050 413191 73062 413194
rect 78250 413191 78262 413194
rect 73050 413145 78262 413191
rect 73050 413142 73062 413145
rect 78250 413142 78262 413145
rect 78314 413142 78326 413194
rect 73434 413030 73446 413082
rect 73498 413079 73510 413082
rect 78362 413079 78374 413082
rect 73498 413033 78374 413079
rect 73498 413030 73510 413033
rect 78362 413030 78374 413033
rect 78426 413030 78438 413082
rect 284218 333510 284230 333562
rect 284282 333559 284294 333562
rect 423882 333559 423894 333562
rect 284282 333513 423894 333559
rect 284282 333510 284294 333513
rect 423882 333510 423894 333513
rect 423946 333510 423958 333562
rect 266522 333398 266534 333450
rect 266586 333447 266598 333450
rect 376282 333447 376294 333450
rect 266586 333401 376294 333447
rect 266586 333398 266598 333401
rect 376282 333398 376294 333401
rect 376346 333398 376358 333450
rect 403386 333398 403398 333450
rect 403450 333447 403462 333450
rect 465546 333447 465558 333450
rect 403450 333401 465558 333447
rect 403450 333398 403462 333401
rect 465546 333398 465558 333401
rect 465610 333398 465622 333450
rect 611034 333398 611046 333450
rect 611098 333447 611110 333450
rect 688090 333447 688102 333450
rect 611098 333401 688102 333447
rect 611098 333398 611110 333401
rect 688090 333398 688102 333401
rect 688154 333398 688166 333450
rect 369674 333286 369686 333338
rect 369738 333335 369750 333338
rect 483802 333335 483814 333338
rect 369738 333289 483814 333335
rect 369738 333286 369750 333289
rect 483802 333286 483814 333289
rect 483866 333286 483878 333338
rect 488394 333286 488406 333338
rect 488458 333335 488470 333338
rect 632426 333335 632438 333338
rect 488458 333289 632438 333335
rect 488458 333286 488470 333289
rect 632426 333286 632438 333289
rect 632490 333286 632502 333338
rect 139178 333174 139190 333226
rect 139242 333223 139254 333226
rect 179834 333223 179846 333226
rect 139242 333177 179846 333223
rect 139242 333174 139254 333177
rect 179834 333174 179846 333177
rect 179898 333174 179910 333226
rect 269098 333174 269110 333226
rect 269162 333223 269174 333226
rect 382106 333223 382118 333226
rect 269162 333177 382118 333223
rect 269162 333174 269174 333177
rect 382106 333174 382118 333177
rect 382170 333174 382182 333226
rect 454794 333174 454806 333226
rect 454858 333223 454870 333226
rect 596698 333223 596710 333226
rect 454858 333177 596710 333223
rect 454858 333174 454870 333177
rect 596698 333174 596710 333177
rect 596762 333174 596774 333226
rect 132570 333062 132582 333114
rect 132634 333111 132646 333114
rect 177706 333111 177718 333114
rect 132634 333065 177718 333111
rect 132634 333062 132646 333065
rect 177706 333062 177718 333065
rect 177770 333062 177782 333114
rect 221386 333062 221398 333114
rect 221450 333111 221462 333114
rect 251626 333111 251638 333114
rect 221450 333065 251638 333111
rect 221450 333062 221462 333065
rect 251626 333062 251638 333065
rect 251690 333062 251702 333114
rect 275370 333062 275382 333114
rect 275434 333111 275446 333114
rect 400698 333111 400710 333114
rect 275434 333065 400710 333111
rect 275434 333062 275446 333065
rect 400698 333062 400710 333065
rect 400762 333062 400774 333114
rect 420858 333062 420870 333114
rect 420922 333111 420934 333114
rect 502058 333111 502070 333114
rect 420922 333065 502070 333111
rect 420922 333062 420934 333065
rect 502058 333062 502070 333065
rect 502122 333062 502134 333114
rect 102666 332950 102678 333002
rect 102730 332999 102742 333002
rect 151946 332999 151958 333002
rect 102730 332953 151958 332999
rect 102730 332950 102742 332953
rect 151946 332950 151958 332953
rect 152010 332950 152022 333002
rect 154410 332950 154422 333002
rect 154474 332999 154486 333002
rect 184986 332999 184998 333002
rect 154474 332953 184998 332999
rect 154474 332950 154486 332953
rect 184986 332950 184998 332953
rect 185050 332950 185062 333002
rect 196074 332950 196086 333002
rect 196138 332999 196150 333002
rect 200218 332999 200230 333002
rect 196138 332953 200230 332999
rect 196138 332950 196150 332953
rect 200218 332950 200230 332953
rect 200282 332950 200294 333002
rect 223626 332950 223638 333002
rect 223690 332999 223702 333002
rect 257562 332999 257574 333002
rect 223690 332953 257574 332999
rect 223690 332950 223702 332953
rect 257562 332950 257574 332953
rect 257626 332950 257638 333002
rect 320058 332950 320070 333002
rect 320122 332999 320134 333002
rect 448298 332999 448310 333002
rect 320122 332953 448310 332999
rect 320122 332950 320134 332953
rect 448298 332950 448310 332953
rect 448362 332950 448374 333002
rect 471146 332950 471158 333002
rect 471210 332999 471222 333002
rect 615290 332999 615302 333002
rect 471210 332953 615302 332999
rect 471210 332950 471222 332953
rect 615290 332950 615302 332953
rect 615354 332950 615366 333002
rect 110618 332838 110630 332890
rect 110682 332887 110694 332890
rect 167962 332887 167974 332890
rect 110682 332841 167974 332887
rect 110682 332838 110694 332841
rect 167962 332838 167974 332841
rect 168026 332838 168038 332890
rect 188010 332838 188022 332890
rect 188074 332887 188086 332890
rect 196634 332887 196646 332890
rect 188074 332841 196646 332887
rect 188074 332838 188086 332841
rect 196634 332838 196646 332841
rect 196698 332838 196710 332890
rect 227210 332838 227222 332890
rect 227274 332887 227286 332890
rect 271450 332887 271462 332890
rect 227274 332841 271462 332887
rect 227274 332838 227286 332841
rect 271450 332838 271462 332841
rect 271514 332838 271526 332890
rect 279738 332838 279750 332890
rect 279802 332887 279814 332890
rect 412570 332887 412582 332890
rect 279802 332841 412582 332887
rect 279802 332838 279814 332841
rect 412570 332838 412582 332841
rect 412634 332838 412646 332890
rect 437546 332838 437558 332890
rect 437610 332887 437622 332890
rect 585498 332887 585510 332890
rect 437610 332841 585510 332887
rect 437610 332838 437622 332841
rect 585498 332838 585510 332841
rect 585562 332838 585574 332890
rect 90794 332726 90806 332778
rect 90858 332775 90870 332778
rect 150602 332775 150614 332778
rect 90858 332729 150614 332775
rect 90858 332726 90870 332729
rect 150602 332726 150614 332729
rect 150666 332726 150678 332778
rect 152394 332726 152406 332778
rect 152458 332775 152470 332778
rect 183530 332775 183542 332778
rect 152458 332729 183542 332775
rect 152458 332726 152470 332729
rect 183530 332726 183542 332729
rect 183594 332726 183606 332778
rect 190138 332726 190150 332778
rect 190202 332775 190214 332778
rect 197866 332775 197878 332778
rect 190202 332729 197878 332775
rect 190202 332726 190214 332729
rect 197866 332726 197878 332729
rect 197930 332726 197942 332778
rect 205370 332726 205382 332778
rect 205434 332775 205446 332778
rect 211866 332775 211878 332778
rect 205434 332729 211878 332775
rect 205434 332726 205446 332729
rect 211866 332726 211878 332729
rect 211930 332726 211942 332778
rect 212090 332726 212102 332778
rect 212154 332775 212166 332778
rect 229786 332775 229798 332778
rect 212154 332729 229798 332775
rect 212154 332726 212166 332729
rect 229786 332726 229798 332729
rect 229850 332726 229862 332778
rect 231578 332726 231590 332778
rect 231642 332775 231654 332778
rect 283434 332775 283446 332778
rect 231642 332729 283446 332775
rect 231642 332726 231654 332729
rect 283434 332726 283446 332729
rect 283498 332726 283510 332778
rect 288474 332726 288486 332778
rect 288538 332775 288550 332778
rect 436426 332775 436438 332778
rect 288538 332729 436438 332775
rect 288538 332726 288550 332729
rect 436426 332726 436438 332729
rect 436490 332726 436502 332778
rect 471370 332726 471382 332778
rect 471434 332775 471446 332778
rect 621226 332775 621238 332778
rect 471434 332729 621238 332775
rect 471434 332726 471446 332729
rect 621226 332726 621238 332729
rect 621290 332726 621302 332778
rect 86874 332614 86886 332666
rect 86938 332663 86950 332666
rect 160234 332663 160246 332666
rect 86938 332617 160246 332663
rect 86938 332614 86950 332617
rect 160234 332614 160246 332617
rect 160298 332614 160310 332666
rect 192154 332614 192166 332666
rect 192218 332663 192230 332666
rect 199546 332663 199558 332666
rect 192218 332617 199558 332663
rect 192218 332614 192230 332617
rect 199546 332614 199558 332617
rect 199610 332614 199622 332666
rect 206826 332614 206838 332666
rect 206890 332663 206902 332666
rect 213882 332663 213894 332666
rect 206890 332617 213894 332663
rect 206890 332614 206902 332617
rect 213882 332614 213894 332617
rect 213946 332614 213958 332666
rect 217466 332614 217478 332666
rect 217530 332663 217542 332666
rect 233706 332663 233718 332666
rect 217530 332617 233718 332663
rect 217530 332614 217542 332617
rect 233706 332614 233718 332617
rect 233770 332614 233782 332666
rect 233930 332614 233942 332666
rect 233994 332663 234006 332666
rect 289370 332663 289382 332666
rect 233994 332617 289382 332663
rect 233994 332614 234006 332617
rect 289370 332614 289382 332617
rect 289434 332614 289446 332666
rect 421306 332614 421318 332666
rect 421370 332663 421382 332666
rect 573514 332663 573526 332666
rect 421370 332617 573526 332663
rect 421370 332614 421382 332617
rect 573514 332614 573526 332617
rect 573578 332614 573590 332666
rect 78810 332502 78822 332554
rect 78874 332551 78886 332554
rect 672298 332551 672310 332554
rect 78874 332505 672310 332551
rect 78874 332502 78886 332505
rect 672298 332502 672310 332505
rect 672362 332502 672374 332554
rect 327226 332390 327238 332442
rect 327290 332439 327302 332442
rect 541706 332439 541718 332442
rect 327290 332393 541718 332439
rect 327290 332390 327302 332393
rect 541706 332390 541718 332393
rect 541770 332390 541782 332442
rect 331482 332278 331494 332330
rect 331546 332327 331558 332330
rect 553690 332327 553702 332330
rect 331546 332281 553702 332327
rect 331546 332278 331558 332281
rect 553690 332278 553702 332281
rect 553754 332278 553766 332330
rect 278954 332166 278966 332218
rect 279018 332215 279030 332218
rect 410554 332215 410566 332218
rect 279018 332169 410566 332215
rect 279018 332166 279030 332169
rect 410554 332166 410566 332169
rect 410618 332166 410630 332218
rect 411338 332166 411350 332218
rect 411402 332215 411414 332218
rect 653034 332215 653046 332218
rect 411402 332169 653046 332215
rect 411402 332166 411414 332169
rect 653034 332166 653046 332169
rect 653098 332166 653110 332218
rect 343802 332054 343814 332106
rect 343866 332103 343878 332106
rect 587402 332103 587414 332106
rect 343866 332057 587414 332103
rect 343866 332054 343878 332057
rect 587402 332054 587414 332057
rect 587466 332054 587478 332106
rect 352538 331942 352550 331994
rect 352602 331991 352614 331994
rect 611258 331991 611270 331994
rect 352602 331945 611270 331991
rect 352602 331942 352614 331945
rect 611258 331942 611270 331945
rect 611322 331942 611334 331994
rect 379306 331830 379318 331882
rect 379370 331879 379382 331882
rect 676890 331879 676902 331882
rect 379370 331833 676902 331879
rect 379370 331830 379382 331833
rect 676890 331830 676902 331833
rect 676954 331830 676966 331882
rect 80042 331718 80054 331770
rect 80106 331767 80118 331770
rect 672410 331767 672422 331770
rect 80106 331721 672422 331767
rect 80106 331718 80118 331721
rect 672410 331718 672422 331721
rect 672474 331718 672486 331770
rect 325994 331606 326006 331658
rect 326058 331655 326070 331658
rect 539802 331655 539814 331658
rect 326058 331609 539814 331655
rect 326058 331606 326070 331609
rect 539802 331606 539814 331609
rect 539866 331606 539878 331658
rect 319834 331494 319846 331546
rect 319898 331543 319910 331546
rect 523898 331543 523910 331546
rect 319898 331497 523910 331543
rect 319898 331494 319910 331497
rect 523898 331494 523910 331497
rect 523962 331494 523974 331546
rect 283322 331382 283334 331434
rect 283386 331431 283398 331434
rect 422538 331431 422550 331434
rect 283386 331385 422550 331431
rect 283386 331382 283398 331385
rect 422538 331382 422550 331385
rect 422602 331382 422614 331434
rect 281194 331270 281206 331322
rect 281258 331319 281270 331322
rect 416602 331319 416614 331322
rect 281258 331273 416614 331319
rect 281258 331270 281270 331273
rect 416602 331270 416614 331273
rect 416666 331270 416678 331322
rect 276826 331158 276838 331210
rect 276890 331207 276902 331210
rect 404618 331207 404630 331210
rect 276890 331161 404630 331207
rect 276890 331158 276902 331161
rect 404618 331158 404630 331161
rect 404682 331158 404694 331210
rect 73210 331046 73222 331098
rect 73274 331046 73286 331098
rect 73225 330871 73271 331046
rect 78250 330871 78262 330874
rect 73225 330825 78262 330871
rect 78250 330822 78262 330825
rect 78314 330822 78326 330874
rect 294298 330822 294310 330874
rect 294362 330871 294374 330874
rect 452330 330871 452342 330874
rect 294362 330825 452342 330871
rect 294362 330822 294374 330825
rect 452330 330822 452342 330825
rect 452394 330822 452406 330874
rect 298666 330710 298678 330762
rect 298730 330759 298742 330762
rect 464202 330759 464214 330762
rect 298730 330713 464214 330759
rect 298730 330710 298742 330713
rect 464202 330710 464214 330713
rect 464266 330710 464278 330762
rect 305162 330598 305174 330650
rect 305226 330647 305238 330650
rect 482122 330647 482134 330650
rect 305226 330601 482134 330647
rect 305226 330598 305238 330601
rect 482122 330598 482134 330601
rect 482186 330598 482198 330650
rect 309530 330486 309542 330538
rect 309594 330535 309606 330538
rect 494106 330535 494118 330538
rect 309594 330489 494118 330535
rect 309594 330486 309606 330489
rect 494106 330486 494118 330489
rect 494170 330486 494182 330538
rect 249386 330374 249398 330426
rect 249450 330423 249462 330426
rect 307290 330423 307302 330426
rect 249450 330377 307302 330423
rect 249450 330374 249462 330377
rect 307290 330374 307302 330377
rect 307354 330374 307366 330426
rect 313898 330374 313910 330426
rect 313962 330423 313974 330426
rect 505978 330423 505990 330426
rect 313962 330377 505990 330423
rect 313962 330374 313974 330377
rect 505978 330374 505990 330377
rect 506042 330374 506054 330426
rect 240202 330262 240214 330314
rect 240266 330311 240278 330314
rect 309306 330311 309318 330314
rect 240266 330265 309318 330311
rect 240266 330262 240278 330265
rect 309306 330262 309318 330265
rect 309370 330262 309382 330314
rect 322634 330262 322646 330314
rect 322698 330311 322710 330314
rect 529834 330311 529846 330314
rect 322698 330265 529846 330311
rect 322698 330262 322710 330265
rect 529834 330262 529846 330265
rect 529898 330262 529910 330314
rect 243226 330150 243238 330202
rect 243290 330199 243302 330202
rect 313226 330199 313238 330202
rect 243290 330153 313238 330199
rect 243290 330150 243302 330153
rect 313226 330150 313238 330153
rect 313290 330150 313302 330202
rect 354778 330150 354790 330202
rect 354842 330199 354854 330202
rect 617306 330199 617318 330202
rect 354842 330153 617318 330199
rect 354842 330150 354854 330153
rect 617306 330150 617318 330153
rect 617370 330150 617382 330202
rect 244010 330038 244022 330090
rect 244074 330087 244086 330090
rect 315242 330087 315254 330090
rect 244074 330041 315254 330087
rect 244074 330038 244086 330041
rect 315242 330038 315254 330041
rect 315306 330038 315318 330090
rect 354554 330038 354566 330090
rect 354618 330087 354630 330090
rect 619210 330087 619222 330090
rect 354618 330041 619222 330087
rect 354618 330038 354630 330041
rect 619210 330038 619222 330041
rect 619274 330038 619286 330090
rect 292058 329926 292070 329978
rect 292122 329975 292134 329978
rect 446394 329975 446406 329978
rect 292122 329929 446406 329975
rect 292122 329926 292134 329929
rect 446394 329926 446406 329929
rect 446458 329926 446470 329978
rect 289930 329814 289942 329866
rect 289994 329863 290006 329866
rect 421754 329863 421766 329866
rect 289994 329817 421766 329863
rect 289994 329814 290006 329817
rect 421754 329814 421766 329817
rect 421818 329814 421830 329866
rect 247706 329142 247718 329194
rect 247770 329191 247782 329194
rect 325210 329191 325222 329194
rect 247770 329145 325222 329191
rect 247770 329142 247782 329145
rect 325210 329142 325222 329145
rect 325274 329142 325286 329194
rect 353882 329142 353894 329194
rect 353946 329191 353958 329194
rect 577546 329191 577558 329194
rect 353946 329145 577558 329191
rect 353946 329142 353958 329145
rect 577546 329142 577558 329145
rect 577610 329142 577622 329194
rect 248490 329030 248502 329082
rect 248554 329079 248566 329082
rect 327114 329079 327126 329082
rect 248554 329033 327126 329079
rect 248554 329030 248566 329033
rect 327114 329030 327126 329033
rect 327178 329030 327190 329082
rect 335290 329030 335302 329082
rect 335354 329079 335366 329082
rect 563658 329079 563670 329082
rect 335354 329033 563670 329079
rect 335354 329030 335366 329033
rect 563658 329030 563670 329033
rect 563722 329030 563734 329082
rect 250618 328918 250630 328970
rect 250682 328967 250694 328970
rect 333050 328967 333062 328970
rect 250682 328921 333062 328967
rect 250682 328918 250694 328921
rect 333050 328918 333062 328921
rect 333114 328918 333126 328970
rect 346714 328918 346726 328970
rect 346778 328967 346790 328970
rect 595354 328967 595366 328970
rect 346778 328921 595366 328967
rect 346778 328918 346790 328921
rect 595354 328918 595366 328921
rect 595418 328918 595430 328970
rect 128538 328806 128550 328858
rect 128602 328855 128614 328858
rect 175466 328855 175478 328858
rect 128602 328809 175478 328855
rect 128602 328806 128614 328809
rect 175466 328806 175478 328809
rect 175530 328806 175542 328858
rect 252858 328806 252870 328858
rect 252922 328855 252934 328858
rect 339098 328855 339110 328858
rect 252922 328809 339110 328855
rect 252922 328806 252934 328809
rect 339098 328806 339110 328809
rect 339162 328806 339174 328858
rect 351194 328806 351206 328858
rect 351258 328855 351270 328858
rect 607338 328855 607350 328858
rect 351258 328809 607350 328855
rect 351258 328806 351270 328809
rect 607338 328806 607350 328809
rect 607402 328806 607414 328858
rect 256442 328694 256454 328746
rect 256506 328743 256518 328746
rect 348954 328743 348966 328746
rect 256506 328697 348966 328743
rect 256506 328694 256518 328697
rect 348954 328694 348966 328697
rect 349018 328694 349030 328746
rect 357690 328694 357702 328746
rect 357754 328743 357766 328746
rect 625258 328743 625270 328746
rect 357754 328697 625270 328743
rect 357754 328694 357766 328697
rect 625258 328694 625270 328697
rect 625322 328694 625334 328746
rect 124618 328582 124630 328634
rect 124682 328631 124694 328634
rect 174794 328631 174806 328634
rect 124682 328585 174806 328631
rect 124682 328582 124694 328585
rect 174794 328582 174806 328585
rect 174858 328582 174870 328634
rect 260810 328582 260822 328634
rect 260874 328631 260886 328634
rect 360938 328631 360950 328634
rect 260874 328585 360950 328631
rect 260874 328582 260886 328585
rect 360938 328582 360950 328585
rect 361002 328582 361014 328634
rect 362170 328582 362182 328634
rect 362234 328631 362246 328634
rect 637130 328631 637142 328634
rect 362234 328585 637142 328631
rect 362234 328582 362246 328585
rect 637130 328582 637142 328585
rect 637194 328582 637206 328634
rect 120586 328470 120598 328522
rect 120650 328519 120662 328522
rect 172554 328519 172566 328522
rect 120650 328473 172566 328519
rect 120650 328470 120662 328473
rect 172554 328470 172566 328473
rect 172618 328470 172630 328522
rect 267418 328470 267430 328522
rect 267482 328519 267494 328522
rect 378858 328519 378870 328522
rect 267482 328473 378870 328519
rect 267482 328470 267494 328473
rect 378858 328470 378870 328473
rect 378922 328470 378934 328522
rect 384682 328470 384694 328522
rect 384746 328519 384758 328522
rect 664906 328519 664918 328522
rect 384746 328473 664918 328519
rect 384746 328470 384758 328473
rect 664906 328470 664918 328473
rect 664970 328470 664982 328522
rect 122490 328358 122502 328410
rect 122554 328407 122566 328410
rect 173338 328407 173350 328410
rect 122554 328361 173350 328407
rect 122554 328358 122566 328361
rect 173338 328358 173350 328361
rect 173402 328358 173414 328410
rect 263050 328358 263062 328410
rect 263114 328407 263126 328410
rect 366874 328407 366886 328410
rect 263114 328361 366886 328407
rect 263114 328358 263126 328361
rect 366874 328358 366886 328361
rect 366938 328358 366950 328410
rect 369562 328358 369574 328410
rect 369626 328407 369638 328410
rect 655050 328407 655062 328410
rect 369626 328361 655062 328407
rect 369626 328358 369638 328361
rect 655050 328358 655062 328361
rect 655114 328358 655126 328410
rect 231018 328246 231030 328298
rect 231082 328295 231094 328298
rect 279402 328295 279414 328298
rect 231082 328249 279414 328295
rect 231082 328246 231094 328249
rect 279402 328246 279414 328249
rect 279466 328246 279478 328298
rect 319050 328246 319062 328298
rect 319114 328295 319126 328298
rect 519866 328295 519878 328298
rect 319114 328249 519878 328295
rect 319114 328246 319126 328249
rect 519866 328246 519878 328249
rect 519930 328246 519942 328298
rect 228778 328134 228790 328186
rect 228842 328183 228854 328186
rect 273466 328183 273478 328186
rect 228842 328137 273478 328183
rect 228842 328134 228854 328137
rect 273466 328134 273478 328137
rect 273530 328134 273542 328186
rect 301690 328134 301702 328186
rect 301754 328183 301766 328186
rect 472154 328183 472166 328186
rect 301754 328137 472166 328183
rect 301754 328134 301766 328137
rect 472154 328134 472166 328137
rect 472218 328134 472230 328186
rect 228106 328022 228118 328074
rect 228170 328071 228182 328074
rect 269546 328071 269558 328074
rect 228170 328025 269558 328071
rect 228170 328022 228182 328025
rect 269546 328022 269558 328025
rect 269610 328022 269622 328074
rect 276154 328022 276166 328074
rect 276218 328071 276230 328074
rect 402602 328071 402614 328074
rect 276218 328025 402614 328071
rect 276218 328022 276230 328025
rect 402602 328022 402614 328025
rect 402666 328022 402678 328074
rect 226650 327910 226662 327962
rect 226714 327959 226726 327962
rect 267530 327959 267542 327962
rect 226714 327913 267542 327959
rect 226714 327910 226726 327913
rect 267530 327910 267542 327913
rect 267594 327910 267606 327962
rect 297210 327910 297222 327962
rect 297274 327959 297286 327962
rect 386026 327959 386038 327962
rect 297274 327913 386038 327959
rect 297274 327910 297286 327913
rect 386026 327910 386038 327913
rect 386090 327910 386102 327962
rect 289258 327462 289270 327514
rect 289322 327511 289334 327514
rect 438442 327511 438454 327514
rect 289322 327465 438454 327511
rect 289322 327462 289334 327465
rect 438442 327462 438454 327465
rect 438506 327462 438518 327514
rect 306730 327350 306742 327402
rect 306794 327399 306806 327402
rect 486154 327399 486166 327402
rect 306794 327353 486166 327399
rect 306794 327350 306806 327353
rect 486154 327350 486166 327353
rect 486218 327350 486230 327402
rect 313338 327238 313350 327290
rect 313402 327287 313414 327290
rect 503962 327287 503974 327290
rect 313402 327241 503974 327287
rect 313402 327238 313414 327241
rect 503962 327238 503974 327241
rect 504026 327238 504038 327290
rect 315466 327126 315478 327178
rect 315530 327175 315542 327178
rect 509898 327175 509910 327178
rect 315530 327129 509910 327175
rect 315530 327126 315542 327129
rect 509898 327126 509910 327129
rect 509962 327126 509974 327178
rect 322074 327014 322086 327066
rect 322138 327063 322150 327066
rect 527818 327063 527830 327066
rect 322138 327017 527830 327063
rect 322138 327014 322150 327017
rect 527818 327014 527830 327017
rect 527882 327014 527894 327066
rect 333050 326902 333062 326954
rect 333114 326951 333126 326954
rect 557610 326951 557622 326954
rect 333114 326905 557622 326951
rect 333114 326902 333126 326905
rect 557610 326902 557622 326905
rect 557674 326902 557686 326954
rect 348282 326790 348294 326842
rect 348346 326839 348358 326842
rect 599386 326839 599398 326842
rect 348346 326793 599398 326839
rect 348346 326790 348358 326793
rect 599386 326790 599398 326793
rect 599450 326790 599462 326842
rect 363626 326678 363638 326730
rect 363690 326727 363702 326730
rect 641050 326727 641062 326730
rect 363690 326681 641062 326727
rect 363690 326678 363702 326681
rect 641050 326678 641062 326681
rect 641114 326678 641126 326730
rect 284890 326566 284902 326618
rect 284954 326615 284966 326618
rect 426458 326615 426470 326618
rect 284954 326569 426470 326615
rect 284954 326566 284966 326569
rect 426458 326566 426470 326569
rect 426522 326566 426534 326618
rect 280410 326454 280422 326506
rect 280474 326503 280486 326506
rect 414586 326503 414598 326506
rect 280474 326457 414598 326503
rect 280474 326454 280486 326457
rect 414586 326454 414598 326457
rect 414650 326454 414662 326506
rect 299786 326342 299798 326394
rect 299850 326391 299862 326394
rect 432506 326391 432518 326394
rect 299850 326345 432518 326391
rect 299850 326342 299862 326345
rect 432506 326342 432518 326345
rect 432570 326342 432582 326394
rect 351978 325782 351990 325834
rect 352042 325831 352054 325834
rect 454682 325831 454694 325834
rect 352042 325785 454694 325831
rect 352042 325782 352054 325785
rect 454682 325782 454694 325785
rect 454746 325782 454758 325834
rect 312554 325670 312566 325722
rect 312618 325719 312630 325722
rect 420858 325719 420870 325722
rect 312618 325673 420870 325719
rect 312618 325670 312630 325673
rect 420858 325670 420870 325673
rect 420922 325670 420934 325722
rect 264506 325558 264518 325610
rect 264570 325607 264582 325610
rect 319722 325607 319734 325610
rect 264570 325561 319734 325607
rect 264570 325558 264582 325561
rect 319722 325558 319734 325561
rect 319786 325558 319798 325610
rect 356346 325558 356358 325610
rect 356410 325607 356422 325610
rect 471370 325607 471382 325610
rect 356410 325561 471382 325607
rect 356410 325558 356422 325561
rect 471370 325558 471382 325561
rect 471434 325558 471446 325610
rect 485482 325558 485494 325610
rect 485546 325607 485558 325610
rect 668602 325607 668614 325610
rect 485546 325561 668614 325607
rect 485546 325558 485558 325561
rect 668602 325558 668614 325561
rect 668666 325558 668678 325610
rect 310426 325446 310438 325498
rect 310490 325495 310502 325498
rect 495562 325495 495574 325498
rect 310490 325449 495574 325495
rect 310490 325446 310502 325449
rect 495562 325446 495574 325449
rect 495626 325446 495638 325498
rect 314794 325334 314806 325386
rect 314858 325383 314870 325386
rect 507322 325383 507334 325386
rect 314858 325337 507334 325383
rect 314858 325334 314870 325337
rect 507322 325334 507334 325337
rect 507386 325334 507398 325386
rect 262266 325222 262278 325274
rect 262330 325271 262342 325274
rect 320170 325271 320182 325274
rect 262330 325225 320182 325271
rect 262330 325222 262342 325225
rect 320170 325222 320182 325225
rect 320234 325222 320246 325274
rect 323530 325222 323542 325274
rect 323594 325271 323606 325274
rect 530842 325271 530854 325274
rect 323594 325225 530854 325271
rect 323594 325222 323606 325225
rect 530842 325222 530854 325225
rect 530906 325222 530918 325274
rect 271786 325110 271798 325162
rect 271850 325159 271862 325162
rect 335066 325159 335078 325162
rect 271850 325113 335078 325159
rect 271850 325110 271862 325113
rect 335066 325110 335078 325113
rect 335130 325110 335142 325162
rect 362730 325110 362742 325162
rect 362794 325159 362806 325162
rect 638362 325159 638374 325162
rect 362794 325113 638374 325159
rect 362794 325110 362806 325113
rect 638362 325110 638374 325113
rect 638426 325110 638438 325162
rect 265962 324998 265974 325050
rect 266026 325047 266038 325050
rect 335178 325047 335190 325050
rect 266026 325001 335190 325047
rect 266026 324998 266038 325001
rect 335178 324998 335190 325001
rect 335242 324998 335254 325050
rect 365082 324998 365094 325050
rect 365146 325047 365158 325050
rect 645082 325047 645094 325050
rect 365146 325001 645094 325047
rect 365146 324998 365158 325001
rect 645082 324998 645094 325001
rect 645146 324998 645158 325050
rect 343242 324886 343254 324938
rect 343306 324935 343318 324938
rect 437546 324935 437558 324938
rect 343306 324889 437558 324935
rect 343306 324886 343318 324889
rect 437546 324886 437558 324889
rect 437610 324886 437622 324938
rect 338874 324774 338886 324826
rect 338938 324823 338950 324826
rect 421306 324823 421318 324826
rect 338938 324777 421318 324823
rect 338938 324774 338950 324777
rect 421306 324774 421318 324777
rect 421370 324774 421382 324826
rect 340890 324662 340902 324714
rect 340954 324711 340966 324714
rect 421082 324711 421094 324714
rect 340954 324665 421094 324711
rect 340954 324662 340966 324665
rect 421082 324662 421094 324665
rect 421146 324662 421158 324714
rect 161354 324214 161366 324266
rect 161418 324263 161430 324266
rect 162586 324263 162598 324266
rect 161418 324217 162598 324263
rect 161418 324214 161430 324217
rect 162586 324214 162598 324217
rect 162650 324214 162662 324266
rect 280634 324214 280646 324266
rect 280698 324263 280710 324266
rect 281922 324263 281934 324266
rect 280698 324217 281934 324263
rect 280698 324214 280710 324217
rect 281922 324214 281934 324217
rect 281986 324214 281998 324266
rect 354554 324214 354566 324266
rect 354618 324263 354630 324266
rect 355506 324263 355518 324266
rect 354618 324217 355518 324263
rect 354618 324214 354630 324217
rect 355506 324214 355518 324217
rect 355570 324214 355582 324266
rect 95722 324102 95734 324154
rect 95786 324151 95798 324154
rect 155194 324151 155206 324154
rect 95786 324105 155206 324151
rect 95786 324102 95798 324105
rect 155194 324102 155206 324105
rect 155258 324102 155270 324154
rect 155418 324102 155430 324154
rect 155482 324151 155494 324154
rect 163202 324151 163214 324154
rect 155482 324105 163214 324151
rect 155482 324102 155494 324105
rect 163202 324102 163214 324105
rect 163266 324102 163278 324154
rect 203354 324102 203366 324154
rect 203418 324151 203430 324154
rect 204642 324151 204654 324154
rect 203418 324105 204654 324151
rect 203418 324102 203430 324105
rect 204642 324102 204654 324105
rect 204706 324102 204718 324154
rect 375218 324102 375230 324154
rect 375282 324151 375294 324154
rect 377850 324151 377862 324154
rect 375282 324105 377862 324151
rect 375282 324102 375294 324105
rect 377850 324102 377862 324105
rect 377914 324102 377926 324154
rect 133690 323990 133702 324042
rect 133754 324039 133766 324042
rect 164658 324039 164670 324042
rect 133754 323993 164670 324039
rect 133754 323990 133766 323993
rect 164658 323990 164670 323993
rect 164722 323990 164734 324042
rect 372306 323990 372318 324042
rect 372370 324039 372382 324042
rect 384682 324039 384694 324042
rect 372370 323993 384694 324039
rect 372370 323990 372382 323993
rect 384682 323990 384694 323993
rect 384746 323990 384758 324042
rect 94042 323878 94054 323930
rect 94106 323927 94118 323930
rect 155306 323927 155318 323930
rect 94106 323881 155318 323927
rect 94106 323878 94118 323881
rect 155306 323878 155318 323881
rect 155370 323878 155382 323930
rect 163874 323927 163886 323930
rect 155433 323881 163886 323927
rect 155194 323766 155206 323818
rect 155258 323815 155270 323818
rect 155433 323815 155479 323881
rect 163874 323878 163886 323881
rect 163938 323878 163950 323930
rect 287074 323878 287086 323930
rect 287138 323927 287150 323930
rect 299786 323927 299798 323930
rect 287138 323881 299798 323927
rect 287138 323878 287150 323881
rect 299786 323878 299798 323881
rect 299850 323878 299862 323930
rect 370066 323878 370078 323930
rect 370130 323927 370142 323930
rect 385466 323927 385478 323930
rect 370130 323881 385478 323927
rect 370130 323878 370142 323881
rect 385466 323878 385478 323881
rect 385530 323878 385542 323930
rect 155258 323769 155479 323815
rect 155258 323766 155270 323769
rect 673194 308807 673206 308810
rect 377305 308761 673206 308807
rect 377305 308698 377351 308761
rect 673194 308758 673206 308761
rect 673258 308758 673270 308810
rect 178042 308646 178054 308698
rect 178106 308695 178118 308698
rect 179666 308695 179678 308698
rect 178106 308649 179678 308695
rect 178106 308646 178118 308649
rect 179666 308646 179678 308649
rect 179730 308646 179742 308698
rect 228386 308646 228398 308698
rect 228450 308695 228462 308698
rect 228450 308649 231862 308695
rect 228450 308646 228462 308649
rect 231816 308583 231862 308649
rect 282314 308646 282326 308698
rect 282378 308695 282390 308698
rect 283826 308695 283838 308698
rect 282378 308649 283838 308695
rect 282378 308646 282390 308649
rect 283826 308646 283838 308649
rect 283890 308646 283902 308698
rect 315914 308646 315926 308698
rect 315978 308695 315990 308698
rect 317426 308695 317438 308698
rect 315978 308649 317438 308695
rect 315978 308646 315990 308649
rect 317426 308646 317438 308649
rect 317490 308646 317502 308698
rect 377290 308646 377302 308698
rect 377354 308646 377366 308698
rect 233818 308583 233830 308586
rect 231816 308537 233830 308583
rect 233818 308534 233830 308537
rect 233882 308534 233894 308586
rect 259522 308583 259534 308586
rect 258809 308537 259534 308583
rect 171434 308422 171446 308474
rect 171498 308471 171510 308474
rect 172946 308471 172958 308474
rect 171498 308425 172958 308471
rect 171498 308422 171510 308425
rect 172946 308422 172958 308425
rect 173010 308422 173022 308474
rect 208506 308422 208518 308474
rect 208570 308471 208582 308474
rect 216178 308471 216190 308474
rect 208570 308425 216190 308471
rect 208570 308422 208582 308425
rect 216178 308422 216190 308425
rect 216242 308422 216254 308474
rect 225362 308422 225374 308474
rect 225426 308471 225438 308474
rect 226762 308471 226774 308474
rect 225426 308425 226774 308471
rect 225426 308422 225438 308425
rect 226762 308422 226774 308425
rect 226826 308422 226838 308474
rect 227826 308422 227838 308474
rect 227890 308471 227902 308474
rect 231802 308471 231814 308474
rect 227890 308425 231814 308471
rect 227890 308422 227902 308425
rect 231802 308422 231814 308425
rect 231866 308422 231878 308474
rect 243562 308422 243574 308474
rect 243626 308471 243638 308474
rect 244850 308471 244862 308474
rect 243626 308425 244862 308471
rect 243626 308422 243638 308425
rect 244850 308422 244862 308425
rect 244914 308422 244926 308474
rect 247034 308422 247046 308474
rect 247098 308471 247110 308474
rect 248546 308471 248558 308474
rect 247098 308425 248558 308471
rect 247098 308422 247110 308425
rect 248546 308422 248558 308425
rect 248610 308422 248622 308474
rect 248714 308422 248726 308474
rect 248778 308471 248790 308474
rect 249778 308471 249790 308474
rect 248778 308425 249790 308471
rect 248778 308422 248790 308425
rect 249778 308422 249790 308425
rect 249842 308422 249854 308474
rect 253642 308422 253654 308474
rect 253706 308471 253718 308474
rect 255266 308471 255278 308474
rect 253706 308425 255278 308471
rect 253706 308422 253718 308425
rect 255266 308422 255278 308425
rect 255330 308422 255342 308474
rect 258809 308362 258855 308537
rect 259522 308534 259534 308537
rect 259586 308534 259598 308586
rect 326498 308534 326510 308586
rect 326562 308583 326574 308586
rect 327450 308583 327462 308586
rect 326562 308537 327462 308583
rect 326562 308534 326574 308537
rect 327450 308534 327462 308537
rect 327514 308534 327526 308586
rect 336074 308422 336086 308474
rect 336138 308471 336150 308474
rect 336914 308471 336926 308474
rect 336138 308425 336926 308471
rect 336138 308422 336150 308425
rect 336914 308422 336926 308425
rect 336978 308422 336990 308474
rect 337754 308422 337766 308474
rect 337818 308471 337830 308474
rect 338706 308471 338718 308474
rect 337818 308425 338718 308471
rect 337818 308422 337830 308425
rect 338706 308422 338718 308425
rect 338770 308422 338782 308474
rect 258794 308310 258806 308362
rect 258858 308310 258870 308362
rect 247930 308198 247942 308250
rect 247994 308247 248006 308250
rect 273914 308247 273926 308250
rect 247994 308201 273926 308247
rect 247994 308198 248006 308201
rect 273914 308198 273926 308201
rect 273978 308198 273990 308250
rect 191818 308086 191830 308138
rect 191882 308135 191894 308138
rect 208842 308135 208854 308138
rect 191882 308089 208854 308135
rect 191882 308086 191894 308089
rect 208842 308086 208854 308089
rect 208906 308086 208918 308138
rect 156202 307974 156214 308026
rect 156266 308023 156278 308026
rect 191594 308023 191606 308026
rect 156266 307977 191606 308023
rect 156266 307974 156278 307977
rect 191594 307974 191606 307977
rect 191658 307974 191670 308026
rect 235050 307974 235062 308026
rect 235114 308023 235126 308026
rect 247146 308023 247158 308026
rect 235114 307977 247158 308023
rect 235114 307974 235126 307977
rect 247146 307974 247158 307977
rect 247210 307974 247222 308026
rect 292506 307974 292518 308026
rect 292570 308023 292582 308026
rect 368218 308023 368230 308026
rect 292570 307977 368230 308023
rect 292570 307974 292582 307977
rect 368218 307974 368230 307977
rect 368282 307974 368294 308026
rect 95722 307862 95734 307914
rect 95786 307911 95798 307914
rect 163146 307911 163158 307914
rect 95786 307865 163158 307911
rect 95786 307862 95798 307865
rect 163146 307862 163158 307865
rect 163210 307862 163222 307914
rect 205146 307862 205158 307914
rect 205210 307911 205222 307914
rect 214890 307911 214902 307914
rect 205210 307865 214902 307911
rect 205210 307862 205222 307865
rect 214890 307862 214902 307865
rect 214954 307862 214966 307914
rect 243114 307862 243126 307914
rect 243178 307911 243190 307914
rect 263946 307911 263958 307914
rect 243178 307865 263958 307911
rect 243178 307862 243190 307865
rect 263946 307862 263958 307865
rect 264010 307862 264022 307914
rect 319274 307862 319286 307914
rect 319338 307911 319350 307914
rect 423322 307911 423334 307914
rect 319338 307865 423334 307911
rect 319338 307862 319350 307865
rect 423322 307862 423334 307865
rect 423386 307862 423398 307914
rect 97402 307750 97414 307802
rect 97466 307799 97478 307802
rect 163706 307799 163718 307802
rect 97466 307753 163718 307799
rect 97466 307750 97478 307753
rect 163706 307750 163718 307753
rect 163770 307750 163782 307802
rect 201562 307750 201574 307802
rect 201626 307799 201638 307802
rect 213098 307799 213110 307802
rect 201626 307753 213110 307799
rect 201626 307750 201638 307753
rect 213098 307750 213110 307753
rect 213162 307750 213174 307802
rect 235722 307750 235734 307802
rect 235786 307799 235798 307802
rect 248602 307799 248614 307802
rect 235786 307753 248614 307799
rect 235786 307750 235798 307753
rect 248602 307750 248614 307753
rect 248666 307750 248678 307802
rect 280298 307750 280310 307802
rect 280362 307799 280374 307802
rect 316586 307799 316598 307802
rect 280362 307753 316598 307799
rect 280362 307750 280374 307753
rect 316586 307750 316598 307753
rect 316650 307750 316662 307802
rect 327450 307750 327462 307802
rect 327514 307799 327526 307802
rect 440234 307799 440246 307802
rect 327514 307753 440246 307799
rect 327514 307750 327526 307753
rect 440234 307750 440246 307753
rect 440298 307750 440310 307802
rect 94266 307638 94278 307690
rect 94330 307687 94342 307690
rect 161914 307687 161926 307690
rect 94330 307641 161926 307687
rect 94330 307638 94342 307641
rect 161914 307638 161926 307641
rect 161978 307638 161990 307690
rect 166394 307638 166406 307690
rect 166458 307687 166470 307690
rect 196522 307687 196534 307690
rect 166458 307641 196534 307687
rect 166458 307638 166470 307641
rect 196522 307638 196534 307641
rect 196586 307638 196598 307690
rect 203354 307638 203366 307690
rect 203418 307687 203430 307690
rect 214330 307687 214342 307690
rect 203418 307641 214342 307687
rect 203418 307638 203430 307641
rect 214330 307638 214342 307641
rect 214394 307638 214406 307690
rect 236954 307638 236966 307690
rect 237018 307687 237030 307690
rect 250506 307687 250518 307690
rect 237018 307641 250518 307687
rect 237018 307638 237030 307641
rect 250506 307638 250518 307641
rect 250570 307638 250582 307690
rect 251626 307638 251638 307690
rect 251690 307687 251702 307690
rect 282202 307687 282214 307690
rect 251690 307641 282214 307687
rect 251690 307638 251702 307641
rect 282202 307638 282214 307641
rect 282266 307638 282278 307690
rect 337530 307638 337542 307690
rect 337594 307687 337606 307690
rect 467786 307687 467798 307690
rect 337594 307641 467798 307687
rect 337594 307638 337606 307641
rect 467786 307638 467798 307641
rect 467850 307638 467862 307690
rect 94042 307526 94054 307578
rect 94106 307575 94118 307578
rect 162474 307575 162486 307578
rect 94106 307529 162486 307575
rect 94106 307526 94118 307529
rect 162474 307526 162486 307529
rect 162538 307526 162550 307578
rect 187450 307575 187462 307578
rect 173016 307529 187462 307575
rect 147802 307414 147814 307466
rect 147866 307463 147878 307466
rect 173016 307463 173062 307529
rect 187450 307526 187462 307529
rect 187514 307526 187526 307578
rect 206714 307526 206726 307578
rect 206778 307575 206790 307578
rect 215562 307575 215574 307578
rect 206778 307529 215574 307575
rect 206778 307526 206790 307529
rect 215562 307526 215574 307529
rect 215626 307526 215638 307578
rect 239418 307526 239430 307578
rect 239482 307575 239494 307578
rect 257002 307575 257014 307578
rect 239482 307529 257014 307575
rect 239482 307526 239494 307529
rect 257002 307526 257014 307529
rect 257066 307526 257078 307578
rect 261930 307526 261942 307578
rect 261994 307575 262006 307578
rect 304042 307575 304054 307578
rect 261994 307529 304054 307575
rect 261994 307526 262006 307529
rect 304042 307526 304054 307529
rect 304106 307526 304118 307578
rect 357690 307526 357702 307578
rect 357754 307575 357766 307578
rect 509786 307575 509798 307578
rect 357754 307529 509798 307575
rect 357754 307526 357766 307529
rect 509786 307526 509798 307529
rect 509850 307526 509862 307578
rect 147866 307417 173062 307463
rect 147866 307414 147878 307417
rect 186778 307414 186790 307466
rect 186842 307463 186854 307466
rect 205818 307463 205830 307466
rect 186842 307417 205830 307463
rect 186842 307414 186854 307417
rect 205818 307414 205830 307417
rect 205882 307414 205894 307466
rect 226650 307414 226662 307466
rect 226714 307463 226726 307466
rect 230234 307463 230246 307466
rect 226714 307417 230246 307463
rect 226714 307414 226726 307417
rect 230234 307414 230246 307417
rect 230298 307414 230310 307466
rect 236394 307414 236406 307466
rect 236458 307463 236470 307466
rect 250282 307463 250294 307466
rect 236458 307417 250294 307463
rect 236458 307414 236470 307417
rect 250282 307414 250294 307417
rect 250346 307414 250358 307466
rect 258346 307414 258358 307466
rect 258410 307463 258422 307466
rect 295978 307463 295990 307466
rect 258410 307417 295990 307463
rect 258410 307414 258422 307417
rect 295978 307414 295990 307417
rect 296042 307414 296054 307466
rect 363850 307414 363862 307466
rect 363914 307463 363926 307466
rect 520874 307463 520886 307466
rect 363914 307417 520886 307463
rect 363914 307414 363926 307417
rect 520874 307414 520886 307417
rect 520938 307414 520950 307466
rect 358362 307302 358374 307354
rect 358426 307351 358438 307354
rect 509898 307351 509910 307354
rect 358426 307305 509910 307351
rect 358426 307302 358438 307305
rect 509898 307302 509910 307305
rect 509962 307302 509974 307354
rect 366090 307190 366102 307242
rect 366154 307239 366166 307242
rect 526810 307239 526822 307242
rect 366154 307193 526822 307239
rect 366154 307190 366166 307193
rect 526810 307190 526822 307193
rect 526874 307190 526886 307242
rect 365642 307078 365654 307130
rect 365706 307127 365718 307130
rect 526586 307127 526598 307130
rect 365706 307081 526598 307127
rect 365706 307078 365718 307081
rect 526586 307078 526598 307081
rect 526650 307078 526662 307130
rect 291274 306966 291286 307018
rect 291338 307015 291350 307018
rect 364634 307015 364646 307018
rect 291338 306969 364646 307015
rect 291338 306966 291350 306969
rect 364634 306966 364646 306969
rect 364698 306966 364710 307018
rect 366874 306966 366886 307018
rect 366938 307015 366950 307018
rect 528266 307015 528278 307018
rect 366938 306969 528278 307015
rect 366938 306966 366950 306969
rect 528266 306966 528278 306969
rect 528330 306966 528342 307018
rect 291834 306854 291846 306906
rect 291898 306903 291910 306906
rect 366202 306903 366214 306906
rect 291898 306857 366214 306903
rect 291898 306854 291910 306857
rect 366202 306854 366214 306857
rect 366266 306854 366278 306906
rect 368106 306854 368118 306906
rect 368170 306903 368182 306906
rect 531626 306903 531638 306906
rect 368170 306857 531638 306903
rect 368170 306854 368182 306857
rect 531626 306854 531638 306857
rect 531690 306854 531702 306906
rect 83738 306742 83750 306794
rect 83802 306791 83814 306794
rect 660986 306791 660998 306794
rect 83802 306745 660998 306791
rect 83802 306742 83814 306745
rect 660986 306742 660998 306745
rect 661050 306742 661062 306794
rect 83626 306630 83638 306682
rect 83690 306679 83702 306682
rect 662666 306679 662678 306682
rect 83690 306633 662678 306679
rect 83690 306630 83702 306633
rect 662666 306630 662678 306633
rect 662730 306630 662742 306682
rect 77242 306518 77254 306570
rect 77306 306567 77318 306570
rect 672298 306567 672310 306570
rect 77306 306521 672310 306567
rect 77306 306518 77318 306521
rect 672298 306518 672310 306521
rect 672362 306518 672374 306570
rect 160010 305846 160022 305898
rect 160074 305895 160086 305898
rect 336858 305895 336870 305898
rect 160074 305849 336870 305895
rect 160074 305846 160086 305849
rect 336858 305846 336870 305849
rect 336922 305846 336934 305898
rect 84746 305734 84758 305786
rect 84810 305783 84822 305786
rect 655946 305783 655958 305786
rect 84810 305737 655958 305783
rect 84810 305734 84822 305737
rect 655946 305734 655958 305737
rect 656010 305734 656022 305786
rect 349178 305622 349190 305674
rect 349242 305671 349254 305674
rect 491306 305671 491318 305674
rect 349242 305625 491318 305671
rect 349242 305622 349254 305625
rect 491306 305622 491318 305625
rect 491370 305622 491382 305674
rect 174794 305510 174806 305562
rect 174858 305559 174870 305562
rect 175354 305559 175366 305562
rect 174858 305513 175366 305559
rect 174858 305510 174870 305513
rect 175354 305510 175366 305513
rect 175418 305510 175430 305562
rect 350970 305510 350982 305562
rect 351034 305559 351046 305562
rect 494666 305559 494678 305562
rect 351034 305513 494678 305559
rect 351034 305510 351046 305513
rect 494666 305510 494678 305513
rect 494730 305510 494742 305562
rect 350410 305398 350422 305450
rect 350474 305447 350486 305450
rect 494890 305447 494902 305450
rect 350474 305401 494902 305447
rect 350474 305398 350486 305401
rect 494890 305398 494902 305401
rect 494954 305398 494966 305450
rect 353434 305286 353446 305338
rect 353498 305335 353510 305338
rect 499706 305335 499718 305338
rect 353498 305289 499718 305335
rect 353498 305286 353510 305289
rect 499706 305286 499718 305289
rect 499770 305286 499782 305338
rect 353994 305174 354006 305226
rect 354058 305223 354070 305226
rect 501386 305223 501398 305226
rect 354058 305177 501398 305223
rect 354058 305174 354070 305177
rect 501386 305174 501398 305177
rect 501450 305174 501462 305226
rect 354666 305062 354678 305114
rect 354730 305111 354742 305114
rect 502282 305111 502294 305114
rect 354730 305065 502294 305111
rect 354730 305062 354742 305065
rect 502282 305062 502294 305065
rect 502346 305062 502358 305114
rect 355898 304950 355910 305002
rect 355962 304999 355974 305002
rect 504746 304999 504758 305002
rect 355962 304953 504758 304999
rect 355962 304950 355974 304953
rect 504746 304950 504758 304953
rect 504810 304950 504822 305002
rect 355226 304838 355238 304890
rect 355290 304887 355302 304890
rect 503962 304887 503974 304890
rect 355290 304841 503974 304887
rect 355290 304838 355302 304841
rect 503962 304838 503974 304841
rect 504026 304838 504038 304890
rect 347386 304726 347398 304778
rect 347450 304775 347462 304778
rect 487946 304775 487958 304778
rect 347450 304729 487958 304775
rect 347450 304726 347462 304729
rect 487946 304726 487958 304729
rect 488010 304726 488022 304778
rect 339994 304614 340006 304666
rect 340058 304663 340070 304666
rect 472042 304663 472054 304666
rect 340058 304617 472054 304663
rect 340058 304614 340070 304617
rect 472042 304614 472054 304617
rect 472106 304614 472118 304666
rect 340666 303942 340678 303994
rect 340730 303991 340742 303994
rect 472826 303991 472838 303994
rect 340730 303945 472838 303991
rect 340730 303942 340742 303945
rect 472826 303942 472838 303945
rect 472890 303942 472902 303994
rect 341898 303830 341910 303882
rect 341962 303879 341974 303882
rect 475402 303879 475414 303882
rect 341962 303833 475414 303879
rect 341962 303830 341974 303833
rect 475402 303830 475414 303833
rect 475466 303830 475478 303882
rect 343018 303718 343030 303770
rect 343082 303767 343094 303770
rect 477866 303767 477878 303770
rect 343082 303721 477878 303767
rect 343082 303718 343094 303721
rect 477866 303718 477878 303721
rect 477930 303718 477942 303770
rect 346154 303606 346166 303658
rect 346218 303655 346230 303658
rect 483802 303655 483814 303658
rect 346218 303609 483814 303655
rect 346218 303606 346230 303609
rect 483802 303606 483814 303609
rect 483866 303606 483878 303658
rect 361386 303494 361398 303546
rect 361450 303543 361462 303546
rect 516506 303543 516518 303546
rect 361450 303497 516518 303543
rect 361450 303494 361462 303497
rect 516506 303494 516518 303497
rect 516570 303494 516582 303546
rect 360154 303382 360166 303434
rect 360218 303431 360230 303434
rect 514826 303431 514838 303434
rect 360218 303385 514838 303431
rect 360218 303382 360230 303385
rect 514826 303382 514838 303385
rect 514890 303382 514902 303434
rect 361946 303270 361958 303322
rect 362010 303319 362022 303322
rect 518186 303319 518198 303322
rect 362010 303273 518198 303319
rect 362010 303270 362022 303273
rect 518186 303270 518198 303273
rect 518250 303270 518262 303322
rect 168746 303158 168758 303210
rect 168810 303207 168822 303210
rect 184426 303207 184438 303210
rect 168810 303161 184438 303207
rect 168810 303158 168822 303161
rect 184426 303158 184438 303161
rect 184490 303158 184502 303210
rect 360714 303158 360726 303210
rect 360778 303207 360790 303210
rect 516730 303207 516742 303210
rect 360778 303161 516742 303207
rect 360778 303158 360790 303161
rect 516730 303158 516742 303161
rect 516794 303158 516806 303210
rect 298218 302262 298230 302314
rect 298282 302311 298294 302314
rect 335850 302311 335862 302314
rect 298282 302265 335862 302311
rect 298282 302262 298294 302265
rect 335850 302262 335862 302265
rect 335914 302262 335926 302314
rect 297434 301702 297446 301754
rect 297498 301751 297510 301754
rect 335066 301751 335078 301754
rect 297498 301705 335078 301751
rect 297498 301702 297510 301705
rect 335066 301702 335078 301705
rect 335130 301702 335142 301754
rect 659306 301702 659318 301754
rect 659370 301751 659382 301754
rect 670730 301751 670742 301754
rect 659370 301705 670742 301751
rect 659370 301702 659382 301705
rect 670730 301702 670742 301705
rect 670794 301702 670806 301754
rect 295866 301590 295878 301642
rect 295930 301639 295942 301642
rect 335290 301639 335302 301642
rect 295930 301593 335302 301639
rect 295930 301590 295942 301593
rect 335290 301590 335302 301593
rect 335354 301590 335366 301642
rect 660986 301590 660998 301642
rect 661050 301639 661062 301642
rect 670954 301639 670966 301642
rect 661050 301593 670966 301639
rect 661050 301590 661062 301593
rect 670954 301590 670966 301593
rect 671018 301590 671030 301642
rect 287466 301478 287478 301530
rect 287530 301527 287542 301530
rect 357802 301527 357814 301530
rect 287530 301481 357814 301527
rect 287530 301478 287542 301481
rect 357802 301478 357814 301481
rect 357866 301478 357878 301530
rect 655946 301478 655958 301530
rect 656010 301527 656022 301530
rect 670282 301527 670294 301530
rect 656010 301481 670294 301527
rect 656010 301478 656022 301481
rect 670282 301478 670294 301481
rect 670346 301478 670358 301530
rect 299450 300470 299462 300522
rect 299514 300519 299526 300522
rect 383002 300519 383014 300522
rect 299514 300473 383014 300519
rect 299514 300470 299526 300473
rect 383002 300470 383014 300473
rect 383066 300470 383078 300522
rect 301018 300358 301030 300410
rect 301082 300407 301094 300410
rect 386362 300407 386374 300410
rect 301082 300361 386374 300407
rect 301082 300358 301094 300361
rect 386362 300358 386374 300361
rect 386426 300358 386438 300410
rect 299226 300246 299238 300298
rect 299290 300295 299302 300298
rect 384682 300295 384694 300298
rect 299290 300249 384694 300295
rect 299290 300246 299302 300249
rect 384682 300246 384694 300249
rect 384746 300246 384758 300298
rect 300794 300134 300806 300186
rect 300858 300183 300870 300186
rect 386922 300183 386934 300186
rect 300858 300137 386934 300183
rect 300858 300134 300870 300137
rect 386922 300134 386934 300137
rect 386986 300134 386998 300186
rect 304154 300022 304166 300074
rect 304218 300071 304230 300074
rect 394762 300071 394774 300074
rect 304218 300025 394774 300071
rect 304218 300022 304230 300025
rect 394762 300022 394774 300025
rect 394826 300022 394838 300074
rect 310874 299910 310886 299962
rect 310938 299959 310950 299962
rect 408650 299959 408662 299962
rect 310938 299913 408662 299959
rect 310938 299910 310950 299913
rect 408650 299910 408662 299913
rect 408714 299910 408726 299962
rect 83290 299798 83302 299850
rect 83354 299847 83366 299850
rect 654490 299847 654502 299850
rect 83354 299801 654502 299847
rect 83354 299798 83366 299801
rect 654490 299798 654502 299801
rect 654554 299798 654566 299850
rect 337530 293974 337542 294026
rect 337594 294023 337606 294026
rect 670394 294023 670406 294026
rect 337594 293977 670406 294023
rect 337594 293974 337606 293977
rect 670394 293974 670406 293977
rect 670458 293974 670470 294026
rect 467002 293862 467014 293914
rect 467066 293911 467078 293914
rect 467786 293911 467798 293914
rect 467066 293865 467798 293911
rect 467066 293862 467078 293865
rect 467786 293862 467798 293865
rect 467850 293862 467862 293914
rect 487162 293862 487174 293914
rect 487226 293911 487238 293914
rect 487946 293911 487958 293914
rect 487226 293865 487958 293911
rect 487226 293862 487238 293865
rect 487946 293862 487958 293865
rect 488010 293862 488022 293914
rect 495786 293862 495798 293914
rect 495850 293911 495862 293914
rect 496346 293911 496358 293914
rect 495850 293865 496358 293911
rect 495850 293862 495862 293865
rect 496346 293862 496358 293865
rect 496410 293862 496422 293914
rect 515722 293862 515734 293914
rect 515786 293911 515798 293914
rect 516730 293911 516742 293914
rect 515786 293865 516742 293911
rect 515786 293862 515798 293865
rect 516730 293862 516742 293865
rect 516794 293862 516806 293914
rect 517514 293862 517526 293914
rect 517578 293911 517590 293914
rect 518186 293911 518198 293914
rect 517578 293865 518198 293911
rect 517578 293862 517590 293865
rect 518186 293862 518198 293865
rect 518250 293862 518262 293914
rect 519082 293526 519094 293578
rect 519146 293575 519158 293578
rect 520538 293575 520550 293578
rect 519146 293529 520550 293575
rect 519146 293526 519158 293529
rect 520538 293526 520550 293529
rect 520602 293526 520614 293578
rect 492202 293414 492214 293466
rect 492266 293463 492278 293466
rect 492986 293463 492998 293466
rect 492266 293417 492998 293463
rect 492266 293414 492278 293417
rect 492986 293414 492998 293417
rect 493050 293414 493062 293466
rect 493994 293414 494006 293466
rect 494058 293463 494070 293466
rect 494890 293463 494902 293466
rect 494058 293417 494902 293463
rect 494058 293414 494070 293417
rect 494890 293414 494902 293417
rect 494954 293414 494966 293466
rect 566010 293414 566022 293466
rect 566074 293463 566086 293466
rect 645418 293463 645430 293466
rect 566074 293417 645430 293463
rect 566074 293414 566086 293417
rect 645418 293414 645430 293417
rect 645482 293414 645494 293466
rect 520762 293302 520774 293354
rect 520826 293351 520838 293354
rect 522330 293351 522342 293354
rect 520826 293305 522342 293351
rect 520826 293302 520838 293305
rect 522330 293302 522342 293305
rect 522394 293351 522406 293354
rect 631418 293351 631430 293354
rect 522394 293305 631430 293351
rect 522394 293302 522406 293305
rect 631418 293302 631430 293305
rect 631482 293302 631494 293354
rect 520538 293190 520550 293242
rect 520602 293239 520614 293242
rect 630970 293239 630982 293242
rect 520602 293193 630982 293239
rect 520602 293190 520614 293193
rect 630970 293190 630982 293193
rect 631034 293190 631046 293242
rect 494890 293078 494902 293130
rect 494954 293127 494966 293130
rect 606218 293127 606230 293130
rect 494954 293081 606230 293127
rect 494954 293078 494966 293081
rect 606218 293078 606230 293081
rect 606282 293078 606294 293130
rect 516730 292966 516742 293018
rect 516794 293015 516806 293018
rect 629514 293015 629526 293018
rect 516794 292969 629526 293015
rect 516794 292966 516806 292969
rect 629514 292966 629526 292969
rect 629578 292966 629590 293018
rect 517514 292854 517526 292906
rect 517578 292903 517590 292906
rect 630522 292903 630534 292906
rect 517578 292857 630534 292903
rect 517578 292854 517590 292857
rect 630522 292854 630534 292857
rect 630586 292854 630598 292906
rect 492986 292742 492998 292794
rect 493050 292791 493062 292794
rect 613498 292791 613510 292794
rect 493050 292745 613510 292791
rect 493050 292742 493062 292745
rect 613498 292742 613510 292745
rect 613562 292742 613574 292794
rect 487162 292630 487174 292682
rect 487226 292679 487238 292682
rect 606330 292679 606342 292682
rect 487226 292633 606342 292679
rect 487226 292630 487238 292633
rect 606330 292630 606342 292633
rect 606394 292630 606406 292682
rect 495786 292518 495798 292570
rect 495850 292567 495862 292570
rect 495850 292521 508391 292567
rect 495850 292518 495862 292521
rect 500826 292406 500838 292458
rect 500890 292455 500902 292458
rect 501386 292455 501398 292458
rect 500890 292409 501398 292455
rect 500890 292406 500902 292409
rect 501386 292406 501398 292409
rect 501450 292455 501462 292458
rect 508218 292455 508230 292458
rect 501450 292409 508230 292455
rect 501450 292406 501462 292409
rect 508218 292406 508230 292409
rect 508282 292406 508294 292458
rect 508345 292455 508391 292521
rect 508554 292518 508566 292570
rect 508618 292567 508630 292570
rect 624250 292567 624262 292570
rect 508618 292521 624262 292567
rect 508618 292518 508630 292521
rect 624250 292518 624262 292521
rect 624314 292518 624326 292570
rect 622346 292455 622358 292458
rect 508345 292409 622358 292455
rect 622346 292406 622358 292409
rect 622410 292406 622422 292458
rect 467002 292294 467014 292346
rect 467066 292343 467078 292346
rect 643962 292343 643974 292346
rect 467066 292297 643974 292343
rect 467066 292294 467078 292297
rect 643962 292294 643974 292297
rect 644026 292294 644038 292346
rect 92474 292182 92486 292234
rect 92538 292231 92550 292234
rect 609802 292231 609814 292234
rect 92538 292185 609814 292231
rect 92538 292182 92550 292185
rect 609802 292182 609814 292185
rect 609866 292182 609878 292234
rect 529162 292070 529174 292122
rect 529226 292119 529238 292122
rect 529946 292119 529958 292122
rect 529226 292073 529958 292119
rect 529226 292070 529238 292073
rect 529946 292070 529958 292073
rect 530010 292070 530022 292122
rect 531066 292070 531078 292122
rect 531130 292119 531142 292122
rect 531626 292119 531638 292122
rect 531130 292073 531638 292119
rect 531130 292070 531142 292073
rect 531626 292070 531638 292073
rect 531690 292070 531702 292122
rect 530842 291958 530854 292010
rect 530906 292007 530918 292010
rect 532410 292007 532422 292010
rect 530906 291961 532422 292007
rect 530906 291958 530918 291961
rect 532410 291958 532422 291961
rect 532474 291958 532486 292010
rect 610810 291958 610822 292010
rect 610874 292007 610886 292010
rect 617978 292007 617990 292010
rect 610874 291961 617990 292007
rect 610874 291958 610886 291961
rect 617978 291958 617990 291961
rect 618042 291958 618054 292010
rect 612378 291846 612390 291898
rect 612442 291895 612454 291898
rect 615738 291895 615750 291898
rect 612442 291849 615750 291895
rect 612442 291846 612454 291849
rect 615738 291846 615750 291849
rect 615802 291846 615814 291898
rect 322522 291734 322534 291786
rect 322586 291783 322598 291786
rect 433402 291783 433414 291786
rect 322586 291737 433414 291783
rect 322586 291734 322598 291737
rect 433402 291734 433414 291737
rect 433466 291734 433478 291786
rect 609914 291734 609926 291786
rect 609978 291783 609990 291786
rect 620666 291783 620678 291786
rect 609978 291737 620678 291783
rect 609978 291734 609990 291737
rect 620666 291734 620678 291737
rect 620730 291734 620742 291786
rect 324090 291622 324102 291674
rect 324154 291671 324166 291674
rect 435194 291671 435206 291674
rect 324154 291625 435206 291671
rect 324154 291622 324166 291625
rect 435194 291622 435206 291625
rect 435258 291622 435270 291674
rect 504746 291622 504758 291674
rect 504810 291671 504822 291674
rect 625706 291671 625718 291674
rect 504810 291625 625718 291671
rect 504810 291622 504822 291625
rect 625706 291622 625718 291625
rect 625770 291622 625782 291674
rect 334506 291510 334518 291562
rect 334570 291559 334582 291562
rect 456026 291559 456038 291562
rect 334570 291513 456038 291559
rect 334570 291510 334582 291513
rect 456026 291510 456038 291513
rect 456090 291510 456102 291562
rect 531066 291510 531078 291562
rect 531130 291559 531142 291562
rect 635338 291559 635350 291562
rect 531130 291513 635350 291559
rect 531130 291510 531142 291513
rect 635338 291510 635350 291513
rect 635402 291510 635414 291562
rect 334618 291398 334630 291450
rect 334682 291447 334694 291450
rect 457370 291447 457382 291450
rect 334682 291401 457382 291447
rect 334682 291398 334694 291401
rect 457370 291398 457382 291401
rect 457434 291398 457446 291450
rect 532410 291398 532422 291450
rect 532474 291447 532486 291450
rect 635786 291447 635798 291450
rect 532474 291401 635798 291447
rect 532474 291398 532486 291401
rect 635786 291398 635798 291401
rect 635850 291398 635862 291450
rect 529162 291286 529174 291338
rect 529226 291335 529238 291338
rect 634778 291335 634790 291338
rect 529226 291289 634790 291335
rect 529226 291286 529238 291289
rect 634778 291286 634790 291289
rect 634842 291286 634854 291338
rect 528266 291174 528278 291226
rect 528330 291223 528342 291226
rect 634330 291223 634342 291226
rect 528330 291177 634342 291223
rect 528330 291174 528342 291177
rect 634330 291174 634342 291177
rect 634394 291174 634406 291226
rect 525802 291062 525814 291114
rect 525866 291111 525878 291114
rect 526810 291111 526822 291114
rect 525866 291065 526822 291111
rect 525866 291062 525878 291065
rect 526810 291062 526822 291065
rect 526874 291111 526886 291114
rect 633882 291111 633894 291114
rect 526874 291065 633894 291111
rect 526874 291062 526886 291065
rect 633882 291062 633894 291065
rect 633946 291062 633958 291114
rect 516506 290950 516518 291002
rect 516570 290999 516582 291002
rect 629962 290999 629974 291002
rect 516570 290953 629974 290999
rect 516570 290950 516582 290953
rect 629962 290950 629974 290953
rect 630026 290950 630038 291002
rect 509898 290838 509910 290890
rect 509962 290887 509974 290890
rect 627610 290887 627622 290890
rect 509962 290841 627622 290887
rect 509962 290838 509974 290841
rect 627610 290838 627622 290841
rect 627674 290838 627686 290890
rect 610698 290726 610710 290778
rect 610762 290775 610774 290778
rect 612714 290775 612726 290778
rect 610762 290729 612726 290775
rect 610762 290726 610774 290729
rect 612714 290726 612726 290729
rect 612778 290726 612790 290778
rect 620666 290726 620678 290778
rect 620730 290775 620742 290778
rect 669834 290775 669846 290778
rect 620730 290729 669846 290775
rect 620730 290726 620742 290729
rect 669834 290726 669846 290729
rect 669898 290726 669910 290778
rect 92586 290614 92598 290666
rect 92650 290663 92662 290666
rect 612378 290663 612390 290666
rect 92650 290617 612390 290663
rect 92650 290614 92662 290617
rect 612378 290614 612390 290617
rect 612442 290614 612454 290666
rect 615738 290614 615750 290666
rect 615802 290663 615814 290666
rect 671290 290663 671302 290666
rect 615802 290617 671302 290663
rect 615802 290614 615814 290617
rect 671290 290614 671302 290617
rect 671354 290614 671366 290666
rect 606330 290502 606342 290554
rect 606394 290551 606406 290554
rect 612490 290551 612502 290554
rect 606394 290505 612502 290551
rect 606394 290502 606406 290505
rect 612490 290502 612502 290505
rect 612554 290502 612566 290554
rect 612826 290502 612838 290554
rect 612890 290551 612902 290554
rect 618986 290551 618998 290554
rect 612890 290505 618998 290551
rect 612890 290502 612902 290505
rect 618986 290502 618998 290505
rect 619050 290502 619062 290554
rect 651130 290502 651142 290554
rect 651194 290551 651206 290554
rect 689322 290551 689334 290554
rect 651194 290505 689334 290551
rect 651194 290502 651206 290505
rect 689322 290502 689334 290505
rect 689386 290502 689398 290554
rect 605770 290390 605782 290442
rect 605834 290439 605846 290442
rect 619434 290439 619446 290442
rect 605834 290393 619446 290439
rect 605834 290390 605846 290393
rect 619434 290390 619446 290393
rect 619498 290390 619510 290442
rect 650234 290390 650246 290442
rect 650298 290439 650310 290442
rect 688202 290439 688214 290442
rect 650298 290393 688214 290439
rect 650298 290390 650310 290393
rect 688202 290390 688214 290393
rect 688266 290390 688278 290442
rect 606106 290278 606118 290330
rect 606170 290327 606182 290330
rect 610810 290327 610822 290330
rect 606170 290281 610822 290327
rect 606170 290278 606182 290281
rect 610810 290278 610822 290281
rect 610874 290278 610886 290330
rect 611034 290278 611046 290330
rect 611098 290327 611110 290330
rect 614730 290327 614742 290330
rect 611098 290281 614742 290327
rect 611098 290278 611110 290281
rect 614730 290278 614742 290281
rect 614794 290278 614806 290330
rect 655946 290278 655958 290330
rect 656010 290327 656022 290330
rect 656010 290281 668663 290327
rect 656010 290278 656022 290281
rect 606330 290166 606342 290218
rect 606394 290215 606406 290218
rect 613162 290215 613174 290218
rect 606394 290169 613174 290215
rect 606394 290166 606406 290169
rect 613162 290166 613174 290169
rect 613226 290166 613238 290218
rect 615178 290166 615190 290218
rect 615242 290215 615254 290218
rect 615626 290215 615638 290218
rect 615242 290169 615638 290215
rect 615242 290166 615254 290169
rect 615626 290166 615638 290169
rect 615690 290166 615702 290218
rect 654042 290166 654054 290218
rect 654106 290215 654118 290218
rect 668154 290215 668166 290218
rect 654106 290169 668166 290215
rect 654106 290166 654118 290169
rect 668154 290166 668166 290169
rect 668218 290166 668230 290218
rect 668617 290215 668663 290281
rect 670058 290278 670070 290330
rect 670122 290327 670134 290330
rect 670730 290327 670742 290330
rect 670122 290281 670742 290327
rect 670122 290278 670134 290281
rect 670730 290278 670742 290281
rect 670794 290278 670806 290330
rect 670282 290215 670294 290218
rect 668617 290169 670294 290215
rect 670282 290166 670294 290169
rect 670346 290166 670358 290218
rect 610810 290054 610822 290106
rect 610874 290103 610886 290106
rect 613722 290103 613734 290106
rect 610874 290057 613734 290103
rect 610874 290054 610886 290057
rect 613722 290054 613734 290057
rect 613786 290054 613798 290106
rect 649674 290054 649686 290106
rect 649738 290103 649750 290106
rect 688874 290103 688886 290106
rect 649738 290057 688886 290103
rect 649738 290054 649750 290057
rect 688874 290054 688886 290057
rect 688938 290054 688950 290106
rect 80378 289942 80390 289994
rect 80442 289991 80454 289994
rect 659754 289991 659766 289994
rect 80442 289945 659766 289991
rect 80442 289942 80454 289945
rect 659754 289942 659766 289945
rect 659818 289942 659830 289994
rect 660314 289942 660326 289994
rect 660378 289991 660390 289994
rect 670954 289991 670966 289994
rect 660378 289945 670966 289991
rect 660378 289942 660390 289945
rect 670954 289942 670966 289945
rect 671018 289942 671030 289994
rect 78698 289830 78710 289882
rect 78762 289879 78774 289882
rect 661210 289879 661222 289882
rect 78762 289833 661222 289879
rect 78762 289830 78774 289833
rect 661210 289830 661222 289833
rect 661274 289830 661286 289882
rect 664570 289830 664582 289882
rect 664634 289879 664646 289882
rect 670618 289879 670630 289882
rect 664634 289833 670630 289879
rect 664634 289830 664646 289833
rect 670618 289830 670630 289833
rect 670682 289830 670694 289882
rect 80154 289718 80166 289770
rect 80218 289767 80230 289770
rect 665578 289767 665590 289770
rect 80218 289721 665590 289767
rect 80218 289718 80230 289721
rect 665578 289718 665590 289721
rect 665642 289718 665654 289770
rect 667930 289767 667942 289770
rect 666936 289721 667942 289767
rect 78698 289606 78710 289658
rect 78762 289655 78774 289658
rect 666936 289655 666982 289721
rect 667930 289718 667942 289721
rect 667994 289718 668006 289770
rect 668938 289718 668950 289770
rect 669002 289767 669014 289770
rect 670282 289767 670294 289770
rect 669002 289721 670294 289767
rect 669002 289718 669014 289721
rect 670282 289718 670294 289721
rect 670346 289718 670358 289770
rect 671850 289718 671862 289770
rect 671914 289767 671926 289770
rect 687418 289767 687430 289770
rect 671914 289721 687430 289767
rect 671914 289718 671926 289721
rect 687418 289718 687430 289721
rect 687482 289718 687494 289770
rect 78762 289609 666982 289655
rect 78762 289606 78774 289609
rect 668154 289606 668166 289658
rect 668218 289655 668230 289658
rect 672186 289655 672198 289658
rect 668218 289609 672198 289655
rect 668218 289606 668230 289609
rect 672186 289606 672198 289609
rect 672250 289606 672262 289658
rect 606330 288822 606342 288874
rect 606394 288871 606406 288874
rect 611370 288871 611382 288874
rect 606394 288825 611382 288871
rect 606394 288822 606406 288825
rect 611370 288822 611382 288825
rect 611434 288822 611446 288874
rect 606218 288710 606230 288762
rect 606282 288759 606294 288762
rect 610810 288759 610822 288762
rect 606282 288713 610822 288759
rect 606282 288710 606294 288713
rect 610810 288710 610822 288713
rect 610874 288710 610886 288762
rect 105802 285574 105814 285626
rect 105866 285623 105878 285626
rect 106474 285623 106486 285626
rect 105866 285577 106486 285623
rect 105866 285574 105878 285577
rect 106474 285574 106486 285577
rect 106538 285574 106550 285626
rect 196858 285574 196870 285626
rect 196922 285623 196934 285626
rect 197418 285623 197430 285626
rect 196922 285577 197430 285623
rect 196922 285574 196934 285577
rect 197418 285574 197430 285577
rect 197482 285574 197494 285626
rect 278842 285574 278854 285626
rect 278906 285623 278918 285626
rect 279402 285623 279414 285626
rect 278906 285577 279414 285623
rect 278906 285574 278918 285577
rect 279402 285574 279414 285577
rect 279466 285574 279478 285626
rect 525802 285574 525814 285626
rect 525866 285623 525878 285626
rect 526586 285623 526598 285626
rect 525866 285577 526598 285623
rect 525866 285574 525878 285577
rect 526586 285574 526598 285577
rect 526650 285574 526662 285626
rect 542602 285574 542614 285626
rect 542666 285623 542678 285626
rect 543274 285623 543286 285626
rect 542666 285577 543286 285623
rect 542666 285574 542678 285577
rect 543274 285574 543286 285577
rect 543338 285574 543350 285626
rect 331034 285014 331046 285066
rect 331098 285063 331110 285066
rect 451658 285063 451670 285066
rect 331098 285017 451670 285063
rect 331098 285014 331110 285017
rect 451658 285014 451670 285017
rect 451722 285014 451734 285066
rect 329354 284902 329366 284954
rect 329418 284951 329430 284954
rect 449194 284951 449206 284954
rect 329418 284905 449206 284951
rect 329418 284902 329430 284905
rect 449194 284902 449206 284905
rect 449258 284902 449270 284954
rect 332826 284790 332838 284842
rect 332890 284839 332902 284842
rect 454234 284839 454246 284842
rect 332890 284793 454246 284839
rect 332890 284790 332902 284793
rect 454234 284790 454246 284793
rect 454298 284790 454310 284842
rect 332938 284678 332950 284730
rect 333002 284727 333014 284730
rect 455578 284727 455590 284730
rect 333002 284681 455590 284727
rect 333002 284678 333014 284681
rect 455578 284678 455590 284681
rect 455642 284678 455654 284730
rect 530842 282774 530854 282826
rect 530906 282823 530918 282826
rect 531738 282823 531750 282826
rect 530906 282777 531750 282823
rect 530906 282774 530918 282777
rect 531738 282774 531750 282777
rect 531802 282774 531814 282826
rect 331370 282102 331382 282154
rect 331434 282151 331446 282154
rect 332154 282151 332166 282154
rect 331434 282105 332166 282151
rect 331434 282102 331446 282105
rect 332154 282102 332166 282105
rect 332218 282102 332230 282154
rect 345146 281878 345158 281930
rect 345210 281927 345222 281930
rect 352426 281927 352438 281930
rect 345210 281881 352438 281927
rect 345210 281878 345222 281881
rect 352426 281878 352438 281881
rect 352490 281878 352502 281930
rect 335290 281766 335302 281818
rect 335354 281815 335366 281818
rect 378746 281815 378758 281818
rect 335354 281769 378758 281815
rect 335354 281766 335366 281769
rect 378746 281766 378758 281769
rect 378810 281766 378822 281818
rect 301690 281654 301702 281706
rect 301754 281703 301766 281706
rect 345370 281703 345382 281706
rect 301754 281657 345382 281703
rect 301754 281654 301766 281657
rect 345370 281654 345382 281657
rect 345434 281654 345446 281706
rect 335066 281542 335078 281594
rect 335130 281591 335142 281594
rect 379978 281591 379990 281594
rect 335130 281545 379990 281591
rect 335130 281542 335142 281545
rect 379978 281542 379990 281545
rect 380042 281542 380054 281594
rect 165610 281430 165622 281482
rect 165674 281479 165686 281482
rect 173114 281479 173126 281482
rect 165674 281433 173126 281479
rect 165674 281430 165686 281433
rect 173114 281430 173126 281433
rect 173178 281430 173190 281482
rect 173898 281430 173910 281482
rect 173962 281479 173974 281482
rect 179834 281479 179846 281482
rect 173962 281433 179846 281479
rect 173962 281430 173974 281433
rect 179834 281430 179846 281433
rect 179898 281430 179910 281482
rect 265738 281430 265750 281482
rect 265802 281479 265814 281482
rect 313338 281479 313350 281482
rect 265802 281433 313350 281479
rect 265802 281430 265814 281433
rect 313338 281430 313350 281433
rect 313402 281430 313414 281482
rect 334618 281430 334630 281482
rect 334682 281479 334694 281482
rect 396666 281479 396678 281482
rect 334682 281433 396678 281479
rect 334682 281430 334694 281433
rect 396666 281430 396678 281433
rect 396730 281430 396742 281482
rect 166058 281318 166070 281370
rect 166122 281367 166134 281370
rect 195066 281367 195078 281370
rect 166122 281321 178103 281367
rect 166122 281318 166134 281321
rect 131450 281206 131462 281258
rect 131514 281255 131526 281258
rect 177930 281255 177942 281258
rect 131514 281209 177942 281255
rect 131514 281206 131526 281209
rect 177930 281206 177942 281209
rect 177994 281206 178006 281258
rect 178057 281255 178103 281321
rect 179736 281321 195078 281367
rect 179736 281255 179782 281321
rect 195066 281318 195078 281321
rect 195130 281318 195142 281370
rect 265514 281318 265526 281370
rect 265578 281367 265590 281370
rect 314682 281367 314694 281370
rect 265578 281321 314694 281367
rect 265578 281318 265590 281321
rect 314682 281318 314694 281321
rect 314746 281318 314758 281370
rect 334394 281318 334406 281370
rect 334458 281367 334470 281370
rect 408202 281367 408214 281370
rect 334458 281321 408214 281367
rect 334458 281318 334470 281321
rect 408202 281318 408214 281321
rect 408266 281318 408278 281370
rect 255546 281255 255558 281258
rect 178057 281209 179782 281255
rect 255337 281209 255558 281255
rect 132794 281094 132806 281146
rect 132858 281143 132870 281146
rect 173898 281143 173910 281146
rect 132858 281097 173910 281143
rect 132858 281094 132870 281097
rect 173898 281094 173910 281097
rect 173962 281094 173974 281146
rect 196634 281143 196646 281146
rect 196536 281097 196646 281143
rect 128314 280982 128326 281034
rect 128378 281031 128390 281034
rect 176474 281031 176486 281034
rect 128378 280985 176486 281031
rect 128378 280982 128390 280985
rect 176474 280982 176486 280985
rect 176538 280982 176550 281034
rect 130890 280870 130902 280922
rect 130954 280919 130966 280922
rect 178266 280919 178278 280922
rect 130954 280873 178278 280919
rect 130954 280870 130966 280873
rect 178266 280870 178278 280873
rect 178330 280870 178342 280922
rect 124170 280758 124182 280810
rect 124234 280807 124246 280810
rect 174682 280807 174694 280810
rect 124234 280761 174694 280807
rect 124234 280758 124246 280761
rect 174682 280758 174694 280761
rect 174746 280758 174758 280810
rect 196536 280807 196582 281097
rect 196634 281094 196646 281097
rect 196698 281094 196710 281146
rect 200106 281094 200118 281146
rect 200170 281094 200182 281146
rect 176601 280761 196582 280807
rect 110394 280646 110406 280698
rect 110458 280646 110470 280698
rect 120586 280646 120598 280698
rect 120650 280695 120662 280698
rect 165610 280695 165622 280698
rect 120650 280649 165622 280695
rect 120650 280646 120662 280649
rect 165610 280646 165622 280649
rect 165674 280646 165686 280698
rect 167850 280646 167862 280698
rect 167914 280646 167926 280698
rect 169194 280646 169206 280698
rect 169258 280646 169270 280698
rect 110409 280583 110455 280646
rect 167865 280583 167911 280646
rect 110409 280537 167911 280583
rect 169209 280583 169255 280646
rect 176601 280583 176647 280761
rect 180730 280646 180742 280698
rect 180794 280695 180806 280698
rect 200121 280695 200167 281094
rect 255337 280919 255383 281209
rect 255546 281206 255558 281209
rect 255610 281206 255622 281258
rect 268874 281206 268886 281258
rect 268938 281255 268950 281258
rect 319834 281255 319846 281258
rect 268938 281209 319846 281255
rect 268938 281206 268950 281209
rect 319834 281206 319846 281209
rect 319898 281206 319910 281258
rect 320058 281206 320070 281258
rect 320122 281255 320134 281258
rect 397898 281255 397910 281258
rect 320122 281209 397910 281255
rect 320122 281206 320134 281209
rect 397898 281206 397910 281209
rect 397962 281206 397974 281258
rect 255434 281094 255446 281146
rect 255498 281094 255510 281146
rect 268986 281094 268998 281146
rect 269050 281143 269062 281146
rect 321066 281143 321078 281146
rect 269050 281097 321078 281143
rect 269050 281094 269062 281097
rect 321066 281094 321078 281097
rect 321130 281094 321142 281146
rect 331930 281094 331942 281146
rect 331994 281143 332006 281146
rect 335178 281143 335190 281146
rect 331994 281097 335190 281143
rect 331994 281094 332006 281097
rect 335178 281094 335190 281097
rect 335242 281094 335254 281146
rect 335514 281094 335526 281146
rect 335578 281143 335590 281146
rect 417162 281143 417174 281146
rect 335578 281097 417174 281143
rect 335578 281094 335590 281097
rect 417162 281094 417174 281097
rect 417226 281094 417238 281146
rect 255449 281031 255495 281094
rect 291162 281031 291174 281034
rect 255449 280985 291174 281031
rect 291162 280982 291174 280985
rect 291226 280982 291238 281034
rect 307514 280982 307526 281034
rect 307578 281031 307590 281034
rect 401482 281031 401494 281034
rect 307578 280985 401494 281031
rect 307578 280982 307590 280985
rect 401482 280982 401494 280985
rect 401546 280982 401558 281034
rect 292282 280919 292294 280922
rect 255337 280873 292294 280919
rect 292282 280870 292294 280873
rect 292346 280870 292358 280922
rect 312666 280870 312678 280922
rect 312730 280919 312742 280922
rect 413018 280919 413030 280922
rect 312730 280873 413030 280919
rect 312730 280870 312742 280873
rect 413018 280870 413030 280873
rect 413082 280870 413094 280922
rect 273018 280758 273030 280810
rect 273082 280807 273094 280810
rect 273082 280761 278902 280807
rect 273082 280758 273094 280761
rect 180794 280649 186502 280695
rect 180794 280646 180806 280649
rect 169209 280537 176647 280583
rect 186456 280583 186502 280649
rect 188136 280649 200167 280695
rect 188136 280583 188182 280649
rect 275594 280646 275606 280698
rect 275658 280646 275670 280698
rect 278856 280695 278902 280761
rect 289706 280758 289718 280810
rect 289770 280807 289782 280810
rect 347722 280807 347734 280810
rect 289770 280761 347734 280807
rect 289770 280758 289782 280761
rect 347722 280758 347734 280761
rect 347786 280758 347798 280810
rect 349416 280761 358647 280807
rect 325882 280695 325894 280698
rect 278856 280649 325894 280695
rect 325882 280646 325894 280649
rect 325946 280646 325958 280698
rect 331930 280646 331942 280698
rect 331994 280646 332006 280698
rect 332154 280646 332166 280698
rect 332218 280695 332230 280698
rect 349416 280695 349462 280761
rect 332218 280649 349462 280695
rect 332218 280646 332230 280649
rect 352426 280646 352438 280698
rect 352490 280646 352502 280698
rect 358474 280695 358486 280698
rect 352776 280649 358486 280695
rect 186456 280537 188182 280583
rect 275609 280583 275655 280646
rect 331945 280583 331991 280646
rect 275609 280537 331991 280583
rect 352441 280583 352487 280646
rect 352776 280583 352822 280649
rect 358474 280646 358486 280649
rect 358538 280646 358550 280698
rect 352441 280537 352822 280583
rect 358601 280583 358647 280761
rect 362730 280758 362742 280810
rect 362794 280807 362806 280810
rect 375498 280807 375510 280810
rect 362794 280761 375510 280807
rect 362794 280758 362806 280761
rect 375498 280758 375510 280761
rect 375562 280758 375574 280810
rect 375625 280761 378023 280807
rect 375625 280583 375671 280761
rect 377850 280646 377862 280698
rect 377914 280646 377926 280698
rect 377977 280695 378023 280761
rect 378074 280758 378086 280810
rect 378138 280807 378150 280810
rect 552682 280807 552694 280810
rect 378138 280761 552694 280807
rect 378138 280758 378150 280761
rect 552682 280758 552694 280761
rect 552746 280758 552758 280810
rect 450202 280695 450214 280698
rect 377977 280649 450214 280695
rect 450202 280646 450214 280649
rect 450266 280646 450278 280698
rect 553578 280646 553590 280698
rect 553642 280646 553654 280698
rect 358601 280537 375671 280583
rect 377865 280583 377911 280646
rect 553593 280583 553639 280646
rect 377865 280537 553639 280583
rect 693242 236742 693254 236794
rect 693306 236791 693318 236794
rect 700522 236791 700534 236794
rect 693306 236745 700534 236791
rect 693306 236742 693318 236745
rect 700522 236742 700534 236745
rect 700586 236742 700598 236794
rect 73434 208070 73446 208122
rect 73498 208119 73510 208122
rect 78250 208119 78262 208122
rect 73498 208073 78262 208119
rect 73498 208070 73510 208073
rect 78250 208070 78262 208073
rect 78314 208070 78326 208122
rect 560186 139862 560198 139914
rect 560250 139911 560262 139914
rect 647882 139911 647894 139914
rect 560250 139865 647894 139911
rect 560250 139862 560262 139865
rect 647882 139862 647894 139865
rect 647946 139862 647958 139914
rect 619770 139750 619782 139802
rect 619834 139799 619846 139802
rect 619834 139753 619942 139799
rect 619834 139750 619846 139753
rect 619896 139687 619942 139753
rect 621562 139750 621574 139802
rect 621626 139799 621638 139802
rect 634330 139799 634342 139802
rect 621626 139753 634342 139799
rect 621626 139750 621638 139753
rect 634330 139750 634342 139753
rect 634394 139750 634406 139802
rect 633658 139687 633670 139690
rect 619896 139641 633670 139687
rect 633658 139638 633670 139641
rect 633722 139638 633734 139690
rect 652586 139687 652598 139690
rect 648905 139641 652598 139687
rect 619546 139526 619558 139578
rect 619610 139575 619622 139578
rect 633210 139575 633222 139578
rect 619610 139529 633222 139575
rect 619610 139526 619622 139529
rect 633210 139526 633222 139529
rect 633274 139526 633286 139578
rect 648905 139466 648951 139641
rect 652586 139638 652598 139641
rect 652650 139638 652662 139690
rect 668714 139638 668726 139690
rect 668778 139687 668790 139690
rect 671514 139687 671526 139690
rect 668778 139641 671526 139687
rect 668778 139638 668790 139641
rect 671514 139638 671526 139641
rect 671578 139638 671590 139690
rect 651914 139575 651926 139578
rect 649129 139529 651926 139575
rect 618986 139414 618998 139466
rect 619050 139463 619062 139466
rect 632090 139463 632102 139466
rect 619050 139417 632102 139463
rect 619050 139414 619062 139417
rect 632090 139414 632102 139417
rect 632154 139414 632166 139466
rect 648890 139414 648902 139466
rect 648954 139414 648966 139466
rect 649129 139354 649175 139529
rect 651914 139526 651926 139529
rect 651978 139526 651990 139578
rect 671626 139575 671638 139578
rect 666936 139529 671638 139575
rect 649226 139414 649238 139466
rect 649290 139463 649302 139466
rect 651690 139463 651702 139466
rect 649290 139417 651702 139463
rect 649290 139414 649302 139417
rect 651690 139414 651702 139417
rect 651754 139414 651766 139466
rect 665802 139414 665814 139466
rect 665866 139463 665878 139466
rect 666936 139463 666982 139529
rect 671626 139526 671638 139529
rect 671690 139526 671702 139578
rect 665866 139417 666982 139463
rect 665866 139414 665878 139417
rect 667146 139414 667158 139466
rect 667210 139463 667222 139466
rect 669498 139463 669510 139466
rect 667210 139417 669510 139463
rect 667210 139414 667222 139417
rect 669498 139414 669510 139417
rect 669562 139414 669574 139466
rect 669834 139414 669846 139466
rect 669898 139463 669910 139466
rect 671290 139463 671302 139466
rect 669898 139417 671302 139463
rect 669898 139414 669910 139417
rect 671290 139414 671302 139417
rect 671354 139414 671366 139466
rect 649114 139302 649126 139354
rect 649178 139302 649190 139354
rect 627498 123559 627510 123562
rect 621576 123513 627510 123559
rect 618538 123062 618550 123114
rect 618602 123111 618614 123114
rect 621576 123111 621622 123513
rect 627498 123510 627510 123513
rect 627562 123510 627574 123562
rect 633098 123510 633110 123562
rect 633162 123559 633174 123562
rect 654714 123559 654726 123562
rect 633162 123513 654726 123559
rect 633162 123510 633174 123513
rect 654714 123510 654726 123513
rect 654778 123510 654790 123562
rect 618602 123065 621622 123111
rect 622473 123401 635062 123447
rect 618602 123062 618614 123065
rect 622473 122999 622519 123401
rect 627498 123286 627510 123338
rect 627562 123335 627574 123338
rect 627562 123289 633382 123335
rect 627562 123286 627574 123289
rect 614856 122953 622519 122999
rect 566010 122838 566022 122890
rect 566074 122887 566086 122890
rect 614856 122887 614902 122953
rect 633336 122887 633382 123289
rect 635016 123223 635062 123401
rect 640953 123401 646822 123447
rect 636906 123286 636918 123338
rect 636970 123286 636982 123338
rect 636921 123223 636967 123286
rect 635016 123177 636967 123223
rect 640953 122887 640999 123401
rect 641162 123286 641174 123338
rect 641226 123286 641238 123338
rect 566074 122841 614902 122887
rect 623593 122841 625095 122887
rect 633336 122841 640999 122887
rect 566074 122838 566086 122841
rect 560186 122726 560198 122778
rect 560250 122775 560262 122778
rect 623593 122775 623639 122841
rect 560250 122729 623639 122775
rect 625049 122775 625095 122841
rect 641177 122775 641223 123286
rect 646776 123223 646822 123401
rect 652362 123335 652374 123338
rect 650136 123289 652374 123335
rect 650136 123223 650182 123289
rect 652362 123286 652374 123289
rect 652426 123286 652438 123338
rect 646776 123177 650182 123223
rect 625049 122729 641223 122775
rect 560250 122726 560262 122729
rect 559402 82182 559414 82234
rect 559466 82231 559478 82234
rect 600506 82231 600518 82234
rect 559466 82185 600518 82231
rect 559466 82182 559478 82185
rect 600506 82182 600518 82185
rect 600570 82182 600582 82234
rect 78026 82070 78038 82122
rect 78090 82119 78102 82122
rect 559514 82119 559526 82122
rect 78090 82073 559526 82119
rect 78090 82070 78102 82073
rect 559514 82070 559526 82073
rect 559578 82070 559590 82122
rect 78250 80950 78262 81002
rect 78314 80999 78326 81002
rect 672074 80999 672086 81002
rect 78314 80953 672086 80999
rect 78314 80950 78326 80953
rect 672074 80950 672086 80953
rect 672138 80950 672150 81002
rect 92362 80838 92374 80890
rect 92426 80887 92438 80890
rect 671962 80887 671974 80890
rect 92426 80841 671974 80887
rect 92426 80838 92438 80841
rect 671962 80838 671974 80841
rect 672026 80838 672038 80890
rect 335962 80726 335974 80778
rect 336026 80775 336038 80778
rect 672970 80775 672982 80778
rect 336026 80729 672982 80775
rect 336026 80726 336038 80729
rect 672970 80726 672982 80729
rect 673034 80726 673046 80778
rect 560298 80614 560310 80666
rect 560362 80663 560374 80666
rect 611706 80663 611718 80666
rect 560362 80617 611718 80663
rect 560362 80614 560374 80617
rect 611706 80614 611718 80617
rect 611770 80614 611782 80666
rect 469130 71766 469142 71818
rect 469194 71815 469206 71818
rect 615290 71815 615302 71818
rect 469194 71769 615302 71815
rect 469194 71766 469206 71769
rect 615290 71766 615302 71769
rect 615354 71766 615366 71818
rect 450986 71654 450998 71706
rect 451050 71703 451062 71706
rect 616634 71703 616646 71706
rect 451050 71657 616646 71703
rect 451050 71654 451062 71657
rect 616634 71654 616646 71657
rect 616698 71654 616710 71706
rect 439898 71542 439910 71594
rect 439962 71591 439974 71594
rect 615962 71591 615974 71594
rect 439962 71545 615974 71591
rect 439962 71542 439974 71545
rect 615962 71542 615974 71545
rect 616026 71542 616038 71594
rect 395882 71430 395894 71482
rect 395946 71479 395958 71482
rect 611930 71479 611942 71482
rect 395946 71433 611942 71479
rect 395946 71430 395958 71433
rect 611930 71430 611942 71433
rect 611994 71430 612006 71482
rect 340890 71318 340902 71370
rect 340954 71367 340966 71370
rect 613274 71367 613286 71370
rect 340954 71321 613286 71367
rect 340954 71318 340966 71321
rect 613274 71318 613286 71321
rect 613338 71318 613350 71370
<< via1 >>
rect 73222 946038 73274 946090
rect 77590 945702 77642 945754
rect 105814 942342 105866 942394
rect 196534 942342 196586 942394
rect 216358 942342 216410 942394
rect 306518 942342 306570 942394
rect 161142 942230 161194 942282
rect 251302 942230 251354 942282
rect 270454 942230 270506 942282
rect 361174 942230 361226 942282
rect 160358 942118 160410 942170
rect 251078 942118 251130 942170
rect 271350 942118 271402 942170
rect 335862 942118 335914 942170
rect 106374 942006 106426 942058
rect 196310 942006 196362 942058
rect 215574 942006 215626 942058
rect 306070 942006 306122 942058
rect 177046 938198 177098 938250
rect 687766 938198 687818 938250
rect 341014 937414 341066 937466
rect 344598 937414 344650 937466
rect 120934 937302 120986 937354
rect 688214 937302 688266 937354
rect 505654 936966 505706 937018
rect 689222 936966 689274 937018
rect 453574 936854 453626 936906
rect 687318 936854 687370 936906
rect 450214 936742 450266 936794
rect 687654 936742 687706 936794
rect 344710 936630 344762 936682
rect 687542 936630 687594 936682
rect 84758 936518 84810 936570
rect 141542 936518 141594 936570
rect 233830 936518 233882 936570
rect 688102 936518 688154 936570
rect 176710 935622 176762 935674
rect 185782 935622 185834 935674
rect 176486 935398 176538 935450
rect 208070 935398 208122 935450
rect 630422 935398 630474 935450
rect 674102 935398 674154 935450
rect 341014 935286 341066 935338
rect 289158 935174 289210 935226
rect 296326 935174 296378 935226
rect 282438 935062 282490 935114
rect 318950 935062 319002 935114
rect 385254 934950 385306 935002
rect 497366 934950 497418 935002
rect 507446 934950 507498 935002
rect 342582 934838 342634 934890
rect 407430 934838 407482 934890
rect 453350 934838 453402 934890
rect 458502 934838 458554 934890
rect 700422 739062 700474 739114
rect 701318 739062 701370 739114
rect 700422 712070 700474 712122
rect 704566 712070 704618 712122
rect 72998 618102 73050 618154
rect 73446 618102 73498 618154
rect 77702 618102 77754 618154
rect 78374 617990 78426 618042
rect 73222 536118 73274 536170
rect 77478 535782 77530 535834
rect 72998 413142 73050 413194
rect 78262 413142 78314 413194
rect 73446 413030 73498 413082
rect 78374 413030 78426 413082
rect 284230 333510 284282 333562
rect 423894 333510 423946 333562
rect 266534 333398 266586 333450
rect 376294 333398 376346 333450
rect 403398 333398 403450 333450
rect 465558 333398 465610 333450
rect 611046 333398 611098 333450
rect 688102 333398 688154 333450
rect 369686 333286 369738 333338
rect 483814 333286 483866 333338
rect 488406 333286 488458 333338
rect 632438 333286 632490 333338
rect 139190 333174 139242 333226
rect 179846 333174 179898 333226
rect 269110 333174 269162 333226
rect 382118 333174 382170 333226
rect 454806 333174 454858 333226
rect 596710 333174 596762 333226
rect 132582 333062 132634 333114
rect 177718 333062 177770 333114
rect 221398 333062 221450 333114
rect 251638 333062 251690 333114
rect 275382 333062 275434 333114
rect 400710 333062 400762 333114
rect 420870 333062 420922 333114
rect 502070 333062 502122 333114
rect 102678 332950 102730 333002
rect 151958 332950 152010 333002
rect 154422 332950 154474 333002
rect 184998 332950 185050 333002
rect 196086 332950 196138 333002
rect 200230 332950 200282 333002
rect 223638 332950 223690 333002
rect 257574 332950 257626 333002
rect 320070 332950 320122 333002
rect 448310 332950 448362 333002
rect 471158 332950 471210 333002
rect 615302 332950 615354 333002
rect 110630 332838 110682 332890
rect 167974 332838 168026 332890
rect 188022 332838 188074 332890
rect 196646 332838 196698 332890
rect 227222 332838 227274 332890
rect 271462 332838 271514 332890
rect 279750 332838 279802 332890
rect 412582 332838 412634 332890
rect 437558 332838 437610 332890
rect 585510 332838 585562 332890
rect 90806 332726 90858 332778
rect 150614 332726 150666 332778
rect 152406 332726 152458 332778
rect 183542 332726 183594 332778
rect 190150 332726 190202 332778
rect 197878 332726 197930 332778
rect 205382 332726 205434 332778
rect 211878 332726 211930 332778
rect 212102 332726 212154 332778
rect 229798 332726 229850 332778
rect 231590 332726 231642 332778
rect 283446 332726 283498 332778
rect 288486 332726 288538 332778
rect 436438 332726 436490 332778
rect 471382 332726 471434 332778
rect 621238 332726 621290 332778
rect 86886 332614 86938 332666
rect 160246 332614 160298 332666
rect 192166 332614 192218 332666
rect 199558 332614 199610 332666
rect 206838 332614 206890 332666
rect 213894 332614 213946 332666
rect 217478 332614 217530 332666
rect 233718 332614 233770 332666
rect 233942 332614 233994 332666
rect 289382 332614 289434 332666
rect 421318 332614 421370 332666
rect 573526 332614 573578 332666
rect 78822 332502 78874 332554
rect 672310 332502 672362 332554
rect 327238 332390 327290 332442
rect 541718 332390 541770 332442
rect 331494 332278 331546 332330
rect 553702 332278 553754 332330
rect 278966 332166 279018 332218
rect 410566 332166 410618 332218
rect 411350 332166 411402 332218
rect 653046 332166 653098 332218
rect 343814 332054 343866 332106
rect 587414 332054 587466 332106
rect 352550 331942 352602 331994
rect 611270 331942 611322 331994
rect 379318 331830 379370 331882
rect 676902 331830 676954 331882
rect 80054 331718 80106 331770
rect 672422 331718 672474 331770
rect 326006 331606 326058 331658
rect 539814 331606 539866 331658
rect 319846 331494 319898 331546
rect 523910 331494 523962 331546
rect 283334 331382 283386 331434
rect 422550 331382 422602 331434
rect 281206 331270 281258 331322
rect 416614 331270 416666 331322
rect 276838 331158 276890 331210
rect 404630 331158 404682 331210
rect 73222 331046 73274 331098
rect 78262 330822 78314 330874
rect 294310 330822 294362 330874
rect 452342 330822 452394 330874
rect 298678 330710 298730 330762
rect 464214 330710 464266 330762
rect 305174 330598 305226 330650
rect 482134 330598 482186 330650
rect 309542 330486 309594 330538
rect 494118 330486 494170 330538
rect 249398 330374 249450 330426
rect 307302 330374 307354 330426
rect 313910 330374 313962 330426
rect 505990 330374 506042 330426
rect 240214 330262 240266 330314
rect 309318 330262 309370 330314
rect 322646 330262 322698 330314
rect 529846 330262 529898 330314
rect 243238 330150 243290 330202
rect 313238 330150 313290 330202
rect 354790 330150 354842 330202
rect 617318 330150 617370 330202
rect 244022 330038 244074 330090
rect 315254 330038 315306 330090
rect 354566 330038 354618 330090
rect 619222 330038 619274 330090
rect 292070 329926 292122 329978
rect 446406 329926 446458 329978
rect 289942 329814 289994 329866
rect 421766 329814 421818 329866
rect 247718 329142 247770 329194
rect 325222 329142 325274 329194
rect 353894 329142 353946 329194
rect 577558 329142 577610 329194
rect 248502 329030 248554 329082
rect 327126 329030 327178 329082
rect 335302 329030 335354 329082
rect 563670 329030 563722 329082
rect 250630 328918 250682 328970
rect 333062 328918 333114 328970
rect 346726 328918 346778 328970
rect 595366 328918 595418 328970
rect 128550 328806 128602 328858
rect 175478 328806 175530 328858
rect 252870 328806 252922 328858
rect 339110 328806 339162 328858
rect 351206 328806 351258 328858
rect 607350 328806 607402 328858
rect 256454 328694 256506 328746
rect 348966 328694 349018 328746
rect 357702 328694 357754 328746
rect 625270 328694 625322 328746
rect 124630 328582 124682 328634
rect 174806 328582 174858 328634
rect 260822 328582 260874 328634
rect 360950 328582 361002 328634
rect 362182 328582 362234 328634
rect 637142 328582 637194 328634
rect 120598 328470 120650 328522
rect 172566 328470 172618 328522
rect 267430 328470 267482 328522
rect 378870 328470 378922 328522
rect 384694 328470 384746 328522
rect 664918 328470 664970 328522
rect 122502 328358 122554 328410
rect 173350 328358 173402 328410
rect 263062 328358 263114 328410
rect 366886 328358 366938 328410
rect 369574 328358 369626 328410
rect 655062 328358 655114 328410
rect 231030 328246 231082 328298
rect 279414 328246 279466 328298
rect 319062 328246 319114 328298
rect 519878 328246 519930 328298
rect 228790 328134 228842 328186
rect 273478 328134 273530 328186
rect 301702 328134 301754 328186
rect 472166 328134 472218 328186
rect 228118 328022 228170 328074
rect 269558 328022 269610 328074
rect 276166 328022 276218 328074
rect 402614 328022 402666 328074
rect 226662 327910 226714 327962
rect 267542 327910 267594 327962
rect 297222 327910 297274 327962
rect 386038 327910 386090 327962
rect 289270 327462 289322 327514
rect 438454 327462 438506 327514
rect 306742 327350 306794 327402
rect 486166 327350 486218 327402
rect 313350 327238 313402 327290
rect 503974 327238 504026 327290
rect 315478 327126 315530 327178
rect 509910 327126 509962 327178
rect 322086 327014 322138 327066
rect 527830 327014 527882 327066
rect 333062 326902 333114 326954
rect 557622 326902 557674 326954
rect 348294 326790 348346 326842
rect 599398 326790 599450 326842
rect 363638 326678 363690 326730
rect 641062 326678 641114 326730
rect 284902 326566 284954 326618
rect 426470 326566 426522 326618
rect 280422 326454 280474 326506
rect 414598 326454 414650 326506
rect 299798 326342 299850 326394
rect 432518 326342 432570 326394
rect 351990 325782 352042 325834
rect 454694 325782 454746 325834
rect 312566 325670 312618 325722
rect 420870 325670 420922 325722
rect 264518 325558 264570 325610
rect 319734 325558 319786 325610
rect 356358 325558 356410 325610
rect 471382 325558 471434 325610
rect 485494 325558 485546 325610
rect 668614 325558 668666 325610
rect 310438 325446 310490 325498
rect 495574 325446 495626 325498
rect 314806 325334 314858 325386
rect 507334 325334 507386 325386
rect 262278 325222 262330 325274
rect 320182 325222 320234 325274
rect 323542 325222 323594 325274
rect 530854 325222 530906 325274
rect 271798 325110 271850 325162
rect 335078 325110 335130 325162
rect 362742 325110 362794 325162
rect 638374 325110 638426 325162
rect 265974 324998 266026 325050
rect 335190 324998 335242 325050
rect 365094 324998 365146 325050
rect 645094 324998 645146 325050
rect 343254 324886 343306 324938
rect 437558 324886 437610 324938
rect 338886 324774 338938 324826
rect 421318 324774 421370 324826
rect 340902 324662 340954 324714
rect 421094 324662 421146 324714
rect 161366 324214 161418 324266
rect 162598 324214 162650 324266
rect 280646 324214 280698 324266
rect 281934 324214 281986 324266
rect 354566 324214 354618 324266
rect 355518 324214 355570 324266
rect 95734 324102 95786 324154
rect 155206 324102 155258 324154
rect 155430 324102 155482 324154
rect 163214 324102 163266 324154
rect 203366 324102 203418 324154
rect 204654 324102 204706 324154
rect 375230 324102 375282 324154
rect 377862 324102 377914 324154
rect 133702 323990 133754 324042
rect 164670 323990 164722 324042
rect 372318 323990 372370 324042
rect 384694 323990 384746 324042
rect 94054 323878 94106 323930
rect 155318 323878 155370 323930
rect 155206 323766 155258 323818
rect 163886 323878 163938 323930
rect 287086 323878 287138 323930
rect 299798 323878 299850 323930
rect 370078 323878 370130 323930
rect 385478 323878 385530 323930
rect 673206 308758 673258 308810
rect 178054 308646 178106 308698
rect 179678 308646 179730 308698
rect 228398 308646 228450 308698
rect 282326 308646 282378 308698
rect 283838 308646 283890 308698
rect 315926 308646 315978 308698
rect 317438 308646 317490 308698
rect 377302 308646 377354 308698
rect 233830 308534 233882 308586
rect 171446 308422 171498 308474
rect 172958 308422 173010 308474
rect 208518 308422 208570 308474
rect 216190 308422 216242 308474
rect 225374 308422 225426 308474
rect 226774 308422 226826 308474
rect 227838 308422 227890 308474
rect 231814 308422 231866 308474
rect 243574 308422 243626 308474
rect 244862 308422 244914 308474
rect 247046 308422 247098 308474
rect 248558 308422 248610 308474
rect 248726 308422 248778 308474
rect 249790 308422 249842 308474
rect 253654 308422 253706 308474
rect 255278 308422 255330 308474
rect 259534 308534 259586 308586
rect 326510 308534 326562 308586
rect 327462 308534 327514 308586
rect 336086 308422 336138 308474
rect 336926 308422 336978 308474
rect 337766 308422 337818 308474
rect 338718 308422 338770 308474
rect 258806 308310 258858 308362
rect 247942 308198 247994 308250
rect 273926 308198 273978 308250
rect 191830 308086 191882 308138
rect 208854 308086 208906 308138
rect 156214 307974 156266 308026
rect 191606 307974 191658 308026
rect 235062 307974 235114 308026
rect 247158 307974 247210 308026
rect 292518 307974 292570 308026
rect 368230 307974 368282 308026
rect 95734 307862 95786 307914
rect 163158 307862 163210 307914
rect 205158 307862 205210 307914
rect 214902 307862 214954 307914
rect 243126 307862 243178 307914
rect 263958 307862 264010 307914
rect 319286 307862 319338 307914
rect 423334 307862 423386 307914
rect 97414 307750 97466 307802
rect 163718 307750 163770 307802
rect 201574 307750 201626 307802
rect 213110 307750 213162 307802
rect 235734 307750 235786 307802
rect 248614 307750 248666 307802
rect 280310 307750 280362 307802
rect 316598 307750 316650 307802
rect 327462 307750 327514 307802
rect 440246 307750 440298 307802
rect 94278 307638 94330 307690
rect 161926 307638 161978 307690
rect 166406 307638 166458 307690
rect 196534 307638 196586 307690
rect 203366 307638 203418 307690
rect 214342 307638 214394 307690
rect 236966 307638 237018 307690
rect 250518 307638 250570 307690
rect 251638 307638 251690 307690
rect 282214 307638 282266 307690
rect 337542 307638 337594 307690
rect 467798 307638 467850 307690
rect 94054 307526 94106 307578
rect 162486 307526 162538 307578
rect 147814 307414 147866 307466
rect 187462 307526 187514 307578
rect 206726 307526 206778 307578
rect 215574 307526 215626 307578
rect 239430 307526 239482 307578
rect 257014 307526 257066 307578
rect 261942 307526 261994 307578
rect 304054 307526 304106 307578
rect 357702 307526 357754 307578
rect 509798 307526 509850 307578
rect 186790 307414 186842 307466
rect 205830 307414 205882 307466
rect 226662 307414 226714 307466
rect 230246 307414 230298 307466
rect 236406 307414 236458 307466
rect 250294 307414 250346 307466
rect 258358 307414 258410 307466
rect 295990 307414 296042 307466
rect 363862 307414 363914 307466
rect 520886 307414 520938 307466
rect 358374 307302 358426 307354
rect 509910 307302 509962 307354
rect 366102 307190 366154 307242
rect 526822 307190 526874 307242
rect 365654 307078 365706 307130
rect 526598 307078 526650 307130
rect 291286 306966 291338 307018
rect 364646 306966 364698 307018
rect 366886 306966 366938 307018
rect 528278 306966 528330 307018
rect 291846 306854 291898 306906
rect 366214 306854 366266 306906
rect 368118 306854 368170 306906
rect 531638 306854 531690 306906
rect 83750 306742 83802 306794
rect 660998 306742 661050 306794
rect 83638 306630 83690 306682
rect 662678 306630 662730 306682
rect 77254 306518 77306 306570
rect 672310 306518 672362 306570
rect 160022 305846 160074 305898
rect 336870 305846 336922 305898
rect 84758 305734 84810 305786
rect 655958 305734 656010 305786
rect 349190 305622 349242 305674
rect 491318 305622 491370 305674
rect 174806 305510 174858 305562
rect 175366 305510 175418 305562
rect 350982 305510 351034 305562
rect 494678 305510 494730 305562
rect 350422 305398 350474 305450
rect 494902 305398 494954 305450
rect 353446 305286 353498 305338
rect 499718 305286 499770 305338
rect 354006 305174 354058 305226
rect 501398 305174 501450 305226
rect 354678 305062 354730 305114
rect 502294 305062 502346 305114
rect 355910 304950 355962 305002
rect 504758 304950 504810 305002
rect 355238 304838 355290 304890
rect 503974 304838 504026 304890
rect 347398 304726 347450 304778
rect 487958 304726 488010 304778
rect 340006 304614 340058 304666
rect 472054 304614 472106 304666
rect 340678 303942 340730 303994
rect 472838 303942 472890 303994
rect 341910 303830 341962 303882
rect 475414 303830 475466 303882
rect 343030 303718 343082 303770
rect 477878 303718 477930 303770
rect 346166 303606 346218 303658
rect 483814 303606 483866 303658
rect 361398 303494 361450 303546
rect 516518 303494 516570 303546
rect 360166 303382 360218 303434
rect 514838 303382 514890 303434
rect 361958 303270 362010 303322
rect 518198 303270 518250 303322
rect 168758 303158 168810 303210
rect 184438 303158 184490 303210
rect 360726 303158 360778 303210
rect 516742 303158 516794 303210
rect 298230 302262 298282 302314
rect 335862 302262 335914 302314
rect 297446 301702 297498 301754
rect 335078 301702 335130 301754
rect 659318 301702 659370 301754
rect 670742 301702 670794 301754
rect 295878 301590 295930 301642
rect 335302 301590 335354 301642
rect 660998 301590 661050 301642
rect 670966 301590 671018 301642
rect 287478 301478 287530 301530
rect 357814 301478 357866 301530
rect 655958 301478 656010 301530
rect 670294 301478 670346 301530
rect 299462 300470 299514 300522
rect 383014 300470 383066 300522
rect 301030 300358 301082 300410
rect 386374 300358 386426 300410
rect 299238 300246 299290 300298
rect 384694 300246 384746 300298
rect 300806 300134 300858 300186
rect 386934 300134 386986 300186
rect 304166 300022 304218 300074
rect 394774 300022 394826 300074
rect 310886 299910 310938 299962
rect 408662 299910 408714 299962
rect 83302 299798 83354 299850
rect 654502 299798 654554 299850
rect 337542 293974 337594 294026
rect 670406 293974 670458 294026
rect 467014 293862 467066 293914
rect 467798 293862 467850 293914
rect 487174 293862 487226 293914
rect 487958 293862 488010 293914
rect 495798 293862 495850 293914
rect 496358 293862 496410 293914
rect 515734 293862 515786 293914
rect 516742 293862 516794 293914
rect 517526 293862 517578 293914
rect 518198 293862 518250 293914
rect 519094 293526 519146 293578
rect 520550 293526 520602 293578
rect 492214 293414 492266 293466
rect 492998 293414 493050 293466
rect 494006 293414 494058 293466
rect 494902 293414 494954 293466
rect 566022 293414 566074 293466
rect 645430 293414 645482 293466
rect 520774 293302 520826 293354
rect 522342 293302 522394 293354
rect 631430 293302 631482 293354
rect 520550 293190 520602 293242
rect 630982 293190 631034 293242
rect 494902 293078 494954 293130
rect 606230 293078 606282 293130
rect 516742 292966 516794 293018
rect 629526 292966 629578 293018
rect 517526 292854 517578 292906
rect 630534 292854 630586 292906
rect 492998 292742 493050 292794
rect 613510 292742 613562 292794
rect 487174 292630 487226 292682
rect 606342 292630 606394 292682
rect 495798 292518 495850 292570
rect 500838 292406 500890 292458
rect 501398 292406 501450 292458
rect 508230 292406 508282 292458
rect 508566 292518 508618 292570
rect 624262 292518 624314 292570
rect 622358 292406 622410 292458
rect 467014 292294 467066 292346
rect 643974 292294 644026 292346
rect 92486 292182 92538 292234
rect 609814 292182 609866 292234
rect 529174 292070 529226 292122
rect 529958 292070 530010 292122
rect 531078 292070 531130 292122
rect 531638 292070 531690 292122
rect 530854 291958 530906 292010
rect 532422 291958 532474 292010
rect 610822 291958 610874 292010
rect 617990 291958 618042 292010
rect 612390 291846 612442 291898
rect 615750 291846 615802 291898
rect 322534 291734 322586 291786
rect 433414 291734 433466 291786
rect 609926 291734 609978 291786
rect 620678 291734 620730 291786
rect 324102 291622 324154 291674
rect 435206 291622 435258 291674
rect 504758 291622 504810 291674
rect 625718 291622 625770 291674
rect 334518 291510 334570 291562
rect 456038 291510 456090 291562
rect 531078 291510 531130 291562
rect 635350 291510 635402 291562
rect 334630 291398 334682 291450
rect 457382 291398 457434 291450
rect 532422 291398 532474 291450
rect 635798 291398 635850 291450
rect 529174 291286 529226 291338
rect 634790 291286 634842 291338
rect 528278 291174 528330 291226
rect 634342 291174 634394 291226
rect 525814 291062 525866 291114
rect 526822 291062 526874 291114
rect 633894 291062 633946 291114
rect 516518 290950 516570 291002
rect 629974 290950 630026 291002
rect 509910 290838 509962 290890
rect 627622 290838 627674 290890
rect 610710 290726 610762 290778
rect 612726 290726 612778 290778
rect 620678 290726 620730 290778
rect 669846 290726 669898 290778
rect 92598 290614 92650 290666
rect 612390 290614 612442 290666
rect 615750 290614 615802 290666
rect 671302 290614 671354 290666
rect 606342 290502 606394 290554
rect 612502 290502 612554 290554
rect 612838 290502 612890 290554
rect 618998 290502 619050 290554
rect 651142 290502 651194 290554
rect 689334 290502 689386 290554
rect 605782 290390 605834 290442
rect 619446 290390 619498 290442
rect 650246 290390 650298 290442
rect 688214 290390 688266 290442
rect 606118 290278 606170 290330
rect 610822 290278 610874 290330
rect 611046 290278 611098 290330
rect 614742 290278 614794 290330
rect 655958 290278 656010 290330
rect 606342 290166 606394 290218
rect 613174 290166 613226 290218
rect 615190 290166 615242 290218
rect 615638 290166 615690 290218
rect 654054 290166 654106 290218
rect 668166 290166 668218 290218
rect 670070 290278 670122 290330
rect 670742 290278 670794 290330
rect 670294 290166 670346 290218
rect 610822 290054 610874 290106
rect 613734 290054 613786 290106
rect 649686 290054 649738 290106
rect 688886 290054 688938 290106
rect 80390 289942 80442 289994
rect 659766 289942 659818 289994
rect 660326 289942 660378 289994
rect 670966 289942 671018 289994
rect 78710 289830 78762 289882
rect 661222 289830 661274 289882
rect 664582 289830 664634 289882
rect 670630 289830 670682 289882
rect 80166 289718 80218 289770
rect 665590 289718 665642 289770
rect 78710 289606 78762 289658
rect 667942 289718 667994 289770
rect 668950 289718 669002 289770
rect 670294 289718 670346 289770
rect 671862 289718 671914 289770
rect 687430 289718 687482 289770
rect 668166 289606 668218 289658
rect 672198 289606 672250 289658
rect 606342 288822 606394 288874
rect 611382 288822 611434 288874
rect 606230 288710 606282 288762
rect 610822 288710 610874 288762
rect 105814 285574 105866 285626
rect 106486 285574 106538 285626
rect 196870 285574 196922 285626
rect 197430 285574 197482 285626
rect 278854 285574 278906 285626
rect 279414 285574 279466 285626
rect 525814 285574 525866 285626
rect 526598 285574 526650 285626
rect 542614 285574 542666 285626
rect 543286 285574 543338 285626
rect 331046 285014 331098 285066
rect 451670 285014 451722 285066
rect 329366 284902 329418 284954
rect 449206 284902 449258 284954
rect 332838 284790 332890 284842
rect 454246 284790 454298 284842
rect 332950 284678 333002 284730
rect 455590 284678 455642 284730
rect 530854 282774 530906 282826
rect 531750 282774 531802 282826
rect 331382 282102 331434 282154
rect 332166 282102 332218 282154
rect 345158 281878 345210 281930
rect 352438 281878 352490 281930
rect 335302 281766 335354 281818
rect 378758 281766 378810 281818
rect 301702 281654 301754 281706
rect 345382 281654 345434 281706
rect 335078 281542 335130 281594
rect 379990 281542 380042 281594
rect 165622 281430 165674 281482
rect 173126 281430 173178 281482
rect 173910 281430 173962 281482
rect 179846 281430 179898 281482
rect 265750 281430 265802 281482
rect 313350 281430 313402 281482
rect 334630 281430 334682 281482
rect 396678 281430 396730 281482
rect 166070 281318 166122 281370
rect 131462 281206 131514 281258
rect 177942 281206 177994 281258
rect 195078 281318 195130 281370
rect 265526 281318 265578 281370
rect 314694 281318 314746 281370
rect 334406 281318 334458 281370
rect 408214 281318 408266 281370
rect 132806 281094 132858 281146
rect 173910 281094 173962 281146
rect 128326 280982 128378 281034
rect 176486 280982 176538 281034
rect 130902 280870 130954 280922
rect 178278 280870 178330 280922
rect 124182 280758 124234 280810
rect 174694 280758 174746 280810
rect 196646 281094 196698 281146
rect 200118 281094 200170 281146
rect 110406 280646 110458 280698
rect 120598 280646 120650 280698
rect 165622 280646 165674 280698
rect 167862 280646 167914 280698
rect 169206 280646 169258 280698
rect 180742 280646 180794 280698
rect 255558 281206 255610 281258
rect 268886 281206 268938 281258
rect 319846 281206 319898 281258
rect 320070 281206 320122 281258
rect 397910 281206 397962 281258
rect 255446 281094 255498 281146
rect 268998 281094 269050 281146
rect 321078 281094 321130 281146
rect 331942 281094 331994 281146
rect 335190 281094 335242 281146
rect 335526 281094 335578 281146
rect 417174 281094 417226 281146
rect 291174 280982 291226 281034
rect 307526 280982 307578 281034
rect 401494 280982 401546 281034
rect 292294 280870 292346 280922
rect 312678 280870 312730 280922
rect 413030 280870 413082 280922
rect 273030 280758 273082 280810
rect 275606 280646 275658 280698
rect 289718 280758 289770 280810
rect 347734 280758 347786 280810
rect 325894 280646 325946 280698
rect 331942 280646 331994 280698
rect 332166 280646 332218 280698
rect 352438 280646 352490 280698
rect 358486 280646 358538 280698
rect 362742 280758 362794 280810
rect 375510 280758 375562 280810
rect 377862 280646 377914 280698
rect 378086 280758 378138 280810
rect 552694 280758 552746 280810
rect 450214 280646 450266 280698
rect 553590 280646 553642 280698
rect 693254 236742 693306 236794
rect 700534 236742 700586 236794
rect 73446 208070 73498 208122
rect 78262 208070 78314 208122
rect 560198 139862 560250 139914
rect 647894 139862 647946 139914
rect 619782 139750 619834 139802
rect 621574 139750 621626 139802
rect 634342 139750 634394 139802
rect 633670 139638 633722 139690
rect 619558 139526 619610 139578
rect 633222 139526 633274 139578
rect 652598 139638 652650 139690
rect 668726 139638 668778 139690
rect 671526 139638 671578 139690
rect 618998 139414 619050 139466
rect 632102 139414 632154 139466
rect 648902 139414 648954 139466
rect 651926 139526 651978 139578
rect 649238 139414 649290 139466
rect 651702 139414 651754 139466
rect 665814 139414 665866 139466
rect 671638 139526 671690 139578
rect 667158 139414 667210 139466
rect 669510 139414 669562 139466
rect 669846 139414 669898 139466
rect 671302 139414 671354 139466
rect 649126 139302 649178 139354
rect 618550 123062 618602 123114
rect 627510 123510 627562 123562
rect 633110 123510 633162 123562
rect 654726 123510 654778 123562
rect 627510 123286 627562 123338
rect 566022 122838 566074 122890
rect 636918 123286 636970 123338
rect 641174 123286 641226 123338
rect 560198 122726 560250 122778
rect 652374 123286 652426 123338
rect 559414 82182 559466 82234
rect 600518 82182 600570 82234
rect 78038 82070 78090 82122
rect 559526 82070 559578 82122
rect 78262 80950 78314 81002
rect 672086 80950 672138 81002
rect 92374 80838 92426 80890
rect 671974 80838 672026 80890
rect 335974 80726 336026 80778
rect 672982 80726 673034 80778
rect 560310 80614 560362 80666
rect 611718 80614 611770 80666
rect 469142 71766 469194 71818
rect 615302 71766 615354 71818
rect 450998 71654 451050 71706
rect 616646 71654 616698 71706
rect 439910 71542 439962 71594
rect 615974 71542 616026 71594
rect 395894 71430 395946 71482
rect 611942 71430 611994 71482
rect 340902 71318 340954 71370
rect 613286 71318 613338 71370
<< metal2 >>
rect 490868 949228 490924 949238
rect 106586 947732 106596 947788
rect 106652 947732 106662 947788
rect 141120 947732 141484 947788
rect 105588 947284 105840 947340
rect 141120 947284 141372 947340
rect 72772 946092 72828 946102
rect 73220 946092 73276 946102
rect 72688 946036 72772 946092
rect 73136 946090 73276 946092
rect 73136 946038 73222 946090
rect 73274 946038 73276 946090
rect 73136 946036 73276 946038
rect 72772 946026 72828 946036
rect 73220 946026 73276 946036
rect 77476 946092 77532 946102
rect 77252 945980 77308 945990
rect 73556 945868 73612 945878
rect 73556 945802 73612 945812
rect 72212 945756 72268 945766
rect 72212 945690 72268 945700
rect 72996 910924 73052 910934
rect 72212 910588 72268 910896
rect 72688 910868 72996 910924
rect 73136 910868 73500 910924
rect 72996 910858 73052 910868
rect 73444 910812 73500 910868
rect 73444 910746 73500 910756
rect 73556 910700 73612 910896
rect 73556 910634 73612 910644
rect 72212 910522 72268 910532
rect 73780 782124 73836 782134
rect 73584 782068 73780 782124
rect 73780 782058 73836 782068
rect 72660 781900 72716 781910
rect 72660 781834 72716 781844
rect 72212 781788 72268 781798
rect 72212 781722 72268 781732
rect 73108 781676 73164 781686
rect 73108 781610 73164 781620
rect 73556 747516 73612 747526
rect 73556 747450 73612 747460
rect 72660 747404 72716 747414
rect 72660 747338 72716 747348
rect 72212 747292 72268 747302
rect 72212 747226 72268 747236
rect 77252 747292 77308 945924
rect 77364 945868 77420 945878
rect 77364 747404 77420 945812
rect 77476 747516 77532 946036
rect 105588 945868 105644 947284
rect 141316 947100 141372 947284
rect 141428 947100 141484 947732
rect 160244 947732 160832 947788
rect 196112 947732 196700 947788
rect 216570 947732 216580 947788
rect 216636 947732 216646 947788
rect 141876 947100 141932 947110
rect 141428 947044 141596 947100
rect 141316 947034 141372 947044
rect 106260 946652 106316 946864
rect 141120 946836 141484 946892
rect 106260 946586 106316 946596
rect 106260 945868 106316 945878
rect 105588 945812 105868 945868
rect 77476 747450 77532 747460
rect 77588 945754 77644 945766
rect 77588 945702 77590 945754
rect 77642 945702 77644 945754
rect 77364 747338 77420 747348
rect 77252 747226 77308 747236
rect 73108 747180 73164 747190
rect 73108 747114 73164 747124
rect 77588 747180 77644 945702
rect 85204 942844 85260 942854
rect 84756 936570 84812 936582
rect 84756 936518 84758 936570
rect 84810 936518 84812 936570
rect 84084 935788 84140 935798
rect 83972 929852 84028 929862
rect 79716 927388 79772 927398
rect 78372 782124 78428 782134
rect 78148 781900 78204 781910
rect 77588 747114 77644 747124
rect 77700 781788 77756 781798
rect 72772 741132 72828 741142
rect 72688 741076 72772 741132
rect 72772 741066 72828 741076
rect 77476 741132 77532 741142
rect 73556 740908 73612 740918
rect 73556 740842 73612 740852
rect 77364 740908 77420 740918
rect 72212 740796 72268 740806
rect 72212 740730 72268 740740
rect 73108 740684 73164 740694
rect 73108 740618 73164 740628
rect 77252 740684 77308 740694
rect 77252 738108 77308 740628
rect 77252 738042 77308 738052
rect 77364 714027 77420 740852
rect 77252 713971 77420 714027
rect 73108 706636 73164 706646
rect 73108 706570 73164 706580
rect 72212 706524 72268 706534
rect 72212 706458 72268 706468
rect 73556 706412 73612 706422
rect 73556 706346 73612 706356
rect 72660 706300 72716 706310
rect 72660 706234 72716 706244
rect 72548 700140 72604 700150
rect 72240 700084 72548 700140
rect 72548 700074 72604 700084
rect 73108 699916 73164 699926
rect 73108 699850 73164 699860
rect 72660 699804 72716 699814
rect 72660 699738 72716 699748
rect 73556 699692 73612 699702
rect 73556 699626 73612 699636
rect 73556 665196 73612 665206
rect 73556 665130 73612 665140
rect 72660 665084 72716 665094
rect 72660 665018 72716 665028
rect 77252 665084 77308 713971
rect 77476 665196 77532 741076
rect 77700 706524 77756 781732
rect 77924 781676 77980 781686
rect 77700 706458 77756 706468
rect 77812 741020 77868 741030
rect 77700 699804 77756 699814
rect 77476 665130 77532 665140
rect 77588 699692 77644 699702
rect 77252 665018 77308 665028
rect 72548 664972 72604 664982
rect 72240 664916 72548 664972
rect 72548 664906 72604 664916
rect 73444 664860 73500 664870
rect 73136 664804 73444 664860
rect 73444 664794 73500 664804
rect 72324 659148 72380 659158
rect 72240 659092 72324 659148
rect 72324 659082 72380 659092
rect 73108 658924 73164 658934
rect 73108 658858 73164 658868
rect 73556 658812 73612 658822
rect 73556 658746 73612 658756
rect 77476 658812 77532 658822
rect 72660 658700 72716 658710
rect 72660 658634 72716 658644
rect 77252 658700 77308 658710
rect 72660 624652 72716 624662
rect 72660 624586 72716 624596
rect 73556 624540 73612 624550
rect 73556 624474 73612 624484
rect 73108 624428 73164 624438
rect 73108 624362 73164 624372
rect 72212 624316 72268 624326
rect 72212 624250 72268 624260
rect 72996 618156 73052 618166
rect 73444 618156 73500 618166
rect 72688 618154 73052 618156
rect 72688 618102 72998 618154
rect 73050 618102 73052 618154
rect 72688 618100 73052 618102
rect 73136 618154 73500 618156
rect 73136 618102 73446 618154
rect 73498 618102 73500 618154
rect 73136 618100 73500 618102
rect 72996 618090 73052 618100
rect 73444 618090 73500 618100
rect 72212 617708 72268 617718
rect 72212 617642 72268 617652
rect 73556 617596 73612 617606
rect 73556 617530 73612 617540
rect 73444 582876 73500 582886
rect 72212 582540 72268 582848
rect 72660 582652 72716 582848
rect 73136 582820 73444 582876
rect 73584 582820 73836 582876
rect 73444 582810 73500 582820
rect 73780 582764 73836 582820
rect 73780 582698 73836 582708
rect 77252 582764 77308 658644
rect 77252 582698 77308 582708
rect 72660 582586 72716 582596
rect 77476 582652 77532 658756
rect 77588 624652 77644 699636
rect 77588 624586 77644 624596
rect 77700 624540 77756 699748
rect 77812 664972 77868 740964
rect 77924 706636 77980 781620
rect 77924 706570 77980 706580
rect 78036 722428 78092 722438
rect 77812 664906 77868 664916
rect 77924 699916 77980 699926
rect 77700 624474 77756 624484
rect 77924 624428 77980 699860
rect 77924 624362 77980 624372
rect 77700 618154 77756 618166
rect 77700 618102 77702 618154
rect 77754 618102 77756 618154
rect 77476 582586 77532 582596
rect 77588 617596 77644 617606
rect 72212 582474 72268 582484
rect 72212 576940 72268 576950
rect 72212 576874 72268 576884
rect 73556 576828 73612 576838
rect 73556 576762 73612 576772
rect 72660 576716 72716 576726
rect 72660 576650 72716 576660
rect 73108 576604 73164 576614
rect 73108 576538 73164 576548
rect 73108 542556 73164 542566
rect 73108 542490 73164 542500
rect 73556 542444 73612 542454
rect 73556 542378 73612 542388
rect 72212 542332 72268 542342
rect 72212 542266 72268 542276
rect 72660 542220 72716 542230
rect 72660 542154 72716 542164
rect 77588 542220 77644 617540
rect 77700 562716 77756 618102
rect 77700 562650 77756 562660
rect 77812 576716 77868 576726
rect 77588 542154 77644 542164
rect 73220 536172 73276 536182
rect 73136 536170 73276 536172
rect 73136 536118 73222 536170
rect 73274 536118 73276 536170
rect 73136 536116 73276 536118
rect 73220 536106 73276 536116
rect 77252 536060 77308 536070
rect 72212 535836 72268 535846
rect 72212 535770 72268 535780
rect 73556 535836 73612 535846
rect 73556 535770 73612 535780
rect 72660 535612 72716 535622
rect 72660 535546 72716 535556
rect 73108 501676 73164 501686
rect 73108 501610 73164 501620
rect 73556 501564 73612 501574
rect 73556 501498 73612 501508
rect 72660 501452 72716 501462
rect 72660 501386 72716 501396
rect 72212 501340 72268 501350
rect 72212 501274 72268 501284
rect 72996 413196 73052 413206
rect 72688 413194 73052 413196
rect 72688 413142 72998 413194
rect 73050 413142 73052 413194
rect 72688 413140 73052 413142
rect 72996 413130 73052 413140
rect 73444 413084 73500 413094
rect 73136 413082 73500 413084
rect 73136 413030 73446 413082
rect 73498 413030 73500 413082
rect 73136 413028 73500 413030
rect 73444 413018 73500 413028
rect 72212 412748 72268 412758
rect 72212 412682 72268 412692
rect 73556 412636 73612 412646
rect 73556 412570 73612 412580
rect 76132 387996 76188 388006
rect 73780 377916 73836 377926
rect 72212 377580 72268 377888
rect 72688 377860 73052 377916
rect 72996 377804 73052 377860
rect 72996 377738 73052 377748
rect 73108 377692 73164 377888
rect 73584 377860 73780 377916
rect 73780 377850 73836 377860
rect 76132 377804 76188 387940
rect 76132 377738 76188 377748
rect 73108 377626 73164 377636
rect 72212 377514 72268 377524
rect 77252 377580 77308 536004
rect 77364 535948 77420 535958
rect 77364 387996 77420 535892
rect 77476 535834 77532 535846
rect 77476 535782 77478 535834
rect 77530 535782 77532 535834
rect 77476 399756 77532 535782
rect 77476 399690 77532 399700
rect 77588 535612 77644 535622
rect 77588 399644 77644 535556
rect 77812 501564 77868 576660
rect 77924 576604 77980 576614
rect 77924 501676 77980 576548
rect 77924 501610 77980 501620
rect 77812 501498 77868 501508
rect 77588 399578 77644 399588
rect 77700 412636 77756 412646
rect 77364 387930 77420 387940
rect 77252 377514 77308 377524
rect 72212 371980 72268 371990
rect 72212 371914 72268 371924
rect 73556 371868 73612 371878
rect 73556 371802 73612 371812
rect 72660 371756 72716 371766
rect 72660 371690 72716 371700
rect 73108 371644 73164 371654
rect 73108 371578 73164 371588
rect 77588 371644 77644 371654
rect 73108 337596 73164 337606
rect 73108 337530 73164 337540
rect 73556 337484 73612 337494
rect 73556 337418 73612 337428
rect 72212 337372 72268 337382
rect 72212 337306 72268 337316
rect 72660 337260 72716 337270
rect 72660 337194 72716 337204
rect 73220 331100 73276 331110
rect 73892 331100 73948 331110
rect 73136 331098 73276 331100
rect 73136 331046 73222 331098
rect 73274 331046 73276 331098
rect 73136 331044 73276 331046
rect 73584 331044 73892 331100
rect 73220 331034 73276 331044
rect 73892 331034 73948 331044
rect 77364 330988 77420 330998
rect 72212 330876 72268 330886
rect 72212 330810 72268 330820
rect 72660 330652 72716 330662
rect 72660 330586 72716 330596
rect 77252 314524 77308 314534
rect 77252 306570 77308 314468
rect 77252 306518 77254 306570
rect 77306 306518 77308 306570
rect 77252 306506 77308 306518
rect 73108 296604 73164 296614
rect 73108 296538 73164 296548
rect 73556 296492 73612 296502
rect 73556 296426 73612 296436
rect 72212 296380 72268 296390
rect 72212 296314 72268 296324
rect 72660 296268 72716 296278
rect 72660 296202 72716 296212
rect 72772 290108 72828 290118
rect 72688 290052 72772 290108
rect 72772 290042 72828 290052
rect 72212 289884 72268 289894
rect 72212 289818 72268 289828
rect 73556 289772 73612 289782
rect 73556 289706 73612 289716
rect 73108 289660 73164 289670
rect 73108 289594 73164 289604
rect 73108 255276 73164 255286
rect 73108 255210 73164 255220
rect 73556 255164 73612 255174
rect 73556 255098 73612 255108
rect 72548 255052 72604 255062
rect 72240 254996 72548 255052
rect 72548 254986 72604 254996
rect 77364 255052 77420 330932
rect 77476 330652 77532 330662
rect 77476 255164 77532 330596
rect 77588 296604 77644 371588
rect 77700 337260 77756 412580
rect 77924 371980 77980 371990
rect 77700 337194 77756 337204
rect 77812 371756 77868 371766
rect 77588 296538 77644 296548
rect 77812 296492 77868 371700
rect 77812 296426 77868 296436
rect 77924 296380 77980 371924
rect 77924 296314 77980 296324
rect 78036 290108 78092 722372
rect 78148 706412 78204 781844
rect 78148 706346 78204 706356
rect 78260 738108 78316 738118
rect 78260 664860 78316 738052
rect 78372 706300 78428 782068
rect 78372 706234 78428 706244
rect 78260 664794 78316 664804
rect 78372 700140 78428 700150
rect 78260 659148 78316 659158
rect 78148 658924 78204 658934
rect 78148 603148 78204 658868
rect 78148 603082 78204 603092
rect 78260 582540 78316 659092
rect 78372 624316 78428 700084
rect 78372 624250 78428 624260
rect 78820 640108 78876 640118
rect 78260 582474 78316 582484
rect 78372 618042 78428 618054
rect 78372 617990 78374 618042
rect 78426 617990 78428 618042
rect 78148 576940 78204 576950
rect 78148 501340 78204 576884
rect 78372 562604 78428 617990
rect 78596 617708 78652 617718
rect 78372 562538 78428 562548
rect 78484 576828 78540 576838
rect 78484 501452 78540 576772
rect 78596 562492 78652 617652
rect 78596 562426 78652 562436
rect 78484 501386 78540 501396
rect 78708 557788 78764 557798
rect 78148 501274 78204 501284
rect 78260 413194 78316 413206
rect 78260 413142 78262 413194
rect 78314 413142 78316 413194
rect 78148 371868 78204 371878
rect 78148 296268 78204 371812
rect 78260 356412 78316 413142
rect 78260 356346 78316 356356
rect 78372 413082 78428 413094
rect 78372 413030 78374 413082
rect 78426 413030 78428 413082
rect 78372 356188 78428 413030
rect 78596 412748 78652 412758
rect 78596 356300 78652 412692
rect 78596 356234 78652 356244
rect 78372 356122 78428 356132
rect 78372 331100 78428 331110
rect 78148 296202 78204 296212
rect 78260 330874 78316 330886
rect 78260 330822 78262 330874
rect 78314 330822 78316 330874
rect 78036 290042 78092 290052
rect 77476 255098 77532 255108
rect 77700 289884 77756 289894
rect 77364 254986 77420 254996
rect 72996 254940 73052 254950
rect 72688 254884 72996 254940
rect 72996 254874 73052 254884
rect 73220 249116 73276 249126
rect 73136 249060 73220 249116
rect 73220 249050 73276 249060
rect 72212 248892 72268 248902
rect 72212 248826 72268 248836
rect 77588 248892 77644 248902
rect 73556 248780 73612 248790
rect 73556 248714 73612 248724
rect 77476 248780 77532 248790
rect 72660 248668 72716 248678
rect 72660 248602 72716 248612
rect 77364 248668 77420 248678
rect 73108 214620 73164 214630
rect 73108 214554 73164 214564
rect 73556 214508 73612 214518
rect 73556 214442 73612 214452
rect 72212 214396 72268 214406
rect 72212 214330 72268 214340
rect 72660 214284 72716 214294
rect 72660 214218 72716 214228
rect 73444 208124 73500 208134
rect 73136 208122 73500 208124
rect 73136 208070 73446 208122
rect 73498 208070 73500 208122
rect 73136 208068 73500 208070
rect 73444 208058 73500 208068
rect 72660 207900 72716 207910
rect 72660 207834 72716 207844
rect 73556 207788 73612 207798
rect 73556 207722 73612 207732
rect 72212 207676 72268 207686
rect 72212 207610 72268 207620
rect 73780 172956 73836 172966
rect 72688 172900 73052 172956
rect 73584 172900 73780 172956
rect 72996 172844 73052 172900
rect 73780 172890 73836 172900
rect 77364 172956 77420 248612
rect 77364 172890 77420 172900
rect 72212 172620 72268 172816
rect 77476 172844 77532 248724
rect 72996 172778 73052 172788
rect 73108 172732 73164 172816
rect 77476 172778 77532 172788
rect 73108 172666 73164 172676
rect 72212 172554 72268 172564
rect 77588 172620 77644 248836
rect 77700 214396 77756 289828
rect 78036 289884 78092 289894
rect 77924 289772 77980 289782
rect 77812 289660 77868 289670
rect 77812 214620 77868 289604
rect 77812 214554 77868 214564
rect 77700 214330 77756 214340
rect 77924 214284 77980 289716
rect 78036 214508 78092 289828
rect 78260 273980 78316 330822
rect 78260 273914 78316 273924
rect 78372 254940 78428 331044
rect 78708 289882 78764 557732
rect 78820 332554 78876 640052
rect 78820 332502 78822 332554
rect 78874 332502 78876 332554
rect 78820 332490 78876 332502
rect 79716 290332 79772 927332
rect 83972 912716 84028 929796
rect 83972 912650 84028 912660
rect 84084 910700 84140 935732
rect 84308 935788 84364 935798
rect 84308 910924 84364 935732
rect 84308 910858 84364 910868
rect 84532 935788 84588 935798
rect 84532 910812 84588 935732
rect 84532 910746 84588 910756
rect 84084 910634 84140 910644
rect 84756 910588 84812 936518
rect 85204 934668 85260 942788
rect 85428 942732 85484 942742
rect 85428 935452 85484 942676
rect 105812 942394 105868 945812
rect 105812 942342 105814 942394
rect 105866 942342 105868 942394
rect 105812 942330 105868 942342
rect 106260 942060 106316 945812
rect 106260 941994 106316 942004
rect 106372 942058 106428 946416
rect 141092 945868 141148 946416
rect 141092 945802 141148 945812
rect 106372 942006 106374 942058
rect 106426 942006 106428 942058
rect 106372 941994 106428 942006
rect 120932 943404 120988 943414
rect 120932 937354 120988 943348
rect 120932 937302 120934 937354
rect 120986 937302 120988 937354
rect 120932 937290 120988 937302
rect 124292 943404 124348 943414
rect 124292 936572 124348 943348
rect 141428 936684 141484 946836
rect 141428 936618 141484 936628
rect 124292 936506 124348 936516
rect 141540 936570 141596 947044
rect 141652 945868 141708 945878
rect 141652 936796 141708 945812
rect 141876 937020 141932 947044
rect 160244 942284 160300 947732
rect 160244 942218 160300 942228
rect 160356 947284 160832 947340
rect 196112 947284 196364 947340
rect 160356 942170 160412 947284
rect 160356 942118 160358 942170
rect 160410 942118 160412 942170
rect 160356 942106 160412 942118
rect 160580 946836 160832 946892
rect 160580 942172 160636 946836
rect 196084 946764 196140 946864
rect 196084 946698 196140 946708
rect 196308 946652 196364 947284
rect 196308 946586 196364 946596
rect 161140 942282 161196 946416
rect 196112 946388 196588 946444
rect 196308 946316 196364 946326
rect 177044 943516 177100 943526
rect 161140 942230 161142 942282
rect 161194 942230 161196 942282
rect 161140 942218 161196 942230
rect 176484 943404 176540 943414
rect 160580 942106 160636 942116
rect 141876 936954 141932 936964
rect 163716 938588 163772 938598
rect 141652 936730 141708 936740
rect 141540 936518 141542 936570
rect 141594 936518 141596 936570
rect 141540 936506 141596 936518
rect 85428 935386 85484 935396
rect 96964 935676 97020 935686
rect 96964 935088 97020 935620
rect 141316 935452 141372 935462
rect 141316 935088 141372 935396
rect 163716 935088 163772 938532
rect 176484 935450 176540 943348
rect 177044 938250 177100 943460
rect 178164 943516 178220 943526
rect 177044 938198 177046 938250
rect 177098 938198 177100 938250
rect 177044 938186 177100 938198
rect 178052 943404 178108 943414
rect 176708 937468 176764 937478
rect 176708 935674 176764 937412
rect 178052 937020 178108 943348
rect 178164 938588 178220 943460
rect 178164 938522 178220 938532
rect 179732 943404 179788 943414
rect 179732 937468 179788 943348
rect 196308 942058 196364 946260
rect 196532 942394 196588 946388
rect 196532 942342 196534 942394
rect 196586 942342 196588 942394
rect 196532 942330 196588 942342
rect 196644 942396 196700 947732
rect 251076 947660 251132 947760
rect 271562 947732 271572 947788
rect 271628 947732 271638 947788
rect 251076 947594 251132 947604
rect 306068 947660 306124 947760
rect 306068 947594 306124 947604
rect 361060 947548 361116 947760
rect 470250 947732 470260 947788
rect 470316 947732 470326 947788
rect 490868 947760 490924 949172
rect 525690 947732 525700 947788
rect 525756 947732 525766 947788
rect 361060 947482 361116 947492
rect 545860 947548 545916 947760
rect 545860 947482 545916 947492
rect 581140 947548 581196 947760
rect 581140 947482 581196 947492
rect 655844 947548 655900 947760
rect 690330 947732 690340 947788
rect 690396 947732 690406 947788
rect 655844 947482 655900 947492
rect 697956 947548 698012 947558
rect 196644 942330 196700 942340
rect 215572 947284 215824 947340
rect 251104 947284 251356 947340
rect 196308 942006 196310 942058
rect 196362 942006 196364 942058
rect 196308 941994 196364 942006
rect 215572 942058 215628 947284
rect 215572 942006 215574 942058
rect 215626 942006 215628 942058
rect 215572 941994 215628 942006
rect 215684 946836 215824 946892
rect 215684 942060 215740 946836
rect 251076 946764 251132 946864
rect 251076 946698 251132 946708
rect 216356 942394 216412 946416
rect 216356 942342 216358 942394
rect 216410 942342 216412 942394
rect 216356 942330 216412 942342
rect 230132 943516 230188 943526
rect 215684 941994 215740 942004
rect 179732 937402 179788 937412
rect 178052 936954 178108 936964
rect 230132 936684 230188 943460
rect 233492 943516 233548 943526
rect 231812 943404 231868 943414
rect 230132 936618 230188 936628
rect 230356 937468 230412 937478
rect 176708 935622 176710 935674
rect 176762 935622 176764 935674
rect 176708 935610 176764 935622
rect 185780 935674 185836 935686
rect 185780 935622 185782 935674
rect 185834 935622 185836 935674
rect 176484 935398 176486 935450
rect 176538 935398 176540 935450
rect 176484 935386 176540 935398
rect 185780 935088 185836 935622
rect 208068 935450 208124 935462
rect 208068 935398 208070 935450
rect 208122 935398 208124 935450
rect 208068 935088 208124 935398
rect 230356 935088 230412 937412
rect 231812 935004 231868 943348
rect 233492 937468 233548 943460
rect 233492 937402 233548 937412
rect 233828 943404 233884 943414
rect 233828 936570 233884 943348
rect 251076 942170 251132 946416
rect 251300 942282 251356 947284
rect 251300 942230 251302 942282
rect 251354 942230 251356 942282
rect 251300 942218 251356 942230
rect 270452 947284 270816 947340
rect 306096 947284 306572 947340
rect 270452 942282 270508 947284
rect 270452 942230 270454 942282
rect 270506 942230 270508 942282
rect 270452 942218 270508 942230
rect 270564 946836 270816 946892
rect 306096 946836 306460 946892
rect 251076 942118 251078 942170
rect 251130 942118 251132 942170
rect 251076 942106 251132 942118
rect 270564 942172 270620 946836
rect 270564 942106 270620 942116
rect 271348 942170 271404 946416
rect 271348 942118 271350 942170
rect 271402 942118 271404 942170
rect 271348 942106 271404 942118
rect 285684 943404 285740 943414
rect 233828 936518 233830 936570
rect 233882 936518 233884 936570
rect 233828 936506 233884 936518
rect 282436 937468 282492 937478
rect 251972 935228 252028 935238
rect 251972 935116 252028 935172
rect 251972 935060 252560 935116
rect 282436 935114 282492 937412
rect 285684 937132 285740 943348
rect 289156 943404 289212 943414
rect 285684 937066 285740 937076
rect 285908 943292 285964 943302
rect 282436 935062 282438 935114
rect 282490 935062 282492 935114
rect 282436 935050 282492 935062
rect 285908 935116 285964 943236
rect 289156 935226 289212 943348
rect 289380 943404 289436 943414
rect 289380 936796 289436 943348
rect 306068 942058 306124 946416
rect 306068 942006 306070 942058
rect 306122 942006 306124 942058
rect 306068 941994 306124 942006
rect 306404 942060 306460 946836
rect 306516 942394 306572 947284
rect 361060 947212 361116 947312
rect 471184 947284 471884 947340
rect 361060 947146 361116 947156
rect 471268 946892 471324 946902
rect 361060 946764 361116 946864
rect 471184 946836 471268 946892
rect 471268 946826 471324 946836
rect 361060 946698 361116 946708
rect 361171 946428 361227 946444
rect 361171 946372 361228 946428
rect 471184 946388 471772 946444
rect 344596 943516 344652 943526
rect 306516 942342 306518 942394
rect 306570 942342 306572 942394
rect 306516 942330 306572 942342
rect 341124 943292 341180 943302
rect 335860 942172 335916 942182
rect 335860 942078 335916 942116
rect 306404 941994 306460 942004
rect 289380 936730 289436 936740
rect 341012 937466 341068 937478
rect 341012 937414 341014 937466
rect 341066 937414 341068 937466
rect 341012 935338 341068 937414
rect 341124 936124 341180 943236
rect 344596 937466 344652 943460
rect 344596 937414 344598 937466
rect 344650 937414 344652 937466
rect 344596 937402 344652 937414
rect 344708 943404 344764 943414
rect 344708 936682 344764 943348
rect 361172 942282 361228 946372
rect 471716 945868 471772 946388
rect 471828 946092 471884 947284
rect 471828 946026 471884 946036
rect 490532 947284 490896 947340
rect 525578 947284 525588 947340
rect 525644 947284 525654 947340
rect 471716 945802 471772 945812
rect 490532 945868 490588 947284
rect 545860 947100 545916 947312
rect 581168 947284 581308 947340
rect 581252 947212 581308 947284
rect 581252 947146 581308 947156
rect 545860 947034 545916 947044
rect 655844 947100 655900 947312
rect 690330 947284 690340 947340
rect 690396 947284 690406 947340
rect 655844 947034 655900 947044
rect 545636 946892 545692 946902
rect 655620 946892 655676 946902
rect 490644 946836 490896 946892
rect 490644 945980 490700 946836
rect 526148 946764 526204 946864
rect 545692 946836 545888 946892
rect 545636 946826 545692 946836
rect 526148 946698 526204 946708
rect 581028 946764 581084 946864
rect 655676 946836 655872 946892
rect 691152 946876 691852 946892
rect 691152 946836 691796 946876
rect 655620 946826 655676 946836
rect 691796 946810 691852 946820
rect 581028 946698 581084 946708
rect 545524 946444 545580 946454
rect 655508 946444 655564 946454
rect 490868 946092 490924 946416
rect 525690 946388 525700 946444
rect 525756 946388 525766 946444
rect 545580 946388 545888 946444
rect 545524 946378 545580 946388
rect 581140 946316 581196 946416
rect 655564 946388 655872 946444
rect 655508 946378 655564 946388
rect 581140 946250 581196 946260
rect 490868 946026 490924 946036
rect 490644 945914 490700 945924
rect 490532 945802 490588 945812
rect 691124 945868 691180 946416
rect 691124 945802 691180 945812
rect 507444 943516 507500 943526
rect 361172 942230 361174 942282
rect 361226 942230 361228 942282
rect 361172 942218 361228 942230
rect 450212 943404 450268 943414
rect 450212 936794 450268 943348
rect 451892 943404 451948 943414
rect 451892 936908 451948 943348
rect 451892 936842 451948 936852
rect 453572 943404 453628 943414
rect 453572 936906 453628 943348
rect 455028 943404 455084 943414
rect 455028 938252 455084 943348
rect 505652 943404 505708 943414
rect 455028 938186 455084 938196
rect 458500 938252 458556 938262
rect 453572 936854 453574 936906
rect 453626 936854 453628 936906
rect 453572 936842 453628 936854
rect 450212 936742 450214 936794
rect 450266 936742 450268 936794
rect 450212 936730 450268 936742
rect 344708 936630 344710 936682
rect 344762 936630 344764 936682
rect 344708 936618 344764 936630
rect 341124 936058 341180 936068
rect 342580 936124 342636 936134
rect 341012 935286 341014 935338
rect 341066 935286 341068 935338
rect 341012 935274 341068 935286
rect 289156 935174 289158 935226
rect 289210 935174 289212 935226
rect 289156 935162 289212 935174
rect 296324 935226 296380 935238
rect 296324 935174 296326 935226
rect 296378 935174 296380 935226
rect 296324 935116 296380 935174
rect 318948 935116 319004 935126
rect 341012 935116 341068 935126
rect 296324 935060 297024 935116
rect 318948 935114 319200 935116
rect 318948 935062 318950 935114
rect 319002 935062 319200 935114
rect 318948 935060 319200 935062
rect 341068 935060 341376 935116
rect 285908 935050 285964 935060
rect 318948 935050 319004 935060
rect 341012 935050 341068 935060
rect 231812 934938 231868 934948
rect 274036 935004 274092 935014
rect 274092 934948 274736 935004
rect 274036 934938 274092 934948
rect 342580 934890 342636 936068
rect 385252 935004 385308 935014
rect 385252 935002 385840 935004
rect 385252 934950 385254 935002
rect 385306 934950 385840 935002
rect 385252 934948 385840 934950
rect 385252 934938 385308 934948
rect 342580 934838 342582 934890
rect 342634 934838 342636 934890
rect 342580 934826 342636 934838
rect 362964 934892 363020 934902
rect 407428 934892 407484 934902
rect 430948 934892 431004 934902
rect 453348 934892 453404 934902
rect 363020 934836 363664 934892
rect 407428 934890 408128 934892
rect 407428 934838 407430 934890
rect 407482 934838 408128 934890
rect 407428 934836 408128 934838
rect 430416 934836 430948 934892
rect 452704 934890 453404 934892
rect 452704 934838 453350 934890
rect 453402 934838 453404 934890
rect 452704 934836 453404 934838
rect 362964 934826 363020 934836
rect 407428 934826 407484 934836
rect 430948 934826 431004 934836
rect 453348 934826 453404 934836
rect 458500 934890 458556 938196
rect 505652 937018 505708 943348
rect 505652 936966 505654 937018
rect 505706 936966 505708 937018
rect 505652 936954 505708 936966
rect 505876 943292 505932 943302
rect 505876 937020 505932 943236
rect 505876 936954 505932 936964
rect 474740 936908 474796 936918
rect 474740 935088 474796 936852
rect 497364 935004 497420 935014
rect 497168 935002 497420 935004
rect 497168 934950 497366 935002
rect 497418 934950 497420 935002
rect 497168 934948 497420 934950
rect 497364 934938 497420 934948
rect 507444 935002 507500 943460
rect 509012 943404 509068 943414
rect 509012 937132 509068 943348
rect 510580 943404 510636 943414
rect 510580 938476 510636 943348
rect 564228 943404 564284 943414
rect 561092 943292 561148 943302
rect 510580 938410 510636 938420
rect 519204 938476 519260 938486
rect 509012 937066 509068 937076
rect 519204 935088 519260 938420
rect 561092 937244 561148 943236
rect 561092 937178 561148 937188
rect 541380 937020 541436 937030
rect 541380 935088 541436 936964
rect 564228 935116 564284 943348
rect 673428 943404 673484 943414
rect 673428 939148 673484 943348
rect 674100 943404 674156 943414
rect 673428 939082 673484 939092
rect 673652 943292 673708 943302
rect 673652 937356 673708 943236
rect 673652 937290 673708 937300
rect 673876 943180 673932 943190
rect 608132 937244 608188 937254
rect 563808 935060 564284 935116
rect 585956 935676 586012 935686
rect 585956 935088 586012 935620
rect 608132 935088 608188 937188
rect 652708 935564 652764 935574
rect 630420 935450 630476 935462
rect 630420 935398 630422 935450
rect 630474 935398 630476 935450
rect 630420 935088 630476 935398
rect 652708 935088 652764 935508
rect 673876 935564 673932 943124
rect 673876 935498 673932 935508
rect 674100 935450 674156 943348
rect 674100 935398 674102 935450
rect 674154 935398 674156 935450
rect 674100 935386 674156 935398
rect 674772 939148 674828 939158
rect 674772 935088 674828 939092
rect 687764 938250 687820 938262
rect 687764 938198 687766 938250
rect 687818 938198 687820 938250
rect 687428 937244 687484 937254
rect 687204 937132 687260 937142
rect 686980 935340 687036 935350
rect 686644 935116 686700 935126
rect 507444 934950 507446 935002
rect 507498 934950 507500 935002
rect 507444 934938 507500 934950
rect 686532 935004 686588 935014
rect 458500 934838 458502 934890
rect 458554 934838 458556 934890
rect 458500 934826 458556 934838
rect 686308 934780 686364 934790
rect 85204 934602 85260 934612
rect 118468 934668 118524 934678
rect 118524 934612 119168 934668
rect 118468 934602 118524 934612
rect 84756 910522 84812 910532
rect 686196 934556 686252 934566
rect 83972 884044 84028 884054
rect 83076 783692 83132 783702
rect 80500 763196 80556 763206
rect 80388 600684 80444 600694
rect 80276 518924 80332 518934
rect 80052 396172 80108 396182
rect 80052 331770 80108 396116
rect 80052 331718 80054 331770
rect 80106 331718 80108 331770
rect 80052 331706 80108 331718
rect 80164 354172 80220 354182
rect 79716 290266 79772 290276
rect 78708 289830 78710 289882
rect 78762 289830 78764 289882
rect 78708 289818 78764 289830
rect 80164 289770 80220 354116
rect 80276 331772 80332 518868
rect 80276 331706 80332 331716
rect 80388 289994 80444 600628
rect 80500 331884 80556 763140
rect 80500 331818 80556 331828
rect 80388 289942 80390 289994
rect 80442 289942 80444 289994
rect 80388 289930 80444 289942
rect 83076 289884 83132 783636
rect 83188 762860 83244 762870
rect 83188 302428 83244 762804
rect 83972 762860 84028 883988
rect 84308 869820 84364 869830
rect 83972 762794 84028 762804
rect 84084 841260 84140 841270
rect 84084 720748 84140 841204
rect 84084 720682 84140 720692
rect 84196 798364 84252 798374
rect 83972 712684 84028 712694
rect 83188 302362 83244 302372
rect 83300 701372 83356 701382
rect 83300 299850 83356 701316
rect 83860 682220 83916 682230
rect 83748 557788 83804 557798
rect 83412 415772 83468 415782
rect 83412 306572 83468 415716
rect 83636 393484 83692 393494
rect 83636 306682 83692 393428
rect 83748 306794 83804 557732
rect 83748 306742 83750 306794
rect 83802 306742 83804 306794
rect 83748 306730 83804 306742
rect 83636 306630 83638 306682
rect 83690 306630 83692 306682
rect 83636 306618 83692 306630
rect 83412 306506 83468 306516
rect 83300 299798 83302 299850
rect 83354 299798 83356 299850
rect 83300 299786 83356 299798
rect 83076 289818 83132 289828
rect 80164 289718 80166 289770
rect 80218 289718 80220 289770
rect 80164 289706 80220 289718
rect 83860 289772 83916 682164
rect 83972 598556 84028 712628
rect 84196 681212 84252 798308
rect 84308 766108 84364 869764
rect 84644 855484 84700 855494
rect 84308 766042 84364 766052
rect 84420 826924 84476 826934
rect 84196 681146 84252 681156
rect 84308 741244 84364 741254
rect 83972 598490 84028 598500
rect 84084 669788 84140 669798
rect 83972 584108 84028 584118
rect 83972 393708 84028 584052
rect 84084 557900 84140 669732
rect 84308 642348 84364 741188
rect 84420 725116 84476 826868
rect 84420 725050 84476 725060
rect 84532 784028 84588 784038
rect 84308 642282 84364 642292
rect 84420 698348 84476 698358
rect 84084 557834 84140 557844
rect 84196 626892 84252 626902
rect 84196 516460 84252 626836
rect 84420 602028 84476 698292
rect 84532 684348 84588 783972
rect 84644 764540 84700 855428
rect 686196 848204 686252 934500
rect 686196 848138 686252 848148
rect 84644 764474 84700 764484
rect 84756 812700 84812 812710
rect 84532 684282 84588 684292
rect 84644 726908 84700 726918
rect 84420 601962 84476 601972
rect 84532 655564 84588 655574
rect 84196 516394 84252 516404
rect 84308 569772 84364 569782
rect 83972 393642 84028 393652
rect 84084 498428 84140 498438
rect 84084 311500 84140 498372
rect 84084 311434 84140 311444
rect 84196 455532 84252 455542
rect 83860 289706 83916 289716
rect 78708 289658 78764 289670
rect 78708 289606 78710 289658
rect 78762 289606 78764 289658
rect 78484 283052 78540 283062
rect 78484 273868 78540 282996
rect 78708 274092 78764 289606
rect 78708 274026 78764 274036
rect 78820 283164 78876 283174
rect 78484 273802 78540 273812
rect 78372 254874 78428 254884
rect 78036 214442 78092 214452
rect 78148 249116 78204 249126
rect 77924 214218 77980 214228
rect 77588 172554 77644 172564
rect 78036 207788 78092 207798
rect 78036 82122 78092 207732
rect 78148 172732 78204 249060
rect 78820 233548 78876 283108
rect 84196 270844 84252 455476
rect 84308 396956 84364 569716
rect 84532 561820 84588 655508
rect 84644 642124 84700 726852
rect 84756 722652 84812 812644
rect 686196 793548 686252 793558
rect 84756 722586 84812 722596
rect 84868 769804 84924 769814
rect 84868 682332 84924 769748
rect 84868 682266 84924 682276
rect 84980 683788 85036 683798
rect 84644 642058 84700 642068
rect 84532 561754 84588 561764
rect 84644 641228 84700 641238
rect 84644 559468 84700 641172
rect 84868 619052 84924 619062
rect 84644 559402 84700 559412
rect 84756 612668 84812 612678
rect 84644 555548 84700 555558
rect 84308 396890 84364 396900
rect 84420 526988 84476 526998
rect 84420 356972 84476 526932
rect 84420 356906 84476 356916
rect 84532 484092 84588 484102
rect 84196 270778 84252 270788
rect 84308 341292 84364 341302
rect 78820 233482 78876 233492
rect 78148 172666 78204 172676
rect 78260 208122 78316 208134
rect 78260 208070 78262 208122
rect 78314 208070 78316 208122
rect 78036 82070 78038 82122
rect 78090 82070 78092 82122
rect 78036 82058 78092 82070
rect 78260 81002 78316 208070
rect 84308 190988 84364 341236
rect 84532 314412 84588 484036
rect 84644 395052 84700 555492
rect 84756 519148 84812 612612
rect 84756 519082 84812 519092
rect 84644 394986 84700 394996
rect 84756 512652 84812 512662
rect 84532 314346 84588 314356
rect 84644 384076 84700 384086
rect 84644 232092 84700 384020
rect 84756 355068 84812 512596
rect 84756 355002 84812 355012
rect 84868 306796 84924 618996
rect 84980 599788 85036 683732
rect 84980 599722 85036 599732
rect 84980 598108 85036 598118
rect 84980 517916 85036 598052
rect 84980 517850 85036 517860
rect 84980 469196 85036 469206
rect 84980 312508 85036 469140
rect 84980 312442 85036 312452
rect 85092 426748 85148 426758
rect 84868 306730 84924 306740
rect 84756 305788 84812 305798
rect 84756 305694 84812 305732
rect 85092 272188 85148 426692
rect 85092 272122 85148 272132
rect 85204 398188 85260 398198
rect 84644 232026 84700 232036
rect 85204 231868 85260 398132
rect 686196 334124 686252 793492
rect 686308 661500 686364 934724
rect 686420 740684 686476 740694
rect 686420 671132 686476 740628
rect 686532 688156 686588 934948
rect 686644 767788 686700 935060
rect 686756 934668 686812 934678
rect 686756 914732 686812 934612
rect 686868 934220 686924 934230
rect 686868 928060 686924 934164
rect 686868 927994 686924 928004
rect 686756 914666 686812 914676
rect 686644 767722 686700 767732
rect 686980 754012 687036 935284
rect 686980 753946 687036 753956
rect 686532 688090 686588 688100
rect 686420 671066 686476 671076
rect 686308 661434 686364 661444
rect 686532 606844 686588 606854
rect 686532 488236 686588 606788
rect 686532 488170 686588 488180
rect 686644 593516 686700 593526
rect 686420 446908 686476 446918
rect 686196 334058 686252 334068
rect 686308 366940 686364 366950
rect 222852 333788 222908 333798
rect 119140 333676 119196 333686
rect 118608 333620 119140 333676
rect 119140 333610 119196 333620
rect 171108 333676 171164 333686
rect 160692 333564 160748 333574
rect 160384 333508 160692 333564
rect 160692 333498 160748 333508
rect 127204 333452 127260 333462
rect 126560 333396 127204 333452
rect 127204 333386 127260 333396
rect 162820 333340 162876 333350
rect 86884 332666 86940 333312
rect 88788 332892 88844 333312
rect 88788 332826 88844 332836
rect 90804 332778 90860 333312
rect 90804 332726 90806 332778
rect 90858 332726 90860 332778
rect 90804 332714 90860 332726
rect 86884 332614 86886 332666
rect 86938 332614 86940 332666
rect 86884 332602 86940 332614
rect 92820 332668 92876 333312
rect 92820 332602 92876 332612
rect 94052 333284 94640 333340
rect 95732 333284 96656 333340
rect 94052 323930 94108 333284
rect 95732 324154 95788 333284
rect 98756 332780 98812 333312
rect 100660 333004 100716 333312
rect 100660 332938 100716 332948
rect 102676 333002 102732 333312
rect 102676 332950 102678 333002
rect 102730 332950 102732 333002
rect 102676 332938 102732 332950
rect 104132 333284 104608 333340
rect 98756 332714 98812 332724
rect 95732 324102 95734 324154
rect 95786 324102 95788 324154
rect 95732 324090 95788 324102
rect 104132 324156 104188 333284
rect 106708 333116 106764 333312
rect 106708 333050 106764 333060
rect 108724 330092 108780 333312
rect 110628 332890 110684 333312
rect 110628 332838 110630 332890
rect 110682 332838 110684 332890
rect 110628 332826 110684 332838
rect 108724 330026 108780 330036
rect 112644 328412 112700 333312
rect 112644 328346 112700 328356
rect 114660 328076 114716 333312
rect 116676 328636 116732 333312
rect 116676 328570 116732 328580
rect 120596 328522 120652 333312
rect 120596 328470 120598 328522
rect 120650 328470 120652 328522
rect 120596 328458 120652 328470
rect 122500 328410 122556 333312
rect 124628 328634 124684 333312
rect 128548 328858 128604 333312
rect 128548 328806 128550 328858
rect 128602 328806 128604 328858
rect 128548 328794 128604 328806
rect 130564 328748 130620 333312
rect 132580 333114 132636 333312
rect 132580 333062 132582 333114
rect 132634 333062 132636 333114
rect 132580 333050 132636 333062
rect 130564 328682 130620 328692
rect 133476 333004 133532 333014
rect 124628 328582 124630 328634
rect 124682 328582 124684 328634
rect 124628 328570 124684 328582
rect 122500 328358 122502 328410
rect 122554 328358 122556 328410
rect 122500 328346 122556 328358
rect 114660 328010 114716 328020
rect 104132 324090 104188 324100
rect 94052 323878 94054 323930
rect 94106 323878 94108 323930
rect 94052 323866 94108 323878
rect 133476 323932 133532 332948
rect 133924 332892 133980 332902
rect 133700 332780 133756 332790
rect 133700 324042 133756 332724
rect 133700 323990 133702 324042
rect 133754 323990 133756 324042
rect 133700 323978 133756 323990
rect 133476 323866 133532 323876
rect 133924 322588 133980 332836
rect 134484 332892 134540 333312
rect 134484 332826 134540 332836
rect 135156 333116 135212 333126
rect 135156 324044 135212 333060
rect 136500 328860 136556 333312
rect 138544 333284 139244 333340
rect 139188 333226 139244 333284
rect 139188 333174 139190 333226
rect 139242 333174 139244 333226
rect 139188 333162 139244 333174
rect 140532 333004 140588 333312
rect 140532 332938 140588 332948
rect 142436 328972 142492 333312
rect 144340 332108 144396 333312
rect 146468 333116 146524 333312
rect 148400 333284 149100 333340
rect 149044 333228 149100 333284
rect 149044 333162 149100 333172
rect 146468 333050 146524 333060
rect 144340 332042 144396 332052
rect 150388 329084 150444 333312
rect 151956 333002 152012 333014
rect 151956 332950 151958 333002
rect 152010 332950 152012 333002
rect 150388 329018 150444 329028
rect 150612 332778 150668 332790
rect 150612 332726 150614 332778
rect 150666 332726 150668 332778
rect 142436 328906 142492 328916
rect 136500 328794 136556 328804
rect 135156 323978 135212 323988
rect 149492 324044 149548 324054
rect 149492 323820 149548 323988
rect 150612 323932 150668 332726
rect 150612 323866 150668 323876
rect 149492 323754 149548 323764
rect 151956 323820 152012 332950
rect 152404 332778 152460 333312
rect 154420 333002 154476 333312
rect 154420 332950 154422 333002
rect 154474 332950 154476 333002
rect 154420 332938 154476 332950
rect 152404 332726 152406 332778
rect 152458 332726 152460 332778
rect 152404 332714 152460 332726
rect 156324 329196 156380 333312
rect 156324 329130 156380 329140
rect 157892 333284 158256 333340
rect 162400 333284 162820 333340
rect 157892 325052 157948 333284
rect 162820 333274 162876 333284
rect 162932 333284 164192 333340
rect 157892 324986 157948 324996
rect 160244 332666 160300 332678
rect 160244 332614 160246 332666
rect 160298 332614 160300 332666
rect 160244 324380 160300 332614
rect 162932 325164 162988 333284
rect 166180 328300 166236 333312
rect 166180 328234 166236 328244
rect 167972 332890 168028 332902
rect 167972 332838 167974 332890
rect 168026 332838 168028 332890
rect 162932 325098 162988 325108
rect 161700 324380 161756 324390
rect 160244 324324 160356 324380
rect 159908 324268 159964 324278
rect 151956 323754 152012 323764
rect 155204 324154 155260 324166
rect 155204 324102 155206 324154
rect 155258 324102 155260 324154
rect 155204 323818 155260 324102
rect 155428 324154 155484 324166
rect 155428 324102 155430 324154
rect 155482 324102 155484 324154
rect 155316 323932 155372 323942
rect 155428 323932 155484 324102
rect 155316 323930 155484 323932
rect 155316 323878 155318 323930
rect 155370 323878 155484 323930
rect 155316 323876 155484 323878
rect 159572 323932 159628 323942
rect 155316 323866 155372 323876
rect 155204 323766 155206 323818
rect 155258 323766 155260 323818
rect 155204 323754 155260 323766
rect 133924 322522 133980 322532
rect 159572 322588 159628 323876
rect 159908 323820 159964 324212
rect 159908 323754 159964 323764
rect 160300 323680 160356 324324
rect 161364 324266 161420 324278
rect 161364 324214 161366 324266
rect 161418 324214 161420 324266
rect 161028 324156 161084 324166
rect 161084 324100 161196 324156
rect 161028 324090 161084 324100
rect 160972 323932 161028 323942
rect 160972 323680 161028 323876
rect 161140 323932 161196 324100
rect 161364 324044 161420 324214
rect 161700 324156 161756 324324
rect 162596 324266 162652 324278
rect 162596 324214 162598 324266
rect 162650 324214 162652 324266
rect 161700 324100 161812 324156
rect 161364 323978 161420 323988
rect 161140 323866 161196 323876
rect 161756 323680 161812 324100
rect 162428 323932 162484 323942
rect 162428 323680 162484 323876
rect 162596 323932 162652 324214
rect 162596 323866 162652 323876
rect 163212 324154 163268 324166
rect 163212 324102 163214 324154
rect 163266 324102 163268 324154
rect 163212 323680 163268 324102
rect 165340 324156 165396 324166
rect 164668 324042 164724 324054
rect 164668 323990 164670 324042
rect 164722 323990 164724 324042
rect 163884 323930 163940 323942
rect 163884 323878 163886 323930
rect 163938 323878 163940 323930
rect 163884 323680 163940 323878
rect 164668 323680 164724 323990
rect 165340 323680 165396 324100
rect 166796 324156 166852 324166
rect 166124 324044 166180 324054
rect 166124 323680 166180 323988
rect 166796 323680 166852 324100
rect 167972 324044 168028 332838
rect 168084 330092 168140 330102
rect 168084 325947 168140 330036
rect 168308 328188 168364 333312
rect 170324 328524 170380 333312
rect 170324 328458 170380 328468
rect 168308 328122 168364 328132
rect 170436 328076 170492 328086
rect 168084 325891 169036 325947
rect 168980 324380 169036 325891
rect 170436 324380 170492 328020
rect 171108 324380 171164 333620
rect 209636 333676 209692 333686
rect 187124 333564 187180 333574
rect 173460 333452 173516 333462
rect 174580 333452 174636 333462
rect 174272 333396 174580 333452
rect 171892 328636 171948 328646
rect 171892 324380 171948 328580
rect 172228 328412 172284 333312
rect 173460 333116 173516 333396
rect 174580 333386 174636 333396
rect 173460 333050 173516 333060
rect 174020 333116 174076 333126
rect 172228 328346 172284 328356
rect 172564 328522 172620 328534
rect 172564 328470 172566 328522
rect 172618 328470 172620 328522
rect 172564 324380 172620 328470
rect 173348 328410 173404 328422
rect 173348 328358 173350 328410
rect 173402 328358 173404 328410
rect 173348 324380 173404 328358
rect 174020 324380 174076 333060
rect 176260 332668 176316 333312
rect 177716 333114 177772 333126
rect 177716 333062 177718 333114
rect 177770 333062 177772 333114
rect 176260 332602 176316 332612
rect 176932 332892 176988 332902
rect 175476 328858 175532 328870
rect 175476 328806 175478 328858
rect 175530 328806 175532 328858
rect 174804 328634 174860 328646
rect 174804 328582 174806 328634
rect 174858 328582 174860 328634
rect 174804 324380 174860 328582
rect 175476 324380 175532 328806
rect 176260 328748 176316 328758
rect 176260 324380 176316 328692
rect 176932 324380 176988 332836
rect 177716 324380 177772 333062
rect 178276 333004 178332 333312
rect 178276 332938 178332 332948
rect 179844 333226 179900 333238
rect 179844 333174 179846 333226
rect 179898 333174 179900 333226
rect 179172 332892 179228 332902
rect 178388 328860 178444 328870
rect 178388 324380 178444 328804
rect 179172 324380 179228 332836
rect 179844 324380 179900 333174
rect 180180 332780 180236 333312
rect 180180 332714 180236 332724
rect 181300 333228 181356 333238
rect 180628 328972 180684 328982
rect 180628 324380 180684 328916
rect 181300 324380 181356 333172
rect 182196 333116 182252 333312
rect 184240 333284 184492 333340
rect 184436 333228 184492 333284
rect 184436 333162 184492 333172
rect 184884 333284 186144 333340
rect 182196 333050 182252 333060
rect 182756 332892 182812 332902
rect 181636 332108 181692 332118
rect 181636 325947 181692 332052
rect 181636 325891 182140 325947
rect 182084 324380 182140 325891
rect 182756 324380 182812 332836
rect 183540 332778 183596 332790
rect 183540 332726 183542 332778
rect 183594 332726 183596 332778
rect 183540 324380 183596 332726
rect 184212 329084 184268 329094
rect 184212 324380 184268 329028
rect 168980 324324 169092 324380
rect 170436 324324 170548 324380
rect 171108 324324 171220 324380
rect 171892 324324 172004 324380
rect 172564 324324 172676 324380
rect 173348 324324 173460 324380
rect 174020 324324 174132 324380
rect 174804 324324 174916 324380
rect 175476 324324 175588 324380
rect 176260 324324 176372 324380
rect 176932 324324 177044 324380
rect 177716 324324 177828 324380
rect 178388 324324 178500 324380
rect 179172 324324 179284 324380
rect 179844 324324 179956 324380
rect 180628 324324 180740 324380
rect 181300 324324 181412 324380
rect 182084 324324 182196 324380
rect 182756 324324 182868 324380
rect 183540 324324 183652 324380
rect 184212 324324 184324 324380
rect 167972 323988 168308 324044
rect 167580 323932 167636 323942
rect 167580 323680 167636 323876
rect 168252 323680 168308 323988
rect 169036 323680 169092 324324
rect 169708 324156 169764 324166
rect 169708 323680 169764 324100
rect 170492 323680 170548 324324
rect 171164 323680 171220 324324
rect 171948 323680 172004 324324
rect 172620 323680 172676 324324
rect 173404 323680 173460 324324
rect 174076 323680 174132 324324
rect 174860 323680 174916 324324
rect 175532 323680 175588 324324
rect 176316 323680 176372 324324
rect 176988 323680 177044 324324
rect 177772 323680 177828 324324
rect 178444 323680 178500 324324
rect 179228 323680 179284 324324
rect 179900 323680 179956 324324
rect 180684 323680 180740 324324
rect 181356 323680 181412 324324
rect 182140 323680 182196 324324
rect 182812 323680 182868 324324
rect 183596 323680 183652 324324
rect 184268 323680 184324 324324
rect 184884 323932 184940 333284
rect 184996 333002 185052 333014
rect 184996 332950 184998 333002
rect 185050 332950 185052 333002
rect 184996 324380 185052 332950
rect 185668 325052 185724 325062
rect 185668 324380 185724 324996
rect 187124 324380 187180 333508
rect 188020 332890 188076 333312
rect 188020 332838 188022 332890
rect 188074 332838 188076 332890
rect 188020 332826 188076 332838
rect 188580 333228 188636 333238
rect 187908 325164 187964 325174
rect 187908 324380 187964 325108
rect 188580 324380 188636 333172
rect 190148 332778 190204 333312
rect 190148 332726 190150 332778
rect 190202 332726 190204 332778
rect 190148 332714 190204 332726
rect 192164 332666 192220 333312
rect 193732 333004 193788 333014
rect 192164 332614 192166 332666
rect 192218 332614 192220 332666
rect 192164 332602 192220 332614
rect 192276 332668 192332 332678
rect 190036 328524 190092 328534
rect 189364 328300 189420 328310
rect 189364 324380 189420 328244
rect 190036 324380 190092 328468
rect 191492 328412 191548 328422
rect 190820 328188 190876 328198
rect 190820 324380 190876 328132
rect 191492 324380 191548 328356
rect 192276 324380 192332 332612
rect 193732 324380 193788 332948
rect 194180 332668 194236 333312
rect 194180 332602 194236 332612
rect 194404 333116 194460 333126
rect 194404 324380 194460 333060
rect 196084 333002 196140 333312
rect 196084 332950 196086 333002
rect 196138 332950 196140 333002
rect 196084 332938 196140 332950
rect 194852 332892 194908 332902
rect 184996 324324 185108 324380
rect 185668 324324 185780 324380
rect 187124 324324 187236 324380
rect 187908 324324 188020 324380
rect 188580 324324 188692 324380
rect 189364 324324 189476 324380
rect 190036 324324 190148 324380
rect 190820 324324 190932 324380
rect 191492 324324 191604 324380
rect 192276 324324 192388 324380
rect 193732 324324 193844 324380
rect 194404 324324 194516 324380
rect 184884 323866 184940 323876
rect 185052 323680 185108 324324
rect 185724 323680 185780 324324
rect 186508 324156 186564 324166
rect 186508 323680 186564 324100
rect 187180 323680 187236 324324
rect 187964 323680 188020 324324
rect 188636 323680 188692 324324
rect 189420 323680 189476 324324
rect 190092 323680 190148 324324
rect 190876 323680 190932 324324
rect 191548 323680 191604 324324
rect 192332 323680 192388 324324
rect 193004 324156 193060 324166
rect 193004 323680 193060 324100
rect 193788 323680 193844 324324
rect 194460 323680 194516 324324
rect 194852 324268 194908 332836
rect 196644 332890 196700 332902
rect 196644 332838 196646 332890
rect 196698 332838 196700 332890
rect 195188 332780 195244 332790
rect 195188 324380 195244 332724
rect 196644 324380 196700 332838
rect 197876 332778 197932 332790
rect 197876 332726 197878 332778
rect 197930 332726 197932 332778
rect 197876 325947 197932 332726
rect 198100 332668 198156 333312
rect 198100 332602 198156 332612
rect 198324 332780 198380 332790
rect 198324 325947 198380 332724
rect 199556 332666 199612 332678
rect 199556 332614 199558 332666
rect 199610 332614 199612 332666
rect 197876 325891 198156 325947
rect 198324 325891 198828 325947
rect 198100 324380 198156 325891
rect 198772 324380 198828 325891
rect 199556 324380 199612 332614
rect 195188 324324 195300 324380
rect 196644 324324 196756 324380
rect 198100 324324 198212 324380
rect 198772 324324 198884 324380
rect 199556 324324 199668 324380
rect 194852 324202 194908 324212
rect 195244 323680 195300 324324
rect 195916 324268 195972 324278
rect 195916 323680 195972 324212
rect 196700 323680 196756 324324
rect 197372 323932 197428 323942
rect 197372 323680 197428 323876
rect 198156 323680 198212 324324
rect 198828 323680 198884 324324
rect 199612 323680 199668 324324
rect 200004 324268 200060 333312
rect 202160 333284 202524 333340
rect 200228 333002 200284 333014
rect 200228 332950 200230 333002
rect 200282 332950 200284 333002
rect 200228 324380 200284 332950
rect 202468 324380 202524 333284
rect 203364 332892 203420 332902
rect 200228 324324 200340 324380
rect 202468 324324 202580 324380
rect 200004 324202 200060 324212
rect 200284 323680 200340 324324
rect 201068 324268 201124 324278
rect 201068 323680 201124 324212
rect 201740 324156 201796 324166
rect 201740 323680 201796 324100
rect 202524 323680 202580 324324
rect 203196 324156 203252 324166
rect 203196 323680 203252 324100
rect 203364 324154 203420 332836
rect 203924 324380 203980 333312
rect 205044 333284 205968 333340
rect 203924 324324 204036 324380
rect 203364 324102 203366 324154
rect 203418 324102 203420 324154
rect 203364 324090 203420 324102
rect 203980 323680 204036 324324
rect 204652 324154 204708 324166
rect 204652 324102 204654 324154
rect 204706 324102 204708 324154
rect 204652 323680 204708 324102
rect 205044 324156 205100 333284
rect 207508 333228 207564 333238
rect 205380 332778 205436 332790
rect 205380 332726 205382 332778
rect 205434 332726 205436 332778
rect 205380 324380 205436 332726
rect 206836 332666 206892 332678
rect 206836 332614 206838 332666
rect 206890 332614 206892 332666
rect 206836 324380 206892 332614
rect 207508 324380 207564 333172
rect 207956 332892 208012 333312
rect 207956 332826 208012 332836
rect 208964 332892 209020 332902
rect 208964 324380 209020 332836
rect 209636 325947 209692 333620
rect 210644 333564 210700 333574
rect 209860 332668 209916 333312
rect 209860 332602 209916 332612
rect 210084 332668 210140 332678
rect 210084 325947 210140 332612
rect 210644 332668 210700 333508
rect 221620 333564 221676 333574
rect 221676 333508 221872 333564
rect 221620 333498 221676 333508
rect 216356 333452 216412 333462
rect 210644 332602 210700 332612
rect 211204 333116 211260 333126
rect 209636 325891 209804 325947
rect 210084 325891 210476 325947
rect 209748 324380 209804 325891
rect 205380 324324 205492 324380
rect 206836 324324 206948 324380
rect 207508 324324 207620 324380
rect 208964 324324 209076 324380
rect 209748 324324 209860 324380
rect 205044 324090 205100 324100
rect 205436 323680 205492 324324
rect 206108 324156 206164 324166
rect 206108 323680 206164 324100
rect 206892 323680 206948 324324
rect 207564 323680 207620 324324
rect 208348 324156 208404 324166
rect 208348 323680 208404 324100
rect 209020 323680 209076 324324
rect 209804 323680 209860 324324
rect 210420 324044 210476 325891
rect 211204 324380 211260 333060
rect 211764 333004 211820 333014
rect 211204 324324 211316 324380
rect 210420 323988 210532 324044
rect 210476 323680 210532 323988
rect 211260 323680 211316 324324
rect 211764 324268 211820 332948
rect 211876 332778 211932 333312
rect 211876 332726 211878 332778
rect 211930 332726 211932 332778
rect 211876 332714 211932 332726
rect 212100 332778 212156 332790
rect 212100 332726 212102 332778
rect 212154 332726 212156 332778
rect 212100 325947 212156 332726
rect 213892 332666 213948 333312
rect 215908 332780 215964 333312
rect 215908 332714 215964 332724
rect 213892 332614 213894 332666
rect 213946 332614 213948 332666
rect 213892 332602 213948 332614
rect 215124 330092 215180 330102
rect 211988 325891 212156 325947
rect 214228 328972 214284 328982
rect 211988 324380 212044 325891
rect 214228 324380 214284 328916
rect 215124 325947 215180 330036
rect 215124 325891 215628 325947
rect 211764 324202 211820 324212
rect 211932 324324 212044 324380
rect 214172 324324 214284 324380
rect 215572 324380 215628 325891
rect 216356 324380 216412 333396
rect 217028 333340 217084 333350
rect 216692 330764 216748 330774
rect 215572 324324 215684 324380
rect 216356 324324 216468 324380
rect 211932 323680 211988 324324
rect 212716 324268 212772 324278
rect 212716 323680 212772 324212
rect 213388 324156 213444 324166
rect 213388 323680 213444 324100
rect 214172 323680 214228 324324
rect 214844 324156 214900 324166
rect 214844 323680 214900 324100
rect 215628 323680 215684 324324
rect 216412 323680 216468 324324
rect 216692 324268 216748 330708
rect 217028 324380 217084 333284
rect 217140 333284 217840 333340
rect 217140 333228 217196 333284
rect 217140 333162 217196 333172
rect 218484 333228 218540 333238
rect 217476 332666 217532 332678
rect 217476 332614 217478 332666
rect 217530 332614 217532 332666
rect 217028 324324 217140 324380
rect 216692 324202 216748 324212
rect 217084 323680 217140 324324
rect 217476 324156 217532 332614
rect 218484 324380 218540 333172
rect 219828 332892 219884 333312
rect 219828 332826 219884 332836
rect 220164 333116 220220 333126
rect 219940 328636 219996 328646
rect 219940 324380 219996 328580
rect 220164 325947 220220 333060
rect 221396 333114 221452 333126
rect 221396 333062 221398 333114
rect 221450 333062 221452 333114
rect 220164 325891 220780 325947
rect 220724 324380 220780 325891
rect 221396 324380 221452 333062
rect 222292 328524 222348 328534
rect 222292 324380 222348 328468
rect 218484 324324 218596 324380
rect 219940 324324 220052 324380
rect 220724 324324 220836 324380
rect 221396 324324 221508 324380
rect 217476 324090 217532 324100
rect 217868 324268 217924 324278
rect 217868 323680 217924 324212
rect 218540 323680 218596 324324
rect 219324 324156 219380 324166
rect 219324 323680 219380 324100
rect 219996 323680 220052 324324
rect 220780 323680 220836 324324
rect 221452 323680 221508 324324
rect 222236 324324 222348 324380
rect 222852 324380 222908 333732
rect 258916 333788 258972 333798
rect 271012 333788 271068 333798
rect 258972 333732 259616 333788
rect 258916 333722 258972 333732
rect 223412 333676 223468 333686
rect 223468 333620 223888 333676
rect 223412 333610 223468 333620
rect 240996 333452 241052 333462
rect 241052 333396 241696 333452
rect 266532 333450 266588 333462
rect 266532 333398 266534 333450
rect 266586 333398 266588 333450
rect 240996 333386 241052 333396
rect 239092 333340 239148 333350
rect 240548 333340 240604 333350
rect 223636 333002 223692 333014
rect 223636 332950 223638 333002
rect 223690 332950 223692 333002
rect 223636 324380 223692 332950
rect 225204 332892 225260 332902
rect 224420 328412 224476 328422
rect 224420 324380 224476 328356
rect 225204 324380 225260 332836
rect 225764 332780 225820 333312
rect 227780 333004 227836 333312
rect 227780 332938 227836 332948
rect 225764 332714 225820 332724
rect 227220 332890 227276 332902
rect 227220 332838 227222 332890
rect 227274 332838 227276 332890
rect 226660 327962 226716 327974
rect 226660 327910 226662 327962
rect 226714 327910 226716 327962
rect 226660 324380 226716 327910
rect 222852 324324 222964 324380
rect 223636 324324 223748 324380
rect 222236 323680 222292 324324
rect 222908 323680 222964 324324
rect 223692 323680 223748 324324
rect 224364 324324 224476 324380
rect 225148 324324 225260 324380
rect 226604 324324 226716 324380
rect 227220 324380 227276 332838
rect 229460 332892 229516 332902
rect 228788 328186 228844 328198
rect 228788 328134 228790 328186
rect 228842 328134 228844 328186
rect 228116 328074 228172 328086
rect 228116 328022 228118 328074
rect 228170 328022 228172 328074
rect 228116 324380 228172 328022
rect 228788 324380 228844 328134
rect 227220 324324 227332 324380
rect 224364 323680 224420 324324
rect 225148 323680 225204 324324
rect 225820 324156 225876 324166
rect 225820 323680 225876 324100
rect 226604 323680 226660 324324
rect 227276 323680 227332 324324
rect 228060 324324 228172 324380
rect 228732 324324 228844 324380
rect 229460 324380 229516 332836
rect 229796 332778 229852 333312
rect 229796 332726 229798 332778
rect 229850 332726 229852 332778
rect 229796 332714 229852 332726
rect 231588 332778 231644 332790
rect 231588 332726 231590 332778
rect 231642 332726 231644 332778
rect 231028 328298 231084 328310
rect 231028 328246 231030 328298
rect 231082 328246 231084 328298
rect 231028 324380 231084 328246
rect 229460 324324 229572 324380
rect 228060 323680 228116 324324
rect 228732 323680 228788 324324
rect 229516 323680 229572 324324
rect 230972 324324 231084 324380
rect 231588 324380 231644 332726
rect 231812 332668 231868 333312
rect 231812 332602 231868 332612
rect 233604 332668 233660 332678
rect 233156 328188 233212 328198
rect 232484 328076 232540 328086
rect 232484 324380 232540 328020
rect 233156 324380 233212 328132
rect 231588 324324 231700 324380
rect 230188 324156 230244 324166
rect 230188 323680 230244 324100
rect 230972 323680 231028 324324
rect 231644 323680 231700 324324
rect 232428 324324 232540 324380
rect 233100 324324 233212 324380
rect 232428 323680 232484 324324
rect 233100 323680 233156 324324
rect 233604 324156 233660 332612
rect 233716 332666 233772 333312
rect 233716 332614 233718 332666
rect 233770 332614 233772 332666
rect 233716 332602 233772 332614
rect 233940 332666 233996 332678
rect 233940 332614 233942 332666
rect 233994 332614 233996 332666
rect 233940 324380 233996 332614
rect 233604 324090 233660 324100
rect 233884 324324 233996 324380
rect 235284 330652 235340 330662
rect 235284 324380 235340 330596
rect 235732 328972 235788 333312
rect 235732 328906 235788 328916
rect 237412 330540 237468 330550
rect 236068 327180 236124 327190
rect 236068 324380 236124 327124
rect 235284 324324 235396 324380
rect 233884 323680 233940 324324
rect 234556 324156 234612 324166
rect 234556 323680 234612 324100
rect 235340 323680 235396 324324
rect 236012 324324 236124 324380
rect 237412 324380 237468 330484
rect 237748 330092 237804 333312
rect 239148 333284 239792 333340
rect 239092 333274 239148 333284
rect 237748 330026 237804 330036
rect 238532 330428 238588 330438
rect 238308 327068 238364 327078
rect 238308 324380 238364 327012
rect 238532 325947 238588 330372
rect 239652 330316 239708 330326
rect 238532 325891 238924 325947
rect 237412 324324 237524 324380
rect 236012 323680 236068 324324
rect 236796 324156 236852 324166
rect 236796 323680 236852 324100
rect 237468 323680 237524 324324
rect 238252 324324 238364 324380
rect 238868 324380 238924 325891
rect 239652 324380 239708 330260
rect 240212 330314 240268 330326
rect 240212 330262 240214 330314
rect 240266 330262 240268 330314
rect 238868 324324 238980 324380
rect 239652 324324 239764 324380
rect 238252 323680 238308 324324
rect 238924 323680 238980 324324
rect 239708 323680 239764 324324
rect 240212 324268 240268 330262
rect 240548 325947 240604 333284
rect 243684 330764 243740 333312
rect 243684 330698 243740 330708
rect 243236 330202 243292 330214
rect 243236 330150 243238 330202
rect 243290 330150 243292 330202
rect 240436 325891 240604 325947
rect 242676 326956 242732 326966
rect 240436 324380 240492 325891
rect 242676 324380 242732 326900
rect 240212 324202 240268 324212
rect 240380 324324 240492 324380
rect 242620 324324 242732 324380
rect 243236 324380 243292 330150
rect 245476 330204 245532 330214
rect 244020 330090 244076 330102
rect 244020 330038 244022 330090
rect 244074 330038 244076 330090
rect 244020 324380 244076 330038
rect 244804 325388 244860 325398
rect 243236 324324 243348 324380
rect 244020 324324 244132 324380
rect 240380 323680 240436 324324
rect 241836 324268 241892 324278
rect 241164 323932 241220 323942
rect 241164 323680 241220 323876
rect 241836 323680 241892 324212
rect 242620 323680 242676 324324
rect 243292 323680 243348 324324
rect 244076 323680 244132 324324
rect 244804 324268 244860 325332
rect 245476 324380 245532 330148
rect 245700 328748 245756 333312
rect 247044 333284 247744 333340
rect 247044 333228 247100 333284
rect 247044 333162 247100 333172
rect 249396 330426 249452 330438
rect 249396 330374 249398 330426
rect 249450 330374 249452 330426
rect 245700 328682 245756 328692
rect 246260 329196 246316 329206
rect 246260 324380 246316 329140
rect 247716 329194 247772 329206
rect 247716 329142 247718 329194
rect 247770 329142 247772 329194
rect 245476 324324 245588 324380
rect 244748 324212 244860 324268
rect 244748 323680 244804 324212
rect 245532 323680 245588 324324
rect 246204 324324 246316 324380
rect 247044 325276 247100 325286
rect 246204 323680 246260 324324
rect 247044 324156 247100 325220
rect 247716 324380 247772 329142
rect 248500 329082 248556 329094
rect 248500 329030 248502 329082
rect 248554 329030 248556 329082
rect 248500 324380 248556 329030
rect 246988 324100 247100 324156
rect 247660 324324 247772 324380
rect 248444 324324 248556 324380
rect 249172 325164 249228 325174
rect 246988 323680 247044 324100
rect 247660 323680 247716 324324
rect 248444 323680 248500 324324
rect 249172 324156 249228 325108
rect 249116 324100 249228 324156
rect 249116 323680 249172 324100
rect 249396 323932 249452 330374
rect 249620 328636 249676 333312
rect 251636 333114 251692 333312
rect 251636 333062 251638 333114
rect 251690 333062 251692 333114
rect 251636 333050 251692 333062
rect 253652 333116 253708 333312
rect 253652 333050 253708 333060
rect 249620 328570 249676 328580
rect 249956 329084 250012 329094
rect 249956 324380 250012 329028
rect 250628 328970 250684 328982
rect 250628 328918 250630 328970
rect 250682 328918 250684 328970
rect 250628 324380 250684 328918
rect 252084 328972 252140 328982
rect 249396 323866 249452 323876
rect 249900 324324 250012 324380
rect 250572 324324 250684 324380
rect 251412 325052 251468 325062
rect 249900 323680 249956 324324
rect 250572 323680 250628 324324
rect 251412 324044 251468 324996
rect 252084 324380 252140 328916
rect 252868 328858 252924 328870
rect 252868 328806 252870 328858
rect 252922 328806 252924 328858
rect 252868 324380 252924 328806
rect 254324 328748 254380 328758
rect 254324 324380 254380 328692
rect 254996 328636 255052 328646
rect 254996 324380 255052 328580
rect 255668 328524 255724 333312
rect 257572 333002 257628 333312
rect 257572 332950 257574 333002
rect 257626 332950 257628 333002
rect 257572 332938 257628 332950
rect 257124 330092 257180 330102
rect 255668 328458 255724 328468
rect 256452 328746 256508 328758
rect 256452 328694 256454 328746
rect 256506 328694 256508 328746
rect 256452 324380 256508 328694
rect 251356 323988 251468 324044
rect 252028 324324 252140 324380
rect 252812 324324 252924 324380
rect 254268 324324 254380 324380
rect 254940 324324 255052 324380
rect 256396 324324 256508 324380
rect 257124 324380 257180 330036
rect 260820 328634 260876 328646
rect 260820 328582 260822 328634
rect 260874 328582 260876 328634
rect 257908 326844 257964 326854
rect 257908 324380 257964 326788
rect 260820 324380 260876 328582
rect 261604 328412 261660 333312
rect 263620 328860 263676 333312
rect 265524 332780 265580 333312
rect 265524 332714 265580 332724
rect 263620 328794 263676 328804
rect 261604 328346 261660 328356
rect 263060 328410 263116 328422
rect 263060 328358 263062 328410
rect 263114 328358 263116 328410
rect 257124 324324 257236 324380
rect 251356 323680 251412 323988
rect 252028 323680 252084 324324
rect 252812 323680 252868 324324
rect 253484 324156 253540 324166
rect 253484 323680 253540 324100
rect 254268 323680 254324 324324
rect 254940 323680 254996 324324
rect 255724 324156 255780 324166
rect 255724 323680 255780 324100
rect 256396 323680 256452 324324
rect 257180 323680 257236 324324
rect 257852 324324 257964 324380
rect 260764 324324 260876 324380
rect 262276 325274 262332 325286
rect 262276 325222 262278 325274
rect 262330 325222 262332 325274
rect 257852 323680 257908 324324
rect 258636 324156 258692 324166
rect 258636 323680 258692 324100
rect 259308 324156 259364 324166
rect 259308 323680 259364 324100
rect 260092 324044 260148 324054
rect 260092 323680 260148 323988
rect 260764 323680 260820 324324
rect 261548 324156 261604 324166
rect 262276 324156 262332 325222
rect 263060 324380 263116 328358
rect 265188 328412 265244 328422
rect 264516 325610 264572 325622
rect 264516 325558 264518 325610
rect 264570 325558 264572 325610
rect 264516 324380 264572 325558
rect 265188 324380 265244 328356
rect 261548 323680 261604 324100
rect 262220 324100 262332 324156
rect 263004 324324 263116 324380
rect 264460 324324 264572 324380
rect 265132 324324 265244 324380
rect 265972 325050 266028 325062
rect 265972 324998 265974 325050
rect 266026 324998 266028 325050
rect 262220 323680 262276 324100
rect 263004 323680 263060 324324
rect 263676 324156 263732 324166
rect 263676 323680 263732 324100
rect 264460 323680 264516 324324
rect 265132 323680 265188 324324
rect 265972 324044 266028 324998
rect 266532 324380 266588 333398
rect 267428 328522 267484 328534
rect 267428 328470 267430 328522
rect 267482 328470 267484 328522
rect 267428 324380 267484 328470
rect 267540 327962 267596 333312
rect 269108 333226 269164 333238
rect 269108 333174 269110 333226
rect 269162 333174 269164 333226
rect 267540 327910 267542 327962
rect 267594 327910 267596 327962
rect 267540 327898 267596 327910
rect 267988 331548 268044 331558
rect 266532 324324 266644 324380
rect 265916 323988 266028 324044
rect 265916 323680 265972 323988
rect 266588 323680 266644 324324
rect 267372 324324 267484 324380
rect 267988 324380 268044 331492
rect 269108 325947 269164 333174
rect 269556 328074 269612 333312
rect 269556 328022 269558 328074
rect 269610 328022 269612 328074
rect 269556 328010 269612 328022
rect 270228 331212 270284 331222
rect 268884 325891 269164 325947
rect 268884 324380 268940 325891
rect 267988 324324 268100 324380
rect 267372 323680 267428 324324
rect 268044 323680 268100 324324
rect 268828 324324 268940 324380
rect 270228 324380 270284 331156
rect 271012 324380 271068 333732
rect 388052 333788 388108 333798
rect 656740 333788 656796 333798
rect 388108 333732 388752 333788
rect 656796 333732 656992 333788
rect 388052 333722 388108 333732
rect 656740 333722 656796 333732
rect 278292 333676 278348 333686
rect 271460 332890 271516 333312
rect 271460 332838 271462 332890
rect 271514 332838 271516 332890
rect 271460 332826 271516 332838
rect 273140 333228 273196 333238
rect 272244 331324 272300 331334
rect 272244 325947 272300 331268
rect 272244 325891 272524 325947
rect 271796 325162 271852 325174
rect 271796 325110 271798 325162
rect 271850 325110 271852 325162
rect 270228 324324 270340 324380
rect 271012 324324 271124 324380
rect 268828 323680 268884 324324
rect 269500 324156 269556 324166
rect 269500 323680 269556 324100
rect 270284 323680 270340 324324
rect 271068 323680 271124 324324
rect 271796 324156 271852 325110
rect 272468 324380 272524 325891
rect 273140 324380 273196 333172
rect 273476 328186 273532 333312
rect 275380 333114 275436 333126
rect 275380 333062 275382 333114
rect 275434 333062 275436 333114
rect 273476 328134 273478 328186
rect 273530 328134 273532 328186
rect 273476 328122 273532 328134
rect 274596 331436 274652 331446
rect 274596 324380 274652 331380
rect 275380 324380 275436 333062
rect 275492 327964 275548 333312
rect 277508 332892 277564 333312
rect 277508 332826 277564 332836
rect 277396 332780 277452 332790
rect 276836 331210 276892 331222
rect 276836 331158 276838 331210
rect 276890 331158 276892 331210
rect 275492 327898 275548 327908
rect 276164 328074 276220 328086
rect 276164 328022 276166 328074
rect 276218 328022 276220 328074
rect 276164 324380 276220 328022
rect 272468 324324 272580 324380
rect 273140 324324 273252 324380
rect 274596 324324 274708 324380
rect 275380 324324 275492 324380
rect 271740 324100 271852 324156
rect 271740 323680 271796 324100
rect 272524 323680 272580 324324
rect 273196 323680 273252 324324
rect 273980 324156 274036 324166
rect 273980 323680 274036 324100
rect 274652 323680 274708 324324
rect 275436 323680 275492 324324
rect 276108 324324 276220 324380
rect 276836 324380 276892 331158
rect 277396 325947 277452 332724
rect 278292 332780 278348 333620
rect 406420 333676 406476 333686
rect 406476 333620 406672 333676
rect 406420 333610 406476 333620
rect 284228 333562 284284 333574
rect 284228 333510 284230 333562
rect 284282 333510 284284 333562
rect 278292 332714 278348 332724
rect 278964 332218 279020 332230
rect 278964 332166 278966 332218
rect 279018 332166 279020 332218
rect 278404 326732 278460 326742
rect 277396 325891 277564 325947
rect 277508 324380 277564 325891
rect 278404 324380 278460 326676
rect 276836 324324 276948 324380
rect 277508 324324 277620 324380
rect 276108 323680 276164 324324
rect 276892 323680 276948 324324
rect 277564 323680 277620 324324
rect 278348 324324 278460 324380
rect 278964 324380 279020 332166
rect 279412 328298 279468 333312
rect 279412 328246 279414 328298
rect 279466 328246 279468 328298
rect 279412 328234 279468 328246
rect 279748 332890 279804 332902
rect 279748 332838 279750 332890
rect 279802 332838 279804 332890
rect 279748 324380 279804 332838
rect 280644 332892 280700 332902
rect 280420 326506 280476 326518
rect 280420 326454 280422 326506
rect 280474 326454 280476 326506
rect 280420 324380 280476 326454
rect 278964 324324 279076 324380
rect 279748 324324 279860 324380
rect 280420 324324 280532 324380
rect 278348 323680 278404 324324
rect 279020 323680 279076 324324
rect 279804 323680 279860 324324
rect 280476 323680 280532 324324
rect 280644 324266 280700 332836
rect 281204 331322 281260 331334
rect 281204 331270 281206 331322
rect 281258 331270 281260 331322
rect 281204 324380 281260 331270
rect 281428 328076 281484 333312
rect 283444 332778 283500 333312
rect 283444 332726 283446 332778
rect 283498 332726 283500 332778
rect 283444 332714 283500 332726
rect 281428 328010 281484 328020
rect 283332 331434 283388 331446
rect 283332 331382 283334 331434
rect 283386 331382 283388 331434
rect 282772 326396 282828 326406
rect 282772 324380 282828 326340
rect 281204 324324 281316 324380
rect 280644 324214 280646 324266
rect 280698 324214 280700 324266
rect 280644 324202 280700 324214
rect 281260 323680 281316 324324
rect 282716 324324 282828 324380
rect 283332 324380 283388 331382
rect 284228 324380 284284 333510
rect 320180 333564 320236 333574
rect 319956 333452 320012 333462
rect 319732 333396 319956 333452
rect 304612 333340 304668 333350
rect 285460 328188 285516 333312
rect 286244 333004 286300 333014
rect 285460 328122 285516 328132
rect 285572 329644 285628 329654
rect 284900 326618 284956 326630
rect 284900 326566 284902 326618
rect 284954 326566 284956 326618
rect 284900 324380 284956 326566
rect 283332 324324 283444 324380
rect 281932 324266 281988 324278
rect 281932 324214 281934 324266
rect 281986 324214 281988 324266
rect 281932 323680 281988 324214
rect 282716 323680 282772 324324
rect 283388 323680 283444 324324
rect 284172 324324 284284 324380
rect 284844 324324 284956 324380
rect 285572 324380 285628 329588
rect 286244 324380 286300 332948
rect 287364 332668 287420 333312
rect 287364 332602 287420 332612
rect 288484 332778 288540 332790
rect 288484 332726 288486 332778
rect 288538 332726 288540 332778
rect 287252 329756 287308 329766
rect 287252 325947 287308 329700
rect 287252 325891 287756 325947
rect 287700 324380 287756 325891
rect 288484 324380 288540 332726
rect 289380 332666 289436 333312
rect 289380 332614 289382 332666
rect 289434 332614 289436 332666
rect 289380 332602 289436 332614
rect 290724 333116 290780 333126
rect 289940 329866 289996 329878
rect 289940 329814 289942 329866
rect 289994 329814 289996 329866
rect 289268 327514 289324 327526
rect 289268 327462 289270 327514
rect 289322 327462 289324 327514
rect 289268 324380 289324 327462
rect 285572 324324 285684 324380
rect 286244 324324 286356 324380
rect 287700 324324 287812 324380
rect 288484 324324 288596 324380
rect 284172 323680 284228 324324
rect 284844 323680 284900 324324
rect 285628 323680 285684 324324
rect 286300 323680 286356 324324
rect 287084 323930 287140 323942
rect 287084 323878 287086 323930
rect 287138 323878 287140 323930
rect 287084 323680 287140 323878
rect 287756 323680 287812 324324
rect 288540 323680 288596 324324
rect 289212 324324 289324 324380
rect 289940 324380 289996 329814
rect 290724 324380 290780 333060
rect 291396 330652 291452 333312
rect 291396 330586 291452 330596
rect 289940 324324 290052 324380
rect 289212 323680 289268 324324
rect 289996 323680 290052 324324
rect 290668 324324 290780 324380
rect 292068 329978 292124 329990
rect 292068 329926 292070 329978
rect 292122 329926 292124 329978
rect 292068 324380 292124 329926
rect 293412 328300 293468 333312
rect 293412 328234 293468 328244
rect 294308 330874 294364 330886
rect 294308 330822 294310 330874
rect 294362 330822 294364 330874
rect 293636 326508 293692 326518
rect 292964 325500 293020 325510
rect 292068 324324 292180 324380
rect 290668 323680 290724 324324
rect 291452 324156 291508 324166
rect 291452 323680 291508 324100
rect 292124 323680 292180 324324
rect 292964 324268 293020 325444
rect 293636 324380 293692 326452
rect 292908 324212 293020 324268
rect 293580 324324 293692 324380
rect 294308 324380 294364 330822
rect 295316 327180 295372 333312
rect 297332 330540 297388 333312
rect 297332 330474 297388 330484
rect 298676 330762 298732 330774
rect 298676 330710 298678 330762
rect 298730 330710 298732 330762
rect 295316 327114 295372 327124
rect 296436 329868 296492 329878
rect 295092 324604 295148 324614
rect 294308 324324 294420 324380
rect 292908 323680 292964 324212
rect 293580 323680 293636 324324
rect 294364 323680 294420 324324
rect 295092 323932 295148 324548
rect 296436 324380 296492 329812
rect 298004 328188 298060 328198
rect 297220 327962 297276 327974
rect 297220 327910 297222 327962
rect 297274 327910 297276 327962
rect 297220 324380 297276 327910
rect 298004 324380 298060 328132
rect 296436 324324 296548 324380
rect 297220 324324 297332 324380
rect 295036 323876 295148 323932
rect 295820 324156 295876 324166
rect 295036 323680 295092 323876
rect 295820 323680 295876 324100
rect 296492 323680 296548 324324
rect 297276 323680 297332 324324
rect 297948 324324 298060 324380
rect 298676 324380 298732 330710
rect 299348 327068 299404 333312
rect 301364 330428 301420 333312
rect 301364 330362 301420 330372
rect 303044 330876 303100 330886
rect 299348 327002 299404 327012
rect 300804 329980 300860 329990
rect 300244 326620 300300 326630
rect 299796 326394 299852 326406
rect 299796 326342 299798 326394
rect 299850 326342 299852 326394
rect 298676 324324 298788 324380
rect 297948 323680 298004 324324
rect 298732 323680 298788 324324
rect 299404 324156 299460 324166
rect 299404 323680 299460 324100
rect 299796 323930 299852 326342
rect 300244 324380 300300 326564
rect 299796 323878 299798 323930
rect 299850 323878 299852 323930
rect 299796 323866 299852 323878
rect 300188 324324 300300 324380
rect 300804 324380 300860 329924
rect 301700 328186 301756 328198
rect 301700 328134 301702 328186
rect 301754 328134 301756 328186
rect 301700 324380 301756 328134
rect 300804 324324 300916 324380
rect 300188 323680 300244 324324
rect 300860 323680 300916 324324
rect 301644 324324 301756 324380
rect 303044 324380 303100 330820
rect 303268 330316 303324 333312
rect 304668 333284 305312 333340
rect 304612 333274 304668 333284
rect 303268 330250 303324 330260
rect 305172 330650 305228 330662
rect 305172 330598 305174 330650
rect 305226 330598 305228 330650
rect 304612 326060 304668 326070
rect 303828 325724 303884 325734
rect 303828 324380 303884 325668
rect 304612 324380 304668 326004
rect 303044 324324 303156 324380
rect 301644 323680 301700 324324
rect 302316 324156 302372 324166
rect 302316 323680 302372 324100
rect 303100 323680 303156 324324
rect 303772 324324 303884 324380
rect 304556 324324 304668 324380
rect 305172 324380 305228 330598
rect 307300 330426 307356 333312
rect 307300 330374 307302 330426
rect 307354 330374 307356 330426
rect 307300 330362 307356 330374
rect 307524 330764 307580 330774
rect 306740 327402 306796 327414
rect 306740 327350 306742 327402
rect 306794 327350 306796 327402
rect 306740 324380 306796 327350
rect 307524 324380 307580 330708
rect 309316 330314 309372 333312
rect 309316 330262 309318 330314
rect 309370 330262 309372 330314
rect 309316 330250 309372 330262
rect 309540 330538 309596 330550
rect 309540 330486 309542 330538
rect 309594 330486 309596 330538
rect 305172 324324 305284 324380
rect 303772 323680 303828 324324
rect 304556 323680 304612 324324
rect 305228 323680 305284 324324
rect 306684 324324 306796 324380
rect 307468 324324 307580 324380
rect 308196 324492 308252 324502
rect 306012 324156 306068 324166
rect 306012 323680 306068 324100
rect 306684 323680 306740 324324
rect 307468 323680 307524 324324
rect 308196 323932 308252 324436
rect 309540 324380 309596 330486
rect 311220 326956 311276 333312
rect 311220 326890 311276 326900
rect 311780 330652 311836 330662
rect 310436 325498 310492 325510
rect 310436 325446 310438 325498
rect 310490 325446 310492 325498
rect 309540 324324 309652 324380
rect 308140 323876 308252 323932
rect 308924 324156 308980 324166
rect 308140 323680 308196 323876
rect 308924 323680 308980 324100
rect 309596 323680 309652 324324
rect 310436 324268 310492 325446
rect 311780 324380 311836 330596
rect 313236 330202 313292 333312
rect 313236 330150 313238 330202
rect 313290 330150 313292 330202
rect 313236 330138 313292 330150
rect 313908 330426 313964 330438
rect 313908 330374 313910 330426
rect 313962 330374 313964 330426
rect 313348 327290 313404 327302
rect 313348 327238 313350 327290
rect 313402 327238 313404 327290
rect 312564 325722 312620 325734
rect 312564 325670 312566 325722
rect 312618 325670 312620 325722
rect 312564 324380 312620 325670
rect 313348 324380 313404 327238
rect 311780 324324 311892 324380
rect 310380 324212 310492 324268
rect 310380 323680 310436 324212
rect 311052 324156 311108 324166
rect 311052 323680 311108 324100
rect 311836 323680 311892 324324
rect 312508 324324 312620 324380
rect 313292 324324 313404 324380
rect 313908 324380 313964 330374
rect 315252 330090 315308 333312
rect 315252 330038 315254 330090
rect 315306 330038 315308 330090
rect 315252 330026 315308 330038
rect 315812 333284 317296 333340
rect 315476 327178 315532 327190
rect 315476 327126 315478 327178
rect 315530 327126 315532 327178
rect 314804 325386 314860 325398
rect 314804 325334 314806 325386
rect 314858 325334 314860 325386
rect 313908 324324 314020 324380
rect 312508 323680 312564 324324
rect 313292 323680 313348 324324
rect 313964 323680 314020 324324
rect 314804 324268 314860 325334
rect 315476 324380 315532 327126
rect 315812 325388 315868 333284
rect 318276 331660 318332 331670
rect 315812 325322 315868 325332
rect 316148 330540 316204 330550
rect 314748 324212 314860 324268
rect 315420 324324 315532 324380
rect 316148 324380 316204 330484
rect 318276 324380 318332 331604
rect 319172 330204 319228 333312
rect 319172 330138 319228 330148
rect 319060 328298 319116 328310
rect 319060 328246 319062 328298
rect 319114 328246 319116 328298
rect 319060 324380 319116 328246
rect 319620 327180 319676 327190
rect 319620 324380 319676 327124
rect 319732 325610 319788 333396
rect 319956 333386 320012 333396
rect 320068 333002 320124 333014
rect 320068 332950 320070 333002
rect 320122 332950 320124 333002
rect 319844 331546 319900 331558
rect 319844 331494 319846 331546
rect 319898 331494 319900 331546
rect 319844 325947 319900 331494
rect 319844 325891 320012 325947
rect 319732 325558 319734 325610
rect 319786 325558 319788 325610
rect 319732 325546 319788 325558
rect 319956 324380 320012 325891
rect 320068 325500 320124 332950
rect 320068 325434 320124 325444
rect 320180 325274 320236 333508
rect 364532 333564 364588 333574
rect 386036 333564 386092 333574
rect 364588 333508 364896 333564
rect 364532 333498 364588 333508
rect 370244 333452 370300 333462
rect 376292 333452 376348 333462
rect 370300 333396 370944 333452
rect 376292 333450 376880 333452
rect 376292 333398 376294 333450
rect 376346 333398 376880 333450
rect 376292 333396 376880 333398
rect 370244 333386 370300 333396
rect 376292 333386 376348 333396
rect 321188 329196 321244 333312
rect 321188 329130 321244 329140
rect 322532 333284 323232 333340
rect 322084 327066 322140 327078
rect 322084 327014 322086 327066
rect 322138 327014 322140 327066
rect 320180 325222 320182 325274
rect 320234 325222 320236 325274
rect 320180 325210 320236 325222
rect 321300 325612 321356 325622
rect 321300 324380 321356 325556
rect 322084 324380 322140 327014
rect 322532 325276 322588 333284
rect 324884 332556 324940 332566
rect 322532 325210 322588 325220
rect 322644 330314 322700 330326
rect 322644 330262 322646 330314
rect 322698 330262 322700 330314
rect 316148 324324 316260 324380
rect 318276 324324 318388 324380
rect 319060 324324 319172 324380
rect 319620 324324 319844 324380
rect 319956 324324 320628 324380
rect 314748 323680 314804 324212
rect 315420 323680 315476 324324
rect 316204 323680 316260 324324
rect 317660 324156 317716 324166
rect 316876 323932 316932 323942
rect 316876 323680 316932 323876
rect 317660 323680 317716 324100
rect 318332 323680 318388 324324
rect 319116 323680 319172 324324
rect 319788 323680 319844 324324
rect 320572 323680 320628 324324
rect 321244 324324 321356 324380
rect 322028 324324 322140 324380
rect 322644 324380 322700 330262
rect 323540 325274 323596 325286
rect 323540 325222 323542 325274
rect 323594 325222 323596 325274
rect 322644 324324 322756 324380
rect 321244 323680 321300 324324
rect 322028 323680 322084 324324
rect 322700 323680 322756 324324
rect 323540 324156 323596 325222
rect 324884 324380 324940 332500
rect 325220 329194 325276 333312
rect 325220 329142 325222 329194
rect 325274 329142 325276 329194
rect 325220 329130 325276 329142
rect 326004 331658 326060 331670
rect 326004 331606 326006 331658
rect 326058 331606 326060 331658
rect 326004 325947 326060 331606
rect 327124 329082 327180 333312
rect 327572 333284 329168 333340
rect 327124 329030 327126 329082
rect 327178 329030 327180 329082
rect 327124 329018 327180 329030
rect 327236 332442 327292 332454
rect 327236 332390 327238 332442
rect 327290 332390 327292 332442
rect 326004 325891 326396 325947
rect 326340 324380 326396 325891
rect 327236 324380 327292 332390
rect 327572 325164 327628 333284
rect 329252 332444 329308 332454
rect 328692 326956 328748 326966
rect 327572 325098 327628 325108
rect 327908 325500 327964 325510
rect 324884 324324 324996 324380
rect 326340 324324 326452 324380
rect 323484 324100 323596 324156
rect 323484 323680 323540 324100
rect 324156 323932 324212 323942
rect 324156 323680 324212 323876
rect 324940 323680 324996 324324
rect 325724 324044 325780 324054
rect 325724 323680 325780 323988
rect 326396 323680 326452 324324
rect 327180 324324 327292 324380
rect 327180 323680 327236 324324
rect 327908 324268 327964 325444
rect 328692 324380 328748 326900
rect 327852 324212 327964 324268
rect 328636 324324 328748 324380
rect 329252 324380 329308 332388
rect 331156 329084 331212 333312
rect 331156 329018 331212 329028
rect 331492 332330 331548 332342
rect 331492 332278 331494 332330
rect 331546 332278 331548 332330
rect 330148 325388 330204 325398
rect 329252 324324 329364 324380
rect 327852 323680 327908 324212
rect 328636 323680 328692 324324
rect 329308 323680 329364 324324
rect 330148 324268 330204 325332
rect 331492 324380 331548 332278
rect 333060 328970 333116 333312
rect 333060 328918 333062 328970
rect 333114 328918 333116 328970
rect 333060 328906 333116 328918
rect 334292 333284 335104 333340
rect 369684 333338 369740 333350
rect 333060 326954 333116 326966
rect 333060 326902 333062 326954
rect 333114 326902 333116 326954
rect 333060 324380 333116 326902
rect 334292 325052 334348 333284
rect 335972 330204 336028 330214
rect 335300 329082 335356 329094
rect 335300 329030 335302 329082
rect 335354 329030 335356 329082
rect 335188 327964 335244 327974
rect 335076 327852 335132 327862
rect 334292 324986 334348 324996
rect 334516 325276 334572 325286
rect 331492 324324 331604 324380
rect 330092 324212 330204 324268
rect 330092 323680 330148 324212
rect 330764 324156 330820 324166
rect 330764 323680 330820 324100
rect 331548 323680 331604 324324
rect 333004 324324 333116 324380
rect 332220 323932 332276 323942
rect 332220 323680 332276 323876
rect 333004 323680 333060 324324
rect 334516 324156 334572 325220
rect 335076 325162 335132 327796
rect 335076 325110 335078 325162
rect 335130 325110 335132 325162
rect 335076 325098 335132 325110
rect 335188 325050 335244 327908
rect 335188 324998 335190 325050
rect 335242 324998 335244 325050
rect 335188 324986 335244 324998
rect 335300 324380 335356 329030
rect 335972 328300 336028 330148
rect 337092 328972 337148 333312
rect 337092 328906 337148 328916
rect 339108 328858 339164 333312
rect 339108 328806 339110 328858
rect 339162 328806 339164 328858
rect 339108 328794 339164 328806
rect 335972 328234 336028 328244
rect 338100 328300 338156 328310
rect 334460 324100 334572 324156
rect 335132 324324 335356 324380
rect 337428 325052 337484 325062
rect 333676 323932 333732 323942
rect 333676 323680 333732 323876
rect 334460 323680 334516 324100
rect 335132 323680 335188 324324
rect 336588 324156 336644 324166
rect 335916 324044 335972 324054
rect 335916 323680 335972 323988
rect 336588 323680 336644 324100
rect 337428 324044 337484 324996
rect 338100 324380 338156 328244
rect 341012 327068 341068 333312
rect 342468 329196 342524 329206
rect 341012 327002 341068 327012
rect 341796 327068 341852 327078
rect 340340 325164 340396 325174
rect 337372 323988 337484 324044
rect 338044 324324 338156 324380
rect 338884 324826 338940 324838
rect 338884 324774 338886 324826
rect 338938 324774 338940 324826
rect 337372 323680 337428 323988
rect 338044 323680 338100 324324
rect 338884 323932 338940 324774
rect 338828 323876 338940 323932
rect 339500 324156 339556 324166
rect 340340 324156 340396 325108
rect 338828 323680 338884 323876
rect 339500 323680 339556 324100
rect 340284 324100 340396 324156
rect 340900 324714 340956 324726
rect 340900 324662 340902 324714
rect 340954 324662 340956 324714
rect 340284 323680 340340 324100
rect 340900 323932 340956 324662
rect 341796 324380 341852 327012
rect 342468 324380 342524 329140
rect 343028 328748 343084 333312
rect 343028 328682 343084 328692
rect 343812 332106 343868 332118
rect 343812 332054 343814 332106
rect 343866 332054 343868 332106
rect 343476 327964 343532 327974
rect 343532 327908 343756 327964
rect 343476 327898 343532 327908
rect 343700 327852 343756 327908
rect 343700 327786 343756 327796
rect 341740 324324 341852 324380
rect 342412 324324 342524 324380
rect 343252 324938 343308 324950
rect 343252 324886 343254 324938
rect 343306 324886 343308 324938
rect 340900 323876 341012 323932
rect 340956 323680 341012 323876
rect 341740 323680 341796 324324
rect 342412 323680 342468 324324
rect 343252 324044 343308 324886
rect 343812 324380 343868 332054
rect 344708 329084 344764 329094
rect 344708 324380 344764 329028
rect 345044 328636 345100 333312
rect 347060 330316 347116 333312
rect 347060 330250 347116 330260
rect 347732 332108 347788 332118
rect 346052 329532 346108 329542
rect 345044 328570 345100 328580
rect 345268 328636 345324 328646
rect 345268 326844 345324 328580
rect 346052 327628 346108 329476
rect 346052 327562 346108 327572
rect 346164 329420 346220 329430
rect 345268 326778 345324 326788
rect 343812 324324 343924 324380
rect 343196 323988 343308 324044
rect 343196 323680 343252 323988
rect 343868 323680 343924 324324
rect 344652 324324 344764 324380
rect 345380 324716 345436 324726
rect 344652 323680 344708 324324
rect 345380 323932 345436 324660
rect 346164 324380 346220 329364
rect 345324 323876 345436 323932
rect 346108 324324 346220 324380
rect 346724 328970 346780 328982
rect 346724 328918 346726 328970
rect 346778 328918 346780 328970
rect 346724 324380 346780 328918
rect 347732 327740 347788 332052
rect 348964 328746 349020 333312
rect 350980 330092 351036 333312
rect 350980 330026 351036 330036
rect 352548 331994 352604 332006
rect 352548 331942 352550 331994
rect 352602 331942 352604 331994
rect 348964 328694 348966 328746
rect 349018 328694 349020 328746
rect 348964 328682 349020 328694
rect 349076 328972 349132 328982
rect 347732 327674 347788 327684
rect 348292 326842 348348 326854
rect 348292 326790 348294 326842
rect 348346 326790 348348 326842
rect 348292 324380 348348 326790
rect 349076 324380 349132 328916
rect 351204 328858 351260 328870
rect 351204 328806 351206 328858
rect 351258 328806 351260 328858
rect 350532 326844 350588 326854
rect 346724 324324 346836 324380
rect 345324 323680 345380 323876
rect 346108 323680 346164 324324
rect 346780 323680 346836 324324
rect 348236 324324 348348 324380
rect 349020 324324 349132 324380
rect 349748 324828 349804 324838
rect 347564 324156 347620 324166
rect 347564 323680 347620 324100
rect 348236 323680 348292 324324
rect 349020 323680 349076 324324
rect 349748 323932 349804 324772
rect 350532 324380 350588 326788
rect 351204 324380 351260 328806
rect 351988 325834 352044 325846
rect 351988 325782 351990 325834
rect 352042 325782 352044 325834
rect 351988 324380 352044 325782
rect 349692 323876 349804 323932
rect 350476 324324 350588 324380
rect 351148 324324 351260 324380
rect 351932 324324 352044 324380
rect 352548 324380 352604 331942
rect 352996 328636 353052 333312
rect 354116 330316 354172 330326
rect 353892 329194 353948 329206
rect 353892 329142 353894 329194
rect 353946 329142 353948 329194
rect 352996 328570 353052 328580
rect 353444 328748 353500 328758
rect 353444 324380 353500 328692
rect 353892 325164 353948 329142
rect 354116 327068 354172 330260
rect 354788 330202 354844 330214
rect 354788 330150 354790 330202
rect 354842 330150 354844 330202
rect 354564 330090 354620 330102
rect 354564 330038 354566 330090
rect 354618 330038 354620 330090
rect 354116 327002 354172 327012
rect 354340 327068 354396 327078
rect 353892 325098 353948 325108
rect 354340 325052 354396 327012
rect 354340 324986 354396 324996
rect 352548 324324 352660 324380
rect 349692 323680 349748 323876
rect 350476 323680 350532 324324
rect 351148 323680 351204 324324
rect 351932 323680 351988 324324
rect 352604 323680 352660 324324
rect 353388 324324 353500 324380
rect 354116 324940 354172 324950
rect 353388 323680 353444 324324
rect 354116 324044 354172 324884
rect 354564 324266 354620 330038
rect 354788 324380 354844 330150
rect 355012 328524 355068 333312
rect 356916 330204 356972 333312
rect 358932 332668 358988 333312
rect 358932 332602 358988 332612
rect 359492 332332 359548 332342
rect 356916 330138 356972 330148
rect 359156 330204 359212 330214
rect 355012 328458 355068 328468
rect 357700 328746 357756 328758
rect 357700 328694 357702 328746
rect 357754 328694 357756 328746
rect 356356 325610 356412 325622
rect 356356 325558 356358 325610
rect 356410 325558 356412 325610
rect 356356 324380 356412 325558
rect 354788 324324 354900 324380
rect 354564 324214 354566 324266
rect 354618 324214 354620 324266
rect 354564 324202 354620 324214
rect 354060 323988 354172 324044
rect 354060 323680 354116 323988
rect 354844 323680 354900 324324
rect 356300 324324 356412 324380
rect 357700 324380 357756 328694
rect 359156 324380 359212 330148
rect 359492 329420 359548 332276
rect 359492 329354 359548 329364
rect 359828 330092 359884 330102
rect 359828 324380 359884 330036
rect 360948 328634 361004 333312
rect 362964 332108 363020 333312
rect 362964 332042 363020 332052
rect 366436 332108 366492 332118
rect 360948 328582 360950 328634
rect 361002 328582 361004 328634
rect 360948 328570 361004 328582
rect 362180 328634 362236 328646
rect 362180 328582 362182 328634
rect 362234 328582 362236 328634
rect 360724 325724 360780 325734
rect 360724 324380 360780 325668
rect 362180 324380 362236 328582
rect 364308 328524 364364 328534
rect 363636 326730 363692 326742
rect 363636 326678 363638 326730
rect 363690 326678 363692 326730
rect 357700 324324 357812 324380
rect 359156 324324 359268 324380
rect 359828 324324 359940 324380
rect 355516 324266 355572 324278
rect 355516 324214 355518 324266
rect 355570 324214 355572 324266
rect 355516 323680 355572 324214
rect 356300 323680 356356 324324
rect 356972 324156 357028 324166
rect 356972 323680 357028 324100
rect 357756 323680 357812 324324
rect 358428 324156 358484 324166
rect 358428 323680 358484 324100
rect 359212 323680 359268 324324
rect 359884 323680 359940 324324
rect 360668 324324 360780 324380
rect 362124 324324 362236 324380
rect 362740 325162 362796 325174
rect 362740 325110 362742 325162
rect 362794 325110 362796 325162
rect 360668 323680 360724 324324
rect 361340 324156 361396 324166
rect 361340 323680 361396 324100
rect 362124 323680 362180 324324
rect 362740 324156 362796 325110
rect 363636 324380 363692 326678
rect 364308 324380 364364 328468
rect 363580 324324 363692 324380
rect 364252 324324 364364 324380
rect 365092 325050 365148 325062
rect 365092 324998 365094 325050
rect 365146 324998 365148 325050
rect 362740 324100 362852 324156
rect 362796 323680 362852 324100
rect 363580 323680 363636 324324
rect 364252 323680 364308 324324
rect 365092 324044 365148 324998
rect 366436 324380 366492 332052
rect 366884 328410 366940 333312
rect 367892 331100 367948 331110
rect 367892 329308 367948 331044
rect 368900 329532 368956 333312
rect 368900 329466 368956 329476
rect 369684 333286 369686 333338
rect 369738 333286 369740 333338
rect 366884 328358 366886 328410
rect 366938 328358 366940 328410
rect 366884 328346 366940 328358
rect 367780 329252 367948 329308
rect 367780 327852 367836 329252
rect 367780 327786 367836 327796
rect 369572 328410 369628 328422
rect 369572 328358 369574 328410
rect 369626 328358 369628 328410
rect 368676 327516 368732 327526
rect 367220 325164 367276 325174
rect 366436 324324 366548 324380
rect 365036 323988 365148 324044
rect 365708 324044 365764 324054
rect 365036 323680 365092 323988
rect 365708 323680 365764 323988
rect 366492 323680 366548 324324
rect 367220 324156 367276 325108
rect 367164 324100 367276 324156
rect 368004 325052 368060 325062
rect 367164 323680 367220 324100
rect 368004 324044 368060 324996
rect 368676 324380 368732 327460
rect 369572 327516 369628 328358
rect 369684 327628 369740 333286
rect 372820 328412 372876 333312
rect 374836 331100 374892 333312
rect 374836 331034 374892 331044
rect 372820 328346 372876 328356
rect 373604 329532 373660 329542
rect 373604 327740 373660 329476
rect 378868 328522 378924 333312
rect 378868 328470 378870 328522
rect 378922 328470 378924 328522
rect 378868 328458 378924 328470
rect 379316 331882 379372 331894
rect 379316 331830 379318 331882
rect 379370 331830 379372 331882
rect 373604 327674 373660 327684
rect 369684 327562 369740 327572
rect 369572 327450 369628 327460
rect 376292 327516 376348 327526
rect 376292 325052 376348 327460
rect 379316 326284 379372 331830
rect 380772 331548 380828 333312
rect 382116 333284 382816 333340
rect 382116 333226 382172 333284
rect 382116 333174 382118 333226
rect 382170 333174 382172 333226
rect 382116 333162 382172 333174
rect 380772 331482 380828 331492
rect 380996 331548 381052 331558
rect 379652 331100 379708 331110
rect 379652 329644 379708 331044
rect 379652 329578 379708 329588
rect 380996 329532 381052 331492
rect 380996 329466 381052 329476
rect 381444 329644 381500 329654
rect 381332 327852 381388 327862
rect 381332 326732 381388 327796
rect 381444 327516 381500 329588
rect 384804 328860 384860 333312
rect 384804 328794 384860 328804
rect 385476 329308 385532 329318
rect 381444 327450 381500 327460
rect 384692 328522 384748 328534
rect 384692 328470 384694 328522
rect 384746 328470 384748 328522
rect 381332 326666 381388 326676
rect 382340 326732 382396 326742
rect 379316 326218 379372 326228
rect 382340 325836 382396 326676
rect 382340 325770 382396 325780
rect 376292 324986 376348 324996
rect 367948 323988 368060 324044
rect 368620 324324 368732 324380
rect 375956 324380 376012 324390
rect 367948 323680 368004 323988
rect 368620 323680 368676 324324
rect 369404 324156 369460 324166
rect 369404 323680 369460 324100
rect 373772 324156 373828 324166
rect 370860 324044 370916 324054
rect 370076 323930 370132 323942
rect 370076 323878 370078 323930
rect 370130 323878 370132 323930
rect 370076 323680 370132 323878
rect 370860 323680 370916 323988
rect 372316 324042 372372 324054
rect 372316 323990 372318 324042
rect 372370 323990 372372 324042
rect 371532 323932 371588 323942
rect 371532 323680 371588 323876
rect 372316 323680 372372 323990
rect 372988 323932 373044 323942
rect 372988 323680 373044 323876
rect 373772 323680 373828 324100
rect 375228 324154 375284 324166
rect 375228 324102 375230 324154
rect 375282 324102 375284 324154
rect 374444 324044 374500 324054
rect 374444 323680 374500 323988
rect 375228 323680 375284 324102
rect 375956 324044 376012 324324
rect 376740 324380 376796 324390
rect 376740 324156 376796 324324
rect 375900 323988 376012 324044
rect 376684 324100 376796 324156
rect 377860 324156 377916 324166
rect 375900 323680 375956 323988
rect 376684 323680 376740 324100
rect 377860 324062 377916 324100
rect 384692 324042 384748 328470
rect 384692 323990 384694 324042
rect 384746 323990 384748 324042
rect 384692 323978 384748 323990
rect 377356 323932 377412 323942
rect 377356 323680 377412 323876
rect 378140 323932 378196 323942
rect 378140 323680 378196 323876
rect 378812 323932 378868 323942
rect 378812 323680 378868 323876
rect 385476 323930 385532 329252
rect 386036 327962 386092 333508
rect 423892 333564 423948 333574
rect 460068 333564 460124 333574
rect 423892 333562 424592 333564
rect 423892 333510 423894 333562
rect 423946 333510 424592 333562
rect 423892 333508 424592 333510
rect 460124 333508 460320 333564
rect 423892 333498 423948 333508
rect 460068 333498 460124 333508
rect 403396 333450 403452 333462
rect 403396 333398 403398 333450
rect 403450 333398 403452 333450
rect 386820 331212 386876 333312
rect 386820 331146 386876 331156
rect 387156 331996 387212 332006
rect 387156 329308 387212 331940
rect 387156 329242 387212 329252
rect 386036 327910 386038 327962
rect 386090 327910 386092 327962
rect 386036 327898 386092 327910
rect 390740 327964 390796 333312
rect 392756 331324 392812 333312
rect 393988 333284 394688 333340
rect 396452 333284 396704 333340
rect 393988 333228 394044 333284
rect 393988 333162 394044 333172
rect 392756 331258 392812 331268
rect 390740 327898 390796 327908
rect 391188 327964 391244 327974
rect 386372 327516 386428 327526
rect 386372 324604 386428 327460
rect 391188 327516 391244 327908
rect 391188 327450 391244 327460
rect 386372 324538 386428 324548
rect 396452 324268 396508 333284
rect 398692 331436 398748 333312
rect 400708 333114 400764 333312
rect 400708 333062 400710 333114
rect 400762 333062 400764 333114
rect 400708 333050 400764 333062
rect 398692 331370 398748 331380
rect 399700 331436 399756 331446
rect 399700 329756 399756 331380
rect 399700 329690 399756 329700
rect 402612 328074 402668 333312
rect 403396 328860 403452 333398
rect 465556 333452 465612 333462
rect 489412 333452 489468 333462
rect 610932 333452 610988 333462
rect 465556 333450 466256 333452
rect 465556 333398 465558 333450
rect 465610 333398 466256 333450
rect 465556 333396 466256 333398
rect 489468 333396 490112 333452
rect 465556 333386 465612 333396
rect 489412 333386 489468 333396
rect 477540 333340 477596 333350
rect 483812 333340 483868 333350
rect 404628 331210 404684 333312
rect 404628 331158 404630 331210
rect 404682 331158 404684 331210
rect 404628 331146 404684 331158
rect 403396 328794 403452 328804
rect 402612 328022 402614 328074
rect 402666 328022 402668 328074
rect 402612 328010 402668 328022
rect 408660 327852 408716 333312
rect 410564 332218 410620 333312
rect 412580 332890 412636 333312
rect 412580 332838 412582 332890
rect 412634 332838 412636 332890
rect 412580 332826 412636 332838
rect 410564 332166 410566 332218
rect 410618 332166 410620 332218
rect 410564 332154 410620 332166
rect 411348 332218 411404 332230
rect 411348 332166 411350 332218
rect 411402 332166 411404 332218
rect 411348 329644 411404 332166
rect 411348 329578 411404 329588
rect 408660 327786 408716 327796
rect 414596 326506 414652 333312
rect 416612 331322 416668 333312
rect 418516 332892 418572 333312
rect 418516 332826 418572 332836
rect 416612 331270 416614 331322
rect 416666 331270 416668 331322
rect 416612 331258 416668 331270
rect 418292 332668 418348 332678
rect 414596 326454 414598 326506
rect 414650 326454 414652 326506
rect 414596 326442 414652 326454
rect 418292 326396 418348 332612
rect 420532 332668 420588 333312
rect 421540 333228 421596 333238
rect 420532 332602 420588 332612
rect 420868 333114 420924 333126
rect 420868 333062 420870 333114
rect 420922 333062 420924 333114
rect 418292 326330 418348 326340
rect 420868 325722 420924 333062
rect 420868 325670 420870 325722
rect 420922 325670 420924 325722
rect 420868 325658 420924 325670
rect 421092 332892 421148 332902
rect 421092 324714 421148 332836
rect 421316 332666 421372 332678
rect 421316 332614 421318 332666
rect 421370 332614 421372 332666
rect 421316 324826 421372 332614
rect 421540 327964 421596 333172
rect 422548 331434 422604 333312
rect 422548 331382 422550 331434
rect 422602 331382 422604 331434
rect 422548 331370 422604 331382
rect 421764 331324 421820 331334
rect 421764 329866 421820 331268
rect 421764 329814 421766 329866
rect 421818 329814 421820 329866
rect 421764 329802 421820 329814
rect 421540 327898 421596 327908
rect 426468 326618 426524 333312
rect 428484 331100 428540 333312
rect 430500 333004 430556 333312
rect 430500 332938 430556 332948
rect 428484 331034 428540 331044
rect 426468 326566 426470 326618
rect 426522 326566 426524 326618
rect 426468 326554 426524 326566
rect 432516 326394 432572 333312
rect 434420 331436 434476 333312
rect 436436 332778 436492 333312
rect 437668 333004 437724 333014
rect 436436 332726 436438 332778
rect 436490 332726 436492 332778
rect 436436 332714 436492 332726
rect 437556 332890 437612 332902
rect 437556 332838 437558 332890
rect 437610 332838 437612 332890
rect 434420 331370 434476 331380
rect 432516 326342 432518 326394
rect 432570 326342 432572 326394
rect 432516 326330 432572 326342
rect 437556 324938 437612 332838
rect 437556 324886 437558 324938
rect 437610 324886 437612 324938
rect 437556 324874 437612 324886
rect 421316 324774 421318 324826
rect 421370 324774 421372 324826
rect 421316 324762 421372 324774
rect 421092 324662 421094 324714
rect 421146 324662 421148 324714
rect 421092 324650 421148 324662
rect 437668 324716 437724 332948
rect 438452 327514 438508 333312
rect 440468 331324 440524 333312
rect 442372 333116 442428 333312
rect 442372 333050 442428 333060
rect 440468 331258 440524 331268
rect 444388 328076 444444 333312
rect 446404 329978 446460 333312
rect 448308 333002 448364 333312
rect 448308 332950 448310 333002
rect 448362 332950 448364 333002
rect 448308 332938 448364 332950
rect 446404 329926 446406 329978
rect 446458 329926 446460 329978
rect 446404 329914 446460 329926
rect 444388 328010 444444 328020
rect 438452 327462 438454 327514
rect 438506 327462 438508 327514
rect 438452 327450 438508 327462
rect 450324 326508 450380 333312
rect 452340 330874 452396 333312
rect 453684 333284 454384 333340
rect 453684 333228 453740 333284
rect 453684 333162 453740 333172
rect 454804 333226 454860 333238
rect 454804 333174 454806 333226
rect 454858 333174 454860 333226
rect 452340 330822 452342 330874
rect 452394 330822 452396 330874
rect 452340 330810 452396 330822
rect 454692 333116 454748 333126
rect 450324 326442 450380 326452
rect 454692 325834 454748 333060
rect 454804 332668 454860 333174
rect 454804 332602 454860 332612
rect 454916 333228 454972 333238
rect 454692 325782 454694 325834
rect 454746 325782 454748 325834
rect 454692 325770 454748 325782
rect 454916 324828 454972 333172
rect 456260 326620 456316 333312
rect 458276 329868 458332 333312
rect 458276 329802 458332 329812
rect 462308 328188 462364 333312
rect 464212 330762 464268 333312
rect 464212 330710 464214 330762
rect 464266 330710 464268 330762
rect 464212 330698 464268 330710
rect 462308 328122 462364 328132
rect 468244 327516 468300 333312
rect 470260 329980 470316 333312
rect 470260 329914 470316 329924
rect 471156 333002 471212 333014
rect 471156 332950 471158 333002
rect 471210 332950 471212 333002
rect 468244 327450 468300 327460
rect 456260 326554 456316 326564
rect 471156 324940 471212 332950
rect 471380 332778 471436 332790
rect 471380 332726 471382 332778
rect 471434 332726 471436 332778
rect 471380 325610 471436 332726
rect 472164 328186 472220 333312
rect 472164 328134 472166 328186
rect 472218 328134 472220 328186
rect 472164 328122 472220 328134
rect 474180 326172 474236 333312
rect 476196 330876 476252 333312
rect 477596 333284 478240 333340
rect 483812 333338 484176 333340
rect 477540 333274 477596 333284
rect 476196 330810 476252 330820
rect 474180 326106 474236 326116
rect 480116 326060 480172 333312
rect 482132 330650 482188 333312
rect 483812 333286 483814 333338
rect 483866 333286 484176 333338
rect 488404 333338 488460 333350
rect 497364 333340 497420 333350
rect 533092 333340 533148 333350
rect 483812 333284 484176 333286
rect 483812 333274 483868 333284
rect 482132 330598 482134 330650
rect 482186 330598 482188 330650
rect 482132 330586 482188 330598
rect 486164 327402 486220 333312
rect 488068 330764 488124 333312
rect 488068 330698 488124 330708
rect 488404 333286 488406 333338
rect 488458 333286 488460 333338
rect 486164 327350 486166 327402
rect 486218 327350 486220 327402
rect 486164 327338 486220 327350
rect 480116 325994 480172 326004
rect 488404 325724 488460 333286
rect 492100 327404 492156 333312
rect 494116 330538 494172 333312
rect 494116 330486 494118 330538
rect 494170 330486 494172 330538
rect 494116 330474 494172 330486
rect 495572 333284 496048 333340
rect 497420 333284 498064 333340
rect 492100 327338 492156 327348
rect 488404 325658 488460 325668
rect 471380 325558 471382 325610
rect 471434 325558 471436 325610
rect 471380 325546 471436 325558
rect 485492 325610 485548 325622
rect 485492 325558 485494 325610
rect 485546 325558 485548 325610
rect 471156 324874 471212 324884
rect 454916 324762 454972 324772
rect 437668 324650 437724 324660
rect 396452 324202 396508 324212
rect 385476 323878 385478 323930
rect 385530 323878 385532 323930
rect 385476 323866 385532 323878
rect 485492 323932 485548 325558
rect 495572 325498 495628 333284
rect 497364 333274 497420 333284
rect 500052 330652 500108 333312
rect 502068 333114 502124 333312
rect 502068 333062 502070 333114
rect 502122 333062 502124 333114
rect 502068 333050 502124 333062
rect 500052 330586 500108 330596
rect 503972 327290 504028 333312
rect 505988 330426 506044 333312
rect 505988 330374 505990 330426
rect 506042 330374 506044 330426
rect 505988 330362 506044 330374
rect 507332 333284 508032 333340
rect 503972 327238 503974 327290
rect 504026 327238 504028 327290
rect 503972 327226 504028 327238
rect 495572 325446 495574 325498
rect 495626 325446 495628 325498
rect 495572 325434 495628 325446
rect 507332 325386 507388 333284
rect 509908 327178 509964 333312
rect 511924 330540 511980 333312
rect 511924 330474 511980 330484
rect 512372 333284 513968 333340
rect 509908 327126 509910 327178
rect 509962 327126 509964 327178
rect 509908 327114 509964 327126
rect 507332 325334 507334 325386
rect 507386 325334 507388 325386
rect 507332 325322 507388 325334
rect 512372 324940 512428 333284
rect 515956 327292 516012 333312
rect 517860 331660 517916 333312
rect 517860 331594 517916 331604
rect 519876 328298 519932 333312
rect 519876 328246 519878 328298
rect 519930 328246 519932 328298
rect 519876 328234 519932 328246
rect 515956 327226 516012 327236
rect 521892 327180 521948 333312
rect 523908 331546 523964 333312
rect 523908 331494 523910 331546
rect 523962 331494 523964 331546
rect 523908 331482 523964 331494
rect 521892 327114 521948 327124
rect 525812 325612 525868 333312
rect 527828 327066 527884 333312
rect 529844 330314 529900 333312
rect 529844 330262 529846 330314
rect 529898 330262 529900 330314
rect 529844 330250 529900 330262
rect 530852 333284 531888 333340
rect 533148 333284 533792 333340
rect 527828 327014 527830 327066
rect 527882 327014 527884 327066
rect 527828 327002 527884 327014
rect 525812 325546 525868 325556
rect 530852 325274 530908 333284
rect 533092 333274 533148 333284
rect 535780 332556 535836 333312
rect 535780 332490 535836 332500
rect 537572 333284 537824 333340
rect 530852 325222 530854 325274
rect 530906 325222 530908 325274
rect 530852 325210 530908 325222
rect 512372 324874 512428 324884
rect 537572 324604 537628 333284
rect 539812 331658 539868 333312
rect 541716 332442 541772 333312
rect 541716 332390 541718 332442
rect 541770 332390 541772 332442
rect 541716 332378 541772 332390
rect 542612 333284 543760 333340
rect 539812 331606 539814 331658
rect 539866 331606 539868 331658
rect 539812 331594 539868 331606
rect 542612 325500 542668 333284
rect 545748 326956 545804 333312
rect 547764 332444 547820 333312
rect 547764 332378 547820 332388
rect 549332 333284 549696 333340
rect 545748 326890 545804 326900
rect 542612 325434 542668 325444
rect 549332 325388 549388 333284
rect 551684 332668 551740 333312
rect 551684 332602 551740 332612
rect 553700 332330 553756 333312
rect 553700 332278 553702 332330
rect 553754 332278 553756 332330
rect 553700 332266 553756 332278
rect 554372 333284 555744 333340
rect 549332 325322 549388 325332
rect 537572 324538 537628 324548
rect 554372 324492 554428 333284
rect 557620 326954 557676 333312
rect 559636 330428 559692 333312
rect 559636 330362 559692 330372
rect 561092 333284 561680 333340
rect 557620 326902 557622 326954
rect 557674 326902 557676 326954
rect 557620 326890 557676 326902
rect 561092 325276 561148 333284
rect 563668 329082 563724 333312
rect 565572 331548 565628 333312
rect 567588 332780 567644 333312
rect 567588 332714 567644 332724
rect 565572 331482 565628 331492
rect 563668 329030 563670 329082
rect 563722 329030 563724 329082
rect 563668 329018 563724 329030
rect 569604 327068 569660 333312
rect 571508 328300 571564 333312
rect 573524 332666 573580 333312
rect 573524 332614 573526 332666
rect 573578 332614 573580 332666
rect 573524 332602 573580 332614
rect 575540 332220 575596 333312
rect 575540 332154 575596 332164
rect 577556 329194 577612 333312
rect 579460 332892 579516 333312
rect 579460 332826 579516 332836
rect 581476 330316 581532 333312
rect 581476 330250 581532 330260
rect 577556 329142 577558 329194
rect 577610 329142 577612 329194
rect 577556 329130 577612 329142
rect 583492 329196 583548 333312
rect 585508 332890 585564 333312
rect 585508 332838 585510 332890
rect 585562 332838 585564 332890
rect 585508 332826 585564 332838
rect 587412 332106 587468 333312
rect 587412 332054 587414 332106
rect 587466 332054 587468 332106
rect 587412 332042 587468 332054
rect 583492 329130 583548 329140
rect 589428 329084 589484 333312
rect 591444 333004 591500 333312
rect 591444 332938 591500 332948
rect 593460 332332 593516 333312
rect 593460 332266 593516 332276
rect 589428 329018 589484 329028
rect 595364 328970 595420 333312
rect 596708 333284 597408 333340
rect 596708 333226 596764 333284
rect 596708 333174 596710 333226
rect 596762 333174 596764 333226
rect 596708 333162 596764 333174
rect 595364 328918 595366 328970
rect 595418 328918 595420 328970
rect 595364 328906 595420 328918
rect 571508 328234 571564 328244
rect 569604 327002 569660 327012
rect 599396 326842 599452 333312
rect 601412 328972 601468 333312
rect 603092 333284 603344 333340
rect 603092 333228 603148 333284
rect 603092 333162 603148 333172
rect 601412 328906 601468 328916
rect 599396 326790 599398 326842
rect 599450 326790 599452 326842
rect 599396 326778 599452 326790
rect 605332 326844 605388 333312
rect 607348 328858 607404 333312
rect 609364 333116 609420 333312
rect 609364 333050 609420 333060
rect 607348 328806 607350 328858
rect 607402 328806 607404 328858
rect 607348 328794 607404 328806
rect 605332 326778 605388 326788
rect 561092 325210 561148 325220
rect 554372 324426 554428 324436
rect 485492 323866 485548 323876
rect 380324 323148 380380 323158
rect 379680 323092 380324 323148
rect 380324 323082 380380 323092
rect 159572 322522 159628 322532
rect 557732 319452 557788 319462
rect 460292 312508 460348 312518
rect 458612 309260 458668 309270
rect 160188 308476 160244 308896
rect 159684 308420 160244 308476
rect 157892 308364 157948 308374
rect 151172 308252 151228 308262
rect 92372 308028 92428 308038
rect 90580 286412 90636 286422
rect 85204 231802 85260 231812
rect 90356 283276 90412 283286
rect 90356 191324 90412 283220
rect 90580 280896 90636 286356
rect 92372 280924 92428 307972
rect 95732 307914 95788 307926
rect 95732 307862 95734 307914
rect 95786 307862 95788 307914
rect 94276 307690 94332 307702
rect 94276 307638 94278 307690
rect 94330 307638 94332 307690
rect 94052 307578 94108 307590
rect 94052 307526 94054 307578
rect 94106 307526 94108 307578
rect 92484 292236 92540 292246
rect 92484 292142 92540 292180
rect 92596 290668 92652 290706
rect 92596 290602 92652 290612
rect 94052 285628 94108 307526
rect 94052 285562 94108 285572
rect 94276 280924 94332 307638
rect 95732 302427 95788 307862
rect 106036 307916 106092 307926
rect 97412 307802 97468 307814
rect 97412 307750 97414 307802
rect 97466 307750 97468 307802
rect 95732 302371 96236 302427
rect 94948 285628 95004 285638
rect 94948 280924 95004 285572
rect 96180 280924 96236 302371
rect 97412 280924 97468 307750
rect 105812 307804 105868 307814
rect 104132 307692 104188 307702
rect 100772 307580 100828 307590
rect 99092 307468 99148 307478
rect 99092 280924 99148 307412
rect 92372 280868 93072 280924
rect 94276 280868 94416 280924
rect 94948 280868 95648 280924
rect 96180 280868 96992 280924
rect 97412 280868 98224 280924
rect 99092 280868 99568 280924
rect 100772 280896 100828 307524
rect 102452 307468 102508 307478
rect 102452 302427 102508 307412
rect 102452 302371 102620 302427
rect 101444 280924 101500 280934
rect 102564 280924 102620 302371
rect 104132 280924 104188 307636
rect 105812 285626 105868 307748
rect 105812 285574 105814 285626
rect 105866 285574 105868 285626
rect 105812 285562 105868 285574
rect 106036 280924 106092 307860
rect 147812 307466 147868 307478
rect 147812 307414 147814 307466
rect 147866 307414 147868 307466
rect 146132 294812 146188 294822
rect 142996 291676 143052 291686
rect 142772 291564 142828 291574
rect 120932 291452 120988 291462
rect 117908 291116 117964 291126
rect 114884 286636 114940 286646
rect 112308 286524 112364 286534
rect 101500 280868 102032 280924
rect 102564 280868 103376 280924
rect 104132 280868 104608 280924
rect 105952 280868 106092 280924
rect 106484 285626 106540 285638
rect 106484 285574 106486 285626
rect 106538 285574 106540 285626
rect 106484 280924 106540 285574
rect 111636 280924 111692 280934
rect 106484 280868 107184 280924
rect 110992 280868 111636 280924
rect 112308 280896 112364 286468
rect 113540 284732 113596 284742
rect 113540 280896 113596 284676
rect 114884 280896 114940 286580
rect 117460 284956 117516 284966
rect 116116 284844 116172 284854
rect 116116 280896 116172 284788
rect 117460 280896 117516 284900
rect 117908 280924 117964 291060
rect 120932 280924 120988 291396
rect 139188 290444 139244 290454
rect 137956 288316 138012 288326
rect 136612 288204 136668 288214
rect 134036 281708 134092 281718
rect 126420 281372 126476 281382
rect 122500 281148 122556 281158
rect 117908 280868 118720 280924
rect 120932 280868 121296 280924
rect 122500 280896 122556 281092
rect 125076 281148 125132 281158
rect 125076 280896 125132 281092
rect 126420 280896 126476 281316
rect 128996 281260 129052 281270
rect 128324 281034 128380 281046
rect 128324 280982 128326 281034
rect 128378 280982 128380 281034
rect 128324 280924 128380 280982
rect 127680 280868 128380 280924
rect 128996 280896 129052 281204
rect 131460 281258 131516 281270
rect 131460 281206 131462 281258
rect 131514 281206 131516 281258
rect 130900 280924 130956 280934
rect 130256 280922 130956 280924
rect 130256 280870 130902 280922
rect 130954 280870 130956 280922
rect 131460 280896 131516 281206
rect 132804 281146 132860 281158
rect 132804 281094 132806 281146
rect 132858 281094 132860 281146
rect 132804 280896 132860 281094
rect 134036 280896 134092 281652
rect 135380 281484 135436 281494
rect 135380 280896 135436 281428
rect 136612 280896 136668 288148
rect 137956 280896 138012 288260
rect 139188 280896 139244 290388
rect 141764 290332 141820 290342
rect 140532 281820 140588 281830
rect 140532 280896 140588 281764
rect 141764 280896 141820 290276
rect 142772 285628 142828 291508
rect 142772 285562 142828 285572
rect 142996 280896 143052 291620
rect 143668 285628 143724 285638
rect 143668 280924 143724 285572
rect 145572 281820 145628 281830
rect 130256 280868 130956 280870
rect 143668 280868 144368 280924
rect 145572 280896 145628 281764
rect 146132 280924 146188 294756
rect 147812 280924 147868 307414
rect 149492 290108 149548 290118
rect 146132 280868 146944 280924
rect 147812 280868 148176 280924
rect 149492 280896 149548 290052
rect 150724 289996 150780 290006
rect 150724 280896 150780 289940
rect 151172 280924 151228 308196
rect 154644 308140 154700 308150
rect 154644 302427 154700 308084
rect 156212 308026 156268 308038
rect 156212 307974 156214 308026
rect 156266 307974 156268 308026
rect 156212 302427 156268 307974
rect 154644 302371 155148 302427
rect 156212 302371 156380 302427
rect 152852 291788 152908 291798
rect 152852 280924 152908 291732
rect 154644 280924 154700 280934
rect 151172 280868 151984 280924
rect 152852 280868 153328 280924
rect 154560 280868 154644 280924
rect 155092 280924 155148 302371
rect 156324 280924 156380 302371
rect 157892 280924 157948 308308
rect 159684 286412 159740 308420
rect 160748 308364 160804 308896
rect 161308 308364 161364 308896
rect 161980 308364 162036 308896
rect 162540 308364 162596 308896
rect 163212 308364 163268 308896
rect 163772 308364 163828 308896
rect 164444 308588 164500 308896
rect 164444 308522 164500 308532
rect 164836 308700 164892 308710
rect 159684 286346 159740 286356
rect 159908 308308 160804 308364
rect 161252 308308 161364 308364
rect 161924 308308 162036 308364
rect 162484 308308 162596 308364
rect 163156 308308 163268 308364
rect 163716 308308 163828 308364
rect 159908 281932 159964 308308
rect 161252 308028 161308 308308
rect 161252 307962 161308 307972
rect 161924 307690 161980 308308
rect 161924 307638 161926 307690
rect 161978 307638 161980 307690
rect 161924 307626 161980 307638
rect 162484 307578 162540 308308
rect 162484 307526 162486 307578
rect 162538 307526 162540 307578
rect 162484 307514 162540 307526
rect 163044 308028 163100 308038
rect 160020 305900 160076 305910
rect 160020 305806 160076 305844
rect 159908 281866 159964 281876
rect 160244 290220 160300 290230
rect 160244 280924 160300 290164
rect 162260 288092 162316 288102
rect 155092 280868 155904 280924
rect 156324 280868 157136 280924
rect 157892 280868 158480 280924
rect 159712 280868 160300 280924
rect 160580 280924 160636 280934
rect 160636 280868 160944 280924
rect 162260 280896 162316 288036
rect 163044 280924 163100 307972
rect 163156 307914 163212 308308
rect 163156 307862 163158 307914
rect 163210 307862 163212 307914
rect 163156 307850 163212 307862
rect 163716 307802 163772 308308
rect 163716 307750 163718 307802
rect 163770 307750 163772 307802
rect 163716 307738 163772 307750
rect 163044 280868 163520 280924
rect 164836 280896 164892 308644
rect 165004 308364 165060 308896
rect 165564 308588 165620 308896
rect 165564 308522 165620 308532
rect 166236 308476 166292 308896
rect 166236 308410 166292 308420
rect 166796 308364 166852 308896
rect 167468 308364 167524 308896
rect 168028 308700 168084 308896
rect 164948 308308 165060 308364
rect 166740 308308 166852 308364
rect 167412 308308 167524 308364
rect 167972 308644 168084 308700
rect 164948 307580 165004 308308
rect 166404 307690 166460 307702
rect 166404 307638 166406 307690
rect 166458 307638 166460 307690
rect 164948 307514 165004 307524
rect 165396 307580 165452 307590
rect 165396 288316 165452 307524
rect 166404 302427 166460 307638
rect 166740 307692 166796 308308
rect 167412 307916 167468 308308
rect 167412 307850 167468 307860
rect 167972 307804 168028 308644
rect 167972 307738 168028 307748
rect 168084 308476 168140 308486
rect 166740 307626 166796 307636
rect 166404 302371 166684 302427
rect 165396 288250 165452 288260
rect 165620 281482 165676 281494
rect 165620 281430 165622 281482
rect 165674 281430 165676 281482
rect 101444 280858 101500 280868
rect 111636 280858 111692 280868
rect 130900 280858 130956 280868
rect 154644 280858 154700 280868
rect 160580 280858 160636 280868
rect 109060 280812 109116 280822
rect 124180 280812 124236 280822
rect 108528 280756 109060 280812
rect 123872 280810 124236 280812
rect 123872 280758 124182 280810
rect 124234 280758 124236 280810
rect 123872 280756 124236 280758
rect 109060 280746 109116 280756
rect 124180 280746 124236 280756
rect 92260 280700 92316 280710
rect 110404 280700 110460 280710
rect 120596 280700 120652 280710
rect 91840 280644 92260 280700
rect 109760 280698 110460 280700
rect 109760 280646 110406 280698
rect 110458 280646 110460 280698
rect 109760 280644 110460 280646
rect 120064 280698 120652 280700
rect 120064 280646 120598 280698
rect 120650 280646 120652 280698
rect 120064 280644 120652 280646
rect 92260 280634 92316 280644
rect 110404 280634 110460 280644
rect 120596 280634 120652 280644
rect 165620 280698 165676 281430
rect 166068 281370 166124 281382
rect 166068 281318 166070 281370
rect 166122 281318 166124 281370
rect 166068 280896 166124 281318
rect 166628 280924 166684 302371
rect 168084 282267 168140 308420
rect 168700 308364 168756 308896
rect 169260 308476 169316 308896
rect 169932 308476 169988 308896
rect 169260 308410 169316 308420
rect 169652 308420 169988 308476
rect 167860 282211 168140 282267
rect 168196 308308 168756 308364
rect 166628 280868 167440 280924
rect 165620 280646 165622 280698
rect 165674 280646 165676 280698
rect 165620 280634 165676 280646
rect 167860 280698 167916 282211
rect 168196 280924 168252 308308
rect 168756 303210 168812 303222
rect 168756 303158 168758 303210
rect 168810 303158 168812 303210
rect 168756 290332 168812 303158
rect 168756 290266 168812 290276
rect 169652 281036 169708 308420
rect 170492 308364 170548 308896
rect 171052 308364 171108 308896
rect 169876 308308 170548 308364
rect 170996 308308 171108 308364
rect 171332 308476 171388 308486
rect 169764 305676 169820 305686
rect 169764 284732 169820 305620
rect 169876 286524 169932 308308
rect 170996 305676 171052 308308
rect 170996 305610 171052 305620
rect 169876 286458 169932 286468
rect 171332 284844 171388 308420
rect 171444 308474 171500 308486
rect 171444 308422 171446 308474
rect 171498 308422 171500 308474
rect 171444 284956 171500 308422
rect 171724 308364 171780 308896
rect 172284 308476 172340 308896
rect 172284 308410 172340 308420
rect 172956 308474 173012 308896
rect 172956 308422 172958 308474
rect 173010 308422 173012 308474
rect 172956 308410 173012 308422
rect 173124 308476 173180 308486
rect 171668 308308 171780 308364
rect 171556 303212 171612 303222
rect 171556 285627 171612 303156
rect 171668 286636 171724 308308
rect 171668 286570 171724 286580
rect 173012 308028 173068 308038
rect 171556 285571 171724 285627
rect 171444 284890 171500 284900
rect 171332 284778 171388 284788
rect 169764 284666 169820 284676
rect 169652 280970 169708 280980
rect 167972 280868 168252 280924
rect 171668 280924 171724 285571
rect 171668 280868 172480 280924
rect 167972 280812 168028 280868
rect 170548 280812 170604 280822
rect 170016 280756 170548 280812
rect 173012 280812 173068 307972
rect 173124 281482 173180 308420
rect 173516 308364 173572 308896
rect 174188 308476 174244 308896
rect 174188 308410 174244 308420
rect 173236 308308 173572 308364
rect 174748 308364 174804 308896
rect 175420 308364 175476 308896
rect 175980 308364 176036 308896
rect 174748 308308 174972 308364
rect 173236 291900 173292 308308
rect 173236 291834 173292 291844
rect 174692 305676 174748 305686
rect 173124 281430 173126 281482
rect 173178 281430 173180 281482
rect 173124 281418 173180 281430
rect 173908 281482 173964 281494
rect 173908 281430 173910 281482
rect 173962 281430 173964 281482
rect 173908 281146 173964 281430
rect 173908 281094 173910 281146
rect 173962 281094 173964 281146
rect 173908 281082 173964 281094
rect 173012 280756 173824 280812
rect 174692 280810 174748 305620
rect 174804 305562 174860 305574
rect 174804 305510 174806 305562
rect 174858 305510 174860 305562
rect 174804 281148 174860 305510
rect 174916 291452 174972 308308
rect 175364 308308 175476 308364
rect 175924 308308 176036 308364
rect 176372 308476 176428 308486
rect 175364 305562 175420 308308
rect 175924 305676 175980 308308
rect 175924 305610 175980 305620
rect 175364 305510 175366 305562
rect 175418 305510 175420 305562
rect 175364 305498 175420 305510
rect 174916 291386 174972 291396
rect 176372 281596 176428 308420
rect 176540 308364 176596 308896
rect 177212 308476 177268 308896
rect 177212 308410 177268 308420
rect 177772 308364 177828 308896
rect 176540 308308 176652 308364
rect 176148 281540 176428 281596
rect 176484 305676 176540 305686
rect 176148 281372 176204 281540
rect 176148 281306 176204 281316
rect 176372 281372 176428 281382
rect 174804 281082 174860 281092
rect 175700 280924 175756 280934
rect 175056 280868 175700 280924
rect 176372 280896 176428 281316
rect 176484 281034 176540 305620
rect 176596 281260 176652 308308
rect 177716 308308 177828 308364
rect 178052 308698 178108 308710
rect 178052 308646 178054 308698
rect 178106 308646 178108 308698
rect 177716 305676 177772 308308
rect 177716 305610 177772 305620
rect 176596 281194 176652 281204
rect 177940 281260 177996 281270
rect 178052 281260 178108 308646
rect 178444 308364 178500 308896
rect 179004 308364 179060 308896
rect 179676 308698 179732 308896
rect 179676 308646 179678 308698
rect 179730 308646 179732 308698
rect 179676 308634 179732 308646
rect 178164 308308 178500 308364
rect 178724 308308 179060 308364
rect 179732 308476 179788 308486
rect 178164 282044 178220 308308
rect 178724 290667 178780 308308
rect 178164 281978 178220 281988
rect 178276 290611 178780 290667
rect 177940 281258 178108 281260
rect 177940 281206 177942 281258
rect 177994 281206 178108 281258
rect 177940 281204 178108 281206
rect 177940 281194 177996 281204
rect 176484 280982 176486 281034
rect 176538 280982 176540 281034
rect 176484 280970 176540 280982
rect 177940 281036 177996 281046
rect 177940 280924 177996 280980
rect 177632 280868 177996 280924
rect 178276 280922 178332 290611
rect 179732 281932 179788 308420
rect 180236 308364 180292 308896
rect 180908 308476 180964 308896
rect 180908 308410 180964 308420
rect 179732 281866 179788 281876
rect 179844 308308 180292 308364
rect 181468 308364 181524 308896
rect 182028 308476 182084 308896
rect 182028 308410 182084 308420
rect 182700 308364 182756 308896
rect 183092 308476 183148 308486
rect 183260 308476 183316 308896
rect 183148 308420 183316 308476
rect 183092 308410 183148 308420
rect 183932 308364 183988 308896
rect 184492 308364 184548 308896
rect 181468 308308 181580 308364
rect 179844 281482 179900 308308
rect 179844 281430 179846 281482
rect 179898 281430 179900 281482
rect 179844 281418 179900 281430
rect 181524 281484 181580 308308
rect 182644 308308 182756 308364
rect 183204 308308 183988 308364
rect 184436 308308 184548 308364
rect 184884 308476 184940 308486
rect 182644 307580 182700 308308
rect 182644 307514 182700 307524
rect 183204 281596 183260 308308
rect 183204 281530 183260 281540
rect 183428 307580 183484 307590
rect 181524 281418 181580 281428
rect 182756 281484 182812 281494
rect 180180 281260 180236 281270
rect 178276 280870 178278 280922
rect 178330 280870 178332 280922
rect 178948 281148 179004 281158
rect 178948 280896 179004 281092
rect 180180 280896 180236 281204
rect 180740 280924 180796 280934
rect 181636 280924 181692 280934
rect 175700 280858 175756 280868
rect 178276 280858 178332 280870
rect 181440 280868 181636 280924
rect 182756 280896 182812 281428
rect 183428 280924 183484 307524
rect 184436 303210 184492 308308
rect 184436 303158 184438 303210
rect 184490 303158 184492 303210
rect 184436 303146 184492 303158
rect 184772 307692 184828 307702
rect 184772 280924 184828 307636
rect 184884 281820 184940 308420
rect 185164 308364 185220 308896
rect 185724 308364 185780 308896
rect 186396 308476 186452 308896
rect 186396 308410 186452 308420
rect 186956 308364 187012 308896
rect 187516 308364 187572 308896
rect 184996 308308 185220 308364
rect 185444 308308 185780 308364
rect 186676 308308 187012 308364
rect 187460 308308 187572 308364
rect 188188 308364 188244 308896
rect 188748 308364 188804 308896
rect 189420 308364 189476 308896
rect 189980 308364 190036 308896
rect 190652 308374 190708 308896
rect 188188 308308 188300 308364
rect 184996 291676 185052 308308
rect 184996 291610 185052 291620
rect 185444 291564 185500 308308
rect 185444 291498 185500 291508
rect 186564 307916 186620 307926
rect 186564 285628 186620 307860
rect 186676 294812 186732 308308
rect 187460 307578 187516 308308
rect 187460 307526 187462 307578
rect 187514 307526 187516 307578
rect 187460 307514 187516 307526
rect 186676 294746 186732 294756
rect 186788 307466 186844 307478
rect 186788 307414 186790 307466
rect 186842 307414 186844 307466
rect 186564 285562 186620 285572
rect 184884 281754 184940 281764
rect 186788 280924 186844 307414
rect 188132 303324 188188 303334
rect 183428 280868 184016 280924
rect 184772 280868 185360 280924
rect 186592 280868 186844 280924
rect 187236 285628 187292 285638
rect 187236 280924 187292 285572
rect 188132 285627 188188 303268
rect 188244 290108 188300 308308
rect 188244 290042 188300 290052
rect 188356 308308 188804 308364
rect 189364 308308 189476 308364
rect 189924 308308 190036 308364
rect 190596 308364 190708 308374
rect 191212 308364 191268 308896
rect 190652 308308 190708 308364
rect 191156 308308 191268 308364
rect 191492 308588 191548 308598
rect 188356 289996 188412 308308
rect 189364 308252 189420 308308
rect 189364 308186 189420 308196
rect 189924 291788 189980 308308
rect 190596 308298 190652 308308
rect 191156 308140 191212 308308
rect 191492 308252 191548 308532
rect 191884 308476 191940 308896
rect 192444 308588 192500 308896
rect 192444 308522 192500 308532
rect 191492 308186 191548 308196
rect 191604 308420 191940 308476
rect 191156 308074 191212 308084
rect 191604 308026 191660 308420
rect 193004 308364 193060 308896
rect 193676 308588 193732 308896
rect 193676 308522 193732 308532
rect 194236 308364 194292 308896
rect 194908 308476 194964 308896
rect 195468 308700 195524 308896
rect 195468 308634 195524 308644
rect 194908 308410 194964 308420
rect 196140 308364 196196 308896
rect 196700 308588 196756 308896
rect 191604 307974 191606 308026
rect 191658 307974 191660 308026
rect 191604 307962 191660 307974
rect 191716 308308 193060 308364
rect 193284 308308 194292 308364
rect 195076 308308 196196 308364
rect 196532 308532 196756 308588
rect 191604 307804 191660 307814
rect 189924 291722 189980 291732
rect 190036 307468 190092 307478
rect 188356 289930 188412 289940
rect 188132 285571 188412 285627
rect 188356 280924 188412 285571
rect 190036 280924 190092 307412
rect 191604 280924 191660 307748
rect 191716 290220 191772 308308
rect 191828 308138 191884 308150
rect 191828 308086 191830 308138
rect 191882 308086 191884 308138
rect 191828 302427 191884 308086
rect 191828 302371 192220 302427
rect 191716 290154 191772 290164
rect 192164 280924 192220 302371
rect 193284 288092 193340 308308
rect 193396 308140 193452 308150
rect 193396 302427 193452 308084
rect 194964 307916 195020 307926
rect 193396 302371 193564 302427
rect 193284 288026 193340 288036
rect 193508 280924 193564 302371
rect 194964 280924 195020 307860
rect 195076 281370 195132 308308
rect 196532 307690 196588 308532
rect 197372 308476 197428 308896
rect 196532 307638 196534 307690
rect 196586 307638 196588 307690
rect 196532 307626 196588 307638
rect 196644 308420 197428 308476
rect 195076 281318 195078 281370
rect 195130 281318 195132 281370
rect 195076 281306 195132 281318
rect 196532 282156 196588 282166
rect 196532 280924 196588 282100
rect 196644 281146 196700 308420
rect 197932 308364 197988 308896
rect 198492 308364 198548 308896
rect 196980 308308 197988 308364
rect 198324 308308 198548 308364
rect 198660 308700 198716 308710
rect 196868 308252 196924 308262
rect 196868 285626 196924 308196
rect 196868 285574 196870 285626
rect 196922 285574 196924 285626
rect 196868 285562 196924 285574
rect 196644 281094 196646 281146
rect 196698 281094 196700 281146
rect 196644 281082 196700 281094
rect 196980 281036 197036 308308
rect 196980 280970 197036 280980
rect 197428 285626 197484 285638
rect 197428 285574 197430 285626
rect 197482 285574 197484 285626
rect 197428 280924 197484 285574
rect 198324 281036 198380 308308
rect 198324 280970 198380 280980
rect 198660 280924 198716 308644
rect 199164 308364 199220 308896
rect 199724 308364 199780 308896
rect 199108 308308 199220 308364
rect 199668 308308 199780 308364
rect 199892 308700 199948 308710
rect 199108 303212 199164 308308
rect 199668 308028 199724 308308
rect 199668 307962 199724 307972
rect 199108 303146 199164 303156
rect 199892 280924 199948 308644
rect 200004 308476 200060 308486
rect 200004 281148 200060 308420
rect 200396 308364 200452 308896
rect 200956 308476 201012 308896
rect 200956 308410 201012 308420
rect 200004 281082 200060 281092
rect 200116 308308 200452 308364
rect 201628 308364 201684 308896
rect 201796 308476 201852 308486
rect 201628 308308 201740 308364
rect 200116 281146 200172 308308
rect 200116 281094 200118 281146
rect 200170 281094 200172 281146
rect 200116 281082 200172 281094
rect 201572 307802 201628 307814
rect 201572 307750 201574 307802
rect 201626 307750 201628 307802
rect 201572 280924 201628 307750
rect 201684 281372 201740 308308
rect 201684 281306 201740 281316
rect 201796 281260 201852 308420
rect 202188 308364 202244 308896
rect 202860 308476 202916 308896
rect 203420 308588 203476 308896
rect 203420 308522 203476 308532
rect 202860 308410 202916 308420
rect 203980 308364 204036 308896
rect 204652 308364 204708 308896
rect 202020 308308 202244 308364
rect 203476 308308 204036 308364
rect 204596 308308 204708 308364
rect 205212 308364 205268 308896
rect 205884 308364 205940 308896
rect 206444 308374 206500 308896
rect 207116 308476 207172 308896
rect 207116 308410 207172 308420
rect 205212 308308 205324 308364
rect 202020 281596 202076 308308
rect 203364 307690 203420 307702
rect 203364 307638 203366 307690
rect 203418 307638 203420 307690
rect 203364 283948 203420 307638
rect 203476 302427 203532 308308
rect 204596 307580 204652 308308
rect 204596 307514 204652 307524
rect 205156 307914 205212 307926
rect 205156 307862 205158 307914
rect 205210 307862 205212 307914
rect 203476 302371 203868 302427
rect 203364 283892 203756 283948
rect 202020 281530 202076 281540
rect 201796 281194 201852 281204
rect 203588 281036 203644 281046
rect 203588 280924 203644 280980
rect 187236 280868 187936 280924
rect 188356 280868 189168 280924
rect 190036 280868 190512 280924
rect 191604 280868 191744 280924
rect 192164 280868 192976 280924
rect 193508 280868 194320 280924
rect 194964 280868 195552 280924
rect 196532 280868 196896 280924
rect 197428 280868 198128 280924
rect 198660 280868 199472 280924
rect 199892 280868 200704 280924
rect 201572 280868 201936 280924
rect 203280 280868 203644 280924
rect 203700 280924 203756 283892
rect 203812 281484 203868 302371
rect 203812 281418 203868 281428
rect 205156 280924 205212 307862
rect 205268 307692 205324 308308
rect 205268 307626 205324 307636
rect 205828 308308 205940 308364
rect 206388 308364 206500 308374
rect 207676 308364 207732 308896
rect 208348 308364 208404 308896
rect 206444 308308 206500 308364
rect 207620 308308 207732 308364
rect 208292 308308 208404 308364
rect 208516 308474 208572 308486
rect 208516 308422 208518 308474
rect 208570 308422 208572 308474
rect 205828 307466 205884 308308
rect 206388 308298 206444 308308
rect 205828 307414 205830 307466
rect 205882 307414 205884 307466
rect 205828 307402 205884 307414
rect 206724 307578 206780 307590
rect 206724 307526 206726 307578
rect 206778 307526 206780 307578
rect 206724 280924 206780 307526
rect 207620 307468 207676 308308
rect 208292 307804 208348 308308
rect 208292 307738 208348 307748
rect 208404 308028 208460 308038
rect 207620 307402 207676 307412
rect 208404 285628 208460 307972
rect 208404 285562 208460 285572
rect 208516 280924 208572 308422
rect 208908 308364 208964 308896
rect 209468 308364 209524 308896
rect 210140 308364 210196 308896
rect 210700 308476 210756 308896
rect 210700 308410 210756 308420
rect 211372 308364 211428 308896
rect 211932 308700 211988 308896
rect 211932 308634 211988 308644
rect 212604 308588 212660 308896
rect 212604 308522 212660 308532
rect 213164 308364 213220 308896
rect 208852 308308 208964 308364
rect 209412 308308 209524 308364
rect 210084 308308 210196 308364
rect 211316 308308 211428 308364
rect 213108 308308 213220 308364
rect 213444 308588 213500 308598
rect 208852 308138 208908 308308
rect 208852 308086 208854 308138
rect 208906 308086 208908 308138
rect 208852 308074 208908 308086
rect 209412 308140 209468 308308
rect 209412 308074 209468 308084
rect 210084 307916 210140 308308
rect 211316 308252 211372 308308
rect 211316 308186 211372 308196
rect 210084 307850 210140 307860
rect 213108 307802 213164 308308
rect 213108 307750 213110 307802
rect 213162 307750 213164 307802
rect 213108 307738 213164 307750
rect 210084 307692 210140 307702
rect 203700 280868 204512 280924
rect 205156 280868 205856 280924
rect 206724 280868 207088 280924
rect 208432 280868 208572 280924
rect 208964 285628 209020 285638
rect 208964 280924 209020 285572
rect 210084 280924 210140 307636
rect 211876 307580 211932 307590
rect 211876 280924 211932 307524
rect 208964 280868 209664 280924
rect 210084 280868 210896 280924
rect 211876 280868 212240 280924
rect 213444 280896 213500 308532
rect 213836 308364 213892 308896
rect 214396 308364 214452 308896
rect 214956 308364 215012 308896
rect 213556 308308 213892 308364
rect 214340 308308 214452 308364
rect 214900 308308 215012 308364
rect 215124 308476 215180 308486
rect 213556 281036 213612 308308
rect 214340 307690 214396 308308
rect 214900 307914 214956 308308
rect 214900 307862 214902 307914
rect 214954 307862 214956 307914
rect 214900 307850 214956 307862
rect 214340 307638 214342 307690
rect 214394 307638 214396 307690
rect 214340 307626 214396 307638
rect 213668 307468 213724 307478
rect 213668 302427 213724 307412
rect 215124 302427 215180 308420
rect 215628 308364 215684 308896
rect 216188 308474 216244 308896
rect 216860 308588 216916 308896
rect 216188 308422 216190 308474
rect 216242 308422 216244 308474
rect 216188 308410 216244 308422
rect 216804 308532 216916 308588
rect 215572 308308 215684 308364
rect 215572 307578 215628 308308
rect 216804 308028 216860 308532
rect 216804 307962 216860 307972
rect 216916 308364 216972 308374
rect 217420 308364 217476 308896
rect 218092 308364 218148 308896
rect 218652 308588 218708 308896
rect 218652 308522 218708 308532
rect 218820 308588 218876 308598
rect 215572 307526 215574 307578
rect 215626 307526 215628 307578
rect 215572 307514 215628 307526
rect 213668 302371 214060 302427
rect 215124 302371 215292 302427
rect 213556 280970 213612 280980
rect 214004 280924 214060 302371
rect 215236 280924 215292 302371
rect 216916 280924 216972 308308
rect 217364 308308 217476 308364
rect 218036 308308 218148 308364
rect 217364 307692 217420 308308
rect 217364 307626 217420 307636
rect 218036 307580 218092 308308
rect 218036 307514 218092 307524
rect 218596 307692 218652 307702
rect 218596 285628 218652 307636
rect 218596 285562 218652 285572
rect 218820 280924 218876 308532
rect 219212 308364 219268 308896
rect 219884 308476 219940 308896
rect 219884 308410 219940 308420
rect 220276 308700 220332 308710
rect 219156 308308 219268 308364
rect 219156 307468 219212 308308
rect 219156 307402 219212 307412
rect 220276 302427 220332 308644
rect 220444 308374 220500 308896
rect 221116 308588 221172 308896
rect 221116 308522 221172 308532
rect 220388 308364 220500 308374
rect 221676 308364 221732 308896
rect 222348 308700 222404 308896
rect 222348 308634 222404 308644
rect 222908 308364 222964 308896
rect 223580 308364 223636 308896
rect 224140 308364 224196 308896
rect 220444 308308 220500 308364
rect 221620 308308 221732 308364
rect 221844 308308 222964 308364
rect 223412 308308 223636 308364
rect 223860 308308 224196 308364
rect 224700 308364 224756 308896
rect 225372 308474 225428 308896
rect 225372 308422 225374 308474
rect 225426 308422 225428 308474
rect 225372 308410 225428 308422
rect 225932 308476 225988 308896
rect 225932 308410 225988 308420
rect 226604 308364 226660 308896
rect 226772 308474 226828 308486
rect 226772 308422 226774 308474
rect 226826 308422 226828 308474
rect 224700 308308 225148 308364
rect 226604 308308 226716 308364
rect 220388 308298 220444 308308
rect 221620 307692 221676 308308
rect 221620 307626 221676 307636
rect 220276 302371 220444 302427
rect 214004 280868 214816 280924
rect 215236 280868 216048 280924
rect 216916 280868 217392 280924
rect 218624 280868 218876 280924
rect 219268 285628 219324 285638
rect 219268 280924 219324 285572
rect 220388 280924 220444 302371
rect 221844 280924 221900 308308
rect 223412 280924 223468 308308
rect 223860 302427 223916 308308
rect 225092 302427 225148 308308
rect 226660 307466 226716 308308
rect 226660 307414 226662 307466
rect 226714 307414 226716 307466
rect 226660 307402 226716 307414
rect 223860 302371 224252 302427
rect 225092 302371 225596 302427
rect 224196 280924 224252 302371
rect 225540 280924 225596 302371
rect 226772 280924 226828 308422
rect 227164 308364 227220 308896
rect 227836 308474 227892 308896
rect 228396 308698 228452 308896
rect 228396 308646 228398 308698
rect 228450 308646 228452 308698
rect 228396 308634 228452 308646
rect 227836 308422 227838 308474
rect 227890 308422 227892 308474
rect 227836 308410 227892 308422
rect 228452 308476 228508 308486
rect 227164 308308 227276 308364
rect 227220 307468 227276 308308
rect 227220 307402 227276 307412
rect 228452 280924 228508 308420
rect 229068 308364 229124 308896
rect 229628 308364 229684 308896
rect 230188 308476 230244 308896
rect 230188 308410 230244 308420
rect 230860 308364 230916 308896
rect 231420 308588 231476 308896
rect 232092 308700 232148 308896
rect 232092 308634 232148 308644
rect 231420 308522 231476 308532
rect 231812 308474 231868 308486
rect 231812 308422 231814 308474
rect 231866 308422 231868 308474
rect 229068 308308 229180 308364
rect 229628 308308 229740 308364
rect 230860 308308 230972 308364
rect 229124 307580 229180 308308
rect 229684 308252 229740 308308
rect 229684 308186 229740 308196
rect 230916 308140 230972 308308
rect 230916 308074 230972 308084
rect 229124 307514 229180 307524
rect 230132 307468 230188 307478
rect 230132 285628 230188 307412
rect 230132 285562 230188 285572
rect 230244 307466 230300 307478
rect 230244 307414 230246 307466
rect 230298 307414 230300 307466
rect 230244 280924 230300 307414
rect 231812 302427 231868 308422
rect 232652 308364 232708 308896
rect 233324 308364 233380 308896
rect 233884 308812 233940 308896
rect 233884 308756 233996 308812
rect 233828 308586 233884 308598
rect 233828 308534 233830 308586
rect 233882 308534 233884 308586
rect 232652 308308 232764 308364
rect 233324 308308 233436 308364
rect 232708 307468 232764 308308
rect 233380 307916 233436 308308
rect 233380 307850 233436 307860
rect 232708 307402 232764 307412
rect 231812 302371 231980 302427
rect 219268 280868 219968 280924
rect 220388 280868 221200 280924
rect 221844 280868 222432 280924
rect 223412 280868 223776 280924
rect 224196 280868 225008 280924
rect 225540 280868 226352 280924
rect 226772 280868 227584 280924
rect 228452 280868 228928 280924
rect 230160 280868 230300 280924
rect 230692 285628 230748 285638
rect 230692 280924 230748 285572
rect 231924 280924 231980 302371
rect 233828 280924 233884 308534
rect 233940 307692 233996 308756
rect 234556 308374 234612 308896
rect 234556 308364 234668 308374
rect 235116 308364 235172 308896
rect 234556 308308 234612 308364
rect 234612 308298 234668 308308
rect 235060 308308 235172 308364
rect 235676 308364 235732 308896
rect 236348 308364 236404 308896
rect 236908 308364 236964 308896
rect 237580 308588 237636 308896
rect 237580 308522 237636 308532
rect 237076 308476 237132 308486
rect 235676 308308 235788 308364
rect 236348 308308 236460 308364
rect 236908 308308 237020 308364
rect 235060 308026 235116 308308
rect 235060 307974 235062 308026
rect 235114 307974 235116 308026
rect 235060 307962 235116 307974
rect 235284 308252 235340 308262
rect 233940 307626 233996 307636
rect 235172 307580 235228 307590
rect 235172 280924 235228 307524
rect 235284 302427 235340 308196
rect 235732 307802 235788 308308
rect 235732 307750 235734 307802
rect 235786 307750 235788 307802
rect 235732 307738 235788 307750
rect 236404 307466 236460 308308
rect 236964 307690 237020 308308
rect 237076 308028 237132 308420
rect 238140 308364 238196 308896
rect 237076 307962 237132 307972
rect 237188 308308 238196 308364
rect 238532 308476 238588 308486
rect 236964 307638 236966 307690
rect 237018 307638 237020 307690
rect 236964 307626 237020 307638
rect 236404 307414 236406 307466
rect 236458 307414 236460 307466
rect 236404 307402 236460 307414
rect 235284 302371 235788 302427
rect 235732 280924 235788 302371
rect 237188 281148 237244 308308
rect 237188 281082 237244 281092
rect 237412 308028 237468 308038
rect 237412 280924 237468 307972
rect 238532 281036 238588 308420
rect 238812 308364 238868 308896
rect 239372 308364 239428 308896
rect 240044 308476 240100 308896
rect 240044 308410 240100 308420
rect 240436 308700 240492 308710
rect 240324 308364 240380 308374
rect 238812 308308 238924 308364
rect 239372 308308 239484 308364
rect 238532 280970 238588 280980
rect 238644 308140 238700 308150
rect 238644 280924 238700 308084
rect 238868 307692 238924 308308
rect 238868 307626 238924 307636
rect 239428 307578 239484 308308
rect 239428 307526 239430 307578
rect 239482 307526 239484 307578
rect 239428 307514 239484 307526
rect 240324 280924 240380 308308
rect 240436 302427 240492 308644
rect 240604 308374 240660 308896
rect 240604 308364 240716 308374
rect 240604 308308 240660 308364
rect 241164 308364 241220 308896
rect 241836 308476 241892 308896
rect 242396 308588 242452 308896
rect 242396 308522 242452 308532
rect 241836 308410 241892 308420
rect 243068 308364 243124 308896
rect 243628 308700 243684 308896
rect 243628 308644 243740 308700
rect 243572 308474 243628 308486
rect 243572 308422 243574 308474
rect 243626 308422 243628 308474
rect 241164 308308 241276 308364
rect 243068 308308 243180 308364
rect 240660 308298 240716 308308
rect 241220 308140 241276 308308
rect 241220 308074 241276 308084
rect 243124 307914 243180 308308
rect 243124 307862 243126 307914
rect 243178 307862 243180 307914
rect 243124 307850 243180 307862
rect 241892 307468 241948 307478
rect 241892 302427 241948 307412
rect 240436 302371 240940 302427
rect 241892 302371 242172 302427
rect 240884 280924 240940 302371
rect 242116 280924 242172 302371
rect 243572 281036 243628 308422
rect 243684 308252 243740 308644
rect 244300 308364 244356 308896
rect 244860 308474 244916 308896
rect 244860 308422 244862 308474
rect 244914 308422 244916 308474
rect 244860 308410 244916 308422
rect 245532 308364 245588 308896
rect 246092 308364 246148 308896
rect 243684 308186 243740 308196
rect 243796 308308 244356 308364
rect 245364 308308 245588 308364
rect 245812 308308 246148 308364
rect 246652 308364 246708 308896
rect 247324 308700 247380 308896
rect 247324 308634 247380 308644
rect 247044 308474 247100 308486
rect 247044 308422 247046 308474
rect 247098 308422 247100 308474
rect 246652 308308 246764 308364
rect 243572 280970 243628 280980
rect 243684 307916 243740 307926
rect 243684 280924 243740 307860
rect 243796 281596 243852 308308
rect 243796 281530 243852 281540
rect 245252 307580 245308 307590
rect 245252 280924 245308 307524
rect 245364 281932 245420 308308
rect 245812 290667 245868 308308
rect 246708 308028 246764 308308
rect 246708 307962 246764 307972
rect 245364 281866 245420 281876
rect 245588 290611 245868 290667
rect 230692 280868 231392 280924
rect 231924 280868 232736 280924
rect 233828 280868 233968 280924
rect 235172 280868 235312 280924
rect 235732 280868 236544 280924
rect 237412 280868 237888 280924
rect 238644 280868 239120 280924
rect 240324 280868 240464 280924
rect 240884 280868 241696 280924
rect 242116 280868 242928 280924
rect 243684 280868 244272 280924
rect 245252 280868 245504 280924
rect 174692 280758 174694 280810
rect 174746 280758 174748 280810
rect 167972 280746 168028 280756
rect 170548 280746 170604 280756
rect 174692 280746 174748 280758
rect 169204 280700 169260 280710
rect 171332 280700 171388 280710
rect 167860 280646 167862 280698
rect 167914 280646 167916 280698
rect 167860 280634 167916 280646
rect 168672 280698 169260 280700
rect 168672 280646 169206 280698
rect 169258 280646 169260 280698
rect 168672 280644 169260 280646
rect 171248 280644 171332 280700
rect 169204 280634 169260 280644
rect 171332 280634 171388 280644
rect 180740 280698 180796 280868
rect 181636 280858 181692 280868
rect 180740 280646 180742 280698
rect 180794 280646 180796 280698
rect 180740 280634 180796 280646
rect 245588 280700 245644 290611
rect 247044 281820 247100 308422
rect 247884 308364 247940 308896
rect 248556 308474 248612 308896
rect 248556 308422 248558 308474
rect 248610 308422 248612 308474
rect 248556 308410 248612 308422
rect 248724 308474 248780 308486
rect 248724 308422 248726 308474
rect 248778 308422 248780 308474
rect 247884 308308 247996 308364
rect 247940 308250 247996 308308
rect 247940 308198 247942 308250
rect 247994 308198 247996 308250
rect 247940 308186 247996 308198
rect 247156 308026 247212 308038
rect 247156 307974 247158 308026
rect 247210 307974 247212 308026
rect 247156 302427 247212 307974
rect 248612 307802 248668 307814
rect 248612 307750 248614 307802
rect 248666 307750 248668 307802
rect 247156 302371 247324 302427
rect 247044 281754 247100 281764
rect 246148 280924 246204 280934
rect 247268 280924 247324 302371
rect 248612 280924 248668 307750
rect 248724 301644 248780 308422
rect 249116 308364 249172 308896
rect 249788 308474 249844 308896
rect 249788 308422 249790 308474
rect 249842 308422 249844 308474
rect 249788 308410 249844 308422
rect 248724 301578 248780 301588
rect 248948 308308 249172 308364
rect 250348 308364 250404 308896
rect 251020 308364 251076 308896
rect 251580 308364 251636 308896
rect 252140 308364 252196 308896
rect 252812 308364 252868 308896
rect 250348 308308 250460 308364
rect 251020 308308 251132 308364
rect 251580 308308 251692 308364
rect 252140 308308 252364 308364
rect 248948 301532 249004 308308
rect 250404 307580 250460 308308
rect 251076 307916 251132 308308
rect 251076 307850 251132 307860
rect 250404 307514 250460 307524
rect 250516 307690 250572 307702
rect 250516 307638 250518 307690
rect 250570 307638 250572 307690
rect 248948 301466 249004 301476
rect 250292 307466 250348 307478
rect 250292 307414 250294 307466
rect 250346 307414 250348 307466
rect 250292 280924 250348 307414
rect 250516 302427 250572 307638
rect 251636 307690 251692 308308
rect 251636 307638 251638 307690
rect 251690 307638 251692 307690
rect 251636 307626 251692 307638
rect 251972 307804 252028 307814
rect 250516 302371 251132 302427
rect 251076 280924 251132 302371
rect 251972 290667 252028 307748
rect 252084 305676 252140 305686
rect 252084 300076 252140 305620
rect 252308 300188 252364 308308
rect 252756 308308 252868 308364
rect 253372 308364 253428 308896
rect 254044 308700 254100 308896
rect 254044 308634 254100 308644
rect 253652 308474 253708 308486
rect 253652 308422 253654 308474
rect 253706 308422 253708 308474
rect 253372 308308 253484 308364
rect 252756 305676 252812 308308
rect 252756 305610 252812 305620
rect 253428 303548 253484 308308
rect 253428 303482 253484 303492
rect 252308 300122 252364 300132
rect 252084 300010 252140 300020
rect 251972 290611 252476 290667
rect 252420 280924 252476 290611
rect 253652 281484 253708 308422
rect 254604 308364 254660 308896
rect 253876 308308 254660 308364
rect 254772 308700 254828 308710
rect 254772 308364 254828 308644
rect 255276 308474 255332 308896
rect 255276 308422 255278 308474
rect 255330 308422 255332 308474
rect 255276 308410 255332 308422
rect 255836 308364 255892 308896
rect 256508 308364 256564 308896
rect 253876 281708 253932 308308
rect 254772 308298 254828 308308
rect 255444 308308 255892 308364
rect 256228 308308 256564 308364
rect 257068 308364 257124 308896
rect 257628 308700 257684 308896
rect 257628 308634 257684 308644
rect 258300 308364 258356 308896
rect 258860 308588 258916 308896
rect 258860 308532 258972 308588
rect 258692 308476 258748 308486
rect 257068 308308 257180 308364
rect 258300 308308 258412 308364
rect 253876 281642 253932 281652
rect 255332 307692 255388 307702
rect 253652 281418 253708 281428
rect 254436 281148 254492 281158
rect 246204 280868 246848 280924
rect 247268 280868 248080 280924
rect 248612 280868 249424 280924
rect 250292 280868 250656 280924
rect 251076 280868 251888 280924
rect 252420 280868 253232 280924
rect 254436 280896 254492 281092
rect 255332 280924 255388 307636
rect 255444 281146 255500 308308
rect 256228 290667 256284 308308
rect 255556 290611 256284 290667
rect 257012 307578 257068 307590
rect 257012 307526 257014 307578
rect 257066 307526 257068 307578
rect 255556 281258 255612 290611
rect 255556 281206 255558 281258
rect 255610 281206 255612 281258
rect 255556 281194 255612 281206
rect 255444 281094 255446 281146
rect 255498 281094 255500 281146
rect 255444 281082 255500 281094
rect 255332 280868 255808 280924
rect 257012 280896 257068 307526
rect 257124 281148 257180 308308
rect 258356 307466 258412 308308
rect 258356 307414 258358 307466
rect 258410 307414 258412 307466
rect 258356 307402 258412 307414
rect 258692 290667 258748 308420
rect 258804 308362 258860 308374
rect 258804 308310 258806 308362
rect 258858 308310 258860 308362
rect 258804 299852 258860 308310
rect 258916 303660 258972 308532
rect 259532 308586 259588 308896
rect 259532 308534 259534 308586
rect 259586 308534 259588 308586
rect 259532 308522 259588 308534
rect 260092 308364 260148 308896
rect 260764 308476 260820 308896
rect 260764 308410 260820 308420
rect 258916 303594 258972 303604
rect 259028 308308 260148 308364
rect 261324 308364 261380 308896
rect 261996 308364 262052 308896
rect 261324 308308 261436 308364
rect 259028 299964 259084 308308
rect 259028 299898 259084 299908
rect 260596 308140 260652 308150
rect 258804 299786 258860 299796
rect 258692 290611 258860 290667
rect 257124 281082 257180 281092
rect 258804 280924 258860 290611
rect 260596 280924 260652 308084
rect 261380 307804 261436 308308
rect 261380 307738 261436 307748
rect 261940 308308 262052 308364
rect 262276 308588 262332 308598
rect 261940 307578 261996 308308
rect 261940 307526 261942 307578
rect 261994 307526 261996 307578
rect 261940 307514 261996 307526
rect 262052 282156 262108 282166
rect 262052 280924 262108 282100
rect 262276 281260 262332 308532
rect 262556 308588 262612 308896
rect 262556 308522 262612 308532
rect 263116 308364 263172 308896
rect 262388 308308 263172 308364
rect 263620 308588 263676 308598
rect 262388 282156 262444 308308
rect 263620 308140 263676 308532
rect 263788 308476 263844 308896
rect 263788 308410 263844 308420
rect 264348 308364 264404 308896
rect 265020 308364 265076 308896
rect 265580 308700 265636 308896
rect 265580 308644 265692 308700
rect 265524 308476 265580 308486
rect 264348 308308 264460 308364
rect 265020 308308 265132 308364
rect 263620 308074 263676 308084
rect 263956 307914 264012 307926
rect 263956 307862 263958 307914
rect 264010 307862 264012 307914
rect 262388 282090 262444 282100
rect 263508 282156 263564 282166
rect 262276 281204 262668 281260
rect 262612 280924 262668 281204
rect 258804 280868 259616 280924
rect 260596 280868 260848 280924
rect 262052 280868 262192 280924
rect 262612 280868 263424 280924
rect 246148 280858 246204 280868
rect 257684 280812 257740 280822
rect 263508 280812 263564 282100
rect 263956 280924 264012 307862
rect 264404 306460 264460 308308
rect 265076 307356 265132 308308
rect 265076 307290 265132 307300
rect 265412 308252 265468 308262
rect 264404 306394 264460 306404
rect 265412 280924 265468 308196
rect 265524 281370 265580 308420
rect 265636 298396 265692 308644
rect 266252 308364 266308 308896
rect 266812 308476 266868 308896
rect 266812 308410 266868 308420
rect 267484 308364 267540 308896
rect 268044 308476 268100 308896
rect 265636 298330 265692 298340
rect 265748 308308 266308 308364
rect 267204 308308 267540 308364
rect 267652 308420 268100 308476
rect 265748 281482 265804 308308
rect 265748 281430 265750 281482
rect 265802 281430 265804 281482
rect 265748 281418 265804 281430
rect 265524 281318 265526 281370
rect 265578 281318 265580 281370
rect 265524 281306 265580 281318
rect 267204 281372 267260 308308
rect 267652 297387 267708 308420
rect 268604 308364 268660 308896
rect 269276 308364 269332 308896
rect 269836 308364 269892 308896
rect 270508 308700 270564 308896
rect 270508 308644 270620 308700
rect 267428 297331 267708 297387
rect 267988 308308 268660 308364
rect 268884 308308 269332 308364
rect 269556 308308 269892 308364
rect 270452 308476 270508 308486
rect 267204 281306 267260 281316
rect 267316 281596 267372 281606
rect 267428 281596 267484 297331
rect 267988 290667 268044 308308
rect 267540 290611 268044 290667
rect 267540 282044 267596 290611
rect 267540 281978 267596 281988
rect 267540 281596 267596 281606
rect 267428 281540 267540 281596
rect 263956 280868 264768 280924
rect 265412 280868 266000 280924
rect 267316 280896 267372 281540
rect 267540 281530 267596 281540
rect 268884 281258 268940 308308
rect 269556 290667 269612 308308
rect 268884 281206 268886 281258
rect 268938 281206 268940 281258
rect 268884 281194 268940 281206
rect 268996 290611 269612 290667
rect 268996 281146 269052 290611
rect 268996 281094 268998 281146
rect 269050 281094 269052 281146
rect 268996 281082 269052 281094
rect 269892 281932 269948 281942
rect 267876 280924 267932 280934
rect 267932 280868 268576 280924
rect 269892 280896 269948 281876
rect 270452 281260 270508 308420
rect 270564 303436 270620 308644
rect 271068 308364 271124 308896
rect 271740 308476 271796 308896
rect 271740 308410 271796 308420
rect 270564 303370 270620 303380
rect 270900 308308 271124 308364
rect 272300 308364 272356 308896
rect 272860 308364 272916 308896
rect 273532 308364 273588 308896
rect 272300 308308 272412 308364
rect 270900 296604 270956 308308
rect 270900 296538 270956 296548
rect 272132 308028 272188 308038
rect 270452 281194 270508 281204
rect 272132 280924 272188 307972
rect 272356 297836 272412 308308
rect 272356 297770 272412 297780
rect 272468 308308 272916 308364
rect 273028 308308 273588 308364
rect 273812 308588 273868 308598
rect 272468 296492 272524 308308
rect 273028 298060 273084 308308
rect 272468 296426 272524 296436
rect 272580 298004 273084 298060
rect 272132 280868 272384 280924
rect 267876 280858 267932 280868
rect 257740 280756 258384 280812
rect 257684 280746 257740 280756
rect 263508 280746 263564 280756
rect 245588 280634 245644 280644
rect 270452 280700 270508 280710
rect 272580 280700 272636 298004
rect 273028 297836 273084 297846
rect 273028 280810 273084 297780
rect 273812 281036 273868 308532
rect 274092 308364 274148 308896
rect 274764 308588 274820 308896
rect 274764 308522 274820 308532
rect 275324 308364 275380 308896
rect 275996 308364 276052 308896
rect 276556 308364 276612 308896
rect 274036 308308 274148 308364
rect 274260 308308 275380 308364
rect 275604 308308 276052 308364
rect 276276 308308 276612 308364
rect 277228 308364 277284 308896
rect 277788 308476 277844 308896
rect 277788 308420 277900 308476
rect 277228 308308 277340 308364
rect 273924 308250 273980 308262
rect 273924 308198 273926 308250
rect 273978 308198 273980 308250
rect 273924 290667 273980 308198
rect 274036 298172 274092 308308
rect 274260 298508 274316 308308
rect 274260 298442 274316 298452
rect 274036 298106 274092 298116
rect 275604 294812 275660 308308
rect 275604 294746 275660 294756
rect 276276 290667 276332 308308
rect 277284 308252 277340 308308
rect 277284 308186 277340 308196
rect 277844 303212 277900 308420
rect 278348 308364 278404 308896
rect 277844 303146 277900 303156
rect 278068 308308 278404 308364
rect 279020 308364 279076 308896
rect 279580 308588 279636 308896
rect 279580 308522 279636 308532
rect 280252 308364 280308 308896
rect 280812 308476 280868 308896
rect 280812 308410 280868 308420
rect 281484 308364 281540 308896
rect 282044 308364 282100 308896
rect 282324 308698 282380 308710
rect 282324 308646 282326 308698
rect 282378 308646 282380 308698
rect 279020 308308 279132 308364
rect 280252 308308 280364 308364
rect 281484 308308 281596 308364
rect 282044 308308 282156 308364
rect 273924 290611 274204 290667
rect 273812 280970 273868 280980
rect 273252 280924 273308 280934
rect 274148 280924 274204 290611
rect 275604 290611 276332 290667
rect 277172 301532 277228 301542
rect 273308 280868 273728 280924
rect 274148 280868 274960 280924
rect 273252 280858 273308 280868
rect 273028 280758 273030 280810
rect 273082 280758 273084 280810
rect 273028 280746 273084 280758
rect 270508 280644 271152 280700
rect 270452 280634 270508 280644
rect 272580 280634 272636 280644
rect 275604 280698 275660 290611
rect 276276 281820 276332 281830
rect 276276 280896 276332 281764
rect 277172 280924 277228 301476
rect 278068 301532 278124 308308
rect 278068 301466 278124 301476
rect 278852 307580 278908 307590
rect 278852 285626 278908 307524
rect 279076 303324 279132 308308
rect 280308 307802 280364 308308
rect 281540 308028 281596 308308
rect 281540 307962 281596 307972
rect 280308 307750 280310 307802
rect 280362 307750 280364 307802
rect 280308 307738 280364 307750
rect 280644 307916 280700 307926
rect 279076 303258 279132 303268
rect 278852 285574 278854 285626
rect 278906 285574 278908 285626
rect 278852 285562 278908 285574
rect 278964 301644 279020 301654
rect 278964 280924 279020 301588
rect 277172 280868 277536 280924
rect 278880 280868 279020 280924
rect 279412 285626 279468 285638
rect 279412 285574 279414 285626
rect 279466 285574 279468 285626
rect 279412 280924 279468 285574
rect 280644 280924 280700 307860
rect 282100 307580 282156 308308
rect 282100 307514 282156 307524
rect 282212 307690 282268 307702
rect 282212 307638 282214 307690
rect 282266 307638 282268 307690
rect 282212 280924 282268 307638
rect 282324 301868 282380 308646
rect 282716 308476 282772 308896
rect 282716 308420 282828 308476
rect 282772 307468 282828 308420
rect 283276 308364 283332 308896
rect 283836 308698 283892 308896
rect 283836 308646 283838 308698
rect 283890 308646 283892 308698
rect 283836 308634 283892 308646
rect 282772 307402 282828 307412
rect 282996 308308 283332 308364
rect 283892 308476 283948 308486
rect 282996 301980 283052 308308
rect 282996 301914 283052 301924
rect 282324 301802 282380 301812
rect 283892 301756 283948 308420
rect 284508 308364 284564 308896
rect 285068 308476 285124 308896
rect 285068 308410 285124 308420
rect 285572 308476 285628 308486
rect 283892 301690 283948 301700
rect 284228 308308 284564 308364
rect 284228 300524 284284 308308
rect 285572 302092 285628 308420
rect 285740 308364 285796 308896
rect 286300 308364 286356 308896
rect 286972 308476 287028 308896
rect 286972 308410 287028 308420
rect 287364 308476 287420 308486
rect 285740 308308 285852 308364
rect 285572 302026 285628 302036
rect 285796 301644 285852 308308
rect 286020 308308 286356 308364
rect 287252 308364 287308 308374
rect 285796 301578 285852 301588
rect 285908 303548 285964 303558
rect 284228 300458 284284 300468
rect 283892 300188 283948 300198
rect 279412 280868 280112 280924
rect 280644 280868 281344 280924
rect 282212 280868 282688 280924
rect 283892 280896 283948 300132
rect 284452 300076 284508 300086
rect 284452 280924 284508 300020
rect 285908 280924 285964 303492
rect 286020 302204 286076 308308
rect 286020 302138 286076 302148
rect 287252 280924 287308 308308
rect 287364 300300 287420 308420
rect 287532 308364 287588 308896
rect 288204 308364 288260 308896
rect 288764 308476 288820 308896
rect 288764 308410 288820 308420
rect 287476 308308 287588 308364
rect 287924 308308 288260 308364
rect 289324 308364 289380 308896
rect 289996 308364 290052 308896
rect 290556 308364 290612 308896
rect 289324 308308 289436 308364
rect 289996 308308 290108 308364
rect 287476 301530 287532 308308
rect 287476 301478 287478 301530
rect 287530 301478 287532 301530
rect 287476 301466 287532 301478
rect 287924 300412 287980 308308
rect 289380 307244 289436 308308
rect 289380 307178 289436 307188
rect 289716 307468 289772 307478
rect 287924 300346 287980 300356
rect 287364 300234 287420 300244
rect 289044 281708 289100 281718
rect 284452 280868 285264 280924
rect 285908 280868 286496 280924
rect 287252 280868 287840 280924
rect 289044 280896 289100 281652
rect 289716 280810 289772 307412
rect 290052 307132 290108 308308
rect 290052 307066 290108 307076
rect 290500 308308 290612 308364
rect 291228 308364 291284 308896
rect 291788 308364 291844 308896
rect 292292 308476 292348 308486
rect 291228 308308 291340 308364
rect 291788 308308 291900 308364
rect 290500 307020 290556 308308
rect 290500 306954 290556 306964
rect 291284 307018 291340 308308
rect 291284 306966 291286 307018
rect 291338 306966 291340 307018
rect 291284 306954 291340 306966
rect 291844 306906 291900 308308
rect 291844 306854 291846 306906
rect 291898 306854 291900 306906
rect 291844 306842 291900 306854
rect 292292 300636 292348 308420
rect 292460 308364 292516 308896
rect 293020 308364 293076 308896
rect 293692 308476 293748 308896
rect 293692 308410 293748 308420
rect 293972 308700 294028 308710
rect 292460 308308 292572 308364
rect 293020 308308 293132 308364
rect 292516 308026 292572 308308
rect 292516 307974 292518 308026
rect 292570 307974 292572 308026
rect 292516 307962 292572 307974
rect 293076 307692 293132 308308
rect 293076 307626 293132 307636
rect 292292 300570 292348 300580
rect 293972 290667 294028 308644
rect 294084 308476 294140 308486
rect 294252 308476 294308 308896
rect 294252 308420 294364 308476
rect 294084 298284 294140 308420
rect 294308 303548 294364 308420
rect 294812 308364 294868 308896
rect 295484 308476 295540 308896
rect 295484 308410 295540 308420
rect 296044 308364 296100 308896
rect 296716 308588 296772 308896
rect 296716 308522 296772 308532
rect 297276 308364 297332 308896
rect 297948 308364 298004 308896
rect 298508 308364 298564 308896
rect 299180 308364 299236 308896
rect 299740 308364 299796 308896
rect 300300 308364 300356 308896
rect 294308 303482 294364 303492
rect 294532 308308 294868 308364
rect 295764 308308 296100 308364
rect 296212 308308 297332 308364
rect 297444 308308 298004 308364
rect 298228 308308 298564 308364
rect 299012 308308 299236 308364
rect 299460 308308 299796 308364
rect 300244 308308 300356 308364
rect 300804 308476 300860 308486
rect 294532 300636 294588 308308
rect 294532 300570 294588 300580
rect 295764 299628 295820 308308
rect 296212 307692 296268 308308
rect 295876 307636 296268 307692
rect 295876 301642 295932 307636
rect 295876 301590 295878 301642
rect 295930 301590 295932 301642
rect 295876 301578 295932 301590
rect 295988 307466 296044 307478
rect 295988 307414 295990 307466
rect 296042 307414 296044 307466
rect 295764 299562 295820 299572
rect 294084 298218 294140 298228
rect 293972 290611 294700 290667
rect 290388 281484 290444 281494
rect 290388 280896 290444 281428
rect 294196 281148 294252 281158
rect 291172 281034 291228 281046
rect 291172 280982 291174 281034
rect 291226 280982 291228 281034
rect 291172 280924 291228 280982
rect 292292 280924 292348 280934
rect 291172 280868 291648 280924
rect 292292 280922 292880 280924
rect 292292 280870 292294 280922
rect 292346 280870 292880 280922
rect 294196 280896 294252 281092
rect 294644 280924 294700 290611
rect 295988 280924 296044 307414
rect 297332 303660 297388 303670
rect 297332 280924 297388 303604
rect 297444 301754 297500 308308
rect 298228 302314 298284 308308
rect 298228 302262 298230 302314
rect 298282 302262 298284 302314
rect 298228 302250 298284 302262
rect 297444 301702 297446 301754
rect 297498 301702 297500 301754
rect 297444 301690 297500 301702
rect 299012 300636 299068 308308
rect 299012 300570 299068 300580
rect 299236 305676 299292 305686
rect 299236 300298 299292 305620
rect 299460 300522 299516 308308
rect 300244 305676 300300 308308
rect 300244 305610 300300 305620
rect 299460 300470 299462 300522
rect 299514 300470 299516 300522
rect 299460 300458 299516 300470
rect 300692 303772 300748 303782
rect 299236 300246 299238 300298
rect 299290 300246 299292 300298
rect 299236 300234 299292 300246
rect 299796 299964 299852 299974
rect 299012 299852 299068 299862
rect 299012 280924 299068 299796
rect 299796 280924 299852 299908
rect 300692 290667 300748 303716
rect 300804 300186 300860 308420
rect 300972 308364 301028 308896
rect 301532 308476 301588 308896
rect 302204 308588 302260 308896
rect 302204 308522 302260 308532
rect 301532 308410 301588 308420
rect 302596 308476 302652 308486
rect 300972 308308 301084 308364
rect 301028 300410 301084 308308
rect 301700 308028 301756 308038
rect 301028 300358 301030 300410
rect 301082 300358 301084 300410
rect 301028 300346 301084 300358
rect 301476 307580 301532 307590
rect 300804 300134 300806 300186
rect 300858 300134 300860 300186
rect 300804 300122 300860 300134
rect 300692 290611 301084 290667
rect 301028 280924 301084 290611
rect 301476 281484 301532 307524
rect 301700 281706 301756 307972
rect 301700 281654 301702 281706
rect 301754 281654 301756 281706
rect 301700 281642 301756 281654
rect 302372 307916 302428 307926
rect 301476 281418 301532 281428
rect 302372 280924 302428 307860
rect 302596 300636 302652 308420
rect 302764 308364 302820 308896
rect 303436 308364 303492 308896
rect 303996 308476 304052 308896
rect 303996 308410 304052 308420
rect 304164 308476 304220 308486
rect 302764 308308 302876 308364
rect 302596 300570 302652 300580
rect 302708 305676 302764 305686
rect 302708 300076 302764 305620
rect 302820 300636 302876 308308
rect 303380 308308 303492 308364
rect 303380 305676 303436 308308
rect 303380 305610 303436 305620
rect 304052 307578 304108 307590
rect 304052 307526 304054 307578
rect 304106 307526 304108 307578
rect 302820 300570 302876 300580
rect 302708 300010 302764 300020
rect 304052 280924 304108 307526
rect 304164 300074 304220 308420
rect 304668 308364 304724 308896
rect 305228 308476 305284 308896
rect 305228 308410 305284 308420
rect 304164 300022 304166 300074
rect 304218 300022 304220 300074
rect 304164 300010 304220 300022
rect 304276 308308 304724 308364
rect 305788 308364 305844 308896
rect 306460 308364 306516 308896
rect 307020 308700 307076 308896
rect 307020 308634 307076 308644
rect 307524 308476 307580 308486
rect 305788 308308 305900 308364
rect 306460 308308 306572 308364
rect 304276 299964 304332 308308
rect 304276 299898 304332 299908
rect 305732 308140 305788 308150
rect 292292 280868 292880 280870
rect 294644 280868 295456 280924
rect 295988 280868 296800 280924
rect 297332 280868 298032 280924
rect 299012 280868 299376 280924
rect 299796 280868 300608 280924
rect 301028 280868 301840 280924
rect 302372 280868 303184 280924
rect 304052 280868 304416 280924
rect 305732 280896 305788 308084
rect 305844 296716 305900 308308
rect 306516 307580 306572 308308
rect 306516 307514 306572 307524
rect 305844 296650 305900 296660
rect 307524 281034 307580 308420
rect 307692 308364 307748 308896
rect 308252 308476 308308 308896
rect 308924 308588 308980 308896
rect 309484 308700 309540 308896
rect 309484 308634 309540 308644
rect 308924 308522 308980 308532
rect 308252 308410 308308 308420
rect 309204 308476 309260 308486
rect 307636 308308 307748 308364
rect 308084 308364 308140 308374
rect 307636 299852 307692 308308
rect 307636 299786 307692 299796
rect 307860 307468 307916 307478
rect 307524 280982 307526 281034
rect 307578 280982 307580 281034
rect 307524 280970 307580 280982
rect 307860 280924 307916 307412
rect 308084 302427 308140 308308
rect 309092 306460 309148 306470
rect 308084 302371 308252 302427
rect 308196 281708 308252 302371
rect 308196 281642 308252 281652
rect 309092 280924 309148 306404
rect 309204 296828 309260 308420
rect 310156 308374 310212 308896
rect 310716 308476 310772 308896
rect 310716 308410 310772 308420
rect 310884 308476 310940 308486
rect 310156 308364 310268 308374
rect 310156 308308 310212 308364
rect 310212 308298 310268 308308
rect 309204 296762 309260 296772
rect 310772 307356 310828 307366
rect 307860 280868 308336 280924
rect 309092 280868 309568 280924
rect 310772 280896 310828 307300
rect 310884 299962 310940 308420
rect 311276 308364 311332 308896
rect 311948 308476 312004 308896
rect 311948 308410 312004 308420
rect 312508 308476 312564 308896
rect 313180 308588 313236 308896
rect 313180 308522 313236 308532
rect 312508 308410 312564 308420
rect 313740 308364 313796 308896
rect 310884 299910 310886 299962
rect 310938 299910 310940 299962
rect 310884 299898 310940 299910
rect 310996 308308 311332 308364
rect 312676 308308 313796 308364
rect 313908 308588 313964 308598
rect 310996 297276 311052 308308
rect 310996 297210 311052 297220
rect 311332 298396 311388 298406
rect 311332 280924 311388 298340
rect 311332 280868 312144 280924
rect 312676 280922 312732 308308
rect 313908 308140 313964 308532
rect 313908 308074 313964 308084
rect 314244 308476 314300 308486
rect 314244 298396 314300 308420
rect 314412 308364 314468 308896
rect 314972 308364 315028 308896
rect 315644 308476 315700 308896
rect 315644 308410 315700 308420
rect 315924 308698 315980 308710
rect 315924 308646 315926 308698
rect 315978 308646 315980 308698
rect 314412 308308 314524 308364
rect 314972 308308 315084 308364
rect 314244 298330 314300 298340
rect 312676 280870 312678 280922
rect 312730 280870 312732 280922
rect 313348 281482 313404 281494
rect 313348 281430 313350 281482
rect 313402 281430 313404 281482
rect 313348 280896 313404 281430
rect 314468 281148 314524 308308
rect 315028 308028 315084 308308
rect 315028 307962 315084 307972
rect 315924 291676 315980 308646
rect 316204 308588 316260 308896
rect 316204 308522 316260 308532
rect 316764 308364 316820 308896
rect 317436 308698 317492 308896
rect 317436 308646 317438 308698
rect 317490 308646 317492 308698
rect 317436 308634 317492 308646
rect 316036 308308 316820 308364
rect 317492 308476 317548 308486
rect 316036 291900 316092 308308
rect 316036 291834 316092 291844
rect 316596 307802 316652 307814
rect 316596 307750 316598 307802
rect 316650 307750 316652 307802
rect 315924 291610 315980 291620
rect 316596 281820 316652 307750
rect 317492 291564 317548 308420
rect 317996 308364 318052 308896
rect 318668 308476 318724 308896
rect 318668 308410 318724 308420
rect 317716 308308 318052 308364
rect 319228 308364 319284 308896
rect 319900 308476 319956 308896
rect 320460 308588 320516 308896
rect 320460 308522 320516 308532
rect 320964 308588 321020 308598
rect 319900 308410 319956 308420
rect 319228 308308 319340 308364
rect 317716 291788 317772 308308
rect 319284 307914 319340 308308
rect 319284 307862 319286 307914
rect 319338 307862 319340 307914
rect 319284 307850 319340 307862
rect 319956 307580 320012 307590
rect 319956 302427 320012 307524
rect 320852 303436 320908 303446
rect 319956 302371 320124 302427
rect 317716 291722 317772 291732
rect 318276 298508 318332 298518
rect 317492 291498 317548 291508
rect 316596 281754 316652 281764
rect 317268 281596 317324 281606
rect 314468 281082 314524 281092
rect 314692 281370 314748 281382
rect 314692 281318 314694 281370
rect 314746 281318 314748 281370
rect 314692 280896 314748 281318
rect 315924 281372 315980 281382
rect 315924 280896 315980 281316
rect 317268 280896 317324 281540
rect 318276 281372 318332 298452
rect 318276 281306 318332 281316
rect 319844 281258 319900 281270
rect 319844 281206 319846 281258
rect 319898 281206 319900 281258
rect 317828 281036 317884 281046
rect 317828 280924 317884 280980
rect 292292 280858 292348 280868
rect 312676 280858 312732 280870
rect 317828 280868 318528 280924
rect 319844 280896 319900 281206
rect 320068 281258 320124 302371
rect 320852 290667 320908 303380
rect 320964 292236 321020 308532
rect 321132 308364 321188 308896
rect 321692 308588 321748 308896
rect 321692 308522 321748 308532
rect 322252 308364 322308 308896
rect 322924 308476 322980 308896
rect 322924 308420 323036 308476
rect 321132 308308 321244 308364
rect 320964 292170 321020 292180
rect 321188 292236 321244 308308
rect 321188 292170 321244 292180
rect 321412 308308 322308 308364
rect 321412 292236 321468 308308
rect 322980 307580 323036 308420
rect 323484 308364 323540 308896
rect 324156 308700 324212 308896
rect 322980 307514 323036 307524
rect 323092 308308 323540 308364
rect 324100 308644 324212 308700
rect 323092 305788 323148 308308
rect 321412 292170 321468 292180
rect 322532 305732 323148 305788
rect 322532 291786 322588 305732
rect 322532 291734 322534 291786
rect 322586 291734 322588 291786
rect 322532 291722 322588 291734
rect 322868 296604 322924 296614
rect 320852 290611 321580 290667
rect 320068 281206 320070 281258
rect 320122 281206 320124 281258
rect 320068 281194 320124 281206
rect 321076 281146 321132 281158
rect 321076 281094 321078 281146
rect 321130 281094 321132 281146
rect 321076 280896 321132 281094
rect 321524 280924 321580 290611
rect 322868 280924 322924 296548
rect 324100 291674 324156 308644
rect 324100 291622 324102 291674
rect 324154 291622 324156 291674
rect 324100 291610 324156 291622
rect 324212 308476 324268 308486
rect 324212 285404 324268 308420
rect 324716 308364 324772 308896
rect 325388 308476 325444 308896
rect 325948 308476 326004 308896
rect 326508 308586 326564 308896
rect 326508 308534 326510 308586
rect 326562 308534 326564 308586
rect 326508 308522 326564 308534
rect 325948 308420 326060 308476
rect 325388 308410 325444 308420
rect 324436 308308 324772 308364
rect 324436 285516 324492 308308
rect 326004 307916 326060 308420
rect 327180 308364 327236 308896
rect 326004 307850 326060 307860
rect 326340 308308 327236 308364
rect 327460 308586 327516 308598
rect 327460 308534 327462 308586
rect 327514 308534 327516 308586
rect 326340 290667 326396 308308
rect 327460 307802 327516 308534
rect 327740 308364 327796 308896
rect 328412 308364 328468 308896
rect 328972 308364 329028 308896
rect 327740 308308 327852 308364
rect 327460 307750 327462 307802
rect 327514 307750 327516 307802
rect 327460 307738 327516 307750
rect 327684 305676 327740 305686
rect 324436 285450 324492 285460
rect 325892 290611 326396 290667
rect 326676 296492 326732 296502
rect 324212 285338 324268 285348
rect 325892 284844 325948 290611
rect 325892 284778 325948 284788
rect 324884 281260 324940 281270
rect 321524 280868 322336 280924
rect 322868 280868 323680 280924
rect 324884 280896 324940 281204
rect 326676 280924 326732 296436
rect 327684 284956 327740 305620
rect 327796 285068 327852 308308
rect 327908 308308 328468 308364
rect 328916 308308 329028 308364
rect 329364 308476 329420 308486
rect 327908 285292 327964 308308
rect 328916 305676 328972 308308
rect 328916 305610 328972 305620
rect 327908 285226 327964 285236
rect 327796 285002 327852 285012
rect 327684 284890 327740 284900
rect 329364 284954 329420 308420
rect 329644 308364 329700 308896
rect 329588 308308 329700 308364
rect 330204 308374 330260 308896
rect 330876 308476 330932 308896
rect 330876 308410 330932 308420
rect 331044 308476 331100 308486
rect 330204 308364 330316 308374
rect 330204 308308 330260 308364
rect 329364 284902 329366 284954
rect 329418 284902 329420 284954
rect 329364 284890 329420 284902
rect 329476 298172 329532 298182
rect 329476 280924 329532 298116
rect 329588 284956 329644 308308
rect 330260 308298 330316 308308
rect 331044 285066 331100 308420
rect 331436 308364 331492 308896
rect 331996 308476 332052 308896
rect 331996 308410 332052 308420
rect 332668 308476 332724 308896
rect 332668 308410 332724 308420
rect 333228 308364 333284 308896
rect 333900 308364 333956 308896
rect 331044 285014 331046 285066
rect 331098 285014 331100 285066
rect 331044 285002 331100 285014
rect 331380 308308 331492 308364
rect 332836 308308 333284 308364
rect 333620 308308 333956 308364
rect 334460 308364 334516 308896
rect 335132 308364 335188 308896
rect 334460 308308 334572 308364
rect 329588 284890 329644 284900
rect 331380 282154 331436 308308
rect 332724 294812 332780 294822
rect 332724 283948 332780 294756
rect 332836 284842 332892 308308
rect 333620 290667 333676 308308
rect 334516 291562 334572 308308
rect 334516 291510 334518 291562
rect 334570 291510 334572 291562
rect 334516 291498 334572 291510
rect 334628 308308 335188 308364
rect 335692 308364 335748 308896
rect 336084 308474 336140 308486
rect 336084 308422 336086 308474
rect 336138 308422 336140 308474
rect 335692 308308 335804 308364
rect 334628 291450 334684 308308
rect 335748 307804 335804 308308
rect 335748 307738 335804 307748
rect 335860 302316 335916 302326
rect 335860 302222 335916 302260
rect 334628 291398 334630 291450
rect 334682 291398 334684 291450
rect 334628 291386 334684 291398
rect 335076 301754 335132 301766
rect 335076 301702 335078 301754
rect 335130 301702 335132 301754
rect 332836 284790 332838 284842
rect 332890 284790 332892 284842
rect 332836 284778 332892 284790
rect 332948 290611 333676 290667
rect 332948 284730 333004 290611
rect 332948 284678 332950 284730
rect 333002 284678 333004 284730
rect 332948 284666 333004 284678
rect 332724 283892 333116 283948
rect 331380 282102 331382 282154
rect 331434 282102 331436 282154
rect 331380 282090 331436 282102
rect 332164 282154 332220 282166
rect 332164 282102 332166 282154
rect 332218 282102 332220 282154
rect 331940 281146 331996 281158
rect 331940 281094 331942 281146
rect 331994 281094 331996 281146
rect 330932 280924 330988 280934
rect 326676 280868 327488 280924
rect 329476 280868 330064 280924
rect 330988 280868 331296 280924
rect 330932 280858 330988 280868
rect 289716 280758 289718 280810
rect 289770 280758 289772 280810
rect 289716 280746 289772 280758
rect 306404 280812 306460 280822
rect 306460 280756 306992 280812
rect 306404 280746 306460 280756
rect 275604 280646 275606 280698
rect 275658 280646 275660 280698
rect 275604 280634 275660 280646
rect 325892 280700 325948 280710
rect 328132 280700 328188 280710
rect 325892 280698 326256 280700
rect 325892 280646 325894 280698
rect 325946 280646 326256 280698
rect 325892 280644 326256 280646
rect 328188 280644 328832 280700
rect 331940 280698 331996 281094
rect 331940 280646 331942 280698
rect 331994 280646 331996 280698
rect 325892 280634 325948 280644
rect 328132 280634 328188 280644
rect 331940 280634 331996 280646
rect 332164 280698 332220 282102
rect 332612 281372 332668 281382
rect 332612 280896 332668 281316
rect 333060 280924 333116 283892
rect 334404 282156 334460 282166
rect 334404 281370 334460 282100
rect 334628 282156 334684 282166
rect 334628 281482 334684 282100
rect 335076 281594 335132 301702
rect 335300 301642 335356 301654
rect 335300 301590 335302 301642
rect 335354 301590 335356 301642
rect 335300 281818 335356 301590
rect 335748 301532 335804 301542
rect 335412 300524 335468 300534
rect 335412 282044 335468 300468
rect 335412 281978 335468 281988
rect 335524 298396 335580 298406
rect 335300 281766 335302 281818
rect 335354 281766 335356 281818
rect 335300 281754 335356 281766
rect 335076 281542 335078 281594
rect 335130 281542 335132 281594
rect 335076 281530 335132 281542
rect 334628 281430 334630 281482
rect 334682 281430 334684 281482
rect 334628 281418 334684 281430
rect 334404 281318 334406 281370
rect 334458 281318 334460 281370
rect 334404 281306 334460 281318
rect 335188 281146 335244 281158
rect 335188 281094 335190 281146
rect 335242 281094 335244 281146
rect 333060 280868 333872 280924
rect 335188 280896 335244 281094
rect 335524 281146 335580 298340
rect 335748 281372 335804 301476
rect 336084 293132 336140 308422
rect 336364 308476 336420 308896
rect 336364 308410 336420 308420
rect 336924 308474 336980 308896
rect 336924 308422 336926 308474
rect 336978 308422 336980 308474
rect 336924 308410 336980 308422
rect 337092 308700 337148 308710
rect 336084 293066 336140 293076
rect 336420 308252 336476 308262
rect 337092 308252 337148 308644
rect 337484 308364 337540 308896
rect 337764 308474 337820 308486
rect 337764 308422 337766 308474
rect 337818 308422 337820 308474
rect 337484 308308 337596 308364
rect 335748 281306 335804 281316
rect 335524 281094 335526 281146
rect 335578 281094 335580 281146
rect 335524 281082 335580 281094
rect 336420 280896 336476 308196
rect 336980 308196 337148 308252
rect 336644 307692 336700 307702
rect 336644 299740 336700 307636
rect 336644 299674 336700 299684
rect 336756 307580 336812 307590
rect 336756 289996 336812 307524
rect 336868 305898 336924 305910
rect 336868 305846 336870 305898
rect 336922 305846 336924 305898
rect 336868 301532 336924 305846
rect 336868 301466 336924 301476
rect 336980 295036 337036 308196
rect 337540 307690 337596 308308
rect 337540 307638 337542 307690
rect 337594 307638 337596 307690
rect 337540 307626 337596 307638
rect 337204 307468 337260 307478
rect 337092 306908 337148 306918
rect 337092 301644 337148 306852
rect 337092 301578 337148 301588
rect 336980 294970 337036 294980
rect 337204 294924 337260 307412
rect 337204 294858 337260 294868
rect 337652 303212 337708 303222
rect 336756 289930 336812 289940
rect 337540 294026 337596 294038
rect 337540 293974 337542 294026
rect 337594 293974 337596 294026
rect 337540 289212 337596 293974
rect 337540 289146 337596 289156
rect 337652 280924 337708 303156
rect 337764 288092 337820 308422
rect 338156 308364 338212 308896
rect 338716 308474 338772 308896
rect 338716 308422 338718 308474
rect 338770 308422 338772 308474
rect 338716 308410 338772 308422
rect 337988 308308 338212 308364
rect 339388 308364 339444 308896
rect 339948 308364 340004 308896
rect 340620 308364 340676 308896
rect 341180 308700 341236 308896
rect 341180 308634 341236 308644
rect 341852 308364 341908 308896
rect 342412 308364 342468 308896
rect 342972 308364 343028 308896
rect 343644 308700 343700 308896
rect 343644 308634 343700 308644
rect 344204 308364 344260 308896
rect 344876 308364 344932 308896
rect 345436 308364 345492 308896
rect 346108 308364 346164 308896
rect 346668 308364 346724 308896
rect 347340 308364 347396 308896
rect 347900 308364 347956 308896
rect 348460 308364 348516 308896
rect 349132 308364 349188 308896
rect 349692 308364 349748 308896
rect 350364 308364 350420 308896
rect 350924 308364 350980 308896
rect 351596 308364 351652 308896
rect 352156 308364 352212 308896
rect 352828 308364 352884 308896
rect 353388 308364 353444 308896
rect 353948 308364 354004 308896
rect 354620 308364 354676 308896
rect 355180 308364 355236 308896
rect 355852 308364 355908 308896
rect 356412 308700 356468 308896
rect 356412 308634 356468 308644
rect 357084 308364 357140 308896
rect 357644 308364 357700 308896
rect 358316 308364 358372 308896
rect 358876 308364 358932 308896
rect 359436 308364 359492 308896
rect 339388 308308 339500 308364
rect 339948 308308 340060 308364
rect 340620 308308 340732 308364
rect 341852 308308 341964 308364
rect 342412 308308 342524 308364
rect 342972 308308 343084 308364
rect 344204 308308 344316 308364
rect 344876 308308 344988 308364
rect 345436 308308 345548 308364
rect 346108 308308 346220 308364
rect 346668 308308 346780 308364
rect 347340 308308 347452 308364
rect 347900 308308 348012 308364
rect 348460 308308 348572 308364
rect 349132 308308 349244 308364
rect 349692 308308 349804 308364
rect 350364 308308 350476 308364
rect 350924 308308 351036 308364
rect 351596 308308 351708 308364
rect 352156 308308 352268 308364
rect 352828 308308 352940 308364
rect 353388 308308 353500 308364
rect 353948 308308 354060 308364
rect 354620 308308 354732 308364
rect 355180 308308 355292 308364
rect 355852 308308 355964 308364
rect 357084 308308 357196 308364
rect 357644 308308 357756 308364
rect 358316 308308 358428 308364
rect 358876 308308 358988 308364
rect 337988 288316 338044 308308
rect 337988 288250 338044 288260
rect 339332 303324 339388 303334
rect 337764 288026 337820 288036
rect 338996 281372 339052 281382
rect 337652 280868 337792 280924
rect 338996 280896 339052 281316
rect 339332 281260 339388 303268
rect 339444 288204 339500 308308
rect 340004 304666 340060 308308
rect 340004 304614 340006 304666
rect 340058 304614 340060 304666
rect 340004 304602 340060 304614
rect 340676 303994 340732 308308
rect 340676 303942 340678 303994
rect 340730 303942 340732 303994
rect 340676 303930 340732 303942
rect 341908 303882 341964 308308
rect 341908 303830 341910 303882
rect 341962 303830 341964 303882
rect 341908 303818 341964 303830
rect 339444 288138 339500 288148
rect 341796 303548 341852 303558
rect 341572 281708 341628 281718
rect 339332 281204 339612 281260
rect 339556 280924 339612 281204
rect 339556 280868 340368 280924
rect 341572 280896 341628 281652
rect 341796 281708 341852 303492
rect 342468 303100 342524 308308
rect 343028 303770 343084 308308
rect 344260 306348 344316 308308
rect 344932 307692 344988 308308
rect 344932 307626 344988 307636
rect 344260 306282 344316 306292
rect 345492 303884 345548 308308
rect 345492 303818 345548 303828
rect 343028 303718 343030 303770
rect 343082 303718 343084 303770
rect 343028 303706 343084 303718
rect 346164 303658 346220 308308
rect 346724 303772 346780 308308
rect 347396 304778 347452 308308
rect 347396 304726 347398 304778
rect 347450 304726 347452 304778
rect 347396 304714 347452 304726
rect 347956 304780 348012 308308
rect 347956 304714 348012 304724
rect 348516 304668 348572 308308
rect 349188 305674 349244 308308
rect 349188 305622 349190 305674
rect 349242 305622 349244 305674
rect 349188 305610 349244 305622
rect 349748 305676 349804 308308
rect 349748 305610 349804 305620
rect 350420 305450 350476 308308
rect 350980 305562 351036 308308
rect 350980 305510 350982 305562
rect 351034 305510 351036 305562
rect 350980 305498 351036 305510
rect 351652 305564 351708 308308
rect 351652 305498 351708 305508
rect 350420 305398 350422 305450
rect 350474 305398 350476 305450
rect 350420 305386 350476 305398
rect 352212 305452 352268 308308
rect 352212 305386 352268 305396
rect 352884 305340 352940 308308
rect 352884 305274 352940 305284
rect 353444 305338 353500 308308
rect 353444 305286 353446 305338
rect 353498 305286 353500 305338
rect 353444 305274 353500 305286
rect 354004 305226 354060 308308
rect 354004 305174 354006 305226
rect 354058 305174 354060 305226
rect 354004 305162 354060 305174
rect 354676 305114 354732 308308
rect 354676 305062 354678 305114
rect 354730 305062 354732 305114
rect 354676 305050 354732 305062
rect 355236 304890 355292 308308
rect 355908 305002 355964 308308
rect 357140 306460 357196 308308
rect 357700 307578 357756 308308
rect 357700 307526 357702 307578
rect 357754 307526 357756 307578
rect 357700 307514 357756 307526
rect 358372 307354 358428 308308
rect 358372 307302 358374 307354
rect 358426 307302 358428 307354
rect 358372 307290 358428 307302
rect 358932 307356 358988 308308
rect 358932 307290 358988 307300
rect 359380 308308 359492 308364
rect 360108 308364 360164 308896
rect 360668 308364 360724 308896
rect 361340 308364 361396 308896
rect 361900 308364 361956 308896
rect 362572 308476 362628 308896
rect 362572 308410 362628 308420
rect 363132 308476 363188 308896
rect 363132 308410 363188 308420
rect 363804 308364 363860 308896
rect 364364 308364 364420 308896
rect 364924 308364 364980 308896
rect 365596 308364 365652 308896
rect 366156 308364 366212 308896
rect 360108 308308 360220 308364
rect 360668 308308 360780 308364
rect 361340 308308 361452 308364
rect 361900 308308 362012 308364
rect 363804 308308 363916 308364
rect 364364 308308 364476 308364
rect 364924 308308 365036 308364
rect 365596 308308 365708 308364
rect 357140 306394 357196 306404
rect 355908 304950 355910 305002
rect 355962 304950 355964 305002
rect 355908 304938 355964 304950
rect 355236 304838 355238 304890
rect 355290 304838 355292 304890
rect 355236 304826 355292 304838
rect 348516 304602 348572 304612
rect 346724 303706 346780 303716
rect 346164 303606 346166 303658
rect 346218 303606 346220 303658
rect 346164 303594 346220 303606
rect 359380 303660 359436 308308
rect 359380 303594 359436 303604
rect 360164 303434 360220 308308
rect 360164 303382 360166 303434
rect 360218 303382 360220 303434
rect 360164 303370 360220 303382
rect 360724 303210 360780 308308
rect 360724 303158 360726 303210
rect 360778 303158 360780 303210
rect 360724 303146 360780 303158
rect 361172 307244 361228 307254
rect 342468 303034 342524 303044
rect 361172 302427 361228 307188
rect 361396 303546 361452 308308
rect 361396 303494 361398 303546
rect 361450 303494 361452 303546
rect 361396 303482 361452 303494
rect 361956 303322 362012 308308
rect 363860 307466 363916 308308
rect 363860 307414 363862 307466
rect 363914 307414 363916 307466
rect 363860 307402 363916 307414
rect 361956 303270 361958 303322
rect 362010 303270 362012 303322
rect 361956 303258 362012 303270
rect 362852 307132 362908 307142
rect 361172 302371 361340 302427
rect 348516 301980 348572 301990
rect 345156 299628 345212 299638
rect 341796 281642 341852 281652
rect 344148 281932 344204 281942
rect 342804 281596 342860 281606
rect 342804 280896 342860 281540
rect 344148 280896 344204 281876
rect 345156 281930 345212 299572
rect 345156 281878 345158 281930
rect 345210 281878 345212 281930
rect 345156 281866 345212 281878
rect 345380 281706 345436 281718
rect 345380 281654 345382 281706
rect 345434 281654 345436 281706
rect 345380 280896 345436 281654
rect 346724 281484 346780 281494
rect 346724 280896 346780 281428
rect 348516 280924 348572 301924
rect 349748 301868 349804 301878
rect 349748 280924 349804 301812
rect 354900 301868 354956 301878
rect 352772 301756 352828 301766
rect 351764 282044 351820 282054
rect 348516 280868 349328 280924
rect 349748 280868 350560 280924
rect 351764 280896 351820 281988
rect 352436 281930 352492 281942
rect 352436 281878 352438 281930
rect 352490 281878 352492 281930
rect 347732 280812 347788 280822
rect 347732 280810 347984 280812
rect 347732 280758 347734 280810
rect 347786 280758 347984 280810
rect 347732 280756 347984 280758
rect 347732 280746 347788 280756
rect 332164 280646 332166 280698
rect 332218 280646 332220 280698
rect 332164 280634 332220 280646
rect 352436 280698 352492 281878
rect 352772 280924 352828 301700
rect 354340 281708 354396 281718
rect 352772 280868 353136 280924
rect 354340 280896 354396 281652
rect 354900 280924 354956 301812
rect 357812 301530 357868 301542
rect 357812 301478 357814 301530
rect 357866 301478 357868 301530
rect 356132 301420 356188 301430
rect 356132 280924 356188 301364
rect 357812 280924 357868 301478
rect 359492 300412 359548 300422
rect 358484 281484 358540 281494
rect 354900 280868 355712 280924
rect 356132 280868 356944 280924
rect 357812 280868 358288 280924
rect 352436 280646 352438 280698
rect 352490 280646 352492 280698
rect 352436 280634 352492 280646
rect 358484 280698 358540 281428
rect 359492 280896 359548 300356
rect 359940 300300 359996 300310
rect 359940 280924 359996 300244
rect 361284 280924 361340 302371
rect 362740 281484 362796 281494
rect 359940 280868 360752 280924
rect 361284 280868 362096 280924
rect 362740 280810 362796 281428
rect 362852 280924 362908 307076
rect 364420 305116 364476 308308
rect 364420 305050 364476 305060
rect 364532 307020 364588 307030
rect 364532 280924 364588 306964
rect 364644 307018 364700 307030
rect 364644 306966 364646 307018
rect 364698 306966 364700 307018
rect 364644 302427 364700 306966
rect 364980 305228 365036 308308
rect 365652 307130 365708 308308
rect 366100 308308 366212 308364
rect 366828 308364 366884 308896
rect 367388 308364 367444 308896
rect 368060 308364 368116 308896
rect 368620 308476 368676 308896
rect 368620 308410 368676 308420
rect 369292 308364 369348 308896
rect 369852 308700 369908 308896
rect 369852 308634 369908 308644
rect 370412 308364 370468 308896
rect 371084 308812 371140 308896
rect 371028 308756 371140 308812
rect 366828 308308 366940 308364
rect 367388 308308 367500 308364
rect 368060 308308 368172 308364
rect 369292 308308 369404 308364
rect 366100 307242 366156 308308
rect 366100 307190 366102 307242
rect 366154 307190 366156 307242
rect 366100 307178 366156 307190
rect 365652 307078 365654 307130
rect 365706 307078 365708 307130
rect 365652 307066 365708 307078
rect 366884 307018 366940 308308
rect 366884 306966 366886 307018
rect 366938 306966 366940 307018
rect 366884 306954 366940 306966
rect 364980 305162 365036 305172
rect 366212 306906 366268 306918
rect 366212 306854 366214 306906
rect 366266 306854 366268 306906
rect 366212 302427 366268 306854
rect 367444 305004 367500 308308
rect 368116 306906 368172 308308
rect 368116 306854 368118 306906
rect 368170 306854 368172 306906
rect 368116 306842 368172 306854
rect 368228 308026 368284 308038
rect 368228 307974 368230 308026
rect 368282 307974 368284 308026
rect 367444 304938 367500 304948
rect 364644 302371 365148 302427
rect 366212 302371 366492 302427
rect 365092 280924 365148 302371
rect 366436 280924 366492 302371
rect 368228 280924 368284 307974
rect 369348 304892 369404 308308
rect 369348 304826 369404 304836
rect 369684 308308 370468 308364
rect 370916 308700 370972 308710
rect 369572 299740 369628 299750
rect 369572 280924 369628 299684
rect 369684 291452 369740 308308
rect 370916 307580 370972 308644
rect 370916 307514 370972 307524
rect 371028 307020 371084 308756
rect 371644 308364 371700 308896
rect 372316 308364 372372 308896
rect 372876 308364 372932 308896
rect 371644 308308 371756 308364
rect 372316 308308 372428 308364
rect 371700 307244 371756 308308
rect 371700 307178 371756 307188
rect 372372 307132 372428 308308
rect 372372 307066 372428 307076
rect 372820 308308 372932 308364
rect 373548 308364 373604 308896
rect 374108 308364 374164 308896
rect 374780 308364 374836 308896
rect 375340 308364 375396 308896
rect 375900 308364 375956 308896
rect 376572 308364 376628 308896
rect 376964 308588 377020 308598
rect 373548 308308 373660 308364
rect 374108 308308 374220 308364
rect 374780 308308 374892 308364
rect 375340 308308 375452 308364
rect 375900 308308 376012 308364
rect 376572 308308 376684 308364
rect 371028 306954 371084 306964
rect 372820 303996 372876 308308
rect 372820 303930 372876 303940
rect 373604 303436 373660 308308
rect 374164 306908 374220 308308
rect 374164 306842 374220 306852
rect 374836 303548 374892 308308
rect 374836 303482 374892 303492
rect 373604 303370 373660 303380
rect 375396 303324 375452 308308
rect 375396 303258 375452 303268
rect 375956 303212 376012 308308
rect 376628 308140 376684 308308
rect 376628 308074 376684 308084
rect 375956 303146 376012 303156
rect 376964 302427 377020 308532
rect 377132 308476 377188 308896
rect 377300 308700 377356 308710
rect 377300 308606 377356 308644
rect 377132 308410 377188 308420
rect 377412 308364 377468 308374
rect 377804 308364 377860 308896
rect 378084 308476 378140 308486
rect 377804 308308 377916 308364
rect 377412 302427 377468 308308
rect 377860 307468 377916 308308
rect 377860 307402 377916 307412
rect 376964 302371 377244 302427
rect 377412 302371 377580 302427
rect 369684 291386 369740 291396
rect 376628 300524 376684 300534
rect 373604 281596 373660 281606
rect 372260 281260 372316 281270
rect 362852 280868 363328 280924
rect 364532 280868 364672 280924
rect 365092 280868 365904 280924
rect 366436 280868 367248 280924
rect 368228 280868 368480 280924
rect 369572 280868 369824 280924
rect 372260 280896 372316 281204
rect 373604 280896 373660 281540
rect 374612 280924 374668 280934
rect 376628 280924 376684 300468
rect 377188 281596 377244 302371
rect 377188 281530 377244 281540
rect 377524 281484 377580 302371
rect 378084 282267 378140 308420
rect 378364 308364 378420 308896
rect 379036 308476 379092 308896
rect 379680 308868 379820 308924
rect 379036 308410 379092 308420
rect 377524 281418 377580 281428
rect 377860 282211 378140 282267
rect 378196 308308 378420 308364
rect 374668 280868 374864 280924
rect 376628 280868 377440 280924
rect 374612 280858 374668 280868
rect 362740 280758 362742 280810
rect 362794 280758 362796 280810
rect 362740 280746 362796 280758
rect 375508 280812 375564 280822
rect 375508 280810 376208 280812
rect 375508 280758 375510 280810
rect 375562 280758 376208 280810
rect 375508 280756 376208 280758
rect 375508 280746 375564 280756
rect 358484 280646 358486 280698
rect 358538 280646 358540 280698
rect 358484 280634 358540 280646
rect 370468 280700 370524 280710
rect 370524 280644 371056 280700
rect 377860 280698 377916 282211
rect 378084 280812 378140 280822
rect 378196 280812 378252 308308
rect 378756 281818 378812 281830
rect 378756 281766 378758 281818
rect 378810 281766 378812 281818
rect 378756 280896 378812 281766
rect 378084 280810 378252 280812
rect 378084 280758 378086 280810
rect 378138 280758 378252 280810
rect 378084 280756 378252 280758
rect 378084 280746 378140 280756
rect 377860 280646 377862 280698
rect 377914 280646 377916 280698
rect 370468 280634 370524 280644
rect 377860 280634 377916 280646
rect 379764 280700 379820 308868
rect 414932 308028 414988 308038
rect 414932 302427 414988 307972
rect 423332 307914 423388 307926
rect 423332 307862 423334 307914
rect 423386 307862 423388 307914
rect 414932 302371 415100 302427
rect 383012 300522 383068 300534
rect 383012 300470 383014 300522
rect 383066 300470 383068 300522
rect 381780 299740 381836 299750
rect 381220 281820 381276 281830
rect 379988 281594 380044 281606
rect 379988 281542 379990 281594
rect 380042 281542 380044 281594
rect 379988 280896 380044 281542
rect 381220 280896 381276 281764
rect 381780 280924 381836 299684
rect 383012 280924 383068 300470
rect 386372 300410 386428 300422
rect 386372 300358 386374 300410
rect 386426 300358 386428 300410
rect 384692 300298 384748 300310
rect 384692 300246 384694 300298
rect 384746 300246 384748 300298
rect 384692 280924 384748 300246
rect 381780 280868 382592 280924
rect 383012 280868 383824 280924
rect 384692 280868 385168 280924
rect 386372 280896 386428 300358
rect 386932 300186 386988 300198
rect 386932 300134 386934 300186
rect 386986 300134 386988 300186
rect 386932 280924 386988 300134
rect 388164 300188 388220 300198
rect 388164 280924 388220 300132
rect 391524 300076 391580 300086
rect 389732 299740 389788 299750
rect 389732 280924 389788 299684
rect 386932 280868 387744 280924
rect 388164 280868 388976 280924
rect 389732 280868 390320 280924
rect 391524 280896 391580 300020
rect 394772 300074 394828 300086
rect 394772 300022 394774 300074
rect 394826 300022 394828 300074
rect 393316 299964 393372 299974
rect 392756 282156 392812 282166
rect 392756 280896 392812 282100
rect 393316 280924 393372 299908
rect 394772 280924 394828 300022
rect 408660 299962 408716 299974
rect 408660 299910 408662 299962
rect 408714 299910 408716 299962
rect 399812 299852 399868 299862
rect 396676 281482 396732 281494
rect 396676 281430 396678 281482
rect 396730 281430 396732 281482
rect 393316 280868 394128 280924
rect 394772 280868 395360 280924
rect 396676 280896 396732 281430
rect 397908 281258 397964 281270
rect 397908 281206 397910 281258
rect 397962 281206 397964 281258
rect 397908 280896 397964 281206
rect 398580 281036 398636 281046
rect 398580 280924 398636 280980
rect 399812 280924 399868 299796
rect 403508 295036 403564 295046
rect 401492 281034 401548 281046
rect 401492 280982 401494 281034
rect 401546 280982 401548 281034
rect 401492 280924 401548 280982
rect 403508 280924 403564 294980
rect 404852 294924 404908 294934
rect 404852 280924 404908 294868
rect 406868 281372 406924 281382
rect 398580 280868 399280 280924
rect 399812 280868 400512 280924
rect 401492 280868 401744 280924
rect 403508 280868 404320 280924
rect 404852 280868 405664 280924
rect 406868 280896 406924 281316
rect 408212 281370 408268 281382
rect 408212 281318 408214 281370
rect 408266 281318 408268 281370
rect 408212 280896 408268 281318
rect 408660 280924 408716 299910
rect 410676 281820 410732 281830
rect 408660 280868 409472 280924
rect 410676 280896 410732 281764
rect 412020 281708 412076 281718
rect 412020 280896 412076 281652
rect 414596 281148 414652 281158
rect 413028 280924 413084 280934
rect 413028 280922 413280 280924
rect 413028 280870 413030 280922
rect 413082 280870 413280 280922
rect 414596 280896 414652 281092
rect 415044 280924 415100 302371
rect 418292 293244 418348 293254
rect 417172 281146 417228 281158
rect 417172 281094 417174 281146
rect 417226 281094 417228 281146
rect 413028 280868 413280 280870
rect 415044 280868 415856 280924
rect 417172 280896 417228 281094
rect 418292 280924 418348 293188
rect 418964 291900 419020 291910
rect 418964 280924 419020 291844
rect 421652 291788 421708 291798
rect 420196 291676 420252 291686
rect 420196 280924 420252 291620
rect 421652 280924 421708 291732
rect 423332 285628 423388 307862
rect 438452 307916 438508 307926
rect 426692 307468 426748 307478
rect 423332 285562 423388 285572
rect 423444 291564 423500 291574
rect 423444 280924 423500 291508
rect 424116 285628 424172 285638
rect 424116 280924 424172 285572
rect 426132 281596 426188 281606
rect 418292 280868 418432 280924
rect 418964 280868 419776 280924
rect 420196 280868 421008 280924
rect 421652 280868 422240 280924
rect 423444 280868 423584 280924
rect 424116 280868 424816 280924
rect 426132 280896 426188 281540
rect 426692 280924 426748 307412
rect 428820 291900 428876 291910
rect 428596 291788 428652 291798
rect 428596 285628 428652 291732
rect 428596 285562 428652 285572
rect 428820 280924 428876 291844
rect 433412 291786 433468 291798
rect 433412 291734 433414 291786
rect 433466 291734 433468 291786
rect 430388 291564 430444 291574
rect 426692 280868 427392 280924
rect 428736 280868 428876 280924
rect 429268 285628 429324 285638
rect 429268 280924 429324 285572
rect 430388 280924 430444 291508
rect 432516 289996 432572 290006
rect 429268 280868 429968 280924
rect 430388 280868 431200 280924
rect 432516 280896 432572 289940
rect 433412 280924 433468 291734
rect 435204 291674 435260 291686
rect 435204 291622 435206 291674
rect 435258 291622 435260 291674
rect 435204 280924 435260 291622
rect 433412 280868 433776 280924
rect 435120 280868 435260 280924
rect 436324 285180 436380 285190
rect 436324 280896 436380 285124
rect 437668 285068 437724 285078
rect 437668 280896 437724 285012
rect 438452 280924 438508 307860
rect 440244 307802 440300 307814
rect 440244 307750 440246 307802
rect 440298 307750 440300 307802
rect 438452 280868 438928 280924
rect 440244 280896 440300 307750
rect 456036 291562 456092 291574
rect 456036 291510 456038 291562
rect 456090 291510 456092 291562
rect 451668 285066 451724 285078
rect 451668 285014 451670 285066
rect 451722 285014 451724 285066
rect 442708 284956 442764 284966
rect 441476 284844 441532 284854
rect 441476 280896 441532 284788
rect 442708 280896 442764 284900
rect 449204 284954 449260 284966
rect 449204 284902 449206 284954
rect 449258 284902 449260 284954
rect 444052 284620 444108 284630
rect 444052 280896 444108 284564
rect 445284 282156 445340 282166
rect 445284 280896 445340 282100
rect 446628 282156 446684 282166
rect 446628 280896 446684 282100
rect 447860 281484 447916 281494
rect 447860 280896 447916 281428
rect 449204 280896 449260 284902
rect 451668 280896 451724 285014
rect 454244 284842 454300 284854
rect 454244 284790 454246 284842
rect 454298 284790 454300 284842
rect 453012 281260 453068 281270
rect 453012 280896 453068 281204
rect 454244 280896 454300 284790
rect 455588 284730 455644 284742
rect 455588 284678 455590 284730
rect 455642 284678 455644 284730
rect 455588 280896 455644 284678
rect 456036 280924 456092 291510
rect 457380 291450 457436 291462
rect 457380 291398 457382 291450
rect 457434 291398 457436 291450
rect 457380 280924 457436 291398
rect 458612 280924 458668 309204
rect 460292 280924 460348 312452
rect 548436 308140 548492 308150
rect 532420 307804 532476 307814
rect 467796 307690 467852 307702
rect 467796 307638 467798 307690
rect 467850 307638 467852 307690
rect 463764 294812 463820 294822
rect 463764 290780 463820 294756
rect 467012 293914 467068 293926
rect 467012 293862 467014 293914
rect 467066 293862 467068 293914
rect 461748 280924 461804 280934
rect 462644 280924 462700 280934
rect 463764 280924 463820 290724
rect 465332 293132 465388 293142
rect 465332 292348 465388 293076
rect 465332 280924 465388 292292
rect 467012 292346 467068 293862
rect 467796 293914 467852 307638
rect 482916 307692 482972 307702
rect 481236 306348 481292 306358
rect 467796 293862 467798 293914
rect 467850 293862 467852 293914
rect 467796 293850 467852 293862
rect 472052 304666 472108 304678
rect 472052 304614 472054 304666
rect 472106 304614 472108 304666
rect 467012 292294 467014 292346
rect 467066 292294 467068 292346
rect 467012 280924 467068 292294
rect 472052 290332 472108 304614
rect 470932 288428 470988 288438
rect 468580 287308 468636 287318
rect 468580 280924 468636 287252
rect 456036 280868 456848 280924
rect 457380 280868 458192 280924
rect 458612 280868 459424 280924
rect 460292 280868 460656 280924
rect 461804 280868 462000 280924
rect 462700 280868 463232 280924
rect 463764 280868 464576 280924
rect 465332 280868 465808 280924
rect 467012 280868 467152 280924
rect 468384 280868 468636 280924
rect 469140 287308 469196 287318
rect 469140 280924 469196 287252
rect 469140 280868 469728 280924
rect 470932 280896 470988 288372
rect 472052 280924 472108 290276
rect 472836 303994 472892 304006
rect 472836 303942 472838 303994
rect 472890 303942 472892 303994
rect 472836 288092 472892 303942
rect 472836 280924 472892 288036
rect 475412 303882 475468 303894
rect 475412 303830 475414 303882
rect 475466 303830 475468 303882
rect 475412 290556 475468 303830
rect 474516 287308 474572 287318
rect 474516 280924 474572 287252
rect 475412 280924 475468 290500
rect 477876 303770 477932 303782
rect 477876 303718 477878 303770
rect 477930 303718 477932 303770
rect 477876 290332 477932 303718
rect 481236 290444 481292 306292
rect 477876 290266 477932 290276
rect 478660 290332 478716 290342
rect 477876 280924 477932 280934
rect 472052 280868 472192 280924
rect 472836 280868 473536 280924
rect 474516 280868 474768 280924
rect 475412 280868 476112 280924
rect 477344 280868 477876 280924
rect 478660 280896 478716 290276
rect 479556 289324 479612 289334
rect 479556 289100 479612 289268
rect 479556 280924 479612 289044
rect 481236 280924 481292 290388
rect 482916 290556 482972 307636
rect 509796 307578 509852 307590
rect 509796 307526 509798 307578
rect 509850 307526 509852 307578
rect 508116 306460 508172 306470
rect 491316 305674 491372 305686
rect 491316 305622 491318 305674
rect 491370 305622 491372 305674
rect 487956 304778 488012 304790
rect 487956 304726 487958 304778
rect 488010 304726 488012 304778
rect 485492 303772 485548 303782
rect 483812 303658 483868 303670
rect 483812 303606 483814 303658
rect 483866 303606 483868 303658
rect 483812 294140 483868 303606
rect 483812 290667 483868 294084
rect 485492 294028 485548 303716
rect 483812 290611 484316 290667
rect 482916 280924 482972 290500
rect 479556 280868 479920 280924
rect 481152 280868 481292 280924
rect 482496 280868 482972 280924
rect 483028 280924 483084 280934
rect 484260 280924 484316 290611
rect 485492 280924 485548 293972
rect 487172 293914 487228 293926
rect 487172 293862 487174 293914
rect 487226 293862 487228 293914
rect 487172 292682 487228 293862
rect 487956 293914 488012 304726
rect 489636 304780 489692 304790
rect 487956 293862 487958 293914
rect 488010 293862 488012 293914
rect 487956 293850 488012 293862
rect 488852 304668 488908 304678
rect 487172 292630 487174 292682
rect 487226 292630 487228 292682
rect 487172 280924 487228 292630
rect 488852 292908 488908 304612
rect 488852 285628 488908 292852
rect 488852 285562 488908 285572
rect 489076 292684 489132 292694
rect 489076 280924 489132 292628
rect 489636 292684 489692 304724
rect 489636 292618 489692 292628
rect 490644 293916 490700 293926
rect 490644 292908 490700 293860
rect 491316 293916 491372 305622
rect 491316 293850 491372 293860
rect 492996 305676 493052 305686
rect 483084 280868 483728 280924
rect 484260 280868 485072 280924
rect 485492 280868 486304 280924
rect 487172 280868 487648 280924
rect 488880 280868 489132 280924
rect 489524 285628 489580 285638
rect 489524 280924 489580 285572
rect 490644 280924 490700 292852
rect 492212 293466 492268 293478
rect 492212 293414 492214 293466
rect 492266 293414 492268 293466
rect 492212 280924 492268 293414
rect 492996 293466 493052 305620
rect 494676 305562 494732 305574
rect 494676 305510 494678 305562
rect 494730 305510 494732 305562
rect 494676 293692 494732 305510
rect 496356 305564 496412 305574
rect 492996 293414 492998 293466
rect 493050 293414 493052 293466
rect 492996 292794 493052 293414
rect 492996 292742 492998 292794
rect 493050 292742 493052 292794
rect 492996 292730 493052 292742
rect 494004 293466 494060 293478
rect 494004 293414 494006 293466
rect 494058 293414 494060 293466
rect 493892 292348 493948 292358
rect 493892 285628 493948 292292
rect 493892 285562 493948 285572
rect 489524 280868 490224 280924
rect 490644 280868 491456 280924
rect 492212 280868 492688 280924
rect 494004 280896 494060 293414
rect 494676 292348 494732 293636
rect 494900 305450 494956 305462
rect 494900 305398 494902 305450
rect 494954 305398 494956 305450
rect 494900 293466 494956 305398
rect 494900 293414 494902 293466
rect 494954 293414 494956 293466
rect 494900 293130 494956 293414
rect 494900 293078 494902 293130
rect 494954 293078 494956 293130
rect 494900 293066 494956 293078
rect 495796 293914 495852 293926
rect 495796 293862 495798 293914
rect 495850 293862 495852 293914
rect 494676 292282 494732 292292
rect 495796 292570 495852 293862
rect 496356 293914 496412 305508
rect 496356 293862 496358 293914
rect 496410 293862 496412 293914
rect 496356 293850 496412 293862
rect 497252 305452 497308 305462
rect 495796 292518 495798 292570
rect 495850 292518 495852 292570
rect 494564 285628 494620 285638
rect 494564 280924 494620 285572
rect 495796 280924 495852 292518
rect 497252 292572 497308 305396
rect 497252 280924 497308 292516
rect 498932 305340 498988 305350
rect 498932 292796 498988 305284
rect 498932 280924 498988 292740
rect 499716 305338 499772 305350
rect 499716 305286 499718 305338
rect 499770 305286 499772 305338
rect 499716 292348 499772 305286
rect 501396 305226 501452 305238
rect 501396 305174 501398 305226
rect 501450 305174 501452 305226
rect 499716 290667 499772 292292
rect 499604 290611 499772 290667
rect 500836 292458 500892 292470
rect 500836 292406 500838 292458
rect 500890 292406 500892 292458
rect 499604 280924 499660 290611
rect 500836 280924 500892 292406
rect 501396 292458 501452 305174
rect 501396 292406 501398 292458
rect 501450 292406 501452 292458
rect 501396 292394 501452 292406
rect 502292 305114 502348 305126
rect 502292 305062 502294 305114
rect 502346 305062 502348 305114
rect 502292 294364 502348 305062
rect 504756 305002 504812 305014
rect 504756 304950 504758 305002
rect 504810 304950 504812 305002
rect 502292 280924 502348 294308
rect 503972 304890 504028 304902
rect 503972 304838 503974 304890
rect 504026 304838 504028 304890
rect 503972 294252 504028 304838
rect 503972 280924 504028 294196
rect 504756 291674 504812 304950
rect 504756 291622 504758 291674
rect 504810 291622 504812 291674
rect 504756 280924 504812 291622
rect 507332 292236 507388 292246
rect 505988 291564 506044 291574
rect 505988 280924 506044 291508
rect 507332 280924 507388 292180
rect 508116 292236 508172 306404
rect 509012 293916 509068 293926
rect 508564 292570 508620 292582
rect 508564 292518 508566 292570
rect 508618 292518 508620 292570
rect 508228 292460 508284 292470
rect 508564 292460 508620 292518
rect 508228 292458 508620 292460
rect 508228 292406 508230 292458
rect 508282 292406 508620 292458
rect 508228 292404 508620 292406
rect 509012 292572 509068 293860
rect 509796 293916 509852 307526
rect 520884 307466 520940 307478
rect 520884 307414 520886 307466
rect 520938 307414 520940 307466
rect 509796 293850 509852 293860
rect 509908 307354 509964 307366
rect 509908 307302 509910 307354
rect 509962 307302 509964 307354
rect 508228 292394 508284 292404
rect 508116 291788 508172 292180
rect 508116 291722 508172 291732
rect 509012 280924 509068 292516
rect 509908 290890 509964 307302
rect 509908 290838 509910 290890
rect 509962 290838 509964 290890
rect 509908 290667 509964 290838
rect 509796 290611 509964 290667
rect 510692 307356 510748 307366
rect 510692 293020 510748 307300
rect 520548 303996 520604 304006
rect 510692 290667 510748 292964
rect 513156 303660 513212 303670
rect 512372 292796 512428 292806
rect 510692 290611 511196 290667
rect 509796 280924 509852 290611
rect 511140 280924 511196 290611
rect 512372 280924 512428 292740
rect 513156 292796 513212 303604
rect 516516 303546 516572 303558
rect 516516 303494 516518 303546
rect 516570 303494 516572 303546
rect 514836 303434 514892 303446
rect 514836 303382 514838 303434
rect 514890 303382 514892 303434
rect 513156 292730 513212 292740
rect 514052 293916 514108 293926
rect 514052 293020 514108 293860
rect 514836 293916 514892 303382
rect 514836 293850 514892 293860
rect 515732 293914 515788 293926
rect 515732 293862 515734 293914
rect 515786 293862 515788 293914
rect 514052 280924 514108 292964
rect 494564 280868 495264 280924
rect 495796 280868 496608 280924
rect 497252 280868 497840 280924
rect 498932 280868 499184 280924
rect 499604 280868 500416 280924
rect 500836 280868 501648 280924
rect 502292 280868 502992 280924
rect 503972 280868 504224 280924
rect 504756 280868 505568 280924
rect 505988 280868 506800 280924
rect 507332 280868 508144 280924
rect 509012 280868 509376 280924
rect 509796 280868 510608 280924
rect 511140 280868 511952 280924
rect 512372 280868 513184 280924
rect 514052 280868 514528 280924
rect 515732 280896 515788 293862
rect 516516 291002 516572 303494
rect 518196 303322 518252 303334
rect 518196 303270 518198 303322
rect 518250 303270 518252 303322
rect 516740 303210 516796 303222
rect 516740 303158 516742 303210
rect 516794 303158 516796 303210
rect 516740 293914 516796 303158
rect 516740 293862 516742 293914
rect 516794 293862 516796 293914
rect 516740 293018 516796 293862
rect 516740 292966 516742 293018
rect 516794 292966 516796 293018
rect 516740 292954 516796 292966
rect 517524 293914 517580 293926
rect 517524 293862 517526 293914
rect 517578 293862 517580 293914
rect 516516 290950 516518 291002
rect 516570 290950 516572 291002
rect 516516 290667 516572 290950
rect 516292 290611 516572 290667
rect 517524 292906 517580 293862
rect 518196 293914 518252 303270
rect 518196 293862 518198 293914
rect 518250 293862 518252 293914
rect 518196 293850 518252 293862
rect 517524 292854 517526 292906
rect 517578 292854 517580 292906
rect 516292 280924 516348 290611
rect 517524 280924 517580 292854
rect 519092 293578 519148 293590
rect 519092 293526 519094 293578
rect 519146 293526 519148 293578
rect 519092 280924 519148 293526
rect 520548 293578 520604 303940
rect 520548 293526 520550 293578
rect 520602 293526 520604 293578
rect 520548 293242 520604 293526
rect 520548 293190 520550 293242
rect 520602 293190 520604 293242
rect 520548 293178 520604 293190
rect 520772 293354 520828 293366
rect 520772 293302 520774 293354
rect 520826 293302 520828 293354
rect 520772 280924 520828 293302
rect 520884 290667 520940 307414
rect 526820 307242 526876 307254
rect 526820 307190 526822 307242
rect 526874 307190 526876 307242
rect 526596 307130 526652 307142
rect 526596 307078 526598 307130
rect 526650 307078 526652 307130
rect 524916 305228 524972 305238
rect 523236 305116 523292 305126
rect 522340 303772 522396 303782
rect 522340 293354 522396 303716
rect 522340 293302 522342 293354
rect 522394 293302 522396 293354
rect 522340 293290 522396 293302
rect 522676 292236 522732 292246
rect 522676 291116 522732 292180
rect 523236 292236 523292 305060
rect 523236 292170 523292 292180
rect 521332 291004 521388 291014
rect 521332 290667 521388 290948
rect 520884 290611 521388 290667
rect 521332 280924 521388 290611
rect 522676 280924 522732 291060
rect 524132 291228 524188 291238
rect 524132 280924 524188 291172
rect 524916 291228 524972 305172
rect 524916 291162 524972 291172
rect 525924 291564 525980 291574
rect 525812 291114 525868 291126
rect 525812 291062 525814 291114
rect 525866 291062 525868 291114
rect 525812 285626 525868 291062
rect 525812 285574 525814 285626
rect 525866 285574 525868 285626
rect 525812 285562 525868 285574
rect 525924 280924 525980 291508
rect 526596 291564 526652 307078
rect 526596 291498 526652 291508
rect 526820 291114 526876 307190
rect 526820 291062 526822 291114
rect 526874 291062 526876 291114
rect 526820 291050 526876 291062
rect 528276 307018 528332 307030
rect 528276 306966 528278 307018
rect 528330 306966 528332 307018
rect 528276 291226 528332 306966
rect 531636 306906 531692 306918
rect 531636 306854 531638 306906
rect 531690 306854 531692 306906
rect 529956 305004 530012 305014
rect 528276 291174 528278 291226
rect 528330 291174 528332 291226
rect 528276 290667 528332 291174
rect 527828 290611 528332 290667
rect 529172 292122 529228 292134
rect 529172 292070 529174 292122
rect 529226 292070 529228 292122
rect 529172 291338 529228 292070
rect 529956 292122 530012 304948
rect 529956 292070 529958 292122
rect 530010 292070 530012 292122
rect 529956 292058 530012 292070
rect 531076 292122 531132 292134
rect 531076 292070 531078 292122
rect 531130 292070 531132 292122
rect 529172 291286 529174 291338
rect 529226 291286 529228 291338
rect 526596 285626 526652 285638
rect 526596 285574 526598 285626
rect 526650 285574 526652 285626
rect 526596 280924 526652 285574
rect 527828 280924 527884 290611
rect 529172 280924 529228 291286
rect 530852 292010 530908 292022
rect 530852 291958 530854 292010
rect 530906 291958 530908 292010
rect 530852 282826 530908 291958
rect 530852 282774 530854 282826
rect 530906 282774 530908 282826
rect 530852 282762 530908 282774
rect 531076 291562 531132 292070
rect 531636 292122 531692 306854
rect 531636 292070 531638 292122
rect 531690 292070 531692 292122
rect 531636 292058 531692 292070
rect 531076 291510 531078 291562
rect 531130 291510 531132 291562
rect 516292 280868 517104 280924
rect 517524 280868 518336 280924
rect 519092 280868 519680 280924
rect 520772 280868 520912 280924
rect 521332 280868 522144 280924
rect 522676 280868 523488 280924
rect 524132 280868 524720 280924
rect 525924 280868 526064 280924
rect 526596 280868 527296 280924
rect 527828 280868 528640 280924
rect 529172 280868 529872 280924
rect 531076 280896 531132 291510
rect 532420 292010 532476 307748
rect 534212 307580 534268 307590
rect 532420 291958 532422 292010
rect 532474 291958 532476 292010
rect 532420 291450 532476 291958
rect 532420 291398 532422 291450
rect 532474 291398 532476 291450
rect 532420 291386 532476 291398
rect 532532 304892 532588 304902
rect 532532 291340 532588 304836
rect 532532 290667 532588 291284
rect 534212 291676 534268 307524
rect 539252 307132 539308 307142
rect 532532 290611 532924 290667
rect 531748 282826 531804 282838
rect 531748 282774 531750 282826
rect 531802 282774 531804 282826
rect 531748 280924 531804 282774
rect 532868 280924 532924 290611
rect 534212 280924 534268 291620
rect 538356 307020 538412 307030
rect 535892 291452 535948 291462
rect 535892 290892 535948 291396
rect 535892 280924 535948 290836
rect 537572 291452 537628 291462
rect 531748 280868 532448 280924
rect 532868 280868 533680 280924
rect 534212 280868 535024 280924
rect 535892 280868 536256 280924
rect 537572 280896 537628 291396
rect 538356 291452 538412 306964
rect 538356 291386 538412 291396
rect 539252 293468 539308 307076
rect 543396 306908 543452 306918
rect 539252 290667 539308 293412
rect 542612 293916 542668 293926
rect 542612 293132 542668 293860
rect 543396 293916 543452 306852
rect 545076 303548 545132 303558
rect 543396 293850 543452 293860
rect 543508 303436 543564 303446
rect 540932 292236 540988 292246
rect 540932 290892 540988 292180
rect 539252 290611 539420 290667
rect 538244 280924 538300 280934
rect 539364 280924 539420 290611
rect 540932 280924 540988 290836
rect 542612 285626 542668 293076
rect 542612 285574 542614 285626
rect 542666 285574 542668 285626
rect 542612 285562 542668 285574
rect 542724 292236 542780 292246
rect 542724 280924 542780 292180
rect 543508 292236 543564 303380
rect 543508 291564 543564 292180
rect 543508 291498 543564 291508
rect 544404 293916 544460 293926
rect 544404 293244 544460 293860
rect 545076 293916 545132 303492
rect 545076 293850 545132 293860
rect 546756 303324 546812 303334
rect 538300 280868 538832 280924
rect 539364 280868 540176 280924
rect 540932 280868 541408 280924
rect 542640 280868 542780 280924
rect 543284 285626 543340 285638
rect 543284 285574 543286 285626
rect 543338 285574 543340 285626
rect 543284 280924 543340 285574
rect 544404 280924 544460 293188
rect 545972 293356 546028 293366
rect 545972 280924 546028 293300
rect 546756 293356 546812 303268
rect 546756 293290 546812 293300
rect 547652 293468 547708 293478
rect 547652 280924 547708 293412
rect 548436 291676 548492 308084
rect 551012 307468 551068 307478
rect 548548 303212 548604 303222
rect 548548 293468 548604 303156
rect 548548 293402 548604 293412
rect 549556 293916 549612 293926
rect 548436 290667 548492 291620
rect 548324 290611 548492 290667
rect 548324 280924 548380 290611
rect 549556 280924 549612 293860
rect 551012 280924 551068 307412
rect 556724 284732 556780 284742
rect 543284 280868 543984 280924
rect 544404 280868 545216 280924
rect 545972 280868 546560 280924
rect 547652 280868 547792 280924
rect 548324 280868 549136 280924
rect 549556 280868 550368 280924
rect 551012 280868 551600 280924
rect 556724 280896 556780 284676
rect 557732 280924 557788 319396
rect 560196 301644 560252 301654
rect 559076 280924 559132 280934
rect 557732 280868 558096 280924
rect 559132 280868 559328 280924
rect 413028 280858 413084 280868
rect 461748 280858 461804 280868
rect 462644 280858 462700 280868
rect 477876 280858 477932 280868
rect 483028 280858 483084 280868
rect 538244 280858 538300 280868
rect 559076 280858 559132 280868
rect 402388 280812 402444 280822
rect 552692 280812 552748 280822
rect 402444 280756 403088 280812
rect 552692 280810 552944 280812
rect 552692 280758 552694 280810
rect 552746 280758 552944 280810
rect 552692 280756 552944 280758
rect 402388 280746 402444 280756
rect 552692 280746 552748 280756
rect 379764 280634 379820 280644
rect 450212 280700 450268 280710
rect 553588 280700 553644 280710
rect 554820 280700 554876 280710
rect 450212 280698 450464 280700
rect 450212 280646 450214 280698
rect 450266 280646 450464 280698
rect 450212 280644 450464 280646
rect 553588 280698 554176 280700
rect 553588 280646 553590 280698
rect 553642 280646 554176 280698
rect 553588 280644 554176 280646
rect 554876 280644 555520 280700
rect 450212 280634 450268 280644
rect 553588 280634 553644 280644
rect 554820 280634 554876 280644
rect 559636 254380 559692 254390
rect 559636 235228 559692 254324
rect 560084 252028 560140 252038
rect 559636 235162 559692 235172
rect 559748 240268 559804 240278
rect 559748 217980 559804 240212
rect 559972 233884 560028 233894
rect 559748 217914 559804 217924
rect 559860 231644 559916 231654
rect 559860 206220 559916 231588
rect 559972 209132 560028 233828
rect 560084 232764 560140 251972
rect 560084 232698 560140 232708
rect 559972 209066 560028 209076
rect 560084 220444 560140 220454
rect 559860 206154 559916 206164
rect 560084 191436 560140 220388
rect 560084 191370 560140 191380
rect 90356 191258 90412 191268
rect 84308 190922 84364 190932
rect 559412 141708 559468 141718
rect 559412 90747 559468 141652
rect 560196 139914 560252 301588
rect 566020 301532 566076 301542
rect 566020 293466 566076 301476
rect 566020 293414 566022 293466
rect 566074 293414 566076 293466
rect 560420 256620 560476 256630
rect 560420 238476 560476 256564
rect 560868 249676 560924 249686
rect 560644 247548 560700 247558
rect 560532 240716 560588 240726
rect 560532 240268 560588 240660
rect 560532 240202 560588 240212
rect 560420 238410 560476 238420
rect 560420 236236 560476 236246
rect 560420 211596 560476 236180
rect 560644 226268 560700 247492
rect 560868 229180 560924 249620
rect 560868 229114 560924 229124
rect 560980 245308 561036 245318
rect 560644 226202 560700 226212
rect 560868 224812 560924 224822
rect 560644 222572 560700 222582
rect 560532 211596 560588 211606
rect 560420 211540 560532 211596
rect 560532 211530 560588 211540
rect 560420 206668 560476 206678
rect 560308 185724 560364 185734
rect 560308 183036 560364 185668
rect 560308 182970 560364 182980
rect 560420 173852 560476 206612
rect 560644 193900 560700 222516
rect 560868 196812 560924 224756
rect 560980 223356 561036 245252
rect 560980 223290 561036 223300
rect 561876 238476 561932 238486
rect 560868 196746 560924 196756
rect 560980 215740 561036 215750
rect 560644 193834 560700 193844
rect 560868 195244 560924 195254
rect 560756 193004 560812 193014
rect 560644 190764 560700 190774
rect 560532 183036 560588 183046
rect 560532 181692 560588 182980
rect 560532 181626 560588 181636
rect 560420 173786 560476 173796
rect 560420 168028 560476 168038
rect 560196 139862 560198 139914
rect 560250 139862 560252 139914
rect 560196 135660 560252 139862
rect 560196 135594 560252 135604
rect 560308 154364 560364 154374
rect 560196 122778 560252 122790
rect 560196 122726 560198 122778
rect 560250 122726 560252 122778
rect 559412 90691 559580 90747
rect 559412 82234 559468 82246
rect 559412 82182 559414 82234
rect 559466 82182 559468 82234
rect 559412 81676 559468 82182
rect 559524 82122 559580 90691
rect 559524 82070 559526 82122
rect 559578 82070 559580 82122
rect 559524 82058 559580 82070
rect 559412 81610 559468 81620
rect 78260 80950 78262 81002
rect 78314 80950 78316 81002
rect 78260 80938 78316 80950
rect 92372 80892 92428 80902
rect 92372 80798 92428 80836
rect 335972 80780 336028 80790
rect 335972 80686 336028 80724
rect 123508 78988 123564 80304
rect 190596 79100 190652 80304
rect 190596 79034 190652 79044
rect 123508 78922 123564 78932
rect 257796 70588 257852 80304
rect 324884 72156 324940 80304
rect 324884 72090 324940 72100
rect 392084 71820 392140 80304
rect 459172 72044 459228 80304
rect 526372 72156 526428 80304
rect 560196 79100 560252 122726
rect 560308 100380 560364 154308
rect 560420 117516 560476 167972
rect 560644 152796 560700 190708
rect 560756 155708 560812 192948
rect 560868 158620 560924 195188
rect 560980 185052 561036 215684
rect 561876 214508 561932 238420
rect 561876 214442 561932 214452
rect 565236 229404 565292 229414
rect 565236 202076 565292 229348
rect 565236 202010 565292 202020
rect 560980 184986 561036 184996
rect 560868 158554 560924 158564
rect 561876 172620 561932 172630
rect 560756 155642 560812 155652
rect 560644 152730 560700 152740
rect 561876 120428 561932 172564
rect 561876 120362 561932 120372
rect 565236 156716 565292 156726
rect 560532 117516 560588 117526
rect 560420 117460 560532 117516
rect 560532 117450 560588 117460
rect 560308 100314 560364 100324
rect 565236 96236 565292 156660
rect 566020 122890 566076 293414
rect 606116 294140 606172 294150
rect 605780 292684 605836 292694
rect 605780 290442 605836 292628
rect 605780 290390 605782 290442
rect 605834 290390 605836 290442
rect 605780 290378 605836 290390
rect 606116 290330 606172 294084
rect 606228 293130 606284 293142
rect 606228 293078 606230 293130
rect 606282 293078 606284 293130
rect 606228 291900 606284 293078
rect 606228 291834 606284 291844
rect 606340 292682 606396 292694
rect 606340 292630 606342 292682
rect 606394 292630 606396 292682
rect 606340 290554 606396 292630
rect 609812 292348 609868 292358
rect 609812 292234 609868 292292
rect 609812 292182 609814 292234
rect 609866 292182 609868 292234
rect 609812 292170 609868 292182
rect 610820 292010 610876 292022
rect 610820 291958 610822 292010
rect 610874 291958 610876 292010
rect 609924 291786 609980 291798
rect 609924 291734 609926 291786
rect 609978 291734 609980 291786
rect 606340 290502 606342 290554
rect 606394 290502 606396 290554
rect 606340 290490 606396 290502
rect 609812 291004 609868 291014
rect 606116 290278 606118 290330
rect 606170 290278 606172 290330
rect 606116 290266 606172 290278
rect 606340 290220 606396 290230
rect 606340 290126 606396 290164
rect 600516 289212 600572 289222
rect 570500 281260 570556 281270
rect 570388 281036 570444 281046
rect 570276 280812 570332 280822
rect 570276 270284 570332 280756
rect 570388 277116 570444 280980
rect 570388 277050 570444 277060
rect 570500 270396 570556 281204
rect 570500 270330 570556 270340
rect 570276 270218 570332 270228
rect 597156 261212 597212 261222
rect 585396 258860 585452 258870
rect 583716 242956 583772 242966
rect 566916 227052 566972 227062
rect 566916 199164 566972 226996
rect 583716 220220 583772 242900
rect 583716 220154 583772 220164
rect 578676 217980 578732 217990
rect 566916 199098 566972 199108
rect 568596 213500 568652 213510
rect 568596 181468 568652 213444
rect 568596 181402 568652 181412
rect 568708 211148 568764 211158
rect 568708 178556 568764 211092
rect 570612 204428 570668 204438
rect 570500 202076 570556 202086
rect 568708 178490 568764 178500
rect 570276 199836 570332 199846
rect 570276 163884 570332 199780
rect 570276 163818 570332 163828
rect 570388 197596 570444 197606
rect 570388 161308 570444 197540
rect 570500 166796 570556 202020
rect 570612 169708 570668 204372
rect 570612 169642 570668 169652
rect 571956 188524 572012 188534
rect 570500 166730 570556 166740
rect 570388 161242 570444 161252
rect 571956 149548 572012 188468
rect 578676 186508 578732 217924
rect 578676 186442 578732 186452
rect 571956 149482 572012 149492
rect 575316 152124 575372 152134
rect 566020 122838 566022 122890
rect 566074 122838 566076 122890
rect 566020 122826 566076 122838
rect 575316 102508 575372 152068
rect 575316 102442 575372 102452
rect 565236 96170 565292 96180
rect 560308 81900 560364 81910
rect 560308 80666 560364 81844
rect 585396 81676 585452 258804
rect 597156 240380 597212 261156
rect 597156 240314 597212 240324
rect 585396 81610 585452 81620
rect 585620 179340 585676 179350
rect 585620 81228 585676 179284
rect 585844 165788 585900 165798
rect 585844 81340 585900 165732
rect 586068 163436 586124 163446
rect 586068 81452 586124 163380
rect 598836 149884 598892 149894
rect 598836 92428 598892 149828
rect 598836 92362 598892 92372
rect 600516 82234 600572 289156
rect 609812 289212 609868 290948
rect 609812 289146 609868 289156
rect 606340 288874 606396 288886
rect 606340 288822 606342 288874
rect 606394 288822 606396 288874
rect 606228 288762 606284 288774
rect 606228 288710 606230 288762
rect 606282 288710 606284 288762
rect 606228 288092 606284 288710
rect 606340 288204 606396 288822
rect 606340 288138 606396 288148
rect 606228 288026 606284 288036
rect 609924 283164 609980 291734
rect 610708 290778 610764 290790
rect 610708 290726 610710 290778
rect 610762 290726 610764 290778
rect 610708 288316 610764 290726
rect 610820 290330 610876 291958
rect 610820 290278 610822 290330
rect 610874 290278 610876 290330
rect 610820 290266 610876 290278
rect 610820 290106 610876 290118
rect 610820 290054 610822 290106
rect 610874 290054 610876 290106
rect 610820 288762 610876 290054
rect 610932 289996 610988 333396
rect 611044 333450 611100 333462
rect 611044 333398 611046 333450
rect 611098 333398 611100 333450
rect 611044 290330 611100 333398
rect 626612 333340 626668 333350
rect 632436 333340 632492 333350
rect 611268 331994 611324 333312
rect 611268 331942 611270 331994
rect 611322 331942 611324 331994
rect 611268 331930 611324 331942
rect 613284 328748 613340 333312
rect 615300 333002 615356 333312
rect 615300 332950 615302 333002
rect 615354 332950 615356 333002
rect 615300 332938 615356 332950
rect 617316 330202 617372 333312
rect 617316 330150 617318 330202
rect 617370 330150 617372 330202
rect 617316 330138 617372 330150
rect 619220 330090 619276 333312
rect 621236 332778 621292 333312
rect 621236 332726 621238 332778
rect 621290 332726 621292 332778
rect 621236 332714 621292 332726
rect 623252 332668 623308 333312
rect 623252 332602 623308 332612
rect 619220 330038 619222 330090
rect 619274 330038 619276 330090
rect 619220 330026 619276 330038
rect 613284 328682 613340 328692
rect 625268 328746 625324 333312
rect 626668 333284 627200 333340
rect 632436 333338 633136 333340
rect 626612 333274 626668 333284
rect 629188 330204 629244 333312
rect 629188 330138 629244 330148
rect 631204 330092 631260 333312
rect 632436 333286 632438 333338
rect 632490 333286 633136 333338
rect 632436 333284 633136 333286
rect 632436 333274 632492 333284
rect 631204 330026 631260 330036
rect 625268 328694 625270 328746
rect 625322 328694 625324 328746
rect 625268 328682 625324 328694
rect 635124 328636 635180 333312
rect 635124 328570 635180 328580
rect 637140 328634 637196 333312
rect 637140 328582 637142 328634
rect 637194 328582 637196 328634
rect 637140 328570 637196 328582
rect 638372 333284 639184 333340
rect 638372 325162 638428 333284
rect 641060 326730 641116 333312
rect 643076 328524 643132 333312
rect 643076 328458 643132 328468
rect 641060 326678 641062 326730
rect 641114 326678 641116 326730
rect 641060 326666 641116 326678
rect 638372 325110 638374 325162
rect 638426 325110 638428 325162
rect 638372 325098 638428 325110
rect 645092 325050 645148 333312
rect 647108 326732 647164 333312
rect 649012 332108 649068 333312
rect 649012 332042 649068 332052
rect 650132 333284 651056 333340
rect 647108 326666 647164 326676
rect 650132 325164 650188 333284
rect 653044 332218 653100 333312
rect 653044 332166 653046 332218
rect 653098 332166 653100 332218
rect 653044 332154 653100 332166
rect 655060 328410 655116 333312
rect 658980 331996 659036 333312
rect 658980 331930 659036 331940
rect 660996 328860 661052 333312
rect 660996 328794 661052 328804
rect 661892 333284 663040 333340
rect 655060 328358 655062 328410
rect 655114 328358 655116 328410
rect 655060 328346 655116 328358
rect 650132 325098 650188 325108
rect 645092 324998 645094 325050
rect 645146 324998 645148 325050
rect 645092 324986 645148 324998
rect 661892 324940 661948 333284
rect 664916 328522 664972 333312
rect 666932 329196 666988 333312
rect 666932 329130 666988 329140
rect 668612 333284 668976 333340
rect 670292 333284 670992 333340
rect 664916 328470 664918 328522
rect 664970 328470 664972 328522
rect 664916 328458 664972 328470
rect 668612 325610 668668 333284
rect 668612 325558 668614 325610
rect 668666 325558 668668 325610
rect 668612 325546 668668 325558
rect 661892 324874 661948 324884
rect 670292 308812 670348 333284
rect 672308 332556 672364 332566
rect 672308 332462 672364 332500
rect 671300 332108 671356 332118
rect 670292 308746 670348 308756
rect 671076 331996 671132 332006
rect 657636 306796 657692 306806
rect 655956 305786 656012 305798
rect 655956 305734 655958 305786
rect 656010 305734 656012 305786
rect 655956 301530 656012 305734
rect 655956 301478 655958 301530
rect 656010 301478 656012 301530
rect 655956 301466 656012 301478
rect 657636 301532 657692 306740
rect 660996 306794 661052 306806
rect 660996 306742 660998 306794
rect 661050 306742 661052 306794
rect 659316 306684 659372 306694
rect 659316 301754 659372 306628
rect 659316 301702 659318 301754
rect 659370 301702 659372 301754
rect 659316 301690 659372 301702
rect 660996 301642 661052 306742
rect 660996 301590 660998 301642
rect 661050 301590 661052 301642
rect 660996 301578 661052 301590
rect 662676 306682 662732 306694
rect 662676 306630 662678 306682
rect 662730 306630 662732 306682
rect 662676 301644 662732 306630
rect 662676 301578 662732 301588
rect 670628 301756 670684 301766
rect 657636 301466 657692 301476
rect 670292 301530 670348 301542
rect 670292 301478 670294 301530
rect 670346 301478 670348 301530
rect 654500 299850 654556 299862
rect 654500 299798 654502 299850
rect 654554 299798 654556 299850
rect 624708 294364 624764 294374
rect 618548 294028 618604 294038
rect 613508 292794 613564 292806
rect 613508 292742 613510 292794
rect 613562 292742 613564 292794
rect 613508 292124 613564 292742
rect 613508 292058 613564 292068
rect 617988 292010 618044 292022
rect 617988 291958 617990 292010
rect 618042 291958 618044 292010
rect 612388 291898 612444 291910
rect 612388 291846 612390 291898
rect 612442 291846 612444 291898
rect 612388 290666 612444 291846
rect 615748 291898 615804 291910
rect 615748 291846 615750 291898
rect 615802 291846 615804 291898
rect 612388 290614 612390 290666
rect 612442 290614 612444 290666
rect 612388 290602 612444 290614
rect 612500 290948 612892 291004
rect 612500 290554 612556 290948
rect 612500 290502 612502 290554
rect 612554 290502 612556 290554
rect 612500 290490 612556 290502
rect 612724 290778 612780 290790
rect 612724 290726 612726 290778
rect 612778 290726 612780 290778
rect 611044 290278 611046 290330
rect 611098 290278 611100 290330
rect 611044 290266 611100 290278
rect 610932 289930 610988 289940
rect 611044 289940 612332 289996
rect 610820 288710 610822 288762
rect 610874 288710 610876 288762
rect 610820 288698 610876 288710
rect 610708 288250 610764 288260
rect 611044 288204 611100 289940
rect 611380 289828 611884 289884
rect 611380 289660 611436 289828
rect 611380 289594 611436 289604
rect 611828 289520 611884 289828
rect 612276 289520 612332 289940
rect 612724 289520 612780 290726
rect 612836 290554 612892 290948
rect 612836 290502 612838 290554
rect 612890 290502 612892 290554
rect 612836 290490 612892 290502
rect 614404 290668 614460 290678
rect 613172 290218 613228 290230
rect 613172 290166 613174 290218
rect 613226 290166 613228 290218
rect 613172 289520 613228 290166
rect 613732 290106 613788 290118
rect 613732 290054 613734 290106
rect 613786 290054 613788 290106
rect 613732 289520 613788 290054
rect 614180 290108 614236 290118
rect 614180 289520 614236 290052
rect 614404 289996 614460 290612
rect 615748 290666 615804 291846
rect 615748 290614 615750 290666
rect 615802 290614 615804 290666
rect 615748 290602 615804 290614
rect 615412 290556 615468 290566
rect 615300 290444 615356 290454
rect 615076 290388 615300 290444
rect 614740 290332 614796 290342
rect 614740 290238 614796 290276
rect 614852 290220 614908 290230
rect 614404 289940 614684 289996
rect 614628 289520 614684 289940
rect 614852 289884 614908 290164
rect 615076 289884 615132 290388
rect 615300 290378 615356 290388
rect 614852 289828 615132 289884
rect 615188 290218 615244 290230
rect 615188 290166 615190 290218
rect 615242 290166 615244 290218
rect 615188 289520 615244 290166
rect 615412 289884 615468 290500
rect 615636 290556 615692 290566
rect 615636 290218 615692 290500
rect 617092 290556 617148 290566
rect 615636 290166 615638 290218
rect 615690 290166 615692 290218
rect 615636 290154 615692 290166
rect 616084 290444 616140 290454
rect 615412 289828 615692 289884
rect 615636 289520 615692 289828
rect 616084 289520 616140 290388
rect 616532 290220 616588 290230
rect 616532 289520 616588 290164
rect 617092 289520 617148 290500
rect 617540 290108 617596 290118
rect 617540 289520 617596 290052
rect 617988 289520 618044 291958
rect 618548 289520 618604 293972
rect 621908 293692 621964 293702
rect 620900 292124 620956 292134
rect 620676 291786 620732 291798
rect 620676 291734 620678 291786
rect 620730 291734 620732 291786
rect 620676 290778 620732 291734
rect 620676 290726 620678 290778
rect 620730 290726 620732 290778
rect 620676 290714 620732 290726
rect 618996 290554 619052 290566
rect 618996 290502 618998 290554
rect 619050 290502 619052 290554
rect 618996 289520 619052 290502
rect 619444 290442 619500 290454
rect 619444 290390 619446 290442
rect 619498 290390 619500 290442
rect 619444 289520 619500 290390
rect 619892 290444 619948 290454
rect 619892 289520 619948 290388
rect 620452 290220 620508 290230
rect 620452 289520 620508 290164
rect 620900 289520 620956 292068
rect 621348 291900 621404 291910
rect 621348 289520 621404 291844
rect 621908 289520 621964 293636
rect 624260 292570 624316 292582
rect 624260 292518 624262 292570
rect 624314 292518 624316 292570
rect 622356 292458 622412 292470
rect 622356 292406 622358 292458
rect 622410 292406 622412 292458
rect 622356 289520 622412 292406
rect 623812 292460 623868 292470
rect 622804 289772 622860 289782
rect 622804 289520 622860 289716
rect 623252 289772 623308 289782
rect 623252 289520 623308 289716
rect 623812 289520 623868 292404
rect 624260 289520 624316 292518
rect 624708 289520 624764 294308
rect 625268 294252 625324 294262
rect 625268 289520 625324 294196
rect 645428 293466 645484 293478
rect 645428 293414 645430 293466
rect 645482 293414 645484 293466
rect 631428 293354 631484 293366
rect 631428 293302 631430 293354
rect 631482 293302 631484 293354
rect 630980 293242 631036 293254
rect 630980 293190 630982 293242
rect 631034 293190 631036 293242
rect 629524 293018 629580 293030
rect 629524 292966 629526 293018
rect 629578 292966 629580 293018
rect 628628 292796 628684 292806
rect 627172 292572 627228 292582
rect 626612 291788 626668 291798
rect 625716 291674 625772 291686
rect 625716 291622 625718 291674
rect 625770 291622 625772 291674
rect 625716 289520 625772 291622
rect 626164 289772 626220 289782
rect 626164 289520 626220 289716
rect 626612 289520 626668 291732
rect 627172 289520 627228 292516
rect 627620 290890 627676 290902
rect 627620 290838 627622 290890
rect 627674 290838 627676 290890
rect 627620 289520 627676 290838
rect 628068 289772 628124 289782
rect 628068 289520 628124 289716
rect 628628 289520 628684 292740
rect 629076 289772 629132 289782
rect 629076 289520 629132 289716
rect 629524 289520 629580 292966
rect 630532 292906 630588 292918
rect 630532 292854 630534 292906
rect 630586 292854 630588 292906
rect 629972 291002 630028 291014
rect 629972 290950 629974 291002
rect 630026 290950 630028 291002
rect 629972 289520 630028 290950
rect 630532 289520 630588 292854
rect 630980 289520 631036 293190
rect 631428 289520 631484 293302
rect 643972 292346 644028 292358
rect 643972 292294 643974 292346
rect 644026 292294 644028 292346
rect 642068 291676 642124 291686
rect 635348 291562 635404 291574
rect 635348 291510 635350 291562
rect 635402 291510 635404 291562
rect 633332 291340 633388 291350
rect 632884 291228 632940 291238
rect 632436 291116 632492 291126
rect 631988 289772 632044 289782
rect 631988 289520 632044 289716
rect 632436 289520 632492 291060
rect 632884 289520 632940 291172
rect 633332 289520 633388 291284
rect 634788 291338 634844 291350
rect 634788 291286 634790 291338
rect 634842 291286 634844 291338
rect 634340 291226 634396 291238
rect 634340 291174 634342 291226
rect 634394 291174 634396 291226
rect 633892 291114 633948 291126
rect 633892 291062 633894 291114
rect 633946 291062 633948 291114
rect 633892 289520 633948 291062
rect 634340 289520 634396 291174
rect 634788 289520 634844 291286
rect 635348 289520 635404 291510
rect 639604 291564 639660 291574
rect 635796 291450 635852 291462
rect 635796 291398 635798 291450
rect 635850 291398 635852 291450
rect 635796 289520 635852 291398
rect 637700 291452 637756 291462
rect 637252 290556 637308 290566
rect 636244 289772 636300 289782
rect 636244 289520 636300 289716
rect 636692 289772 636748 289782
rect 636692 289520 636748 289716
rect 637252 289520 637308 290500
rect 637700 289520 637756 291396
rect 639156 290892 639212 290902
rect 638148 289772 638204 289782
rect 638148 289520 638204 289716
rect 638708 289772 638764 289782
rect 638708 289520 638764 289716
rect 639156 289520 639212 290836
rect 639604 289520 639660 291508
rect 640052 289772 640108 289782
rect 640052 289520 640108 289716
rect 640612 289772 640668 289782
rect 640612 289520 640668 289716
rect 641060 289772 641116 289782
rect 641060 289520 641116 289716
rect 641508 289772 641564 289782
rect 641508 289520 641564 289716
rect 642068 289520 642124 291620
rect 642964 290780 643020 290790
rect 642740 290108 642796 290118
rect 642516 289772 642572 289782
rect 642516 289520 642572 289716
rect 642740 289772 642796 290052
rect 642740 289706 642796 289716
rect 642964 289520 643020 290724
rect 643524 290556 643580 290566
rect 643524 289520 643580 290500
rect 643972 289520 644028 292294
rect 644868 291004 644924 291014
rect 644420 289772 644476 289782
rect 644420 289520 644476 289716
rect 644868 289520 644924 290948
rect 645428 289520 645484 293414
rect 648788 291676 648844 291686
rect 647332 291564 647388 291574
rect 645876 291452 645932 291462
rect 645876 289520 645932 291396
rect 646884 290108 646940 290118
rect 646884 289520 646940 290052
rect 647332 289520 647388 291508
rect 648228 290220 648284 290230
rect 648228 289520 648284 290164
rect 648788 289520 648844 291620
rect 651140 290554 651196 290566
rect 651140 290502 651142 290554
rect 651194 290502 651196 290554
rect 650244 290442 650300 290454
rect 650244 290390 650246 290442
rect 650298 290390 650300 290442
rect 649684 290106 649740 290118
rect 649684 290054 649686 290106
rect 649738 290054 649740 290106
rect 649684 289520 649740 290054
rect 650244 289520 650300 290390
rect 651140 289520 651196 290502
rect 654052 290218 654108 290230
rect 654052 290166 654054 290218
rect 654106 290166 654108 290218
rect 651588 289884 651644 289894
rect 651588 289520 651644 289828
rect 652596 289884 652652 289894
rect 652596 289520 652652 289828
rect 653044 289772 653100 289782
rect 653044 289520 653100 289716
rect 654052 289520 654108 290166
rect 654500 289520 654556 299798
rect 669396 292012 669452 292022
rect 658868 290668 658924 290678
rect 655956 290330 656012 290342
rect 655956 290278 655958 290330
rect 656010 290278 656012 290330
rect 655508 289772 655564 289782
rect 655508 289520 655564 289716
rect 655956 289520 656012 290278
rect 656964 289996 657020 290006
rect 656964 289520 657020 289940
rect 657412 289884 657468 289894
rect 657412 289520 657468 289828
rect 658308 289772 658364 289782
rect 658308 289520 658364 289716
rect 658868 289520 658924 290612
rect 668388 290556 668444 290566
rect 666036 290444 666092 290454
rect 662676 290220 662732 290230
rect 659764 289994 659820 290006
rect 659764 289942 659766 289994
rect 659818 289942 659820 289994
rect 659764 289520 659820 289942
rect 660324 289994 660380 290006
rect 660324 289942 660326 289994
rect 660378 289942 660380 289994
rect 660324 289520 660380 289942
rect 661220 289882 661276 289894
rect 661220 289830 661222 289882
rect 661274 289830 661276 289882
rect 661220 289520 661276 289830
rect 661668 289772 661724 289782
rect 661668 289520 661724 289716
rect 662676 289520 662732 290164
rect 664132 290108 664188 290118
rect 663124 289884 663180 289894
rect 663124 289520 663180 289828
rect 664132 289520 664188 290052
rect 664580 289882 664636 289894
rect 664580 289830 664582 289882
rect 664634 289830 664636 289882
rect 664580 289520 664636 289830
rect 665588 289770 665644 289782
rect 665588 289718 665590 289770
rect 665642 289718 665644 289770
rect 665588 289520 665644 289718
rect 666036 289520 666092 290388
rect 668164 290218 668220 290230
rect 668164 290166 668166 290218
rect 668218 290166 668220 290218
rect 667156 290108 667212 290118
rect 667156 289884 667212 290052
rect 666932 289828 667212 289884
rect 666932 289772 666988 289828
rect 667268 289772 667324 289782
rect 666932 289706 666988 289716
rect 667044 289716 667268 289772
rect 667044 289520 667100 289716
rect 667268 289706 667324 289716
rect 667492 289772 667548 289782
rect 667492 289520 667548 289716
rect 667940 289770 667996 289782
rect 667940 289718 667942 289770
rect 667994 289718 667996 289770
rect 667940 289520 667996 289718
rect 668164 289658 668220 290166
rect 668164 289606 668166 289658
rect 668218 289606 668220 289658
rect 668164 289594 668220 289606
rect 668388 289520 668444 290500
rect 668948 289770 669004 289782
rect 668948 289718 668950 289770
rect 669002 289718 669004 289770
rect 668948 289520 669004 289718
rect 669396 289520 669452 291956
rect 669844 290778 669900 290790
rect 669844 290726 669846 290778
rect 669898 290726 669900 290778
rect 669844 289520 669900 290726
rect 670068 290668 670124 290678
rect 670068 290330 670124 290612
rect 670068 290278 670070 290330
rect 670122 290278 670124 290330
rect 670068 290266 670124 290278
rect 670292 290218 670348 301478
rect 670292 290166 670294 290218
rect 670346 290166 670348 290218
rect 670292 290154 670348 290166
rect 670404 294026 670460 294038
rect 670404 293974 670406 294026
rect 670458 293974 670460 294026
rect 670292 289884 670348 289894
rect 670292 289770 670348 289828
rect 670292 289718 670294 289770
rect 670346 289718 670348 289770
rect 670292 289706 670348 289718
rect 670404 289520 670460 293974
rect 670628 289882 670684 301700
rect 670740 301754 670796 301766
rect 670740 301702 670742 301754
rect 670794 301702 670796 301754
rect 670740 290330 670796 301702
rect 670740 290278 670742 290330
rect 670794 290278 670796 290330
rect 670740 290266 670796 290278
rect 670964 301642 671020 301654
rect 670964 301590 670966 301642
rect 671018 301590 671020 301642
rect 670964 289994 671020 301590
rect 671076 291564 671132 331940
rect 671076 291498 671132 291508
rect 671188 301644 671244 301654
rect 670964 289942 670966 289994
rect 671018 289942 671020 289994
rect 670964 289930 671020 289942
rect 671188 289996 671244 301588
rect 671300 291452 671356 332052
rect 672196 331884 672252 331894
rect 672084 331772 672140 331782
rect 671524 313292 671580 313302
rect 671524 291676 671580 313236
rect 671524 291610 671580 291620
rect 671300 291386 671356 291396
rect 671188 289930 671244 289940
rect 671300 290666 671356 290678
rect 671300 290614 671302 290666
rect 671354 290614 671356 290666
rect 670628 289830 670630 289882
rect 670682 289830 670684 289882
rect 670628 289818 670684 289830
rect 670852 289772 670908 289782
rect 670852 289520 670908 289716
rect 671300 289520 671356 290614
rect 672084 290220 672140 331716
rect 672084 290154 672140 290164
rect 671860 289770 671916 289782
rect 671860 289718 671862 289770
rect 671914 289718 671916 289770
rect 611380 288876 611436 288886
rect 611380 288782 611436 288820
rect 611044 288138 611100 288148
rect 671860 283836 671916 289718
rect 672196 289658 672252 331828
rect 672420 331770 672476 331782
rect 672420 331718 672422 331770
rect 672474 331718 672476 331770
rect 672308 306570 672364 306582
rect 672308 306518 672310 306570
rect 672362 306518 672364 306570
rect 672308 289884 672364 306518
rect 672420 290332 672476 331718
rect 672868 328412 672924 333312
rect 673652 333284 674912 333340
rect 672868 328346 672924 328356
rect 673204 332668 673260 332678
rect 673204 308810 673260 332612
rect 673652 325052 673708 333284
rect 676900 331882 676956 333312
rect 678916 332668 678972 333312
rect 678916 332602 678972 332612
rect 680372 333284 680848 333340
rect 682052 333284 682864 333340
rect 683732 333284 684880 333340
rect 676900 331830 676902 331882
rect 676954 331830 676956 331882
rect 676900 331818 676956 331830
rect 673652 324986 673708 324996
rect 680372 322588 680428 333284
rect 682052 324044 682108 333284
rect 683732 324156 683788 333284
rect 683732 324090 683788 324100
rect 682052 323978 682108 323988
rect 680372 322522 680428 322532
rect 673204 308758 673206 308810
rect 673258 308758 673260 308810
rect 673204 308746 673260 308758
rect 672420 290266 672476 290276
rect 672308 289818 672364 289828
rect 672196 289606 672198 289658
rect 672250 289606 672252 289658
rect 672196 289594 672252 289606
rect 671860 283770 671916 283780
rect 609924 283098 609980 283108
rect 605556 281596 605612 281606
rect 603876 274764 603932 274774
rect 602308 272524 602364 272534
rect 602196 268044 602252 268054
rect 600628 265692 600684 265702
rect 600628 248780 600684 265636
rect 602196 252140 602252 267988
rect 602308 257068 602364 272468
rect 603876 260428 603932 274708
rect 605556 270396 605612 281540
rect 605556 270330 605612 270340
rect 607236 279356 607292 279366
rect 607236 267148 607292 279300
rect 607236 267082 607292 267092
rect 603876 260362 603932 260372
rect 602308 257002 602364 257012
rect 602196 252074 602252 252084
rect 600628 248714 600684 248724
rect 605556 183932 605612 183942
rect 603876 177100 603932 177110
rect 600628 161196 600684 161206
rect 600628 107548 600684 161140
rect 603876 127708 603932 177044
rect 603876 127642 603932 127652
rect 603988 170268 604044 170278
rect 603988 122668 604044 170212
rect 605556 139468 605612 183876
rect 605556 139402 605612 139412
rect 605668 174860 605724 174870
rect 605668 131068 605724 174804
rect 671748 154588 671804 154598
rect 671748 141148 671804 154532
rect 671860 149996 671916 150006
rect 671860 142156 671916 149940
rect 672756 147644 672812 147654
rect 671860 142090 671916 142100
rect 672196 143052 672252 143062
rect 671748 141082 671804 141092
rect 671972 141596 672028 141606
rect 611716 140140 611772 140150
rect 605668 131002 605724 131012
rect 611492 131852 611548 131862
rect 603988 122602 604044 122612
rect 600628 107482 600684 107492
rect 600516 82182 600518 82234
rect 600570 82182 600572 82234
rect 600516 82170 600572 82182
rect 586068 81386 586124 81396
rect 585844 81274 585900 81284
rect 585620 81162 585676 81172
rect 560308 80614 560310 80666
rect 560362 80614 560364 80666
rect 560308 80602 560364 80614
rect 560196 79034 560252 79044
rect 561876 78988 561932 78998
rect 526372 72090 526428 72100
rect 560980 72156 561036 72166
rect 459172 71978 459228 71988
rect 506772 71932 506828 71942
rect 392084 71754 392140 71764
rect 469140 71818 469196 71830
rect 469140 71766 469142 71818
rect 469194 71766 469196 71818
rect 450996 71706 451052 71718
rect 450996 71654 450998 71706
rect 451050 71654 451052 71706
rect 439908 71594 439964 71606
rect 439908 71542 439910 71594
rect 439962 71542 439964 71594
rect 341684 71484 341740 71494
rect 257796 70522 257852 70532
rect 340900 71370 340956 71382
rect 340900 71318 340902 71370
rect 340954 71318 340956 71370
rect 340900 70252 340956 71318
rect 340890 70196 340956 70252
rect 176182 70140 176238 70150
rect 176182 70074 176238 70084
rect 231182 70140 231238 70150
rect 340890 70112 340946 70196
rect 341684 70140 341740 71428
rect 395892 71482 395948 71494
rect 395892 71430 395894 71482
rect 395946 71430 395948 71482
rect 395892 70252 395948 71430
rect 341064 70084 341740 70140
rect 395890 70196 395948 70252
rect 396036 70588 396092 70598
rect 395890 70112 395946 70196
rect 396036 70112 396092 70532
rect 439908 70140 439964 71542
rect 450996 70476 451052 71654
rect 454580 71708 454636 71718
rect 450996 70420 451092 70476
rect 439315 70084 439964 70140
rect 451036 70112 451092 70420
rect 451181 70140 451237 70150
rect 231182 70074 231238 70084
rect 451181 70074 451237 70084
rect 454580 70140 454636 71652
rect 454580 70074 454636 70084
rect 450890 69804 450946 69814
rect 450890 69738 450946 69748
rect 469140 69804 469196 71766
rect 494287 70140 494343 70150
rect 494287 70074 494343 70084
rect 505890 70140 505946 70150
rect 506772 70140 506828 71876
rect 548548 71820 548604 71830
rect 548548 70700 548604 71764
rect 560980 70700 561036 72100
rect 548548 70644 548630 70700
rect 560980 70644 561092 70700
rect 506210 70084 506828 70140
rect 548432 70140 548488 70150
rect 548574 70112 548630 70644
rect 560890 70588 560946 70598
rect 549287 70364 549343 70374
rect 549287 70112 549343 70308
rect 560890 70112 560946 70532
rect 561036 70112 561092 70644
rect 561876 70140 561932 78932
rect 611492 71596 611548 131796
rect 611716 80666 611772 140084
rect 624036 140140 624092 140150
rect 624036 140074 624092 140084
rect 619108 140028 619164 140038
rect 618884 139916 618940 139926
rect 611716 80614 611718 80666
rect 611770 80614 611772 80666
rect 611716 80602 611772 80614
rect 611492 71530 611548 71540
rect 611940 71482 611996 139664
rect 612164 139636 612640 139692
rect 612164 131852 612220 139636
rect 612164 131786 612220 131796
rect 611940 71430 611942 71482
rect 611994 71430 611996 71482
rect 611940 71418 611996 71430
rect 613284 71370 613340 139664
rect 613956 71484 614012 139664
rect 614628 71708 614684 139664
rect 615300 71818 615356 139664
rect 615300 71766 615302 71818
rect 615354 71766 615356 71818
rect 615300 71754 615356 71766
rect 614628 71642 614684 71652
rect 615972 71594 616028 139664
rect 616644 71706 616700 139664
rect 617316 71932 617372 139664
rect 617316 71866 617372 71876
rect 616644 71654 616646 71706
rect 616698 71654 616700 71706
rect 616644 71642 616700 71654
rect 615972 71542 615974 71594
rect 616026 71542 616028 71594
rect 615972 71530 616028 71542
rect 613956 71418 614012 71428
rect 613284 71318 613286 71370
rect 613338 71318 613340 71370
rect 613284 71306 613340 71318
rect 617988 71036 618044 139664
rect 618436 139636 618688 139692
rect 618324 134652 618380 134662
rect 618324 89964 618380 134596
rect 618436 134428 618492 139636
rect 618436 134362 618492 134372
rect 618548 139468 618604 139478
rect 618548 132747 618604 139412
rect 618324 89898 618380 89908
rect 618436 132691 618604 132747
rect 618436 86268 618492 132691
rect 618436 86202 618492 86212
rect 618548 123114 618604 123126
rect 618548 123062 618550 123114
rect 618602 123062 618604 123114
rect 618548 81340 618604 123062
rect 618660 122668 618716 122678
rect 618660 82572 618716 122612
rect 618884 93772 618940 139860
rect 618996 139466 619052 139478
rect 618996 139414 618998 139466
rect 619050 139414 619052 139466
rect 618996 96236 619052 139414
rect 619108 139468 619164 139972
rect 623364 140028 623420 140038
rect 623364 139962 623420 139972
rect 624708 140028 624764 140038
rect 624708 139962 624764 139972
rect 657076 140028 657132 140038
rect 657076 139962 657132 139972
rect 657748 140028 657804 140038
rect 657748 139962 657804 139972
rect 630756 139916 630812 139926
rect 630756 139850 630812 139860
rect 631428 139916 631484 139926
rect 631428 139850 631484 139860
rect 647892 139916 647948 139926
rect 655732 139916 655788 139926
rect 647892 139914 648368 139916
rect 647892 139862 647894 139914
rect 647946 139888 648368 139914
rect 647946 139862 648396 139888
rect 647892 139860 648396 139862
rect 647892 139850 647948 139860
rect 619780 139802 619836 139814
rect 619780 139750 619782 139802
rect 619834 139750 619836 139802
rect 619108 139402 619164 139412
rect 618996 96170 619052 96180
rect 619108 125468 619164 125478
rect 618884 93706 618940 93716
rect 619108 92540 619164 125412
rect 619108 92474 619164 92484
rect 618660 82506 618716 82516
rect 618548 81274 618604 81284
rect 619332 71148 619388 139664
rect 619556 139578 619612 139590
rect 619556 139526 619558 139578
rect 619610 139526 619612 139578
rect 619556 99036 619612 139526
rect 619780 100604 619836 139750
rect 621572 139802 621628 139814
rect 621572 139750 621574 139802
rect 621626 139750 621628 139802
rect 620032 139636 620508 139692
rect 620704 139636 621180 139692
rect 620452 134540 620508 139636
rect 620452 134474 620508 134484
rect 621124 134428 621180 139636
rect 621348 134652 621404 139664
rect 621460 139468 621516 139478
rect 621572 139468 621628 139750
rect 622692 139804 622748 139814
rect 622692 139738 622748 139748
rect 634340 139804 634396 139814
rect 634340 139802 634816 139804
rect 634340 139750 634342 139802
rect 634394 139750 634816 139802
rect 634340 139748 634816 139750
rect 634340 139738 634396 139748
rect 622020 139692 622076 139702
rect 632772 139692 632828 139702
rect 633668 139692 633724 139702
rect 638820 139692 638876 139702
rect 622020 139626 622076 139636
rect 624932 139636 625408 139692
rect 624932 139580 624988 139636
rect 624932 139514 624988 139524
rect 621516 139412 621628 139468
rect 621460 139402 621516 139412
rect 621348 134586 621404 134596
rect 621124 134362 621180 134372
rect 626052 125916 626108 139664
rect 626052 125850 626108 125860
rect 626724 125132 626780 139664
rect 627396 125244 627452 139664
rect 628068 125916 628124 139664
rect 628068 125850 628124 125860
rect 628740 125916 628796 139664
rect 628740 125850 628796 125860
rect 629412 125356 629468 139664
rect 630084 125468 630140 139664
rect 632100 139466 632156 139664
rect 632772 139626 632828 139636
rect 633220 139636 633472 139692
rect 633668 139690 634144 139692
rect 633668 139638 633670 139690
rect 633722 139638 634144 139690
rect 633668 139636 634144 139638
rect 633220 139578 633276 139636
rect 633668 139626 633724 139636
rect 633220 139526 633222 139578
rect 633274 139526 633276 139578
rect 633220 139514 633276 139526
rect 632100 139414 632102 139466
rect 632154 139414 632156 139466
rect 632100 139402 632156 139414
rect 635460 135436 635516 139664
rect 636132 135660 636188 139664
rect 636132 135594 636188 135604
rect 635460 135370 635516 135380
rect 636804 135212 636860 139664
rect 637476 135324 637532 139664
rect 638148 135548 638204 139664
rect 638820 139626 638876 139636
rect 638148 135482 638204 135492
rect 637476 135258 637532 135268
rect 636804 135146 636860 135156
rect 630084 125402 630140 125412
rect 639492 125468 639548 139664
rect 640164 125580 640220 139664
rect 640836 125692 640892 139664
rect 641508 125916 641564 139664
rect 642292 126812 642348 139664
rect 642292 126746 642348 126756
rect 641508 125850 641564 125860
rect 642964 125804 643020 139664
rect 643636 127596 643692 139664
rect 643636 127530 643692 127540
rect 644308 126924 644364 139664
rect 644980 127036 645036 139664
rect 645652 127260 645708 139664
rect 646324 127484 646380 139664
rect 646324 127418 646380 127428
rect 645652 127194 645708 127204
rect 644980 126970 645036 126980
rect 644308 126858 644364 126868
rect 646996 126028 647052 139664
rect 646996 125962 647052 125972
rect 647668 126028 647724 139664
rect 648340 131628 648396 139860
rect 655732 139850 655788 139860
rect 665140 139916 665196 139926
rect 665140 139850 665196 139860
rect 659092 139804 659148 139814
rect 659092 139738 659148 139748
rect 650692 139692 650748 139702
rect 652596 139692 652652 139702
rect 656404 139692 656460 139702
rect 666484 139692 666540 139702
rect 648900 139466 648956 139478
rect 648900 139414 648902 139466
rect 648954 139414 648956 139466
rect 648900 132076 648956 139414
rect 649012 139468 649068 139664
rect 649460 139636 649712 139692
rect 650020 139636 650384 139692
rect 650748 139636 651056 139692
rect 649012 139402 649068 139412
rect 649236 139466 649292 139478
rect 649236 139414 649238 139466
rect 649290 139414 649292 139466
rect 649124 139354 649180 139366
rect 649124 139302 649126 139354
rect 649178 139302 649180 139354
rect 649124 132188 649180 139302
rect 649236 132300 649292 139414
rect 649460 136332 649516 139636
rect 649460 136266 649516 136276
rect 650020 134876 650076 139636
rect 650692 139626 650748 139636
rect 651700 139466 651756 139664
rect 651924 139636 652400 139692
rect 652596 139690 653072 139692
rect 652596 139638 652598 139690
rect 652650 139638 653072 139690
rect 652596 139636 653072 139638
rect 651924 139578 651980 139636
rect 652596 139626 652652 139636
rect 651924 139526 651926 139578
rect 651978 139526 651980 139578
rect 651924 139514 651980 139526
rect 651700 139414 651702 139466
rect 651754 139414 651756 139466
rect 651700 139402 651756 139414
rect 653716 136332 653772 139664
rect 653716 136266 653772 136276
rect 654388 136108 654444 139664
rect 655060 136220 655116 139664
rect 656404 139626 656460 139636
rect 658420 139468 658476 139664
rect 659792 139636 660044 139692
rect 659988 139580 660044 139636
rect 659988 139514 660044 139524
rect 658420 139402 658476 139412
rect 660436 138012 660492 139664
rect 661136 139636 661612 139692
rect 660436 137946 660492 137956
rect 661556 136892 661612 139636
rect 661780 137788 661836 139664
rect 662452 137900 662508 139664
rect 663152 139636 663516 139692
rect 662452 137834 662508 137844
rect 661780 137722 661836 137732
rect 663460 137004 663516 139636
rect 663796 138796 663852 139664
rect 664468 139020 664524 139664
rect 665812 139466 665868 139664
rect 667828 139692 667884 139702
rect 668724 139692 668780 139702
rect 666484 139626 666540 139636
rect 665812 139414 665814 139466
rect 665866 139414 665868 139466
rect 665812 139402 665868 139414
rect 667156 139466 667212 139664
rect 668528 139690 668780 139692
rect 668528 139638 668726 139690
rect 668778 139638 668780 139690
rect 668528 139636 668780 139638
rect 669200 139636 669676 139692
rect 667828 139626 667884 139636
rect 668724 139626 668780 139636
rect 667156 139414 667158 139466
rect 667210 139414 667212 139466
rect 667156 139402 667212 139414
rect 669508 139466 669564 139478
rect 669508 139414 669510 139466
rect 669562 139414 669564 139466
rect 664468 138954 664524 138964
rect 663796 138730 663852 138740
rect 663460 136938 663516 136948
rect 661556 136826 661612 136836
rect 655060 136154 655116 136164
rect 654388 136042 654444 136052
rect 669508 134988 669564 139414
rect 669620 139468 669676 139636
rect 669620 139402 669676 139412
rect 669844 139466 669900 139664
rect 670544 139636 671020 139692
rect 669844 139414 669846 139466
rect 669898 139414 669900 139466
rect 669844 139402 669900 139414
rect 670964 137787 671020 139636
rect 671524 139690 671580 139702
rect 671524 139638 671526 139690
rect 671578 139638 671580 139690
rect 671300 139466 671356 139478
rect 671300 139414 671302 139466
rect 671354 139414 671356 139466
rect 670964 137731 671244 137787
rect 669508 134922 669564 134932
rect 650020 134810 650076 134820
rect 671188 133196 671244 137731
rect 671094 133140 671244 133196
rect 650122 133084 650178 133094
rect 650122 133018 650178 133028
rect 649572 132748 649628 132758
rect 649478 132692 649572 132748
rect 649572 132682 649628 132692
rect 654378 132636 654434 132646
rect 654378 132570 654434 132580
rect 656394 132636 656450 132646
rect 656394 132570 656450 132580
rect 657972 132636 658028 132646
rect 664580 132636 664636 132646
rect 658028 132580 658550 132636
rect 664150 132580 664580 132636
rect 657972 132570 658028 132580
rect 664580 132570 664636 132580
rect 666922 132636 666978 132646
rect 666922 132570 666978 132580
rect 667594 132636 667650 132646
rect 670180 132636 670236 132646
rect 669750 132580 670180 132636
rect 667594 132570 667650 132580
rect 670180 132570 670236 132580
rect 654836 132524 654892 132534
rect 659652 132524 659708 132534
rect 661994 132524 662050 132534
rect 668266 132524 668322 132534
rect 650692 132468 650934 132524
rect 650692 132412 650748 132468
rect 650692 132346 650748 132356
rect 649236 132234 649292 132244
rect 651578 132300 651634 132496
rect 651578 132234 651634 132244
rect 649124 132122 649180 132132
rect 652250 132188 652306 132496
rect 652250 132122 652306 132132
rect 648900 132010 648956 132020
rect 652922 132076 652978 132496
rect 653604 132198 653660 132524
rect 654892 132468 655078 132524
rect 654836 132458 654892 132468
rect 655722 132300 655778 132496
rect 655722 132234 655778 132244
rect 653594 132188 653660 132198
rect 653650 132132 653660 132188
rect 657178 132188 657234 132496
rect 653594 132122 653650 132132
rect 657178 132122 657234 132132
rect 652922 132010 652978 132020
rect 657850 132076 657906 132496
rect 659222 132468 659652 132524
rect 659894 132468 660156 132524
rect 659652 132458 659708 132468
rect 657850 132010 657906 132020
rect 648340 131562 648396 131572
rect 654724 131628 654780 131638
rect 647668 125962 647724 125972
rect 642964 125738 643020 125748
rect 640836 125626 640892 125636
rect 640164 125514 640220 125524
rect 639492 125402 639548 125412
rect 629412 125290 629468 125300
rect 627396 125178 627452 125188
rect 626724 125066 626780 125076
rect 627508 123562 627564 123574
rect 633108 123564 633164 123574
rect 627508 123510 627510 123562
rect 627562 123510 627564 123562
rect 627284 123452 627340 123462
rect 627284 123386 627340 123396
rect 622132 123340 622188 123350
rect 622132 123274 622188 123284
rect 627508 123338 627564 123510
rect 632464 123562 633164 123564
rect 632464 123510 633110 123562
rect 633162 123510 633164 123562
rect 632464 123508 633164 123510
rect 633108 123498 633164 123508
rect 654724 123562 654780 131572
rect 660100 131516 660156 132468
rect 660650 132300 660706 132496
rect 660650 132234 660706 132244
rect 661322 132188 661378 132496
rect 662694 132468 663292 132524
rect 661994 132458 662050 132468
rect 661322 132122 661378 132132
rect 660100 131450 660156 131460
rect 663236 131404 663292 132468
rect 663460 131852 663516 132524
rect 664822 132468 665196 132524
rect 665494 132468 665980 132524
rect 666166 132468 666652 132524
rect 663460 131786 663516 131796
rect 663236 131338 663292 131348
rect 665140 131068 665196 132468
rect 665924 131964 665980 132468
rect 665924 131898 665980 131908
rect 666596 131740 666652 132468
rect 668266 132458 668322 132468
rect 668938 132076 668994 132496
rect 670422 132468 670908 132524
rect 670852 132300 670908 132468
rect 671300 132300 671356 139414
rect 670852 132244 671356 132300
rect 668938 132010 668994 132020
rect 671524 132076 671580 139638
rect 671524 132010 671580 132020
rect 671636 139578 671692 139590
rect 671636 139526 671638 139578
rect 671690 139526 671692 139578
rect 666596 131674 666652 131684
rect 671636 131740 671692 139526
rect 671636 131674 671692 131684
rect 665140 131002 665196 131012
rect 655396 127260 655452 127270
rect 655172 127036 655228 127046
rect 654724 123510 654726 123562
rect 654778 123510 654780 123562
rect 654724 123498 654780 123510
rect 654948 125244 655004 125254
rect 627508 123286 627510 123338
rect 627562 123286 627564 123338
rect 627508 123274 627564 123286
rect 636916 123340 636972 123350
rect 641172 123340 641228 123378
rect 636916 123338 637616 123340
rect 636916 123286 636918 123338
rect 636970 123286 637616 123338
rect 636916 123284 637616 123286
rect 636916 123274 636972 123284
rect 641172 123274 641228 123284
rect 642740 123340 642796 123350
rect 642740 123274 642796 123284
rect 647892 123340 647948 123350
rect 647892 123274 647948 123284
rect 652372 123340 652428 123350
rect 652372 123338 653072 123340
rect 652372 123286 652374 123338
rect 652426 123286 653072 123338
rect 652372 123284 653072 123286
rect 652372 123274 652428 123284
rect 654948 116620 655004 125188
rect 654948 116554 655004 116564
rect 655060 125132 655116 125142
rect 655060 115052 655116 125076
rect 655060 114986 655116 114996
rect 619780 100538 619836 100548
rect 620564 100716 620620 100726
rect 620564 100492 620620 100660
rect 625380 100716 625436 100726
rect 623364 100492 623420 100502
rect 620564 100436 620816 100492
rect 625380 100492 625436 100660
rect 647556 100716 647612 100726
rect 628628 100492 628684 100502
rect 625380 100436 625968 100492
rect 623364 100426 623420 100436
rect 628628 100426 628684 100436
rect 631204 100492 631260 100502
rect 647556 100492 647612 100660
rect 646912 100436 647612 100492
rect 649572 100492 649628 100502
rect 631204 100426 631260 100436
rect 649572 100426 649628 100436
rect 652148 100492 652204 100502
rect 652148 100426 652204 100436
rect 633780 100044 633836 100054
rect 633780 99978 633836 99988
rect 635796 100044 635852 100054
rect 639044 100044 639100 100054
rect 635852 99988 636496 100044
rect 635796 99978 635852 99988
rect 639044 99978 639100 99988
rect 641732 100044 641788 100054
rect 644980 100044 645036 100054
rect 644336 99988 644980 100044
rect 641732 99978 641788 99988
rect 644980 99978 645036 99988
rect 619556 98970 619612 98980
rect 655172 92316 655228 126980
rect 655284 126924 655340 126934
rect 655284 109676 655340 126868
rect 655396 110236 655452 127204
rect 655396 110170 655452 110180
rect 655956 126700 656012 126710
rect 655284 109610 655340 109620
rect 655172 92250 655228 92260
rect 655956 85596 656012 126644
rect 670180 123564 670236 123574
rect 670180 123498 670236 123508
rect 655956 85530 656012 85540
rect 671972 80890 672028 141540
rect 671972 80838 671974 80890
rect 672026 80838 672028 80890
rect 628068 80668 628124 80678
rect 628068 80602 628124 80612
rect 645092 80668 645148 80678
rect 645092 80602 645148 80612
rect 671972 74508 672028 80838
rect 671972 74442 672028 74452
rect 672084 140812 672140 140822
rect 672084 81002 672140 140756
rect 672196 83468 672252 142996
rect 672196 83402 672252 83412
rect 672084 80950 672086 81002
rect 672138 80950 672140 81002
rect 672084 74284 672140 80950
rect 672084 74218 672140 74228
rect 672756 74060 672812 147588
rect 673540 142716 673596 142726
rect 673540 94108 673596 142660
rect 673540 94042 673596 94052
rect 686308 90748 686364 366884
rect 686420 176428 686476 446852
rect 686420 176362 686476 176372
rect 686532 353612 686588 353622
rect 686532 90860 686588 353556
rect 686644 334012 686700 593460
rect 686868 513996 686924 514006
rect 686644 333946 686700 333956
rect 686756 473788 686812 473798
rect 686756 218428 686812 473732
rect 686868 262220 686924 513940
rect 686868 262154 686924 262164
rect 686980 336028 687036 336038
rect 686756 218362 686812 218372
rect 686980 132748 687036 335972
rect 687204 274540 687260 937076
rect 687316 936906 687372 936918
rect 687316 936854 687318 936906
rect 687370 936854 687372 936906
rect 687316 281484 687372 936854
rect 687428 289770 687484 937188
rect 687652 936794 687708 936806
rect 687652 936742 687654 936794
rect 687706 936742 687708 936794
rect 687428 289718 687430 289770
rect 687482 289718 687484 289770
rect 687428 289706 687484 289718
rect 687540 936682 687596 936694
rect 687540 936630 687542 936682
rect 687594 936630 687596 936682
rect 687540 289212 687596 936630
rect 687652 289772 687708 936742
rect 687764 313292 687820 938198
rect 688212 937356 688268 937366
rect 688212 937262 688268 937300
rect 688996 937244 689052 937254
rect 688436 937020 688492 937030
rect 688212 936796 688268 936806
rect 687876 936684 687932 936694
rect 687876 331996 687932 936628
rect 687988 936572 688044 936582
rect 687988 332108 688044 936516
rect 688100 936570 688156 936582
rect 688100 936518 688102 936570
rect 688154 936518 688156 936570
rect 688100 333450 688156 936518
rect 688100 333398 688102 333450
rect 688154 333398 688156 333450
rect 688100 333386 688156 333398
rect 688212 333452 688268 936740
rect 688212 333386 688268 333396
rect 688324 672812 688380 672822
rect 687988 332042 688044 332052
rect 687876 331930 687932 331940
rect 687764 313226 687820 313236
rect 688212 290444 688268 290454
rect 688212 290350 688268 290388
rect 687652 289706 687708 289716
rect 687540 289146 687596 289156
rect 687316 281418 687372 281428
rect 687204 274474 687260 274484
rect 688324 260764 688380 672756
rect 688436 267708 688492 936964
rect 688884 936460 688940 936470
rect 688884 290106 688940 936404
rect 688996 672812 689052 937188
rect 688996 672746 689052 672756
rect 689220 937018 689276 937030
rect 689220 936966 689222 937018
rect 689274 936966 689276 937018
rect 688996 580748 689052 580758
rect 688996 334236 689052 580692
rect 689108 394156 689164 394166
rect 689108 336028 689164 394100
rect 689108 335962 689164 335972
rect 688996 334170 689052 334180
rect 688884 290054 688886 290106
rect 688938 290054 688940 290106
rect 688884 290042 688940 290054
rect 689220 269948 689276 936966
rect 695380 935564 695436 935574
rect 694820 934892 694876 934902
rect 694708 934780 694764 934790
rect 693812 934556 693868 934566
rect 691348 910812 691404 910822
rect 689556 910588 689612 910598
rect 689332 290556 689388 290566
rect 689332 290462 689388 290500
rect 689220 269882 689276 269892
rect 688436 267642 688492 267652
rect 688324 260698 688380 260708
rect 689556 249228 689612 910532
rect 691236 908572 691292 908582
rect 689556 249162 689612 249172
rect 689668 824908 689724 824918
rect 689668 235340 689724 824852
rect 689780 739228 689836 739238
rect 689780 242284 689836 739172
rect 689780 242218 689836 242228
rect 689892 695548 689948 695558
rect 689668 235274 689724 235284
rect 689892 228396 689948 695492
rect 689892 228330 689948 228340
rect 690004 651868 690060 651878
rect 690004 221564 690060 651812
rect 690004 221498 690060 221508
rect 690116 566188 690172 566198
rect 690116 207676 690172 566132
rect 690116 207610 690172 207620
rect 690228 524188 690284 524198
rect 690228 200732 690284 524132
rect 691236 253820 691292 908516
rect 691348 900844 691404 910756
rect 691348 900778 691404 900788
rect 693028 860748 693084 860758
rect 691236 253754 691292 253764
rect 692916 822556 692972 822566
rect 692916 239932 692972 822500
rect 693028 806988 693084 860692
rect 693812 823004 693868 934500
rect 693812 822938 693868 822948
rect 694484 934332 694540 934342
rect 693028 806922 693084 806932
rect 693028 780780 693084 780790
rect 693028 719852 693084 780724
rect 693028 719786 693084 719796
rect 694484 609756 694540 934276
rect 694596 873628 694652 873638
rect 694596 736092 694652 873572
rect 694596 736026 694652 736036
rect 694484 609690 694540 609700
rect 694596 607516 694652 607526
rect 693140 500780 693196 500790
rect 692916 239866 692972 239876
rect 693028 420812 693084 420822
rect 690228 200666 690284 200676
rect 693028 179788 693084 420756
rect 693140 265804 693196 500724
rect 693140 265738 693196 265748
rect 693252 460796 693308 460806
rect 693252 236794 693308 460740
rect 693252 236742 693254 236794
rect 693306 236742 693308 236794
rect 693252 236730 693308 236742
rect 694596 219212 694652 607460
rect 694708 566860 694764 934724
rect 694820 822108 694876 934836
rect 694820 822042 694876 822052
rect 695156 934444 695212 934454
rect 694708 566794 694764 566804
rect 694820 693084 694876 693094
rect 694596 219146 694652 219156
rect 694708 564508 694764 564518
rect 694708 212268 694764 564452
rect 694820 334124 694876 693028
rect 695156 607964 695212 934388
rect 695156 607898 695212 607908
rect 694820 334058 694876 334068
rect 694932 566748 694988 566758
rect 694932 307020 694988 566692
rect 695380 522060 695436 935508
rect 697956 925148 698012 947492
rect 697956 925082 698012 925092
rect 700532 934668 700588 934678
rect 700532 908124 700588 934612
rect 705012 927276 705068 927286
rect 703892 927164 703948 927174
rect 705012 927164 705068 927220
rect 703948 927108 704416 927164
rect 705012 927108 705312 927164
rect 703892 927098 703948 927108
rect 704836 926380 704892 926390
rect 704836 926314 704892 926324
rect 705732 926380 705788 926390
rect 705732 926314 705788 926324
rect 700532 908058 700588 908068
rect 699188 891548 699244 891558
rect 696276 887068 696332 887078
rect 696276 736988 696332 887012
rect 696276 736922 696332 736932
rect 698740 840588 698796 840598
rect 698740 720188 698796 840532
rect 699188 752556 699244 891492
rect 700196 891436 700252 891446
rect 699748 891324 699804 891334
rect 699412 890652 699468 890662
rect 699188 752490 699244 752500
rect 699300 805532 699356 805542
rect 698740 720122 698796 720132
rect 699300 712124 699356 805476
rect 699412 752556 699468 890596
rect 699748 806428 699804 891268
rect 700084 838348 700140 838358
rect 699972 823116 700028 823126
rect 699748 806362 699804 806372
rect 699860 821884 699916 821894
rect 699412 752490 699468 752500
rect 699524 805420 699580 805430
rect 699524 712236 699580 805364
rect 699524 712170 699580 712180
rect 699748 804972 699804 804982
rect 699300 712058 699356 712068
rect 699748 710556 699804 804916
rect 699860 720300 699916 821828
rect 699860 720234 699916 720244
rect 699972 719068 700028 823060
rect 700084 720412 700140 838292
rect 700196 755692 700252 891380
rect 704388 891324 704444 891856
rect 704836 891548 704892 891856
rect 704836 891482 704892 891492
rect 705284 891436 705340 891856
rect 705284 891370 705340 891380
rect 705572 891828 705760 891884
rect 704388 891258 704444 891268
rect 705572 890652 705628 891828
rect 705572 890586 705628 890596
rect 704388 840588 704444 840598
rect 704388 840522 704444 840532
rect 704836 840364 704892 840374
rect 704836 840298 704892 840308
rect 705284 840364 705340 840374
rect 705284 840298 705340 840308
rect 705732 840364 705788 840374
rect 705732 840298 705788 840308
rect 700644 838348 700700 838358
rect 700644 823116 700700 838292
rect 700644 823050 700700 823060
rect 701428 824788 701484 824798
rect 701428 819980 701484 824732
rect 701428 819914 701484 819924
rect 704388 805420 704444 805840
rect 704388 805354 704444 805364
rect 700196 755626 700252 755636
rect 701316 805308 701372 805318
rect 700084 720346 700140 720356
rect 700420 739114 700476 739126
rect 700420 739062 700422 739114
rect 700474 739062 700476 739114
rect 699972 719002 700028 719012
rect 700420 712122 700476 739062
rect 701316 739114 701372 805252
rect 704836 805308 704892 805840
rect 705284 805532 705340 805840
rect 705284 805466 705340 805476
rect 705572 805812 705760 805868
rect 704836 805242 704892 805252
rect 705572 804972 705628 805812
rect 705572 804906 705628 804916
rect 704388 755692 704444 755702
rect 704388 755104 704444 755636
rect 705124 755132 705180 755142
rect 705180 755076 705312 755132
rect 705124 755066 705180 755076
rect 704836 754460 704892 754470
rect 704836 754394 704892 754404
rect 705732 754460 705788 754470
rect 705732 754394 705788 754404
rect 701316 739062 701318 739114
rect 701370 739062 701372 739114
rect 701316 739050 701372 739062
rect 704388 720412 704444 720422
rect 704388 720346 704444 720356
rect 704836 720300 704892 720310
rect 704836 720234 704892 720244
rect 705284 720188 705340 720198
rect 705284 720122 705340 720132
rect 700420 712070 700422 712122
rect 700474 712070 700476 712122
rect 700420 712058 700476 712070
rect 700644 719852 700700 719862
rect 699748 710490 699804 710500
rect 700644 697116 700700 719796
rect 705572 719796 705760 719852
rect 705572 719068 705628 719796
rect 705572 719002 705628 719012
rect 705012 712236 705068 712246
rect 703892 712124 703948 712134
rect 704564 712124 704620 712134
rect 705012 712124 705068 712180
rect 703948 712068 704416 712124
rect 704564 712122 704864 712124
rect 704564 712070 704566 712122
rect 704618 712070 704864 712122
rect 704564 712068 704864 712070
rect 705012 712068 705312 712124
rect 703892 712058 703948 712068
rect 704564 712058 704620 712068
rect 705732 711452 705788 711462
rect 705732 711386 705788 711396
rect 700644 697050 700700 697060
rect 701540 697116 701596 697126
rect 701540 695788 701596 697060
rect 701540 695722 701596 695732
rect 704388 676508 704444 676816
rect 704836 676620 704892 676816
rect 704836 676554 704892 676564
rect 704388 676442 704444 676452
rect 705284 676396 705340 676816
rect 705284 676330 705340 676340
rect 705732 676284 705788 676816
rect 705684 676228 705788 676284
rect 705684 675500 705740 676228
rect 705684 675434 705740 675444
rect 700532 671132 700588 671142
rect 700532 652764 700588 671076
rect 704676 669116 704732 669126
rect 704732 669060 704864 669116
rect 704676 669050 704732 669060
rect 704388 668556 704444 668566
rect 704388 668490 704444 668500
rect 705284 668556 705340 668566
rect 705284 668490 705340 668500
rect 705732 668444 705788 668454
rect 705732 668378 705788 668388
rect 700532 652698 700588 652708
rect 704388 633612 704444 633808
rect 704388 633546 704444 633556
rect 704836 633500 704892 633808
rect 704836 633434 704892 633444
rect 705284 633388 705340 633808
rect 705284 633322 705340 633332
rect 705732 633388 705788 633808
rect 705732 633322 705788 633332
rect 704388 626556 704444 626566
rect 704388 626192 704444 626500
rect 705284 626332 705340 626342
rect 705284 626192 705340 626276
rect 705732 626332 705788 626342
rect 705732 626192 705788 626276
rect 704836 625436 704892 625446
rect 704836 625370 704892 625380
rect 704388 590268 704444 590800
rect 704836 590492 704892 590800
rect 704836 590426 704892 590436
rect 705284 590380 705340 590800
rect 705284 590314 705340 590324
rect 705732 590268 705788 590800
rect 704388 590202 704444 590212
rect 705684 590212 705788 590268
rect 705684 589820 705740 590212
rect 705684 589754 705740 589764
rect 704836 583324 704892 583334
rect 704836 583184 704892 583268
rect 704004 582876 704060 582886
rect 705284 582876 705340 582886
rect 704060 582820 704416 582876
rect 704004 582810 704060 582820
rect 705284 582810 705340 582820
rect 705732 582428 705788 582438
rect 705732 582362 705788 582372
rect 705012 547932 705068 547942
rect 704388 547708 704444 547904
rect 704564 547876 704864 547932
rect 705068 547876 705312 547932
rect 705572 547876 705760 547932
rect 704564 547820 704620 547876
rect 705012 547866 705068 547876
rect 704564 547754 704620 547764
rect 704388 547642 704444 547652
rect 705572 543452 705628 547876
rect 705572 543386 705628 543396
rect 704564 540204 704620 540214
rect 704416 540148 704564 540204
rect 704564 540138 704620 540148
rect 704676 540092 704732 540102
rect 705124 540092 705180 540102
rect 704732 540036 704864 540092
rect 705180 540036 705312 540092
rect 704676 540026 704732 540036
rect 705124 540026 705180 540036
rect 705732 539420 705788 539430
rect 705732 539354 705788 539364
rect 695380 521994 695436 522004
rect 696276 521500 696332 521510
rect 695156 351820 695212 351830
rect 695156 334236 695212 351764
rect 695156 334170 695212 334180
rect 695380 349132 695436 349142
rect 695380 334012 695436 349076
rect 695380 333946 695436 333956
rect 694932 306954 694988 306964
rect 695156 306572 695212 306582
rect 694708 212202 694764 212212
rect 694820 266252 694876 266262
rect 693028 179722 693084 179732
rect 694596 180236 694652 180246
rect 694596 166124 694652 180180
rect 694820 180012 694876 266196
rect 694820 179946 694876 179956
rect 694932 223244 694988 223254
rect 694932 173068 694988 223188
rect 695044 220556 695100 220566
rect 695044 177660 695100 220500
rect 695156 191548 695212 306516
rect 696276 205324 696332 521444
rect 704388 504588 704444 504896
rect 704388 504522 704444 504532
rect 704836 504476 704892 504896
rect 704836 504410 704892 504420
rect 705284 504364 705340 504896
rect 705284 504298 705340 504308
rect 705572 504868 705760 504924
rect 705572 504140 705628 504868
rect 705572 504074 705628 504084
rect 700532 488012 700588 488022
rect 700532 350028 700588 487956
rect 704564 368172 704620 368182
rect 704620 368116 704864 368172
rect 704564 368106 704620 368116
rect 704004 367836 704060 367846
rect 705284 367836 705340 367846
rect 704060 367780 704416 367836
rect 704004 367770 704060 367780
rect 705284 367770 705340 367780
rect 705732 367388 705788 367398
rect 705732 367322 705788 367332
rect 700532 349962 700588 349972
rect 704836 333116 704892 333126
rect 704836 333050 704892 333060
rect 705012 332892 705068 332902
rect 704388 332668 704444 332864
rect 705068 332836 705312 332892
rect 705572 332836 705760 332892
rect 705012 332826 705068 332836
rect 705572 332780 705628 332836
rect 705572 332714 705628 332724
rect 704388 332602 704444 332612
rect 704004 325164 704060 325174
rect 705124 325164 705180 325174
rect 704060 325108 704416 325164
rect 705180 325108 705312 325164
rect 704004 325098 704060 325108
rect 705124 325098 705180 325108
rect 704564 325052 704620 325062
rect 704620 324996 704864 325052
rect 704564 324986 704620 324996
rect 705732 324380 705788 324390
rect 705732 324314 705788 324324
rect 704676 289884 704732 289894
rect 704416 289828 704676 289884
rect 705012 289884 705068 289894
rect 704676 289818 704732 289828
rect 704836 289436 704892 289856
rect 705068 289828 705312 289884
rect 705572 289828 705760 289884
rect 705012 289818 705068 289828
rect 704836 289370 704892 289380
rect 705572 289100 705628 289828
rect 705572 289034 705628 289044
rect 704676 282156 704732 282166
rect 704416 282100 704676 282156
rect 704676 282090 704732 282100
rect 705012 282044 705068 282054
rect 705068 281988 705312 282044
rect 705012 281978 705068 281988
rect 704836 281932 704892 281942
rect 704836 281866 704892 281876
rect 705732 281372 705788 281382
rect 705732 281306 705788 281316
rect 696276 205258 696332 205268
rect 697956 263564 698012 263574
rect 695156 191482 695212 191492
rect 697956 184604 698012 263508
rect 704676 246876 704732 246886
rect 704416 246820 704676 246876
rect 704676 246810 704732 246820
rect 704788 246820 704864 246876
rect 704564 239148 704620 239158
rect 704416 239092 704564 239148
rect 704788 239148 704844 246820
rect 705284 246316 705340 246848
rect 705284 246250 705340 246260
rect 705684 246820 705760 246876
rect 705684 239148 705740 246820
rect 704788 239092 704864 239148
rect 705684 239092 705760 239148
rect 704564 239082 704620 239092
rect 705284 238476 705340 238486
rect 705284 238410 705340 238420
rect 700532 236794 700588 236806
rect 700532 236742 700534 236794
rect 700586 236742 700588 236794
rect 700532 222796 700588 236742
rect 700532 222730 700588 222740
rect 704388 203308 704444 203840
rect 704836 203532 704892 203840
rect 704836 203466 704892 203476
rect 705284 203420 705340 203840
rect 705732 203644 705788 203840
rect 705732 203578 705788 203588
rect 705284 203354 705340 203364
rect 704388 203242 704444 203252
rect 704564 196252 704620 196262
rect 703892 196140 703948 196150
rect 704564 196140 704620 196196
rect 703948 196084 704416 196140
rect 704564 196084 704864 196140
rect 703892 196074 703948 196084
rect 705012 196028 705068 196038
rect 705068 195972 705312 196028
rect 705012 195962 705068 195972
rect 705732 195468 705788 195478
rect 705732 195402 705788 195412
rect 697956 184538 698012 184548
rect 695044 177594 695100 177604
rect 694932 173002 694988 173012
rect 694596 166058 694652 166068
rect 694708 163884 694764 163894
rect 686980 132682 687036 132692
rect 694596 156940 694652 156950
rect 694596 91532 694652 156884
rect 694708 134540 694764 163828
rect 705012 160860 705068 160870
rect 704388 160300 704444 160832
rect 704836 160412 704892 160832
rect 705068 160804 705312 160860
rect 705572 160804 705760 160860
rect 705012 160794 705068 160804
rect 704836 160346 704892 160356
rect 704388 160234 704444 160244
rect 705572 159740 705628 160804
rect 705572 159674 705628 159684
rect 700532 159180 700588 159190
rect 700532 137228 700588 159124
rect 704388 152796 704444 152806
rect 704388 152730 704444 152740
rect 705284 152796 705340 152806
rect 705284 152730 705340 152740
rect 704836 152572 704892 152582
rect 704836 152506 704892 152516
rect 705732 152460 705788 152470
rect 705732 152394 705788 152404
rect 707896 152180 707952 152236
rect 707896 151900 707952 151956
rect 700532 137162 700588 137172
rect 694708 134474 694764 134484
rect 704836 118076 704892 118086
rect 704836 118010 704892 118020
rect 704676 117852 704732 117862
rect 704416 117796 704676 117852
rect 704676 117786 704732 117796
rect 705012 117796 705312 117852
rect 705572 117796 705760 117852
rect 705012 117628 705068 117796
rect 705572 117740 705628 117796
rect 705572 117674 705628 117684
rect 705012 117562 705068 117572
rect 704004 110124 704060 110134
rect 705012 110124 705068 110134
rect 704060 110068 704416 110124
rect 705068 110068 705312 110124
rect 704004 110058 704060 110068
rect 705012 110058 705068 110068
rect 704564 110012 704620 110022
rect 704620 109956 704864 110012
rect 704564 109946 704620 109956
rect 705732 109452 705788 109462
rect 705732 109386 705788 109396
rect 694596 91466 694652 91476
rect 686532 90794 686588 90804
rect 686308 90682 686364 90692
rect 672756 73994 672812 74004
rect 672980 83468 673036 83478
rect 672980 80778 673036 83412
rect 672980 80726 672982 80778
rect 673034 80726 673036 80778
rect 672980 73948 673036 80726
rect 704388 74172 704444 74816
rect 704836 74284 704892 74816
rect 705284 74508 705340 74816
rect 705284 74442 705340 74452
rect 704836 74218 704892 74228
rect 705732 74172 705788 74816
rect 704340 74116 704444 74172
rect 705684 74116 705788 74172
rect 704340 74060 704396 74116
rect 704340 73994 704396 74004
rect 672980 73882 673036 73892
rect 705684 73948 705740 74116
rect 705684 73882 705740 73892
rect 619332 71082 619388 71092
rect 617988 70970 618044 70980
rect 561210 70084 561932 70140
rect 505890 70074 505946 70084
rect 548432 70074 548488 70084
rect 469140 69738 469196 69748
rect 506036 69804 506092 69814
rect 506036 69738 506092 69748
<< via2 >>
rect 490868 949172 490924 949228
rect 106596 947732 106652 947788
rect 72772 946036 72828 946092
rect 77476 946036 77532 946092
rect 77252 945924 77308 945980
rect 73556 945812 73612 945868
rect 72212 945700 72268 945756
rect 72996 910868 73052 910924
rect 73444 910756 73500 910812
rect 73556 910644 73612 910700
rect 72212 910532 72268 910588
rect 73780 782068 73836 782124
rect 72660 781844 72716 781900
rect 72212 781732 72268 781788
rect 73108 781620 73164 781676
rect 73556 747460 73612 747516
rect 72660 747348 72716 747404
rect 72212 747236 72268 747292
rect 77364 945812 77420 945868
rect 141316 947044 141372 947100
rect 216580 947732 216636 947788
rect 106260 946596 106316 946652
rect 77476 747460 77532 747516
rect 77364 747348 77420 747404
rect 77252 747236 77308 747292
rect 73108 747124 73164 747180
rect 85204 942788 85260 942844
rect 84084 935732 84140 935788
rect 83972 929796 84028 929852
rect 79716 927332 79772 927388
rect 78372 782068 78428 782124
rect 78148 781844 78204 781900
rect 77588 747124 77644 747180
rect 77700 781732 77756 781788
rect 72772 741076 72828 741132
rect 77476 741076 77532 741132
rect 73556 740852 73612 740908
rect 77364 740852 77420 740908
rect 72212 740740 72268 740796
rect 73108 740628 73164 740684
rect 77252 740628 77308 740684
rect 77252 738052 77308 738108
rect 73108 706580 73164 706636
rect 72212 706468 72268 706524
rect 73556 706356 73612 706412
rect 72660 706244 72716 706300
rect 72548 700084 72604 700140
rect 73108 699860 73164 699916
rect 72660 699748 72716 699804
rect 73556 699636 73612 699692
rect 73556 665140 73612 665196
rect 72660 665028 72716 665084
rect 77924 781620 77980 781676
rect 77700 706468 77756 706524
rect 77812 740964 77868 741020
rect 77700 699748 77756 699804
rect 77476 665140 77532 665196
rect 77588 699636 77644 699692
rect 77252 665028 77308 665084
rect 72548 664916 72604 664972
rect 73444 664804 73500 664860
rect 72324 659092 72380 659148
rect 73108 658868 73164 658924
rect 73556 658756 73612 658812
rect 77476 658756 77532 658812
rect 72660 658644 72716 658700
rect 77252 658644 77308 658700
rect 72660 624596 72716 624652
rect 73556 624484 73612 624540
rect 73108 624372 73164 624428
rect 72212 624260 72268 624316
rect 72212 617652 72268 617708
rect 73556 617540 73612 617596
rect 73444 582820 73500 582876
rect 73780 582708 73836 582764
rect 77252 582708 77308 582764
rect 72660 582596 72716 582652
rect 77588 624596 77644 624652
rect 77924 706580 77980 706636
rect 78036 722372 78092 722428
rect 77812 664916 77868 664972
rect 77924 699860 77980 699916
rect 77700 624484 77756 624540
rect 77924 624372 77980 624428
rect 77476 582596 77532 582652
rect 77588 617540 77644 617596
rect 72212 582484 72268 582540
rect 72212 576884 72268 576940
rect 73556 576772 73612 576828
rect 72660 576660 72716 576716
rect 73108 576548 73164 576604
rect 73108 542500 73164 542556
rect 73556 542388 73612 542444
rect 72212 542276 72268 542332
rect 72660 542164 72716 542220
rect 77700 562660 77756 562716
rect 77812 576660 77868 576716
rect 77588 542164 77644 542220
rect 77252 536004 77308 536060
rect 72212 535780 72268 535836
rect 73556 535780 73612 535836
rect 72660 535556 72716 535612
rect 73108 501620 73164 501676
rect 73556 501508 73612 501564
rect 72660 501396 72716 501452
rect 72212 501284 72268 501340
rect 72212 412692 72268 412748
rect 73556 412580 73612 412636
rect 76132 387940 76188 387996
rect 72996 377748 73052 377804
rect 73780 377860 73836 377916
rect 76132 377748 76188 377804
rect 73108 377636 73164 377692
rect 72212 377524 72268 377580
rect 77364 535892 77420 535948
rect 77476 399700 77532 399756
rect 77588 535556 77644 535612
rect 77924 576548 77980 576604
rect 77924 501620 77980 501676
rect 77812 501508 77868 501564
rect 77588 399588 77644 399644
rect 77700 412580 77756 412636
rect 77364 387940 77420 387996
rect 77252 377524 77308 377580
rect 72212 371924 72268 371980
rect 73556 371812 73612 371868
rect 72660 371700 72716 371756
rect 73108 371588 73164 371644
rect 77588 371588 77644 371644
rect 73108 337540 73164 337596
rect 73556 337428 73612 337484
rect 72212 337316 72268 337372
rect 72660 337204 72716 337260
rect 73892 331044 73948 331100
rect 77364 330932 77420 330988
rect 72212 330820 72268 330876
rect 72660 330596 72716 330652
rect 77252 314468 77308 314524
rect 73108 296548 73164 296604
rect 73556 296436 73612 296492
rect 72212 296324 72268 296380
rect 72660 296212 72716 296268
rect 72772 290052 72828 290108
rect 72212 289828 72268 289884
rect 73556 289716 73612 289772
rect 73108 289604 73164 289660
rect 73108 255220 73164 255276
rect 73556 255108 73612 255164
rect 72548 254996 72604 255052
rect 77476 330596 77532 330652
rect 77924 371924 77980 371980
rect 77700 337204 77756 337260
rect 77812 371700 77868 371756
rect 77588 296548 77644 296604
rect 77812 296436 77868 296492
rect 77924 296324 77980 296380
rect 78148 706356 78204 706412
rect 78260 738052 78316 738108
rect 78372 706244 78428 706300
rect 78260 664804 78316 664860
rect 78372 700084 78428 700140
rect 78260 659092 78316 659148
rect 78148 658868 78204 658924
rect 78148 603092 78204 603148
rect 78372 624260 78428 624316
rect 78820 640052 78876 640108
rect 78260 582484 78316 582540
rect 78148 576884 78204 576940
rect 78596 617652 78652 617708
rect 78372 562548 78428 562604
rect 78484 576772 78540 576828
rect 78596 562436 78652 562492
rect 78484 501396 78540 501452
rect 78708 557732 78764 557788
rect 78148 501284 78204 501340
rect 78148 371812 78204 371868
rect 78260 356356 78316 356412
rect 78596 412692 78652 412748
rect 78596 356244 78652 356300
rect 78372 356132 78428 356188
rect 78372 331044 78428 331100
rect 78148 296212 78204 296268
rect 78036 290052 78092 290108
rect 77476 255108 77532 255164
rect 77700 289828 77756 289884
rect 77364 254996 77420 255052
rect 72996 254884 73052 254940
rect 73220 249060 73276 249116
rect 72212 248836 72268 248892
rect 77588 248836 77644 248892
rect 73556 248724 73612 248780
rect 77476 248724 77532 248780
rect 72660 248612 72716 248668
rect 77364 248612 77420 248668
rect 73108 214564 73164 214620
rect 73556 214452 73612 214508
rect 72212 214340 72268 214396
rect 72660 214228 72716 214284
rect 72660 207844 72716 207900
rect 73556 207732 73612 207788
rect 72212 207620 72268 207676
rect 73780 172900 73836 172956
rect 77364 172900 77420 172956
rect 72996 172788 73052 172844
rect 77476 172788 77532 172844
rect 73108 172676 73164 172732
rect 72212 172564 72268 172620
rect 78036 289828 78092 289884
rect 77924 289716 77980 289772
rect 77812 289604 77868 289660
rect 77812 214564 77868 214620
rect 77700 214340 77756 214396
rect 78260 273924 78316 273980
rect 83972 912660 84028 912716
rect 84308 935732 84364 935788
rect 84308 910868 84364 910924
rect 84532 935732 84588 935788
rect 84532 910756 84588 910812
rect 84084 910644 84140 910700
rect 85428 942676 85484 942732
rect 106260 945812 106316 945868
rect 106260 942004 106316 942060
rect 141092 945812 141148 945868
rect 120932 943348 120988 943404
rect 124292 943348 124348 943404
rect 141428 936628 141484 936684
rect 124292 936516 124348 936572
rect 141876 947044 141932 947100
rect 141652 945812 141708 945868
rect 160244 942228 160300 942284
rect 196084 946708 196140 946764
rect 196308 946596 196364 946652
rect 196308 946260 196364 946316
rect 177044 943460 177100 943516
rect 176484 943348 176540 943404
rect 160580 942116 160636 942172
rect 141876 936964 141932 937020
rect 163716 938532 163772 938588
rect 141652 936740 141708 936796
rect 85428 935396 85484 935452
rect 96964 935620 97020 935676
rect 141316 935396 141372 935452
rect 178164 943460 178220 943516
rect 178052 943348 178108 943404
rect 176708 937412 176764 937468
rect 178164 938532 178220 938588
rect 179732 943348 179788 943404
rect 271572 947732 271628 947788
rect 251076 947604 251132 947660
rect 306068 947604 306124 947660
rect 470260 947732 470316 947788
rect 525700 947732 525756 947788
rect 361060 947492 361116 947548
rect 545860 947492 545916 947548
rect 581140 947492 581196 947548
rect 690340 947732 690396 947788
rect 655844 947492 655900 947548
rect 697956 947492 698012 947548
rect 196644 942340 196700 942396
rect 251076 946708 251132 946764
rect 230132 943460 230188 943516
rect 215684 942004 215740 942060
rect 179732 937412 179788 937468
rect 178052 936964 178108 937020
rect 233492 943460 233548 943516
rect 231812 943348 231868 943404
rect 230132 936628 230188 936684
rect 230356 937412 230412 937468
rect 233492 937412 233548 937468
rect 233828 943348 233884 943404
rect 270564 942116 270620 942172
rect 285684 943348 285740 943404
rect 282436 937412 282492 937468
rect 251972 935172 252028 935228
rect 289156 943348 289212 943404
rect 285684 937076 285740 937132
rect 285908 943236 285964 943292
rect 289380 943348 289436 943404
rect 361060 947156 361116 947212
rect 471268 946836 471324 946892
rect 361060 946708 361116 946764
rect 344596 943460 344652 943516
rect 341124 943236 341180 943292
rect 335860 942170 335916 942172
rect 335860 942118 335862 942170
rect 335862 942118 335914 942170
rect 335914 942118 335916 942170
rect 335860 942116 335916 942118
rect 306404 942004 306460 942060
rect 289380 936740 289436 936796
rect 344708 943348 344764 943404
rect 471828 946036 471884 946092
rect 525588 947284 525644 947340
rect 471716 945812 471772 945868
rect 581252 947156 581308 947212
rect 545860 947044 545916 947100
rect 690340 947284 690396 947340
rect 655844 947044 655900 947100
rect 545636 946836 545692 946892
rect 526148 946708 526204 946764
rect 655620 946836 655676 946892
rect 691796 946820 691852 946876
rect 581028 946708 581084 946764
rect 525700 946388 525756 946444
rect 545524 946388 545580 946444
rect 655508 946388 655564 946444
rect 581140 946260 581196 946316
rect 490868 946036 490924 946092
rect 490644 945924 490700 945980
rect 490532 945812 490588 945868
rect 691124 945812 691180 945868
rect 507444 943460 507500 943516
rect 450212 943348 450268 943404
rect 451892 943348 451948 943404
rect 451892 936852 451948 936908
rect 453572 943348 453628 943404
rect 455028 943348 455084 943404
rect 505652 943348 505708 943404
rect 455028 938196 455084 938252
rect 458500 938196 458556 938252
rect 341124 936068 341180 936124
rect 342580 936068 342636 936124
rect 285908 935060 285964 935116
rect 341012 935060 341068 935116
rect 231812 934948 231868 935004
rect 274036 934948 274092 935004
rect 362964 934836 363020 934892
rect 430948 934836 431004 934892
rect 505876 943236 505932 943292
rect 505876 936964 505932 937020
rect 474740 936852 474796 936908
rect 509012 943348 509068 943404
rect 510580 943348 510636 943404
rect 564228 943348 564284 943404
rect 561092 943236 561148 943292
rect 510580 938420 510636 938476
rect 519204 938420 519260 938476
rect 509012 937076 509068 937132
rect 561092 937188 561148 937244
rect 541380 936964 541436 937020
rect 673428 943348 673484 943404
rect 674100 943348 674156 943404
rect 673428 939092 673484 939148
rect 673652 943236 673708 943292
rect 673652 937300 673708 937356
rect 673876 943124 673932 943180
rect 608132 937188 608188 937244
rect 585956 935620 586012 935676
rect 652708 935508 652764 935564
rect 673876 935508 673932 935564
rect 674772 939092 674828 939148
rect 687428 937188 687484 937244
rect 687204 937076 687260 937132
rect 686980 935284 687036 935340
rect 686644 935060 686700 935116
rect 686532 934948 686588 935004
rect 686308 934724 686364 934780
rect 85204 934612 85260 934668
rect 118468 934612 118524 934668
rect 84756 910532 84812 910588
rect 686196 934500 686252 934556
rect 83972 883988 84028 884044
rect 83076 783636 83132 783692
rect 80500 763140 80556 763196
rect 80388 600628 80444 600684
rect 80276 518868 80332 518924
rect 80052 396116 80108 396172
rect 80164 354116 80220 354172
rect 79716 290276 79772 290332
rect 80276 331716 80332 331772
rect 80500 331828 80556 331884
rect 83188 762804 83244 762860
rect 84308 869764 84364 869820
rect 83972 762804 84028 762860
rect 84084 841204 84140 841260
rect 84084 720692 84140 720748
rect 84196 798308 84252 798364
rect 83972 712628 84028 712684
rect 83188 302372 83244 302428
rect 83300 701316 83356 701372
rect 83860 682164 83916 682220
rect 83748 557732 83804 557788
rect 83412 415716 83468 415772
rect 83636 393428 83692 393484
rect 83412 306516 83468 306572
rect 83076 289828 83132 289884
rect 84644 855428 84700 855484
rect 84308 766052 84364 766108
rect 84420 826868 84476 826924
rect 84196 681156 84252 681212
rect 84308 741188 84364 741244
rect 83972 598500 84028 598556
rect 84084 669732 84140 669788
rect 83972 584052 84028 584108
rect 84420 725060 84476 725116
rect 84532 783972 84588 784028
rect 84308 642292 84364 642348
rect 84420 698292 84476 698348
rect 84084 557844 84140 557900
rect 84196 626836 84252 626892
rect 686196 848148 686252 848204
rect 84644 764484 84700 764540
rect 84756 812644 84812 812700
rect 84532 684292 84588 684348
rect 84644 726852 84700 726908
rect 84420 601972 84476 602028
rect 84532 655508 84588 655564
rect 84196 516404 84252 516460
rect 84308 569716 84364 569772
rect 83972 393652 84028 393708
rect 84084 498372 84140 498428
rect 84084 311444 84140 311500
rect 84196 455476 84252 455532
rect 83860 289716 83916 289772
rect 78484 282996 78540 283052
rect 78708 274036 78764 274092
rect 78820 283108 78876 283164
rect 78484 273812 78540 273868
rect 78372 254884 78428 254940
rect 78036 214452 78092 214508
rect 78148 249060 78204 249116
rect 77924 214228 77980 214284
rect 77588 172564 77644 172620
rect 78036 207732 78092 207788
rect 686196 793492 686252 793548
rect 84756 722596 84812 722652
rect 84868 769748 84924 769804
rect 84868 682276 84924 682332
rect 84980 683732 85036 683788
rect 84644 642068 84700 642124
rect 84532 561764 84588 561820
rect 84644 641172 84700 641228
rect 84868 618996 84924 619052
rect 84644 559412 84700 559468
rect 84756 612612 84812 612668
rect 84644 555492 84700 555548
rect 84308 396900 84364 396956
rect 84420 526932 84476 526988
rect 84420 356916 84476 356972
rect 84532 484036 84588 484092
rect 84196 270788 84252 270844
rect 84308 341236 84364 341292
rect 78820 233492 78876 233548
rect 78148 172676 78204 172732
rect 84756 519092 84812 519148
rect 84644 394996 84700 395052
rect 84756 512596 84812 512652
rect 84532 314356 84588 314412
rect 84644 384020 84700 384076
rect 84756 355012 84812 355068
rect 84980 599732 85036 599788
rect 84980 598052 85036 598108
rect 84980 517860 85036 517916
rect 84980 469140 85036 469196
rect 84980 312452 85036 312508
rect 85092 426692 85148 426748
rect 84868 306740 84924 306796
rect 84756 305786 84812 305788
rect 84756 305734 84758 305786
rect 84758 305734 84810 305786
rect 84810 305734 84812 305786
rect 84756 305732 84812 305734
rect 85092 272132 85148 272188
rect 85204 398132 85260 398188
rect 84644 232036 84700 232092
rect 686420 740628 686476 740684
rect 686756 934612 686812 934668
rect 686868 934164 686924 934220
rect 686868 928004 686924 928060
rect 686756 914676 686812 914732
rect 686644 767732 686700 767788
rect 686980 753956 687036 754012
rect 686532 688100 686588 688156
rect 686420 671076 686476 671132
rect 686308 661444 686364 661500
rect 686532 606788 686588 606844
rect 686532 488180 686588 488236
rect 686644 593460 686700 593516
rect 686420 446852 686476 446908
rect 686196 334068 686252 334124
rect 686308 366884 686364 366940
rect 222852 333732 222908 333788
rect 119140 333620 119196 333676
rect 171108 333620 171164 333676
rect 160692 333508 160748 333564
rect 127204 333396 127260 333452
rect 88788 332836 88844 332892
rect 92820 332612 92876 332668
rect 100660 332948 100716 333004
rect 98756 332724 98812 332780
rect 106708 333060 106764 333116
rect 108724 330036 108780 330092
rect 112644 328356 112700 328412
rect 116676 328580 116732 328636
rect 130564 328692 130620 328748
rect 133476 332948 133532 333004
rect 114660 328020 114716 328076
rect 104132 324100 104188 324156
rect 133924 332836 133980 332892
rect 133700 332724 133756 332780
rect 133476 323876 133532 323932
rect 134484 332836 134540 332892
rect 135156 333060 135212 333116
rect 140532 332948 140588 333004
rect 149044 333172 149100 333228
rect 146468 333060 146524 333116
rect 144340 332052 144396 332108
rect 150388 329028 150444 329084
rect 142436 328916 142492 328972
rect 136500 328804 136556 328860
rect 135156 323988 135212 324044
rect 149492 323988 149548 324044
rect 150612 323876 150668 323932
rect 149492 323764 149548 323820
rect 156324 329140 156380 329196
rect 162820 333284 162876 333340
rect 157892 324996 157948 325052
rect 166180 328244 166236 328300
rect 162932 325108 162988 325164
rect 159908 324212 159964 324268
rect 151956 323764 152012 323820
rect 159572 323876 159628 323932
rect 133924 322532 133980 322588
rect 159908 323764 159964 323820
rect 161700 324324 161756 324380
rect 161028 324100 161084 324156
rect 160972 323876 161028 323932
rect 161364 323988 161420 324044
rect 161140 323876 161196 323932
rect 162428 323876 162484 323932
rect 162596 323876 162652 323932
rect 165340 324100 165396 324156
rect 166796 324100 166852 324156
rect 166124 323988 166180 324044
rect 168084 330036 168140 330092
rect 170324 328468 170380 328524
rect 168308 328132 168364 328188
rect 170436 328020 170492 328076
rect 209636 333620 209692 333676
rect 187124 333508 187180 333564
rect 173460 333396 173516 333452
rect 174580 333396 174636 333452
rect 171892 328580 171948 328636
rect 173460 333060 173516 333116
rect 174020 333060 174076 333116
rect 172228 328356 172284 328412
rect 176260 332612 176316 332668
rect 176932 332836 176988 332892
rect 176260 328692 176316 328748
rect 178276 332948 178332 333004
rect 179172 332836 179228 332892
rect 178388 328804 178444 328860
rect 180180 332724 180236 332780
rect 181300 333172 181356 333228
rect 180628 328916 180684 328972
rect 184436 333172 184492 333228
rect 182196 333060 182252 333116
rect 182756 332836 182812 332892
rect 181636 332052 181692 332108
rect 184212 329028 184268 329084
rect 167580 323876 167636 323932
rect 169708 324100 169764 324156
rect 185668 324996 185724 325052
rect 188580 333172 188636 333228
rect 187908 325108 187964 325164
rect 193732 332948 193788 333004
rect 192276 332612 192332 332668
rect 190036 328468 190092 328524
rect 189364 328244 189420 328300
rect 191492 328356 191548 328412
rect 190820 328132 190876 328188
rect 194180 332612 194236 332668
rect 194404 333060 194460 333116
rect 194852 332836 194908 332892
rect 184884 323876 184940 323932
rect 186508 324100 186564 324156
rect 193004 324100 193060 324156
rect 195188 332724 195244 332780
rect 198100 332612 198156 332668
rect 198324 332724 198380 332780
rect 194852 324212 194908 324268
rect 195916 324212 195972 324268
rect 197372 323876 197428 323932
rect 203364 332836 203420 332892
rect 200004 324212 200060 324268
rect 201068 324212 201124 324268
rect 201740 324100 201796 324156
rect 203196 324100 203252 324156
rect 207508 333172 207564 333228
rect 207956 332836 208012 332892
rect 208964 332836 209020 332892
rect 210644 333508 210700 333564
rect 209860 332612 209916 332668
rect 210084 332612 210140 332668
rect 221620 333508 221676 333564
rect 216356 333396 216412 333452
rect 210644 332612 210700 332668
rect 211204 333060 211260 333116
rect 205044 324100 205100 324156
rect 206108 324100 206164 324156
rect 208348 324100 208404 324156
rect 211764 332948 211820 333004
rect 215908 332724 215964 332780
rect 215124 330036 215180 330092
rect 214228 328916 214284 328972
rect 211764 324212 211820 324268
rect 217028 333284 217084 333340
rect 216692 330708 216748 330764
rect 212716 324212 212772 324268
rect 213388 324100 213444 324156
rect 214844 324100 214900 324156
rect 217140 333172 217196 333228
rect 218484 333172 218540 333228
rect 216692 324212 216748 324268
rect 219828 332836 219884 332892
rect 220164 333060 220220 333116
rect 219940 328580 219996 328636
rect 222292 328468 222348 328524
rect 217476 324100 217532 324156
rect 217868 324212 217924 324268
rect 219324 324100 219380 324156
rect 258916 333732 258972 333788
rect 271012 333732 271068 333788
rect 223412 333620 223468 333676
rect 240996 333396 241052 333452
rect 225204 332836 225260 332892
rect 224420 328356 224476 328412
rect 227780 332948 227836 333004
rect 225764 332724 225820 332780
rect 229460 332836 229516 332892
rect 225820 324100 225876 324156
rect 231812 332612 231868 332668
rect 233604 332612 233660 332668
rect 233156 328132 233212 328188
rect 232484 328020 232540 328076
rect 230188 324100 230244 324156
rect 233604 324100 233660 324156
rect 235284 330596 235340 330652
rect 235732 328916 235788 328972
rect 237412 330484 237468 330540
rect 236068 327124 236124 327180
rect 234556 324100 234612 324156
rect 239092 333284 239148 333340
rect 240548 333284 240604 333340
rect 237748 330036 237804 330092
rect 238532 330372 238588 330428
rect 238308 327012 238364 327068
rect 239652 330260 239708 330316
rect 236796 324100 236852 324156
rect 243684 330708 243740 330764
rect 242676 326900 242732 326956
rect 240212 324212 240268 324268
rect 245476 330148 245532 330204
rect 244804 325332 244860 325388
rect 241836 324212 241892 324268
rect 241164 323876 241220 323932
rect 247044 333172 247100 333228
rect 245700 328692 245756 328748
rect 246260 329140 246316 329196
rect 247044 325220 247100 325276
rect 249172 325108 249228 325164
rect 253652 333060 253708 333116
rect 249620 328580 249676 328636
rect 249956 329028 250012 329084
rect 252084 328916 252140 328972
rect 249396 323876 249452 323932
rect 251412 324996 251468 325052
rect 254324 328692 254380 328748
rect 254996 328580 255052 328636
rect 257124 330036 257180 330092
rect 255668 328468 255724 328524
rect 257908 326788 257964 326844
rect 265524 332724 265580 332780
rect 263620 328804 263676 328860
rect 261604 328356 261660 328412
rect 253484 324100 253540 324156
rect 255724 324100 255780 324156
rect 258636 324100 258692 324156
rect 259308 324100 259364 324156
rect 260092 323988 260148 324044
rect 265188 328356 265244 328412
rect 261548 324100 261604 324156
rect 263676 324100 263732 324156
rect 267988 331492 268044 331548
rect 270228 331156 270284 331212
rect 388052 333732 388108 333788
rect 656740 333732 656796 333788
rect 278292 333620 278348 333676
rect 273140 333172 273196 333228
rect 272244 331268 272300 331324
rect 269500 324100 269556 324156
rect 274596 331380 274652 331436
rect 277508 332836 277564 332892
rect 277396 332724 277452 332780
rect 275492 327908 275548 327964
rect 273980 324100 274036 324156
rect 406420 333620 406476 333676
rect 278292 332724 278348 332780
rect 278404 326676 278460 326732
rect 280644 332836 280700 332892
rect 281428 328020 281484 328076
rect 282772 326340 282828 326396
rect 320180 333508 320236 333564
rect 319956 333396 320012 333452
rect 286244 332948 286300 333004
rect 285460 328132 285516 328188
rect 285572 329588 285628 329644
rect 287364 332612 287420 332668
rect 287252 329700 287308 329756
rect 290724 333060 290780 333116
rect 291396 330596 291452 330652
rect 293412 328244 293468 328300
rect 293636 326452 293692 326508
rect 292964 325444 293020 325500
rect 291452 324100 291508 324156
rect 297332 330484 297388 330540
rect 295316 327124 295372 327180
rect 296436 329812 296492 329868
rect 295092 324548 295148 324604
rect 298004 328132 298060 328188
rect 295820 324100 295876 324156
rect 301364 330372 301420 330428
rect 303044 330820 303100 330876
rect 299348 327012 299404 327068
rect 300804 329924 300860 329980
rect 300244 326564 300300 326620
rect 299404 324100 299460 324156
rect 304612 333284 304668 333340
rect 303268 330260 303324 330316
rect 304612 326004 304668 326060
rect 303828 325668 303884 325724
rect 302316 324100 302372 324156
rect 307524 330708 307580 330764
rect 308196 324436 308252 324492
rect 306012 324100 306068 324156
rect 311220 326900 311276 326956
rect 311780 330596 311836 330652
rect 308924 324100 308980 324156
rect 311052 324100 311108 324156
rect 318276 331604 318332 331660
rect 315812 325332 315868 325388
rect 316148 330484 316204 330540
rect 319172 330148 319228 330204
rect 319620 327124 319676 327180
rect 320068 325444 320124 325500
rect 364532 333508 364588 333564
rect 386036 333508 386092 333564
rect 370244 333396 370300 333452
rect 321188 329140 321244 329196
rect 321300 325556 321356 325612
rect 324884 332500 324940 332556
rect 322532 325220 322588 325276
rect 317660 324100 317716 324156
rect 316876 323876 316932 323932
rect 329252 332388 329308 332444
rect 328692 326900 328748 326956
rect 327572 325108 327628 325164
rect 327908 325444 327964 325500
rect 324156 323876 324212 323932
rect 325724 323988 325780 324044
rect 331156 329028 331212 329084
rect 330148 325332 330204 325388
rect 335972 330148 336028 330204
rect 335188 327908 335244 327964
rect 335076 327796 335132 327852
rect 334292 324996 334348 325052
rect 334516 325220 334572 325276
rect 330764 324100 330820 324156
rect 332220 323876 332276 323932
rect 337092 328916 337148 328972
rect 335972 328244 336028 328300
rect 338100 328244 338156 328300
rect 337428 324996 337484 325052
rect 333676 323876 333732 323932
rect 336588 324100 336644 324156
rect 335916 323988 335972 324044
rect 342468 329140 342524 329196
rect 341012 327012 341068 327068
rect 341796 327012 341852 327068
rect 340340 325108 340396 325164
rect 339500 324100 339556 324156
rect 343028 328692 343084 328748
rect 343476 327908 343532 327964
rect 343700 327796 343756 327852
rect 344708 329028 344764 329084
rect 347060 330260 347116 330316
rect 347732 332052 347788 332108
rect 346052 329476 346108 329532
rect 345044 328580 345100 328636
rect 345268 328580 345324 328636
rect 346052 327572 346108 327628
rect 346164 329364 346220 329420
rect 345268 326788 345324 326844
rect 345380 324660 345436 324716
rect 350980 330036 351036 330092
rect 349076 328916 349132 328972
rect 347732 327684 347788 327740
rect 350532 326788 350588 326844
rect 349748 324772 349804 324828
rect 347564 324100 347620 324156
rect 354116 330260 354172 330316
rect 352996 328580 353052 328636
rect 353444 328692 353500 328748
rect 354116 327012 354172 327068
rect 354340 327012 354396 327068
rect 353892 325108 353948 325164
rect 354340 324996 354396 325052
rect 354116 324884 354172 324940
rect 358932 332612 358988 332668
rect 359492 332276 359548 332332
rect 356916 330148 356972 330204
rect 359156 330148 359212 330204
rect 355012 328468 355068 328524
rect 359492 329364 359548 329420
rect 359828 330036 359884 330092
rect 362964 332052 363020 332108
rect 366436 332052 366492 332108
rect 360724 325668 360780 325724
rect 364308 328468 364364 328524
rect 356972 324100 357028 324156
rect 358428 324100 358484 324156
rect 361340 324100 361396 324156
rect 367892 331044 367948 331100
rect 368900 329476 368956 329532
rect 367780 327796 367836 327852
rect 368676 327460 368732 327516
rect 367220 325108 367276 325164
rect 365708 323988 365764 324044
rect 368004 324996 368060 325052
rect 374836 331044 374892 331100
rect 372820 328356 372876 328412
rect 373604 329476 373660 329532
rect 373604 327684 373660 327740
rect 369684 327572 369740 327628
rect 369572 327460 369628 327516
rect 376292 327460 376348 327516
rect 380772 331492 380828 331548
rect 380996 331492 381052 331548
rect 379652 331044 379708 331100
rect 379652 329588 379708 329644
rect 380996 329476 381052 329532
rect 381444 329588 381500 329644
rect 381332 327796 381388 327852
rect 384804 328804 384860 328860
rect 385476 329252 385532 329308
rect 381444 327460 381500 327516
rect 381332 326676 381388 326732
rect 382340 326676 382396 326732
rect 379316 326228 379372 326284
rect 382340 325780 382396 325836
rect 376292 324996 376348 325052
rect 375956 324324 376012 324380
rect 369404 324100 369460 324156
rect 373772 324100 373828 324156
rect 370860 323988 370916 324044
rect 371532 323876 371588 323932
rect 372988 323876 373044 323932
rect 374444 323988 374500 324044
rect 376740 324324 376796 324380
rect 377860 324154 377916 324156
rect 377860 324102 377862 324154
rect 377862 324102 377914 324154
rect 377914 324102 377916 324154
rect 377860 324100 377916 324102
rect 377356 323876 377412 323932
rect 378140 323876 378196 323932
rect 378812 323876 378868 323932
rect 460068 333508 460124 333564
rect 386820 331156 386876 331212
rect 387156 331940 387212 331996
rect 387156 329252 387212 329308
rect 393988 333172 394044 333228
rect 392756 331268 392812 331324
rect 390740 327908 390796 327964
rect 391188 327908 391244 327964
rect 386372 327460 386428 327516
rect 391188 327460 391244 327516
rect 386372 324548 386428 324604
rect 398692 331380 398748 331436
rect 399700 331380 399756 331436
rect 399700 329700 399756 329756
rect 489412 333396 489468 333452
rect 610932 333396 610988 333452
rect 403396 328804 403452 328860
rect 411348 329588 411404 329644
rect 408660 327796 408716 327852
rect 418516 332836 418572 332892
rect 418292 332612 418348 332668
rect 421540 333172 421596 333228
rect 420532 332612 420588 332668
rect 418292 326340 418348 326396
rect 421092 332836 421148 332892
rect 421764 331268 421820 331324
rect 421540 327908 421596 327964
rect 430500 332948 430556 333004
rect 428484 331044 428540 331100
rect 437668 332948 437724 333004
rect 434420 331380 434476 331436
rect 442372 333060 442428 333116
rect 440468 331268 440524 331324
rect 444388 328020 444444 328076
rect 453684 333172 453740 333228
rect 454692 333060 454748 333116
rect 450324 326452 450380 326508
rect 454804 332612 454860 332668
rect 454916 333172 454972 333228
rect 458276 329812 458332 329868
rect 462308 328132 462364 328188
rect 470260 329924 470316 329980
rect 468244 327460 468300 327516
rect 456260 326564 456316 326620
rect 477540 333284 477596 333340
rect 476196 330820 476252 330876
rect 474180 326116 474236 326172
rect 488068 330708 488124 330764
rect 480116 326004 480172 326060
rect 497364 333284 497420 333340
rect 492100 327348 492156 327404
rect 488404 325668 488460 325724
rect 471156 324884 471212 324940
rect 454916 324772 454972 324828
rect 437668 324660 437724 324716
rect 396452 324212 396508 324268
rect 500052 330596 500108 330652
rect 511924 330484 511980 330540
rect 517860 331604 517916 331660
rect 515956 327236 516012 327292
rect 521892 327124 521948 327180
rect 533092 333284 533148 333340
rect 525812 325556 525868 325612
rect 535780 332500 535836 332556
rect 512372 324884 512428 324940
rect 547764 332388 547820 332444
rect 545748 326900 545804 326956
rect 542612 325444 542668 325500
rect 551684 332612 551740 332668
rect 549332 325332 549388 325388
rect 537572 324548 537628 324604
rect 559636 330372 559692 330428
rect 567588 332724 567644 332780
rect 565572 331492 565628 331548
rect 575540 332164 575596 332220
rect 579460 332836 579516 332892
rect 581476 330260 581532 330316
rect 583492 329140 583548 329196
rect 591444 332948 591500 333004
rect 593460 332276 593516 332332
rect 589428 329028 589484 329084
rect 571508 328244 571564 328300
rect 569604 327012 569660 327068
rect 603092 333172 603148 333228
rect 601412 328916 601468 328972
rect 609364 333060 609420 333116
rect 605332 326788 605388 326844
rect 561092 325220 561148 325276
rect 554372 324436 554428 324492
rect 485492 323876 485548 323932
rect 380324 323092 380380 323148
rect 159572 322532 159628 322588
rect 557732 319396 557788 319452
rect 460292 312452 460348 312508
rect 458612 309204 458668 309260
rect 157892 308308 157948 308364
rect 151172 308196 151228 308252
rect 92372 307972 92428 308028
rect 90580 286356 90636 286412
rect 85204 231812 85260 231868
rect 90356 283220 90412 283276
rect 92484 292234 92540 292236
rect 92484 292182 92486 292234
rect 92486 292182 92538 292234
rect 92538 292182 92540 292234
rect 92484 292180 92540 292182
rect 92596 290666 92652 290668
rect 92596 290614 92598 290666
rect 92598 290614 92650 290666
rect 92650 290614 92652 290666
rect 92596 290612 92652 290614
rect 94052 285572 94108 285628
rect 106036 307860 106092 307916
rect 94948 285572 95004 285628
rect 105812 307748 105868 307804
rect 104132 307636 104188 307692
rect 100772 307524 100828 307580
rect 99092 307412 99148 307468
rect 102452 307412 102508 307468
rect 146132 294756 146188 294812
rect 142996 291620 143052 291676
rect 142772 291508 142828 291564
rect 120932 291396 120988 291452
rect 117908 291060 117964 291116
rect 114884 286580 114940 286636
rect 112308 286468 112364 286524
rect 101444 280868 101500 280924
rect 111636 280868 111692 280924
rect 113540 284676 113596 284732
rect 117460 284900 117516 284956
rect 116116 284788 116172 284844
rect 139188 290388 139244 290444
rect 137956 288260 138012 288316
rect 136612 288148 136668 288204
rect 134036 281652 134092 281708
rect 126420 281316 126476 281372
rect 122500 281092 122556 281148
rect 125076 281092 125132 281148
rect 128996 281204 129052 281260
rect 135380 281428 135436 281484
rect 141764 290276 141820 290332
rect 140532 281764 140588 281820
rect 142772 285572 142828 285628
rect 143668 285572 143724 285628
rect 145572 281764 145628 281820
rect 149492 290052 149548 290108
rect 150724 289940 150780 289996
rect 154644 308084 154700 308140
rect 152852 291732 152908 291788
rect 154644 280868 154700 280924
rect 164444 308532 164500 308588
rect 164836 308644 164892 308700
rect 159684 286356 159740 286412
rect 161252 307972 161308 308028
rect 163044 307972 163100 308028
rect 160020 305898 160076 305900
rect 160020 305846 160022 305898
rect 160022 305846 160074 305898
rect 160074 305846 160076 305898
rect 160020 305844 160076 305846
rect 159908 281876 159964 281932
rect 160244 290164 160300 290220
rect 162260 288036 162316 288092
rect 160580 280868 160636 280924
rect 165564 308532 165620 308588
rect 166236 308420 166292 308476
rect 164948 307524 165004 307580
rect 165396 307524 165452 307580
rect 167412 307860 167468 307916
rect 167972 307748 168028 307804
rect 168084 308420 168140 308476
rect 166740 307636 166796 307692
rect 165396 288260 165452 288316
rect 109060 280756 109116 280812
rect 92260 280644 92316 280700
rect 169260 308420 169316 308476
rect 168756 290276 168812 290332
rect 171332 308420 171388 308476
rect 169764 305620 169820 305676
rect 170996 305620 171052 305676
rect 169876 286468 169932 286524
rect 172284 308420 172340 308476
rect 173124 308420 173180 308476
rect 171556 303156 171612 303212
rect 171668 286580 171724 286636
rect 173012 307972 173068 308028
rect 171444 284900 171500 284956
rect 171332 284788 171388 284844
rect 169764 284676 169820 284732
rect 169652 280980 169708 281036
rect 167972 280756 168028 280812
rect 170548 280756 170604 280812
rect 174188 308420 174244 308476
rect 173236 291844 173292 291900
rect 174692 305620 174748 305676
rect 176372 308420 176428 308476
rect 175924 305620 175980 305676
rect 174916 291396 174972 291452
rect 177212 308420 177268 308476
rect 176484 305620 176540 305676
rect 176148 281316 176204 281372
rect 176372 281316 176428 281372
rect 174804 281092 174860 281148
rect 175700 280868 175756 280924
rect 177716 305620 177772 305676
rect 176596 281204 176652 281260
rect 179732 308420 179788 308476
rect 178164 281988 178220 282044
rect 177940 280980 177996 281036
rect 180908 308420 180964 308476
rect 179732 281876 179788 281932
rect 182028 308420 182084 308476
rect 183092 308420 183148 308476
rect 184884 308420 184940 308476
rect 182644 307524 182700 307580
rect 183204 281540 183260 281596
rect 183428 307524 183484 307580
rect 181524 281428 181580 281484
rect 182756 281428 182812 281484
rect 180180 281204 180236 281260
rect 178948 281092 179004 281148
rect 180740 280868 180796 280924
rect 181636 280868 181692 280924
rect 184772 307636 184828 307692
rect 186396 308420 186452 308476
rect 184996 291620 185052 291676
rect 185444 291508 185500 291564
rect 186564 307860 186620 307916
rect 186676 294756 186732 294812
rect 186564 285572 186620 285628
rect 184884 281764 184940 281820
rect 188132 303268 188188 303324
rect 187236 285572 187292 285628
rect 188244 290052 188300 290108
rect 190596 308308 190652 308364
rect 191492 308532 191548 308588
rect 189364 308196 189420 308252
rect 192444 308532 192500 308588
rect 191492 308196 191548 308252
rect 191156 308084 191212 308140
rect 193676 308532 193732 308588
rect 195468 308644 195524 308700
rect 194908 308420 194964 308476
rect 191604 307748 191660 307804
rect 189924 291732 189980 291788
rect 190036 307412 190092 307468
rect 188356 289940 188412 289996
rect 191716 290164 191772 290220
rect 193396 308084 193452 308140
rect 194964 307860 195020 307916
rect 193284 288036 193340 288092
rect 196532 282100 196588 282156
rect 198660 308644 198716 308700
rect 196868 308196 196924 308252
rect 196980 280980 197036 281036
rect 198324 280980 198380 281036
rect 199892 308644 199948 308700
rect 199668 307972 199724 308028
rect 199108 303156 199164 303212
rect 200004 308420 200060 308476
rect 200956 308420 201012 308476
rect 200004 281092 200060 281148
rect 201796 308420 201852 308476
rect 201684 281316 201740 281372
rect 203420 308532 203476 308588
rect 202860 308420 202916 308476
rect 207116 308420 207172 308476
rect 204596 307524 204652 307580
rect 202020 281540 202076 281596
rect 201796 281204 201852 281260
rect 203588 280980 203644 281036
rect 203812 281428 203868 281484
rect 205268 307636 205324 307692
rect 206388 308308 206444 308364
rect 208292 307748 208348 307804
rect 208404 307972 208460 308028
rect 207620 307412 207676 307468
rect 208404 285572 208460 285628
rect 210700 308420 210756 308476
rect 211932 308644 211988 308700
rect 212604 308532 212660 308588
rect 213444 308532 213500 308588
rect 209412 308084 209468 308140
rect 211316 308196 211372 308252
rect 210084 307860 210140 307916
rect 210084 307636 210140 307692
rect 208964 285572 209020 285628
rect 211876 307524 211932 307580
rect 215124 308420 215180 308476
rect 213668 307412 213724 307468
rect 216804 307972 216860 308028
rect 218652 308532 218708 308588
rect 218820 308532 218876 308588
rect 216916 308308 216972 308364
rect 213556 280980 213612 281036
rect 217364 307636 217420 307692
rect 218036 307524 218092 307580
rect 218596 307636 218652 307692
rect 218596 285572 218652 285628
rect 219884 308420 219940 308476
rect 220276 308644 220332 308700
rect 219156 307412 219212 307468
rect 221116 308532 221172 308588
rect 222348 308644 222404 308700
rect 220388 308308 220444 308364
rect 225932 308420 225988 308476
rect 221620 307636 221676 307692
rect 219268 285572 219324 285628
rect 228452 308420 228508 308476
rect 227220 307412 227276 307468
rect 230188 308420 230244 308476
rect 232092 308644 232148 308700
rect 231420 308532 231476 308588
rect 229684 308196 229740 308252
rect 230916 308084 230972 308140
rect 229124 307524 229180 307580
rect 230132 307412 230188 307468
rect 230132 285572 230188 285628
rect 233380 307860 233436 307916
rect 232708 307412 232764 307468
rect 230692 285572 230748 285628
rect 234612 308308 234668 308364
rect 237580 308532 237636 308588
rect 237076 308420 237132 308476
rect 235284 308196 235340 308252
rect 233940 307636 233996 307692
rect 235172 307524 235228 307580
rect 237076 307972 237132 308028
rect 238532 308420 238588 308476
rect 237188 281092 237244 281148
rect 237412 307972 237468 308028
rect 240044 308420 240100 308476
rect 240436 308644 240492 308700
rect 238532 280980 238588 281036
rect 238644 308084 238700 308140
rect 238868 307636 238924 307692
rect 240324 308308 240380 308364
rect 240660 308308 240716 308364
rect 242396 308532 242452 308588
rect 241836 308420 241892 308476
rect 241220 308084 241276 308140
rect 241892 307412 241948 307468
rect 243684 308196 243740 308252
rect 247324 308644 247380 308700
rect 243572 280980 243628 281036
rect 243684 307860 243740 307916
rect 243796 281540 243852 281596
rect 245252 307524 245308 307580
rect 246708 307972 246764 308028
rect 245364 281876 245420 281932
rect 171332 280644 171388 280700
rect 247044 281764 247100 281820
rect 248724 301588 248780 301644
rect 251076 307860 251132 307916
rect 250404 307524 250460 307580
rect 248948 301476 249004 301532
rect 251972 307748 252028 307804
rect 252084 305620 252140 305676
rect 254044 308644 254100 308700
rect 252756 305620 252812 305676
rect 253428 303492 253484 303548
rect 252308 300132 252364 300188
rect 252084 300020 252140 300076
rect 254772 308644 254828 308700
rect 254772 308308 254828 308364
rect 257628 308644 257684 308700
rect 258692 308420 258748 308476
rect 253876 281652 253932 281708
rect 255332 307636 255388 307692
rect 253652 281428 253708 281484
rect 254436 281092 254492 281148
rect 246148 280868 246204 280924
rect 260764 308420 260820 308476
rect 258916 303604 258972 303660
rect 259028 299908 259084 299964
rect 260596 308084 260652 308140
rect 258804 299796 258860 299852
rect 257124 281092 257180 281148
rect 261380 307748 261436 307804
rect 262276 308532 262332 308588
rect 262052 282100 262108 282156
rect 262556 308532 262612 308588
rect 263620 308532 263676 308588
rect 263788 308420 263844 308476
rect 265524 308420 265580 308476
rect 263620 308084 263676 308140
rect 262388 282100 262444 282156
rect 263508 282100 263564 282156
rect 265076 307300 265132 307356
rect 265412 308196 265468 308252
rect 264404 306404 264460 306460
rect 266812 308420 266868 308476
rect 265636 298340 265692 298396
rect 270452 308420 270508 308476
rect 267204 281316 267260 281372
rect 267316 281540 267372 281596
rect 267540 281988 267596 282044
rect 267540 281540 267596 281596
rect 269892 281876 269948 281932
rect 267876 280868 267932 280924
rect 271740 308420 271796 308476
rect 270564 303380 270620 303436
rect 270900 296548 270956 296604
rect 272132 307972 272188 308028
rect 270452 281204 270508 281260
rect 272356 297780 272412 297836
rect 273812 308532 273868 308588
rect 272468 296436 272524 296492
rect 257684 280756 257740 280812
rect 263508 280756 263564 280812
rect 245588 280644 245644 280700
rect 273028 297780 273084 297836
rect 274764 308532 274820 308588
rect 274260 298452 274316 298508
rect 274036 298116 274092 298172
rect 275604 294756 275660 294812
rect 277284 308196 277340 308252
rect 277844 303156 277900 303212
rect 279580 308532 279636 308588
rect 280812 308420 280868 308476
rect 273812 280980 273868 281036
rect 277172 301476 277228 301532
rect 273252 280868 273308 280924
rect 270452 280644 270508 280700
rect 272580 280644 272636 280700
rect 276276 281764 276332 281820
rect 278068 301476 278124 301532
rect 278852 307524 278908 307580
rect 281540 307972 281596 308028
rect 280644 307860 280700 307916
rect 279076 303268 279132 303324
rect 278964 301588 279020 301644
rect 282100 307524 282156 307580
rect 282772 307412 282828 307468
rect 283892 308420 283948 308476
rect 282996 301924 283052 301980
rect 282324 301812 282380 301868
rect 285068 308420 285124 308476
rect 285572 308420 285628 308476
rect 283892 301700 283948 301756
rect 286972 308420 287028 308476
rect 287364 308420 287420 308476
rect 285572 302036 285628 302092
rect 287252 308308 287308 308364
rect 285796 301588 285852 301644
rect 285908 303492 285964 303548
rect 284228 300468 284284 300524
rect 283892 300132 283948 300188
rect 284452 300020 284508 300076
rect 286020 302148 286076 302204
rect 288764 308420 288820 308476
rect 289380 307188 289436 307244
rect 289716 307412 289772 307468
rect 287924 300356 287980 300412
rect 287364 300244 287420 300300
rect 289044 281652 289100 281708
rect 290052 307076 290108 307132
rect 292292 308420 292348 308476
rect 290500 306964 290556 307020
rect 293692 308420 293748 308476
rect 293972 308644 294028 308700
rect 293076 307636 293132 307692
rect 292292 300580 292348 300636
rect 294084 308420 294140 308476
rect 295484 308420 295540 308476
rect 296716 308532 296772 308588
rect 294308 303492 294364 303548
rect 300804 308420 300860 308476
rect 294532 300580 294588 300636
rect 295764 299572 295820 299628
rect 294084 298228 294140 298284
rect 290388 281428 290444 281484
rect 294196 281092 294252 281148
rect 297332 303604 297388 303660
rect 299012 300580 299068 300636
rect 299236 305620 299292 305676
rect 300244 305620 300300 305676
rect 300692 303716 300748 303772
rect 299796 299908 299852 299964
rect 299012 299796 299068 299852
rect 302204 308532 302260 308588
rect 301532 308420 301588 308476
rect 302596 308420 302652 308476
rect 301700 307972 301756 308028
rect 301476 307524 301532 307580
rect 302372 307860 302428 307916
rect 301476 281428 301532 281484
rect 303996 308420 304052 308476
rect 304164 308420 304220 308476
rect 302596 300580 302652 300636
rect 302708 305620 302764 305676
rect 303380 305620 303436 305676
rect 302820 300580 302876 300636
rect 302708 300020 302764 300076
rect 305228 308420 305284 308476
rect 307020 308644 307076 308700
rect 307524 308420 307580 308476
rect 304276 299908 304332 299964
rect 305732 308084 305788 308140
rect 306516 307524 306572 307580
rect 305844 296660 305900 296716
rect 309484 308644 309540 308700
rect 308924 308532 308980 308588
rect 308252 308420 308308 308476
rect 309204 308420 309260 308476
rect 308084 308308 308140 308364
rect 307636 299796 307692 299852
rect 307860 307412 307916 307468
rect 309092 306404 309148 306460
rect 308196 281652 308252 281708
rect 310716 308420 310772 308476
rect 310884 308420 310940 308476
rect 310212 308308 310268 308364
rect 309204 296772 309260 296828
rect 310772 307300 310828 307356
rect 311948 308420 312004 308476
rect 313180 308532 313236 308588
rect 312508 308420 312564 308476
rect 313908 308532 313964 308588
rect 310996 297220 311052 297276
rect 311332 298340 311388 298396
rect 313908 308084 313964 308140
rect 314244 308420 314300 308476
rect 315644 308420 315700 308476
rect 314244 298340 314300 298396
rect 315028 307972 315084 308028
rect 316204 308532 316260 308588
rect 317492 308420 317548 308476
rect 316036 291844 316092 291900
rect 315924 291620 315980 291676
rect 318668 308420 318724 308476
rect 320460 308532 320516 308588
rect 320964 308532 321020 308588
rect 319900 308420 319956 308476
rect 319956 307524 320012 307580
rect 320852 303380 320908 303436
rect 317716 291732 317772 291788
rect 318276 298452 318332 298508
rect 317492 291508 317548 291564
rect 316596 281764 316652 281820
rect 317268 281540 317324 281596
rect 314468 281092 314524 281148
rect 315924 281316 315980 281372
rect 318276 281316 318332 281372
rect 317828 280980 317884 281036
rect 321692 308532 321748 308588
rect 320964 292180 321020 292236
rect 321188 292180 321244 292236
rect 322980 307524 323036 307580
rect 321412 292180 321468 292236
rect 322868 296548 322924 296604
rect 324212 308420 324268 308476
rect 325388 308420 325444 308476
rect 326004 307860 326060 307916
rect 327684 305620 327740 305676
rect 324436 285460 324492 285516
rect 326676 296436 326732 296492
rect 324212 285348 324268 285404
rect 325892 284788 325948 284844
rect 324884 281204 324940 281260
rect 329364 308420 329420 308476
rect 328916 305620 328972 305676
rect 327908 285236 327964 285292
rect 327796 285012 327852 285068
rect 327684 284900 327740 284956
rect 330876 308420 330932 308476
rect 331044 308420 331100 308476
rect 330260 308308 330316 308364
rect 329476 298116 329532 298172
rect 331996 308420 332052 308476
rect 332668 308420 332724 308476
rect 329588 284900 329644 284956
rect 332724 294756 332780 294812
rect 335748 307748 335804 307804
rect 335860 302314 335916 302316
rect 335860 302262 335862 302314
rect 335862 302262 335914 302314
rect 335914 302262 335916 302314
rect 335860 302260 335916 302262
rect 330932 280868 330988 280924
rect 306404 280756 306460 280812
rect 328132 280644 328188 280700
rect 332612 281316 332668 281372
rect 334404 282100 334460 282156
rect 334628 282100 334684 282156
rect 335748 301476 335804 301532
rect 335412 300468 335468 300524
rect 335412 281988 335468 282044
rect 335524 298340 335580 298396
rect 336364 308420 336420 308476
rect 337092 308644 337148 308700
rect 336084 293076 336140 293132
rect 336420 308196 336476 308252
rect 335748 281316 335804 281372
rect 336644 307636 336700 307692
rect 336644 299684 336700 299740
rect 336756 307524 336812 307580
rect 336868 301476 336924 301532
rect 337204 307412 337260 307468
rect 337092 306852 337148 306908
rect 337092 301588 337148 301644
rect 336980 294980 337036 295036
rect 337204 294868 337260 294924
rect 337652 303156 337708 303212
rect 336756 289940 336812 289996
rect 337540 289156 337596 289212
rect 341180 308644 341236 308700
rect 343644 308644 343700 308700
rect 356412 308644 356468 308700
rect 337988 288260 338044 288316
rect 339332 303268 339388 303324
rect 337764 288036 337820 288092
rect 338996 281316 339052 281372
rect 339444 288148 339500 288204
rect 341796 303492 341852 303548
rect 341572 281652 341628 281708
rect 344932 307636 344988 307692
rect 344260 306292 344316 306348
rect 345492 303828 345548 303884
rect 347956 304724 348012 304780
rect 349748 305620 349804 305676
rect 351652 305508 351708 305564
rect 352212 305396 352268 305452
rect 352884 305284 352940 305340
rect 358932 307300 358988 307356
rect 362572 308420 362628 308476
rect 363132 308420 363188 308476
rect 357140 306404 357196 306460
rect 348516 304612 348572 304668
rect 346724 303716 346780 303772
rect 359380 303604 359436 303660
rect 361172 307188 361228 307244
rect 342468 303044 342524 303100
rect 362852 307076 362908 307132
rect 348516 301924 348572 301980
rect 345156 299572 345212 299628
rect 341796 281652 341852 281708
rect 344148 281876 344204 281932
rect 342804 281540 342860 281596
rect 346724 281428 346780 281484
rect 349748 301812 349804 301868
rect 354900 301812 354956 301868
rect 352772 301700 352828 301756
rect 351764 281988 351820 282044
rect 354340 281652 354396 281708
rect 356132 301364 356188 301420
rect 359492 300356 359548 300412
rect 358484 281428 358540 281484
rect 359940 300244 359996 300300
rect 362740 281428 362796 281484
rect 364420 305060 364476 305116
rect 364532 306964 364588 307020
rect 368620 308420 368676 308476
rect 369852 308644 369908 308700
rect 364980 305172 365036 305228
rect 367444 304948 367500 305004
rect 369348 304836 369404 304892
rect 370916 308644 370972 308700
rect 369572 299684 369628 299740
rect 370916 307524 370972 307580
rect 371700 307188 371756 307244
rect 372372 307076 372428 307132
rect 376964 308532 377020 308588
rect 371028 306964 371084 307020
rect 372820 303940 372876 303996
rect 374164 306852 374220 306908
rect 374836 303492 374892 303548
rect 373604 303380 373660 303436
rect 375396 303268 375452 303324
rect 376628 308084 376684 308140
rect 375956 303156 376012 303212
rect 377300 308698 377356 308700
rect 377300 308646 377302 308698
rect 377302 308646 377354 308698
rect 377354 308646 377356 308698
rect 377300 308644 377356 308646
rect 377132 308420 377188 308476
rect 377412 308308 377468 308364
rect 378084 308420 378140 308476
rect 377860 307412 377916 307468
rect 369684 291396 369740 291452
rect 376628 300468 376684 300524
rect 373604 281540 373660 281596
rect 372260 281204 372316 281260
rect 377188 281540 377244 281596
rect 379036 308420 379092 308476
rect 377524 281428 377580 281484
rect 374612 280868 374668 280924
rect 370468 280644 370524 280700
rect 414932 307972 414988 308028
rect 381780 299684 381836 299740
rect 381220 281764 381276 281820
rect 388164 300132 388220 300188
rect 391524 300020 391580 300076
rect 389732 299684 389788 299740
rect 393316 299908 393372 299964
rect 392756 282100 392812 282156
rect 399812 299796 399868 299852
rect 398580 280980 398636 281036
rect 403508 294980 403564 295036
rect 404852 294868 404908 294924
rect 406868 281316 406924 281372
rect 410676 281764 410732 281820
rect 412020 281652 412076 281708
rect 414596 281092 414652 281148
rect 418292 293188 418348 293244
rect 418964 291844 419020 291900
rect 421652 291732 421708 291788
rect 420196 291620 420252 291676
rect 438452 307860 438508 307916
rect 426692 307412 426748 307468
rect 423332 285572 423388 285628
rect 423444 291508 423500 291564
rect 424116 285572 424172 285628
rect 426132 281540 426188 281596
rect 428820 291844 428876 291900
rect 428596 291732 428652 291788
rect 428596 285572 428652 285628
rect 430388 291508 430444 291564
rect 429268 285572 429324 285628
rect 432516 289940 432572 289996
rect 436324 285124 436380 285180
rect 437668 285012 437724 285068
rect 442708 284900 442764 284956
rect 441476 284788 441532 284844
rect 444052 284564 444108 284620
rect 445284 282100 445340 282156
rect 446628 282100 446684 282156
rect 447860 281428 447916 281484
rect 453012 281204 453068 281260
rect 548436 308084 548492 308140
rect 532420 307748 532476 307804
rect 463764 294756 463820 294812
rect 463764 290724 463820 290780
rect 465332 293076 465388 293132
rect 465332 292292 465388 292348
rect 482916 307636 482972 307692
rect 481236 306292 481292 306348
rect 472052 290276 472108 290332
rect 470932 288372 470988 288428
rect 468580 287252 468636 287308
rect 461748 280868 461804 280924
rect 462644 280868 462700 280924
rect 469140 287252 469196 287308
rect 472836 288036 472892 288092
rect 475412 290500 475468 290556
rect 474516 287252 474572 287308
rect 481236 290388 481292 290444
rect 477876 290276 477932 290332
rect 478660 290276 478716 290332
rect 477876 280868 477932 280924
rect 479556 289268 479612 289324
rect 479556 289044 479612 289100
rect 508116 306404 508172 306460
rect 485492 303716 485548 303772
rect 483812 294084 483868 294140
rect 485492 293972 485548 294028
rect 482916 290500 482972 290556
rect 489636 304724 489692 304780
rect 488852 304612 488908 304668
rect 488852 292852 488908 292908
rect 488852 285572 488908 285628
rect 489076 292628 489132 292684
rect 489636 292628 489692 292684
rect 490644 293860 490700 293916
rect 491316 293860 491372 293916
rect 492996 305620 493052 305676
rect 490644 292852 490700 292908
rect 483028 280868 483084 280924
rect 489524 285572 489580 285628
rect 496356 305508 496412 305564
rect 494676 293636 494732 293692
rect 493892 292292 493948 292348
rect 493892 285572 493948 285628
rect 494676 292292 494732 292348
rect 497252 305396 497308 305452
rect 494564 285572 494620 285628
rect 497252 292516 497308 292572
rect 498932 305284 498988 305340
rect 498932 292740 498988 292796
rect 499716 292292 499772 292348
rect 502292 294308 502348 294364
rect 503972 294196 504028 294252
rect 507332 292180 507388 292236
rect 505988 291508 506044 291564
rect 509012 293860 509068 293916
rect 509796 293860 509852 293916
rect 509012 292516 509068 292572
rect 508116 292180 508172 292236
rect 508116 291732 508172 291788
rect 510692 307300 510748 307356
rect 520548 303940 520604 303996
rect 510692 292964 510748 293020
rect 513156 303604 513212 303660
rect 512372 292740 512428 292796
rect 513156 292740 513212 292796
rect 514052 293860 514108 293916
rect 514836 293860 514892 293916
rect 514052 292964 514108 293020
rect 524916 305172 524972 305228
rect 523236 305060 523292 305116
rect 522340 303716 522396 303772
rect 522676 292180 522732 292236
rect 523236 292180 523292 292236
rect 522676 291060 522732 291116
rect 521332 290948 521388 291004
rect 524132 291172 524188 291228
rect 524916 291172 524972 291228
rect 525924 291508 525980 291564
rect 526596 291508 526652 291564
rect 529956 304948 530012 305004
rect 534212 307524 534268 307580
rect 532532 304836 532588 304892
rect 532532 291284 532588 291340
rect 539252 307076 539308 307132
rect 534212 291620 534268 291676
rect 538356 306964 538412 307020
rect 535892 291396 535948 291452
rect 535892 290836 535948 290892
rect 537572 291396 537628 291452
rect 538356 291396 538412 291452
rect 543396 306852 543452 306908
rect 539252 293412 539308 293468
rect 542612 293860 542668 293916
rect 545076 303492 545132 303548
rect 543396 293860 543452 293916
rect 543508 303380 543564 303436
rect 542612 293076 542668 293132
rect 540932 292180 540988 292236
rect 540932 290836 540988 290892
rect 542724 292180 542780 292236
rect 543508 292180 543564 292236
rect 543508 291508 543564 291564
rect 544404 293860 544460 293916
rect 545076 293860 545132 293916
rect 546756 303268 546812 303324
rect 544404 293188 544460 293244
rect 538244 280868 538300 280924
rect 545972 293300 546028 293356
rect 546756 293300 546812 293356
rect 547652 293412 547708 293468
rect 551012 307412 551068 307468
rect 548548 303156 548604 303212
rect 548548 293412 548604 293468
rect 549556 293860 549612 293916
rect 548436 291620 548492 291676
rect 556724 284676 556780 284732
rect 560196 301588 560252 301644
rect 559076 280868 559132 280924
rect 402388 280756 402444 280812
rect 379764 280644 379820 280700
rect 554820 280644 554876 280700
rect 559636 254324 559692 254380
rect 560084 251972 560140 252028
rect 559636 235172 559692 235228
rect 559748 240212 559804 240268
rect 559972 233828 560028 233884
rect 559748 217924 559804 217980
rect 559860 231588 559916 231644
rect 560084 232708 560140 232764
rect 559972 209076 560028 209132
rect 560084 220388 560140 220444
rect 559860 206164 559916 206220
rect 560084 191380 560140 191436
rect 90356 191268 90412 191324
rect 84308 190932 84364 190988
rect 559412 141652 559468 141708
rect 566020 301476 566076 301532
rect 560420 256564 560476 256620
rect 560868 249620 560924 249676
rect 560644 247492 560700 247548
rect 560532 240660 560588 240716
rect 560532 240212 560588 240268
rect 560420 238420 560476 238476
rect 560420 236180 560476 236236
rect 560868 229124 560924 229180
rect 560980 245252 561036 245308
rect 560644 226212 560700 226268
rect 560868 224756 560924 224812
rect 560644 222516 560700 222572
rect 560532 211540 560588 211596
rect 560420 206612 560476 206668
rect 560308 185668 560364 185724
rect 560308 182980 560364 183036
rect 560980 223300 561036 223356
rect 561876 238420 561932 238476
rect 560868 196756 560924 196812
rect 560980 215684 561036 215740
rect 560644 193844 560700 193900
rect 560868 195188 560924 195244
rect 560756 192948 560812 193004
rect 560644 190708 560700 190764
rect 560532 182980 560588 183036
rect 560532 181636 560588 181692
rect 560420 173796 560476 173852
rect 560420 167972 560476 168028
rect 560196 135604 560252 135660
rect 560308 154308 560364 154364
rect 559412 81620 559468 81676
rect 92372 80890 92428 80892
rect 92372 80838 92374 80890
rect 92374 80838 92426 80890
rect 92426 80838 92428 80890
rect 92372 80836 92428 80838
rect 335972 80778 336028 80780
rect 335972 80726 335974 80778
rect 335974 80726 336026 80778
rect 336026 80726 336028 80778
rect 335972 80724 336028 80726
rect 190596 79044 190652 79100
rect 123508 78932 123564 78988
rect 324884 72100 324940 72156
rect 561876 214452 561932 214508
rect 565236 229348 565292 229404
rect 565236 202020 565292 202076
rect 560980 184996 561036 185052
rect 560868 158564 560924 158620
rect 561876 172564 561932 172620
rect 560756 155652 560812 155708
rect 560644 152740 560700 152796
rect 561876 120372 561932 120428
rect 565236 156660 565292 156716
rect 560532 117460 560588 117516
rect 560308 100324 560364 100380
rect 606116 294084 606172 294140
rect 605780 292628 605836 292684
rect 606228 291844 606284 291900
rect 609812 292292 609868 292348
rect 609812 290948 609868 291004
rect 606340 290218 606396 290220
rect 606340 290166 606342 290218
rect 606342 290166 606394 290218
rect 606394 290166 606396 290218
rect 606340 290164 606396 290166
rect 600516 289156 600572 289212
rect 570500 281204 570556 281260
rect 570388 280980 570444 281036
rect 570276 280756 570332 280812
rect 570388 277060 570444 277116
rect 570500 270340 570556 270396
rect 570276 270228 570332 270284
rect 597156 261156 597212 261212
rect 585396 258804 585452 258860
rect 583716 242900 583772 242956
rect 566916 226996 566972 227052
rect 583716 220164 583772 220220
rect 578676 217924 578732 217980
rect 566916 199108 566972 199164
rect 568596 213444 568652 213500
rect 568596 181412 568652 181468
rect 568708 211092 568764 211148
rect 570612 204372 570668 204428
rect 570500 202020 570556 202076
rect 568708 178500 568764 178556
rect 570276 199780 570332 199836
rect 570276 163828 570332 163884
rect 570388 197540 570444 197596
rect 570612 169652 570668 169708
rect 571956 188468 572012 188524
rect 570500 166740 570556 166796
rect 570388 161252 570444 161308
rect 578676 186452 578732 186508
rect 571956 149492 572012 149548
rect 575316 152068 575372 152124
rect 575316 102452 575372 102508
rect 565236 96180 565292 96236
rect 560308 81844 560364 81900
rect 597156 240324 597212 240380
rect 585396 81620 585452 81676
rect 585620 179284 585676 179340
rect 585844 165732 585900 165788
rect 586068 163380 586124 163436
rect 598836 149828 598892 149884
rect 598836 92372 598892 92428
rect 609812 289156 609868 289212
rect 606340 288148 606396 288204
rect 606228 288036 606284 288092
rect 623252 332612 623308 332668
rect 613284 328692 613340 328748
rect 626612 333284 626668 333340
rect 629188 330148 629244 330204
rect 631204 330036 631260 330092
rect 635124 328580 635180 328636
rect 643076 328468 643132 328524
rect 649012 332052 649068 332108
rect 647108 326676 647164 326732
rect 658980 331940 659036 331996
rect 660996 328804 661052 328860
rect 650132 325108 650188 325164
rect 666932 329140 666988 329196
rect 661892 324884 661948 324940
rect 672308 332554 672364 332556
rect 672308 332502 672310 332554
rect 672310 332502 672362 332554
rect 672362 332502 672364 332554
rect 672308 332500 672364 332502
rect 671300 332052 671356 332108
rect 670292 308756 670348 308812
rect 671076 331940 671132 331996
rect 657636 306740 657692 306796
rect 659316 306628 659372 306684
rect 662676 301588 662732 301644
rect 670628 301700 670684 301756
rect 657636 301476 657692 301532
rect 624708 294308 624764 294364
rect 618548 293972 618604 294028
rect 613508 292068 613564 292124
rect 610932 289940 610988 289996
rect 610708 288260 610764 288316
rect 611380 289604 611436 289660
rect 614404 290612 614460 290668
rect 614180 290052 614236 290108
rect 615412 290500 615468 290556
rect 615300 290388 615356 290444
rect 614740 290330 614796 290332
rect 614740 290278 614742 290330
rect 614742 290278 614794 290330
rect 614794 290278 614796 290330
rect 614740 290276 614796 290278
rect 614852 290164 614908 290220
rect 615636 290500 615692 290556
rect 617092 290500 617148 290556
rect 616084 290388 616140 290444
rect 616532 290164 616588 290220
rect 617540 290052 617596 290108
rect 621908 293636 621964 293692
rect 620900 292068 620956 292124
rect 619892 290388 619948 290444
rect 620452 290164 620508 290220
rect 621348 291844 621404 291900
rect 623812 292404 623868 292460
rect 622804 289716 622860 289772
rect 623252 289716 623308 289772
rect 625268 294196 625324 294252
rect 628628 292740 628684 292796
rect 627172 292516 627228 292572
rect 626612 291732 626668 291788
rect 626164 289716 626220 289772
rect 628068 289716 628124 289772
rect 629076 289716 629132 289772
rect 642068 291620 642124 291676
rect 633332 291284 633388 291340
rect 632884 291172 632940 291228
rect 632436 291060 632492 291116
rect 631988 289716 632044 289772
rect 639604 291508 639660 291564
rect 637700 291396 637756 291452
rect 637252 290500 637308 290556
rect 636244 289716 636300 289772
rect 636692 289716 636748 289772
rect 639156 290836 639212 290892
rect 638148 289716 638204 289772
rect 638708 289716 638764 289772
rect 640052 289716 640108 289772
rect 640612 289716 640668 289772
rect 641060 289716 641116 289772
rect 641508 289716 641564 289772
rect 642964 290724 643020 290780
rect 642740 290052 642796 290108
rect 642516 289716 642572 289772
rect 642740 289716 642796 289772
rect 643524 290500 643580 290556
rect 644868 290948 644924 291004
rect 644420 289716 644476 289772
rect 648788 291620 648844 291676
rect 647332 291508 647388 291564
rect 645876 291396 645932 291452
rect 646884 290052 646940 290108
rect 648228 290164 648284 290220
rect 651588 289828 651644 289884
rect 652596 289828 652652 289884
rect 653044 289716 653100 289772
rect 669396 291956 669452 292012
rect 658868 290612 658924 290668
rect 655508 289716 655564 289772
rect 656964 289940 657020 289996
rect 657412 289828 657468 289884
rect 658308 289716 658364 289772
rect 668388 290500 668444 290556
rect 666036 290388 666092 290444
rect 662676 290164 662732 290220
rect 661668 289716 661724 289772
rect 664132 290052 664188 290108
rect 663124 289828 663180 289884
rect 667156 290052 667212 290108
rect 666932 289716 666988 289772
rect 667268 289716 667324 289772
rect 667492 289716 667548 289772
rect 670068 290612 670124 290668
rect 670292 289828 670348 289884
rect 671076 291508 671132 291564
rect 671188 301588 671244 301644
rect 672196 331828 672252 331884
rect 672084 331716 672140 331772
rect 671524 313236 671580 313292
rect 671524 291620 671580 291676
rect 671300 291396 671356 291452
rect 671188 289940 671244 289996
rect 670852 289716 670908 289772
rect 672084 290164 672140 290220
rect 611380 288874 611436 288876
rect 611380 288822 611382 288874
rect 611382 288822 611434 288874
rect 611434 288822 611436 288874
rect 611380 288820 611436 288822
rect 611044 288148 611100 288204
rect 672868 328356 672924 328412
rect 673204 332612 673260 332668
rect 678916 332612 678972 332668
rect 673652 324996 673708 325052
rect 683732 324100 683788 324156
rect 682052 323988 682108 324044
rect 680372 322532 680428 322588
rect 672420 290276 672476 290332
rect 672308 289828 672364 289884
rect 671860 283780 671916 283836
rect 609924 283108 609980 283164
rect 605556 281540 605612 281596
rect 603876 274708 603932 274764
rect 602308 272468 602364 272524
rect 602196 267988 602252 268044
rect 600628 265636 600684 265692
rect 605556 270340 605612 270396
rect 607236 279300 607292 279356
rect 607236 267092 607292 267148
rect 603876 260372 603932 260428
rect 602308 257012 602364 257068
rect 602196 252084 602252 252140
rect 600628 248724 600684 248780
rect 605556 183876 605612 183932
rect 603876 177044 603932 177100
rect 600628 161140 600684 161196
rect 603876 127652 603932 127708
rect 603988 170212 604044 170268
rect 605556 139412 605612 139468
rect 605668 174804 605724 174860
rect 671748 154532 671804 154588
rect 671860 149940 671916 149996
rect 672756 147588 672812 147644
rect 671860 142100 671916 142156
rect 672196 142996 672252 143052
rect 671748 141092 671804 141148
rect 671972 141540 672028 141596
rect 611716 140084 611772 140140
rect 605668 131012 605724 131068
rect 611492 131796 611548 131852
rect 603988 122612 604044 122668
rect 600628 107492 600684 107548
rect 586068 81396 586124 81452
rect 585844 81284 585900 81340
rect 585620 81172 585676 81228
rect 560196 79044 560252 79100
rect 561876 78932 561932 78988
rect 526372 72100 526428 72156
rect 560980 72100 561036 72156
rect 459172 71988 459228 72044
rect 506772 71876 506828 71932
rect 392084 71764 392140 71820
rect 341684 71428 341740 71484
rect 257796 70532 257852 70588
rect 176182 70084 176238 70140
rect 231182 70084 231238 70140
rect 396036 70532 396092 70588
rect 454580 71652 454636 71708
rect 451181 70084 451237 70140
rect 454580 70084 454636 70140
rect 450890 69748 450946 69804
rect 494287 70084 494343 70140
rect 548548 71764 548604 71820
rect 505890 70084 505946 70140
rect 548432 70084 548488 70140
rect 560890 70532 560946 70588
rect 549287 70308 549343 70364
rect 624036 140084 624092 140140
rect 619108 139972 619164 140028
rect 618884 139860 618940 139916
rect 611492 71540 611548 71596
rect 612164 131796 612220 131852
rect 614628 71652 614684 71708
rect 617316 71876 617372 71932
rect 613956 71428 614012 71484
rect 618324 134596 618380 134652
rect 618436 134372 618492 134428
rect 618548 139412 618604 139468
rect 618324 89908 618380 89964
rect 618436 86212 618492 86268
rect 618660 122612 618716 122668
rect 623364 139972 623420 140028
rect 624708 139972 624764 140028
rect 657076 139972 657132 140028
rect 657748 139972 657804 140028
rect 630756 139860 630812 139916
rect 631428 139860 631484 139916
rect 619108 139412 619164 139468
rect 618996 96180 619052 96236
rect 619108 125412 619164 125468
rect 618884 93716 618940 93772
rect 619108 92484 619164 92540
rect 618660 82516 618716 82572
rect 618548 81284 618604 81340
rect 620452 134484 620508 134540
rect 622692 139748 622748 139804
rect 622020 139636 622076 139692
rect 624932 139524 624988 139580
rect 621460 139412 621516 139468
rect 621348 134596 621404 134652
rect 621124 134372 621180 134428
rect 626052 125860 626108 125916
rect 628068 125860 628124 125916
rect 628740 125860 628796 125916
rect 632772 139636 632828 139692
rect 636132 135604 636188 135660
rect 635460 135380 635516 135436
rect 638820 139636 638876 139692
rect 638148 135492 638204 135548
rect 637476 135268 637532 135324
rect 636804 135156 636860 135212
rect 630084 125412 630140 125468
rect 642292 126756 642348 126812
rect 641508 125860 641564 125916
rect 643636 127540 643692 127596
rect 646324 127428 646380 127484
rect 645652 127204 645708 127260
rect 644980 126980 645036 127036
rect 644308 126868 644364 126924
rect 646996 125972 647052 126028
rect 655732 139860 655788 139916
rect 665140 139860 665196 139916
rect 659092 139748 659148 139804
rect 650692 139636 650748 139692
rect 649012 139412 649068 139468
rect 649460 136276 649516 136332
rect 653716 136276 653772 136332
rect 656404 139636 656460 139692
rect 659988 139524 660044 139580
rect 658420 139412 658476 139468
rect 660436 137956 660492 138012
rect 662452 137844 662508 137900
rect 661780 137732 661836 137788
rect 666484 139636 666540 139692
rect 667828 139636 667884 139692
rect 664468 138964 664524 139020
rect 663796 138740 663852 138796
rect 663460 136948 663516 137004
rect 661556 136836 661612 136892
rect 655060 136164 655116 136220
rect 654388 136052 654444 136108
rect 669620 139412 669676 139468
rect 669508 134932 669564 134988
rect 650020 134820 650076 134876
rect 650122 133028 650178 133084
rect 649572 132692 649628 132748
rect 654378 132580 654434 132636
rect 656394 132580 656450 132636
rect 657972 132580 658028 132636
rect 664580 132580 664636 132636
rect 666922 132580 666978 132636
rect 667594 132580 667650 132636
rect 670180 132580 670236 132636
rect 650692 132356 650748 132412
rect 649236 132244 649292 132300
rect 651578 132244 651634 132300
rect 649124 132132 649180 132188
rect 652250 132132 652306 132188
rect 648900 132020 648956 132076
rect 654836 132468 654892 132524
rect 655722 132244 655778 132300
rect 653594 132132 653650 132188
rect 657178 132132 657234 132188
rect 652922 132020 652978 132076
rect 659652 132468 659708 132524
rect 657850 132020 657906 132076
rect 648340 131572 648396 131628
rect 654724 131572 654780 131628
rect 647668 125972 647724 126028
rect 642964 125748 643020 125804
rect 640836 125636 640892 125692
rect 640164 125524 640220 125580
rect 639492 125412 639548 125468
rect 629412 125300 629468 125356
rect 627396 125188 627452 125244
rect 626724 125076 626780 125132
rect 627284 123396 627340 123452
rect 622132 123284 622188 123340
rect 660650 132244 660706 132300
rect 661994 132468 662050 132524
rect 661322 132132 661378 132188
rect 660100 131460 660156 131516
rect 663460 131796 663516 131852
rect 663236 131348 663292 131404
rect 665924 131908 665980 131964
rect 668266 132468 668322 132524
rect 668938 132020 668994 132076
rect 671524 132020 671580 132076
rect 666596 131684 666652 131740
rect 671636 131684 671692 131740
rect 665140 131012 665196 131068
rect 655396 127204 655452 127260
rect 655172 126980 655228 127036
rect 654948 125188 655004 125244
rect 641172 123338 641228 123340
rect 641172 123286 641174 123338
rect 641174 123286 641226 123338
rect 641226 123286 641228 123338
rect 641172 123284 641228 123286
rect 642740 123284 642796 123340
rect 647892 123284 647948 123340
rect 654948 116564 655004 116620
rect 655060 125076 655116 125132
rect 655060 114996 655116 115052
rect 619780 100548 619836 100604
rect 620564 100660 620620 100716
rect 625380 100660 625436 100716
rect 623364 100436 623420 100492
rect 647556 100660 647612 100716
rect 628628 100436 628684 100492
rect 631204 100436 631260 100492
rect 649572 100436 649628 100492
rect 652148 100436 652204 100492
rect 633780 99988 633836 100044
rect 635796 99988 635852 100044
rect 639044 99988 639100 100044
rect 641732 99988 641788 100044
rect 644980 99988 645036 100044
rect 619556 98980 619612 99036
rect 655284 126868 655340 126924
rect 655396 110180 655452 110236
rect 655956 126644 656012 126700
rect 655284 109620 655340 109676
rect 655172 92260 655228 92316
rect 670180 123508 670236 123564
rect 655956 85540 656012 85596
rect 628068 80612 628124 80668
rect 645092 80612 645148 80668
rect 671972 74452 672028 74508
rect 672084 140756 672140 140812
rect 672196 83412 672252 83468
rect 672084 74228 672140 74284
rect 673540 142660 673596 142716
rect 673540 94052 673596 94108
rect 686420 176372 686476 176428
rect 686532 353556 686588 353612
rect 686868 513940 686924 513996
rect 686644 333956 686700 334012
rect 686756 473732 686812 473788
rect 686868 262164 686924 262220
rect 686980 335972 687036 336028
rect 686756 218372 686812 218428
rect 688212 937354 688268 937356
rect 688212 937302 688214 937354
rect 688214 937302 688266 937354
rect 688266 937302 688268 937354
rect 688212 937300 688268 937302
rect 688996 937188 689052 937244
rect 688436 936964 688492 937020
rect 688212 936740 688268 936796
rect 687876 936628 687932 936684
rect 687988 936516 688044 936572
rect 688212 333396 688268 333452
rect 688324 672756 688380 672812
rect 687988 332052 688044 332108
rect 687876 331940 687932 331996
rect 687764 313236 687820 313292
rect 688212 290442 688268 290444
rect 688212 290390 688214 290442
rect 688214 290390 688266 290442
rect 688266 290390 688268 290442
rect 688212 290388 688268 290390
rect 687652 289716 687708 289772
rect 687540 289156 687596 289212
rect 687316 281428 687372 281484
rect 687204 274484 687260 274540
rect 688884 936404 688940 936460
rect 688996 672756 689052 672812
rect 688996 580692 689052 580748
rect 689108 394100 689164 394156
rect 689108 335972 689164 336028
rect 688996 334180 689052 334236
rect 695380 935508 695436 935564
rect 694820 934836 694876 934892
rect 694708 934724 694764 934780
rect 693812 934500 693868 934556
rect 691348 910756 691404 910812
rect 689556 910532 689612 910588
rect 689332 290554 689388 290556
rect 689332 290502 689334 290554
rect 689334 290502 689386 290554
rect 689386 290502 689388 290554
rect 689332 290500 689388 290502
rect 689220 269892 689276 269948
rect 688436 267652 688492 267708
rect 688324 260708 688380 260764
rect 691236 908516 691292 908572
rect 689556 249172 689612 249228
rect 689668 824852 689724 824908
rect 689780 739172 689836 739228
rect 689780 242228 689836 242284
rect 689892 695492 689948 695548
rect 689668 235284 689724 235340
rect 689892 228340 689948 228396
rect 690004 651812 690060 651868
rect 690004 221508 690060 221564
rect 690116 566132 690172 566188
rect 690116 207620 690172 207676
rect 690228 524132 690284 524188
rect 691348 900788 691404 900844
rect 693028 860692 693084 860748
rect 691236 253764 691292 253820
rect 692916 822500 692972 822556
rect 693812 822948 693868 823004
rect 694484 934276 694540 934332
rect 693028 806932 693084 806988
rect 693028 780724 693084 780780
rect 693028 719796 693084 719852
rect 694596 873572 694652 873628
rect 694596 736036 694652 736092
rect 694484 609700 694540 609756
rect 694596 607460 694652 607516
rect 693140 500724 693196 500780
rect 692916 239876 692972 239932
rect 693028 420756 693084 420812
rect 690228 200676 690284 200732
rect 693140 265748 693196 265804
rect 693252 460740 693308 460796
rect 694820 822052 694876 822108
rect 695156 934388 695212 934444
rect 694708 566804 694764 566860
rect 694820 693028 694876 693084
rect 694596 219156 694652 219212
rect 694708 564452 694764 564508
rect 695156 607908 695212 607964
rect 694820 334068 694876 334124
rect 694932 566692 694988 566748
rect 697956 925092 698012 925148
rect 700532 934612 700588 934668
rect 705012 927220 705068 927276
rect 703892 927108 703948 927164
rect 704836 926324 704892 926380
rect 705732 926324 705788 926380
rect 700532 908068 700588 908124
rect 699188 891492 699244 891548
rect 696276 887012 696332 887068
rect 696276 736932 696332 736988
rect 698740 840532 698796 840588
rect 700196 891380 700252 891436
rect 699748 891268 699804 891324
rect 699412 890596 699468 890652
rect 699188 752500 699244 752556
rect 699300 805476 699356 805532
rect 698740 720132 698796 720188
rect 700084 838292 700140 838348
rect 699972 823060 700028 823116
rect 699748 806372 699804 806428
rect 699860 821828 699916 821884
rect 699412 752500 699468 752556
rect 699524 805364 699580 805420
rect 699524 712180 699580 712236
rect 699748 804916 699804 804972
rect 699300 712068 699356 712124
rect 699860 720244 699916 720300
rect 704836 891492 704892 891548
rect 705284 891380 705340 891436
rect 704388 891268 704444 891324
rect 705572 890596 705628 890652
rect 704388 840532 704444 840588
rect 704836 840308 704892 840364
rect 705284 840308 705340 840364
rect 705732 840308 705788 840364
rect 700644 838292 700700 838348
rect 700644 823060 700700 823116
rect 701428 824732 701484 824788
rect 701428 819924 701484 819980
rect 704388 805364 704444 805420
rect 700196 755636 700252 755692
rect 701316 805252 701372 805308
rect 700084 720356 700140 720412
rect 699972 719012 700028 719068
rect 705284 805476 705340 805532
rect 704836 805252 704892 805308
rect 705572 804916 705628 804972
rect 704388 755636 704444 755692
rect 705124 755076 705180 755132
rect 704836 754404 704892 754460
rect 705732 754404 705788 754460
rect 704388 720356 704444 720412
rect 704836 720244 704892 720300
rect 705284 720132 705340 720188
rect 700644 719796 700700 719852
rect 699748 710500 699804 710556
rect 705572 719012 705628 719068
rect 705012 712180 705068 712236
rect 703892 712068 703948 712124
rect 705732 711396 705788 711452
rect 700644 697060 700700 697116
rect 701540 697060 701596 697116
rect 701540 695732 701596 695788
rect 704836 676564 704892 676620
rect 704388 676452 704444 676508
rect 705284 676340 705340 676396
rect 705684 675444 705740 675500
rect 700532 671076 700588 671132
rect 704676 669060 704732 669116
rect 704388 668500 704444 668556
rect 705284 668500 705340 668556
rect 705732 668388 705788 668444
rect 700532 652708 700588 652764
rect 704388 633556 704444 633612
rect 704836 633444 704892 633500
rect 705284 633332 705340 633388
rect 705732 633332 705788 633388
rect 704388 626500 704444 626556
rect 705284 626276 705340 626332
rect 705732 626276 705788 626332
rect 704836 625380 704892 625436
rect 704836 590436 704892 590492
rect 705284 590324 705340 590380
rect 704388 590212 704444 590268
rect 705684 589764 705740 589820
rect 704836 583268 704892 583324
rect 704004 582820 704060 582876
rect 705284 582820 705340 582876
rect 705732 582372 705788 582428
rect 705012 547876 705068 547932
rect 704564 547764 704620 547820
rect 704388 547652 704444 547708
rect 705572 543396 705628 543452
rect 704564 540148 704620 540204
rect 704676 540036 704732 540092
rect 705124 540036 705180 540092
rect 705732 539364 705788 539420
rect 695380 522004 695436 522060
rect 696276 521444 696332 521500
rect 695156 351764 695212 351820
rect 695156 334180 695212 334236
rect 695380 349076 695436 349132
rect 695380 333956 695436 334012
rect 694932 306964 694988 307020
rect 695156 306516 695212 306572
rect 694708 212212 694764 212268
rect 694820 266196 694876 266252
rect 693028 179732 693084 179788
rect 694596 180180 694652 180236
rect 694820 179956 694876 180012
rect 694932 223188 694988 223244
rect 695044 220500 695100 220556
rect 704388 504532 704444 504588
rect 704836 504420 704892 504476
rect 705284 504308 705340 504364
rect 705572 504084 705628 504140
rect 700532 487956 700588 488012
rect 704564 368116 704620 368172
rect 704004 367780 704060 367836
rect 705284 367780 705340 367836
rect 705732 367332 705788 367388
rect 700532 349972 700588 350028
rect 704836 333060 704892 333116
rect 705012 332836 705068 332892
rect 705572 332724 705628 332780
rect 704388 332612 704444 332668
rect 704004 325108 704060 325164
rect 705124 325108 705180 325164
rect 704564 324996 704620 325052
rect 705732 324324 705788 324380
rect 704676 289828 704732 289884
rect 705012 289828 705068 289884
rect 704836 289380 704892 289436
rect 705572 289044 705628 289100
rect 704676 282100 704732 282156
rect 705012 281988 705068 282044
rect 704836 281876 704892 281932
rect 705732 281316 705788 281372
rect 696276 205268 696332 205324
rect 697956 263508 698012 263564
rect 695156 191492 695212 191548
rect 704676 246820 704732 246876
rect 704564 239092 704620 239148
rect 705284 246260 705340 246316
rect 705284 238420 705340 238476
rect 700532 222740 700588 222796
rect 704836 203476 704892 203532
rect 705732 203588 705788 203644
rect 705284 203364 705340 203420
rect 704388 203252 704444 203308
rect 704564 196196 704620 196252
rect 703892 196084 703948 196140
rect 705012 195972 705068 196028
rect 705732 195412 705788 195468
rect 697956 184548 698012 184604
rect 695044 177604 695100 177660
rect 694932 173012 694988 173068
rect 694596 166068 694652 166124
rect 694708 163828 694764 163884
rect 686980 132692 687036 132748
rect 694596 156884 694652 156940
rect 705012 160804 705068 160860
rect 704836 160356 704892 160412
rect 704388 160244 704444 160300
rect 705572 159684 705628 159740
rect 700532 159124 700588 159180
rect 704388 152740 704444 152796
rect 705284 152740 705340 152796
rect 704836 152516 704892 152572
rect 705732 152404 705788 152460
rect 700532 137172 700588 137228
rect 694708 134484 694764 134540
rect 704836 118020 704892 118076
rect 704676 117796 704732 117852
rect 705572 117684 705628 117740
rect 705012 117572 705068 117628
rect 704004 110068 704060 110124
rect 705012 110068 705068 110124
rect 704564 109956 704620 110012
rect 705732 109396 705788 109452
rect 694596 91476 694652 91532
rect 686532 90804 686588 90860
rect 686308 90692 686364 90748
rect 672756 74004 672812 74060
rect 672980 83412 673036 83468
rect 705284 74452 705340 74508
rect 704836 74228 704892 74284
rect 704340 74004 704396 74060
rect 672980 73892 673036 73948
rect 705684 73892 705740 73948
rect 619332 71092 619388 71148
rect 617988 70980 618044 71036
rect 469140 69748 469196 69804
rect 506036 69748 506092 69804
<< metal3 >>
rect 470250 949172 470260 949228
rect 470316 949172 490868 949228
rect 490924 949172 490934 949228
rect 106558 947732 106596 947788
rect 106652 947732 106662 947788
rect 216542 947732 216580 947788
rect 216636 947732 216646 947788
rect 271534 947732 271572 947788
rect 271628 947732 271638 947788
rect 470222 947732 470260 947788
rect 470316 947732 470326 947788
rect 525662 947732 525700 947788
rect 525756 947732 525766 947788
rect 690302 947732 690340 947788
rect 690396 947732 690406 947788
rect 251066 947604 251076 947660
rect 251132 947604 251188 947660
rect 251244 947604 251254 947660
rect 306030 947604 306068 947660
rect 306124 947604 306134 947660
rect 361050 947492 361060 947548
rect 361116 947492 361396 947548
rect 361452 947492 361462 947548
rect 545822 947492 545860 947548
rect 545916 947492 545926 947548
rect 581102 947492 581140 947548
rect 581196 947492 581206 947548
rect 655806 947492 655844 947548
rect 655900 947492 655910 947548
rect 697918 947492 697956 947548
rect 698012 947492 698022 947548
rect 525550 947284 525588 947340
rect 525644 947284 525654 947340
rect 690302 947284 690340 947340
rect 690396 947284 690406 947340
rect 361050 947156 361060 947212
rect 361116 947156 361284 947212
rect 361340 947156 361350 947212
rect 581214 947156 581252 947212
rect 581308 947156 581318 947212
rect 141306 947044 141316 947100
rect 141372 947044 141876 947100
rect 141932 947044 141942 947100
rect 545822 947044 545860 947100
rect 545916 947044 545926 947100
rect 655806 947044 655844 947100
rect 655900 947044 655910 947100
rect 471230 946836 471268 946892
rect 471324 946836 471334 946892
rect 545598 946836 545636 946892
rect 545692 946836 545702 946892
rect 655582 946836 655620 946892
rect 655676 946836 655686 946892
rect 691786 946820 691796 946876
rect 691852 946820 692916 946876
rect 692972 946820 692982 946876
rect 196046 946708 196084 946764
rect 196140 946708 196150 946764
rect 251038 946708 251076 946764
rect 251132 946708 251142 946764
rect 361050 946708 361060 946764
rect 361116 946708 361172 946764
rect 361228 946708 361238 946764
rect 526110 946708 526148 946764
rect 526204 946708 526214 946764
rect 580990 946708 581028 946764
rect 581084 946708 581094 946764
rect 106250 946596 106260 946652
rect 106316 946596 106326 946652
rect 196298 946596 196308 946652
rect 196364 946596 196374 946652
rect 72762 946036 72772 946092
rect 72828 946036 77476 946092
rect 77532 946036 77542 946092
rect 75450 945924 75460 945980
rect 75516 945924 77252 945980
rect 77308 945924 77318 945980
rect 106260 945868 106316 946596
rect 196308 946316 196364 946596
rect 525662 946388 525700 946444
rect 525756 946388 525766 946444
rect 545486 946388 545524 946444
rect 545580 946388 545590 946444
rect 655470 946388 655508 946444
rect 655564 946388 655574 946444
rect 196298 946260 196308 946316
rect 196364 946260 196374 946316
rect 581102 946260 581140 946316
rect 581196 946260 581206 946316
rect 471818 946036 471828 946092
rect 471884 946036 490868 946092
rect 490924 946036 490934 946092
rect 471258 945924 471268 945980
rect 471324 945924 490644 945980
rect 490700 945924 490710 945980
rect 73546 945812 73556 945868
rect 73612 945812 77364 945868
rect 77420 945812 77430 945868
rect 106250 945812 106260 945868
rect 106316 945812 106326 945868
rect 141082 945812 141092 945868
rect 141148 945812 141652 945868
rect 141708 945812 141718 945868
rect 471706 945812 471716 945868
rect 471772 945812 490532 945868
rect 490588 945812 490598 945868
rect 691114 945812 691124 945868
rect 691180 945812 704004 945868
rect 704060 945812 704070 945868
rect 72202 945700 72212 945756
rect 72268 945700 75460 945756
rect 75516 945700 75526 945756
rect 121764 943404 121820 944048
rect 122212 943404 122268 944048
rect 123108 943964 123164 944048
rect 123556 943964 123612 944048
rect 123108 943908 123612 943964
rect 124004 943404 124060 944048
rect 124452 943404 124508 944048
rect 120922 943348 120932 943404
rect 120988 943348 121820 943404
rect 121930 943348 121940 943404
rect 121996 943348 122268 943404
rect 122378 943348 122388 943404
rect 122444 943348 124060 943404
rect 124282 943348 124292 943404
rect 124348 943348 124508 943404
rect 124900 942844 124956 944048
rect 176764 943516 176820 944048
rect 176764 943460 177044 943516
rect 177100 943460 177110 943516
rect 177212 943404 177268 944048
rect 178108 943964 178164 944048
rect 178556 943964 178612 944048
rect 178108 943908 178612 943964
rect 179004 943516 179060 944048
rect 178154 943460 178164 943516
rect 178220 943460 179060 943516
rect 179452 943404 179508 944048
rect 179900 943404 179956 944048
rect 231764 943516 231820 944048
rect 230122 943460 230132 943516
rect 230188 943460 231820 943516
rect 232212 943404 232268 944048
rect 233108 943964 233164 944048
rect 233556 943964 233612 944048
rect 233108 943908 233612 943964
rect 234004 943516 234060 944048
rect 233482 943460 233492 943516
rect 233548 943460 234060 943516
rect 234452 943404 234508 944048
rect 176474 943348 176484 943404
rect 176540 943348 177268 943404
rect 178042 943348 178052 943404
rect 178108 943348 179508 943404
rect 179722 943348 179732 943404
rect 179788 943348 179956 943404
rect 231802 943348 231812 943404
rect 231868 943348 232268 943404
rect 233818 943348 233828 943404
rect 233884 943348 234508 943404
rect 234900 943292 234956 944048
rect 286764 943404 286820 944048
rect 285674 943348 285684 943404
rect 285740 943348 286820 943404
rect 287212 943292 287268 944048
rect 288108 943964 288164 944048
rect 288556 943964 288612 944048
rect 288108 943908 288612 943964
rect 289004 943404 289060 944048
rect 289452 943404 289508 944048
rect 289900 943404 289956 944048
rect 341764 943404 341820 944048
rect 289004 943348 289156 943404
rect 289212 943348 289222 943404
rect 289370 943348 289380 943404
rect 289436 943348 289508 943404
rect 289818 943348 289828 943404
rect 289884 943348 289956 943404
rect 341226 943348 341236 943404
rect 341292 943348 341820 943404
rect 342212 943292 342268 944048
rect 343108 943964 343164 944048
rect 343556 943964 343612 944048
rect 343108 943908 343612 943964
rect 344004 943404 344060 944048
rect 342682 943348 342692 943404
rect 342748 943348 344060 943404
rect 344452 943404 344508 944048
rect 344900 943516 344956 944048
rect 344586 943460 344596 943516
rect 344652 943460 344956 943516
rect 451764 943404 451820 944048
rect 452212 943404 452268 944048
rect 453108 943964 453164 944048
rect 453556 943964 453612 944048
rect 453108 943908 453612 943964
rect 454004 943516 454060 944048
rect 454004 943460 454244 943516
rect 454300 943460 454310 943516
rect 454452 943404 454508 944048
rect 344452 943348 344708 943404
rect 344764 943348 344774 943404
rect 450202 943348 450212 943404
rect 450268 943348 451820 943404
rect 451882 943348 451892 943404
rect 451948 943348 452268 943404
rect 453562 943348 453572 943404
rect 453628 943348 454508 943404
rect 454900 943404 454956 944048
rect 506764 943404 506820 944048
rect 454900 943348 455028 943404
rect 455084 943348 455094 943404
rect 505642 943348 505652 943404
rect 505708 943348 506820 943404
rect 507212 943292 507268 944048
rect 508108 943964 508164 944048
rect 508556 943964 508612 944048
rect 508108 943908 508612 943964
rect 509004 943516 509060 944048
rect 507434 943460 507444 943516
rect 507500 943460 509060 943516
rect 509452 943404 509508 944048
rect 509002 943348 509012 943404
rect 509068 943348 509508 943404
rect 509900 943404 509956 944048
rect 561764 943404 561820 944048
rect 509900 943348 510580 943404
rect 510636 943348 510646 943404
rect 561306 943348 561316 943404
rect 561372 943348 561820 943404
rect 562212 943292 562268 944048
rect 563108 943964 563164 944048
rect 563556 943964 563612 944048
rect 563108 943908 563612 943964
rect 564004 943404 564060 944048
rect 564004 943348 564228 943404
rect 564284 943348 564294 943404
rect 233482 943236 233492 943292
rect 233548 943236 234956 943292
rect 285898 943236 285908 943292
rect 285964 943236 287268 943292
rect 341114 943236 341124 943292
rect 341180 943236 342268 943292
rect 505866 943236 505876 943292
rect 505932 943236 507268 943292
rect 561082 943236 561092 943292
rect 561148 943236 562268 943292
rect 564452 943292 564508 944048
rect 564900 943404 564956 944048
rect 671764 943404 671820 944048
rect 564890 943348 564900 943404
rect 564956 943348 564966 943404
rect 670282 943348 670292 943404
rect 670348 943348 671820 943404
rect 672212 943404 672268 944048
rect 673108 943964 673164 944048
rect 673556 943964 673612 944048
rect 673108 943908 673612 943964
rect 674004 943404 674060 944048
rect 672212 943348 673428 943404
rect 673484 943348 673494 943404
rect 674004 943348 674100 943404
rect 674156 943348 674166 943404
rect 674452 943292 674508 944048
rect 564452 943236 565012 943292
rect 565068 943236 565078 943292
rect 673642 943236 673652 943292
rect 673708 943236 674508 943292
rect 674900 943180 674956 944048
rect 673866 943124 673876 943180
rect 673932 943124 674956 943180
rect 85194 942788 85204 942844
rect 85260 942788 124956 942844
rect 85418 942676 85428 942732
rect 85484 942676 121940 942732
rect 121996 942676 122006 942732
rect 85418 942564 85428 942620
rect 85484 942564 122388 942620
rect 122444 942564 122454 942620
rect 106586 942340 106596 942396
rect 106652 942340 196644 942396
rect 196700 942340 196710 942396
rect 216570 942340 216580 942396
rect 216636 942340 306068 942396
rect 306124 942340 306134 942396
rect 334282 942340 334292 942396
rect 334348 942340 361172 942396
rect 361228 942340 361238 942396
rect 160234 942228 160244 942284
rect 160300 942228 251188 942284
rect 251244 942228 251254 942284
rect 271562 942228 271572 942284
rect 271628 942228 361396 942284
rect 361452 942228 361462 942284
rect 160570 942116 160580 942172
rect 160636 942116 251076 942172
rect 251132 942116 251142 942172
rect 270554 942116 270564 942172
rect 270620 942116 334292 942172
rect 334348 942116 334358 942172
rect 335850 942116 335860 942172
rect 335916 942116 361284 942172
rect 361340 942116 361350 942172
rect 106250 942004 106260 942060
rect 106316 942004 196084 942060
rect 196140 942004 196150 942060
rect 215674 942004 215684 942060
rect 215740 942004 306404 942060
rect 306460 942004 306470 942060
rect 673418 939092 673428 939148
rect 673484 939092 674772 939148
rect 674828 939092 674838 939148
rect 163706 938532 163716 938588
rect 163772 938532 178164 938588
rect 178220 938532 178230 938588
rect 510570 938420 510580 938476
rect 510636 938420 519204 938476
rect 519260 938420 519270 938476
rect 455018 938196 455028 938252
rect 455084 938196 458500 938252
rect 458556 938196 458566 938252
rect 176698 937412 176708 937468
rect 176764 937412 179732 937468
rect 179788 937412 179798 937468
rect 230346 937412 230356 937468
rect 230412 937412 233492 937468
rect 233548 937412 233558 937468
rect 282398 937412 282436 937468
rect 282492 937412 282502 937468
rect 673642 937300 673652 937356
rect 673708 937300 687708 937356
rect 688174 937300 688212 937356
rect 688268 937300 688278 937356
rect 687652 937244 687708 937300
rect 561082 937188 561092 937244
rect 561148 937188 608132 937244
rect 608188 937188 608198 937244
rect 687390 937188 687428 937244
rect 687484 937188 687494 937244
rect 687652 937188 688996 937244
rect 689052 937188 689062 937244
rect 285646 937076 285684 937132
rect 285740 937076 285750 937132
rect 509002 937076 509012 937132
rect 509068 937076 687204 937132
rect 687260 937076 687270 937132
rect 141838 936964 141876 937020
rect 141932 936964 141942 937020
rect 178042 936964 178052 937020
rect 178108 936964 178724 937020
rect 178780 936964 178790 937020
rect 505866 936964 505876 937020
rect 505932 936964 541380 937020
rect 541436 936964 541446 937020
rect 688398 936964 688436 937020
rect 688492 936964 688502 937020
rect 451882 936852 451892 936908
rect 451948 936852 474740 936908
rect 474796 936852 474806 936908
rect 141614 936740 141652 936796
rect 141708 936740 141718 936796
rect 289370 936740 289380 936796
rect 289436 936740 688212 936796
rect 688268 936740 688278 936796
rect 141390 936628 141428 936684
rect 141484 936628 141494 936684
rect 230122 936628 230132 936684
rect 230188 936628 687876 936684
rect 687932 936628 687942 936684
rect 124282 936516 124292 936572
rect 124348 936516 666987 936572
rect 687950 936516 687988 936572
rect 688044 936516 688054 936572
rect 666931 936348 666987 936516
rect 688846 936404 688884 936460
rect 688940 936404 688950 936460
rect 666931 936292 689332 936348
rect 689388 936292 689398 936348
rect 341114 936068 341124 936124
rect 341180 936068 342580 936124
rect 342636 936068 342646 936124
rect 84046 935732 84084 935788
rect 84140 935732 84150 935788
rect 84270 935732 84308 935788
rect 84364 935732 84374 935788
rect 84494 935732 84532 935788
rect 84588 935732 84598 935788
rect 85418 935620 85428 935676
rect 85484 935620 96964 935676
rect 97020 935620 97030 935676
rect 585946 935620 585956 935676
rect 586012 935620 587524 935676
rect 587580 935620 587590 935676
rect 652698 935508 652708 935564
rect 652764 935508 673876 935564
rect 673932 935508 673942 935564
rect 695342 935508 695380 935564
rect 695436 935508 695446 935564
rect 85418 935396 85428 935452
rect 85484 935396 141316 935452
rect 141372 935396 141382 935452
rect 686970 935284 686980 935340
rect 687036 935284 694260 935340
rect 694316 935284 694326 935340
rect 233482 935172 233492 935228
rect 233548 935172 251972 935228
rect 252028 935172 252038 935228
rect 285898 935060 285908 935116
rect 285964 935060 341012 935116
rect 341068 935060 341078 935116
rect 686634 935060 686644 935116
rect 686700 935060 694036 935116
rect 694092 935060 694102 935116
rect 231802 934948 231812 935004
rect 231868 934948 274036 935004
rect 274092 934948 274102 935004
rect 686522 934948 686532 935004
rect 686588 934948 694932 935004
rect 694988 934948 694998 935004
rect 341002 934836 341012 934892
rect 341068 934836 362964 934892
rect 363020 934836 363030 934892
rect 430938 934836 430948 934892
rect 431004 934836 458500 934892
rect 458556 934836 458566 934892
rect 686298 934836 686308 934892
rect 686364 934836 694820 934892
rect 694876 934836 694886 934892
rect 686298 934724 686308 934780
rect 686364 934724 694708 934780
rect 694764 934724 694774 934780
rect 85194 934612 85204 934668
rect 85260 934612 118468 934668
rect 118524 934612 118534 934668
rect 686746 934612 686756 934668
rect 686812 934612 700532 934668
rect 700588 934612 700598 934668
rect 686186 934500 686196 934556
rect 686252 934500 693812 934556
rect 693868 934500 693878 934556
rect 686970 934388 686980 934444
rect 687036 934388 695156 934444
rect 695212 934388 695222 934444
rect 686746 934276 686756 934332
rect 686812 934276 694484 934332
rect 694540 934276 694550 934332
rect 686858 934164 686868 934220
rect 686924 934164 700532 934220
rect 700588 934164 700598 934220
rect 75936 929900 76132 929956
rect 76188 929900 76198 929956
rect 83738 929796 83748 929852
rect 83804 929796 83972 929852
rect 84028 929796 84038 929852
rect 75936 929452 76356 929508
rect 76412 929452 76422 929508
rect 75992 929004 76132 929060
rect 76188 929004 76198 929060
rect 75936 928556 76188 928612
rect 76132 928164 76188 928556
rect 75936 928108 76188 928164
rect 686858 928004 686868 928060
rect 686924 928004 686934 928060
rect 686868 927472 686924 928004
rect 78922 927332 78932 927388
rect 78988 927332 79716 927388
rect 79772 927332 79782 927388
rect 75936 927212 76244 927268
rect 76300 927212 76310 927268
rect 703994 927220 704004 927276
rect 704060 927220 705012 927276
rect 705068 927220 705078 927276
rect 703854 927108 703892 927164
rect 703948 927108 703958 927164
rect 84634 926884 84644 926940
rect 84700 926884 85120 926940
rect 75936 926764 76356 926820
rect 76412 926764 76422 926820
rect 704778 926324 704788 926380
rect 704892 926324 704902 926380
rect 705674 926324 705684 926380
rect 705788 926324 705798 926380
rect 697722 925092 697732 925148
rect 697788 925092 697956 925148
rect 698012 925092 698022 925148
rect 686746 914676 686756 914732
rect 686812 914676 686822 914732
rect 686756 914144 686812 914676
rect 83962 912660 83972 912716
rect 84028 912660 85120 912716
rect 701316 911180 702016 911236
rect 701316 911148 701372 911180
rect 690451 911092 701372 911148
rect 72986 910868 72996 910924
rect 73052 910868 84308 910924
rect 84364 910868 84374 910924
rect 73434 910756 73444 910812
rect 73500 910756 84532 910812
rect 84588 910756 84598 910812
rect 73546 910644 73556 910700
rect 73612 910644 84084 910700
rect 84140 910644 84150 910700
rect 690451 910588 690507 911092
rect 691338 910756 691348 910812
rect 691404 910788 701484 910812
rect 691404 910756 702016 910788
rect 701428 910732 702016 910756
rect 72202 910532 72212 910588
rect 72268 910532 84756 910588
rect 84812 910532 84822 910588
rect 689546 910532 689556 910588
rect 689612 910532 690507 910588
rect 701876 909836 702016 909892
rect 701876 909444 701932 909836
rect 701876 909388 702016 909444
rect 700522 908964 700532 909020
rect 700588 908996 701372 909020
rect 700588 908964 702016 908996
rect 701316 908940 702016 908964
rect 691226 908516 691236 908572
rect 691292 908548 701372 908572
rect 691292 908516 702016 908548
rect 701316 908492 702016 908516
rect 700522 908068 700532 908124
rect 700588 908100 701372 908124
rect 700588 908068 702016 908100
rect 701316 908044 702016 908068
rect 686896 900788 691348 900844
rect 691404 900788 691414 900844
rect 85092 897148 85148 898352
rect 76010 897092 76020 897148
rect 76076 897092 85148 897148
rect 699178 891492 699188 891548
rect 699244 891492 704836 891548
rect 704892 891492 704902 891548
rect 700186 891380 700196 891436
rect 700252 891380 705284 891436
rect 705340 891380 705350 891436
rect 699738 891268 699748 891324
rect 699804 891268 704388 891324
rect 704444 891268 704454 891324
rect 699402 890596 699412 890652
rect 699468 890596 705572 890652
rect 705628 890596 705638 890652
rect 686868 887068 686924 887376
rect 686868 887012 696276 887068
rect 696332 887012 696342 887068
rect 83962 883988 83972 884044
rect 84028 883988 85120 884044
rect 686868 873628 686924 874048
rect 686868 873572 694596 873628
rect 694652 873572 694662 873628
rect 84298 869764 84308 869820
rect 84364 869764 85120 869820
rect 686896 860692 693028 860748
rect 693084 860692 693094 860748
rect 84634 855428 84644 855484
rect 84700 855428 85120 855484
rect 686186 848148 686196 848204
rect 686252 848148 686262 848204
rect 686196 847504 686252 848148
rect 84074 841204 84084 841260
rect 84140 841204 85120 841260
rect 698730 840532 698740 840588
rect 698796 840532 704388 840588
rect 704444 840532 704454 840588
rect 704778 840308 704788 840364
rect 704892 840308 704902 840364
rect 705114 840308 705124 840364
rect 705180 840308 705284 840364
rect 705340 840308 705350 840364
rect 705674 840308 705684 840364
rect 705788 840308 705798 840364
rect 700074 838292 700084 838348
rect 700140 838292 700420 838348
rect 700476 838292 700486 838348
rect 700606 838292 700644 838348
rect 700700 838292 700710 838348
rect 686298 834820 686308 834876
rect 686364 834820 686374 834876
rect 686308 834176 686364 834820
rect 84410 826868 84420 826924
rect 84476 826868 85120 826924
rect 701316 825180 702016 825236
rect 701316 824908 701372 825180
rect 689658 824852 689668 824908
rect 689724 824852 701372 824908
rect 701418 824732 701428 824788
rect 701484 824732 702016 824788
rect 701876 823836 702016 823892
rect 701876 823444 701932 823836
rect 701876 823388 702016 823444
rect 699962 823060 699972 823116
rect 700028 823060 700644 823116
rect 700700 823060 700710 823116
rect 693802 822948 693812 823004
rect 693868 822996 701372 823004
rect 693868 822948 702016 822996
rect 701316 822940 702016 822948
rect 692906 822500 692916 822556
rect 692972 822548 701372 822556
rect 692972 822500 702016 822548
rect 701316 822492 702016 822500
rect 694810 822052 694820 822108
rect 694876 822100 701372 822108
rect 694876 822052 702016 822100
rect 701316 822044 702016 822052
rect 699850 821828 699860 821884
rect 699916 821828 701316 821884
rect 701372 821828 701382 821884
rect 686868 819980 686924 820736
rect 686868 819924 701428 819980
rect 701484 819924 701494 819980
rect 84746 812644 84756 812700
rect 84812 812644 85120 812700
rect 686634 807716 686644 807772
rect 686700 807716 686710 807772
rect 686644 807520 686700 807716
rect 693018 806932 693028 806988
rect 693084 806932 700532 806988
rect 700588 806932 700598 806988
rect 699738 806372 699748 806428
rect 699804 806372 702267 806428
rect 702211 806316 702267 806372
rect 702211 806260 703892 806316
rect 703948 806260 703958 806316
rect 699290 805476 699300 805532
rect 699356 805476 705284 805532
rect 705340 805476 705350 805532
rect 699514 805364 699524 805420
rect 699580 805364 704388 805420
rect 704444 805364 704454 805420
rect 701306 805252 701316 805308
rect 701372 805252 704836 805308
rect 704892 805252 704902 805308
rect 699738 804916 699748 804972
rect 699804 804916 705572 804972
rect 705628 804916 705638 804972
rect 84186 798308 84196 798364
rect 84252 798308 85120 798364
rect 686196 793548 686252 794080
rect 686186 793492 686196 793548
rect 686252 793492 686262 793548
rect 84522 783972 84532 784028
rect 84588 783972 85120 784028
rect 76346 783636 76356 783692
rect 76412 783636 83076 783692
rect 83132 783636 83142 783692
rect 73770 782068 73780 782124
rect 73836 782068 78372 782124
rect 78428 782068 78438 782124
rect 72650 781844 72660 781900
rect 72716 781844 78148 781900
rect 78204 781844 78214 781900
rect 72202 781732 72212 781788
rect 72268 781732 77700 781788
rect 77756 781732 77766 781788
rect 73098 781620 73108 781676
rect 73164 781620 77924 781676
rect 77980 781620 77990 781676
rect 686896 780724 693028 780780
rect 693084 780724 693094 780780
rect 84858 769748 84868 769804
rect 84924 769748 85120 769804
rect 686634 767732 686644 767788
rect 686700 767732 686710 767788
rect 686644 767536 686700 767732
rect 83738 766052 83748 766108
rect 83804 766052 84308 766108
rect 84364 766052 84374 766108
rect 75936 765900 76132 765956
rect 76188 765900 76198 765956
rect 75936 765452 76132 765508
rect 76188 765452 76198 765508
rect 75992 765004 76244 765060
rect 76300 765004 76310 765060
rect 75936 764556 76188 764612
rect 76132 764164 76188 764556
rect 84606 764484 84644 764540
rect 84700 764484 84710 764540
rect 75936 764108 76188 764164
rect 75936 763212 76244 763268
rect 76300 763212 76310 763268
rect 80462 763140 80500 763196
rect 80556 763140 80566 763196
rect 75936 762764 76132 762820
rect 76188 762764 76198 762820
rect 82282 762804 82292 762860
rect 82348 762804 83188 762860
rect 83244 762804 83254 762860
rect 83738 762804 83748 762860
rect 83804 762804 83972 762860
rect 84028 762804 84038 762860
rect 700186 755636 700196 755692
rect 700252 755636 704388 755692
rect 704444 755636 704454 755692
rect 84746 755412 84756 755468
rect 84812 755412 85120 755468
rect 703882 755076 703892 755132
rect 703948 755076 705124 755132
rect 705180 755076 705190 755132
rect 704778 754404 704788 754460
rect 704892 754404 704902 754460
rect 705674 754404 705684 754460
rect 705788 754404 705798 754460
rect 686868 754012 686924 754096
rect 686868 753956 686980 754012
rect 687036 753956 687046 754012
rect 699150 752500 699188 752556
rect 699244 752500 699254 752556
rect 699402 752500 699412 752556
rect 699468 752500 700420 752556
rect 700476 752500 700486 752556
rect 73546 747460 73556 747516
rect 73612 747460 77476 747516
rect 77532 747460 77542 747516
rect 72650 747348 72660 747404
rect 72716 747348 77364 747404
rect 77420 747348 77430 747404
rect 72202 747236 72212 747292
rect 72268 747236 77252 747292
rect 77308 747236 77318 747292
rect 73098 747124 73108 747180
rect 73164 747124 77588 747180
rect 77644 747124 77654 747180
rect 84298 741188 84308 741244
rect 84364 741188 85120 741244
rect 72762 741076 72772 741132
rect 72828 741076 77476 741132
rect 77532 741076 77542 741132
rect 75450 740964 75460 741020
rect 75516 740964 77812 741020
rect 77868 740964 77878 741020
rect 73546 740852 73556 740908
rect 73612 740852 77364 740908
rect 77420 740852 77430 740908
rect 72202 740740 72212 740796
rect 72268 740740 75460 740796
rect 75516 740740 75526 740796
rect 686420 740684 686476 740768
rect 73098 740628 73108 740684
rect 73164 740628 77252 740684
rect 77308 740628 77318 740684
rect 686410 740628 686420 740684
rect 686476 740628 686486 740684
rect 701316 739228 702016 739236
rect 689770 739172 689780 739228
rect 689836 739180 702016 739228
rect 689836 739172 701372 739180
rect 701316 738780 702016 738788
rect 700522 738724 700532 738780
rect 700588 738732 702016 738780
rect 700588 738724 701372 738732
rect 77242 738052 77252 738108
rect 77308 738052 78260 738108
rect 78316 738052 78326 738108
rect 701876 737836 702016 737892
rect 701876 737444 701932 737836
rect 701876 737388 702016 737444
rect 701316 736988 702016 736996
rect 696266 736932 696276 736988
rect 696332 736940 702016 736988
rect 696332 736932 701372 736940
rect 701316 736492 702016 736548
rect 701316 736428 701372 736492
rect 690451 736372 701372 736428
rect 690451 735868 690507 736372
rect 701428 736092 702016 736100
rect 694586 736036 694596 736092
rect 694652 736044 702016 736092
rect 694652 736036 701484 736044
rect 689546 735812 689556 735868
rect 689612 735812 690507 735868
rect 686868 728084 686980 728140
rect 687036 728084 687046 728140
rect 686868 727552 686924 728084
rect 84634 726852 84644 726908
rect 84700 726852 85120 726908
rect 84410 725060 84420 725116
rect 84476 725060 84644 725116
rect 84700 725060 84710 725116
rect 75936 724900 76132 724956
rect 76188 724900 76198 724956
rect 75936 724452 76524 724508
rect 76468 724444 76524 724452
rect 76468 724388 77140 724444
rect 77196 724388 77206 724444
rect 75992 724004 76468 724060
rect 76524 724004 76534 724060
rect 75936 723556 76188 723612
rect 76132 723164 76188 723556
rect 75936 723108 76188 723164
rect 84634 722596 84644 722652
rect 84700 722596 84756 722652
rect 84812 722596 84822 722652
rect 77242 722372 77252 722428
rect 77308 722372 78036 722428
rect 78092 722372 78102 722428
rect 75936 722212 76132 722268
rect 76188 722212 76198 722268
rect 75936 721764 76356 721820
rect 76412 721764 76422 721820
rect 83738 720692 83748 720748
rect 83804 720692 84084 720748
rect 84140 720692 84150 720748
rect 700074 720356 700084 720412
rect 700140 720356 704388 720412
rect 704444 720356 704454 720412
rect 699850 720244 699860 720300
rect 699916 720244 704836 720300
rect 704892 720244 704902 720300
rect 698730 720132 698740 720188
rect 698796 720132 705284 720188
rect 705340 720132 705350 720188
rect 693018 719796 693028 719852
rect 693084 719796 700644 719852
rect 700700 719796 700710 719852
rect 699962 719012 699972 719068
rect 700028 719012 705572 719068
rect 705628 719012 705638 719068
rect 686868 714028 686924 714112
rect 686858 713972 686868 714028
rect 686924 713972 686934 714028
rect 83962 712628 83972 712684
rect 84028 712628 85120 712684
rect 699514 712180 699524 712236
rect 699580 712180 705012 712236
rect 705068 712180 705078 712236
rect 699290 712068 699300 712124
rect 699356 712068 703892 712124
rect 703948 712068 703958 712124
rect 705674 711396 705684 711452
rect 705788 711396 705798 711452
rect 699738 710500 699748 710556
rect 699804 710500 700420 710556
rect 700476 710500 700486 710556
rect 73098 706580 73108 706636
rect 73164 706580 77924 706636
rect 77980 706580 77990 706636
rect 72202 706468 72212 706524
rect 72268 706468 77700 706524
rect 77756 706468 77766 706524
rect 73546 706356 73556 706412
rect 73612 706356 78148 706412
rect 78204 706356 78214 706412
rect 72650 706244 72660 706300
rect 72716 706244 78372 706300
rect 78428 706244 78438 706300
rect 686746 701428 686756 701484
rect 686812 701428 686822 701484
rect 76346 701316 76356 701372
rect 76412 701316 83300 701372
rect 83356 701316 83366 701372
rect 686756 700896 686812 701428
rect 72538 700084 72548 700140
rect 72604 700084 78372 700140
rect 78428 700084 78438 700140
rect 73098 699860 73108 699916
rect 73164 699860 77924 699916
rect 77980 699860 77990 699916
rect 72650 699748 72660 699804
rect 72716 699748 77700 699804
rect 77756 699748 77766 699804
rect 73546 699636 73556 699692
rect 73612 699636 77588 699692
rect 77644 699636 77654 699692
rect 84410 698292 84420 698348
rect 84476 698292 85120 698348
rect 700634 697060 700644 697116
rect 700700 697060 701540 697116
rect 701596 697060 701606 697116
rect 701316 696180 702016 696236
rect 701316 695548 701372 696180
rect 701530 695732 701540 695788
rect 701596 695732 702016 695788
rect 689882 695492 689892 695548
rect 689948 695492 701372 695548
rect 701876 694836 702016 694892
rect 701876 694444 701932 694836
rect 701876 694388 702016 694444
rect 701316 693980 702016 693996
rect 694586 693924 694596 693980
rect 694652 693940 702016 693980
rect 694652 693924 701372 693940
rect 701316 693532 702016 693548
rect 694586 693476 694596 693532
rect 694652 693492 702016 693532
rect 694652 693476 701372 693492
rect 701316 693084 702016 693100
rect 694810 693028 694820 693084
rect 694876 693044 702016 693084
rect 694876 693028 701372 693044
rect 686522 688100 686532 688156
rect 686588 688100 686598 688156
rect 686532 687568 686588 688100
rect 84522 684292 84532 684348
rect 84588 684292 84644 684348
rect 84700 684292 84710 684348
rect 75936 683900 76132 683956
rect 76188 683900 76198 683956
rect 85092 683788 85148 684096
rect 84970 683732 84980 683788
rect 85036 683732 85148 683788
rect 75936 683452 76132 683508
rect 76188 683452 76198 683508
rect 75992 683004 76468 683060
rect 76524 683004 76534 683060
rect 75936 682556 76188 682612
rect 76132 682164 76188 682556
rect 84830 682276 84868 682332
rect 84924 682276 84934 682332
rect 82282 682164 82292 682220
rect 82348 682164 83860 682220
rect 83916 682164 83926 682220
rect 75936 682108 76188 682164
rect 75936 681212 76132 681268
rect 76188 681212 76198 681268
rect 83738 681156 83748 681212
rect 83804 681156 84196 681212
rect 84252 681156 84262 681212
rect 75936 680764 76132 680820
rect 76188 680764 76198 680820
rect 702090 676564 702100 676620
rect 702156 676564 704836 676620
rect 704892 676564 704902 676620
rect 704378 676452 704388 676508
rect 704444 676452 705236 676508
rect 705292 676452 705302 676508
rect 704442 676340 704452 676396
rect 704508 676340 705284 676396
rect 705340 676340 705350 676396
rect 701754 675444 701764 675500
rect 701820 675444 705684 675500
rect 705740 675444 705750 675500
rect 686532 673708 686588 674128
rect 686522 673652 686532 673708
rect 686588 673652 686598 673708
rect 688314 672756 688324 672812
rect 688380 672756 688996 672812
rect 689052 672756 689062 672812
rect 686410 671076 686420 671132
rect 686476 671076 700532 671132
rect 700588 671076 700598 671132
rect 84074 669732 84084 669788
rect 84140 669732 85120 669788
rect 702090 669060 702100 669116
rect 702156 669060 704676 669116
rect 704732 669060 704742 669116
rect 704378 668500 704388 668556
rect 704444 668500 704452 668556
rect 704508 668500 704518 668556
rect 705226 668500 705236 668556
rect 705340 668500 705350 668556
rect 705674 668388 705684 668444
rect 705788 668388 705798 668444
rect 73546 665140 73556 665196
rect 73612 665140 77476 665196
rect 77532 665140 77542 665196
rect 72650 665028 72660 665084
rect 72716 665028 77252 665084
rect 77308 665028 77318 665084
rect 72538 664916 72548 664972
rect 72604 664916 77812 664972
rect 77868 664916 77878 664972
rect 73434 664804 73444 664860
rect 73500 664804 78260 664860
rect 78316 664804 78326 664860
rect 686298 661444 686308 661500
rect 686364 661444 686374 661500
rect 686308 660912 686364 661444
rect 72314 659092 72324 659148
rect 72380 659092 78260 659148
rect 78316 659092 78326 659148
rect 73098 658868 73108 658924
rect 73164 658868 78148 658924
rect 78204 658868 78214 658924
rect 73546 658756 73556 658812
rect 73612 658756 77476 658812
rect 77532 658756 77542 658812
rect 72650 658644 72660 658700
rect 72716 658644 77252 658700
rect 77308 658644 77318 658700
rect 84522 655508 84532 655564
rect 84588 655508 85120 655564
rect 701418 653180 701428 653236
rect 701484 653180 702016 653236
rect 701316 652764 702016 652788
rect 700522 652708 700532 652764
rect 700588 652732 702016 652764
rect 700588 652708 701372 652732
rect 689994 651812 690004 651868
rect 690060 651812 701428 651868
rect 701484 651812 701494 651868
rect 701876 651836 702016 651892
rect 701876 651444 701932 651836
rect 701876 651388 702016 651444
rect 701316 650972 702016 650996
rect 694026 650916 694036 650972
rect 694092 650940 702016 650972
rect 694092 650916 701372 650940
rect 701316 650524 702016 650548
rect 694698 650468 694708 650524
rect 694764 650492 702016 650524
rect 694764 650468 701372 650492
rect 701316 650076 702016 650100
rect 694250 650020 694260 650076
rect 694316 650044 702016 650076
rect 694316 650020 701372 650044
rect 686410 648116 686420 648172
rect 686476 648116 686486 648172
rect 686420 647584 686476 648116
rect 75936 642900 76132 642956
rect 76188 642900 76198 642956
rect 75936 642460 76524 642508
rect 75936 642452 77140 642460
rect 76468 642404 77140 642452
rect 77196 642404 77206 642460
rect 83738 642292 83748 642348
rect 83804 642292 84308 642348
rect 84364 642292 84374 642348
rect 84634 642068 84644 642124
rect 84700 642068 84756 642124
rect 84812 642068 84822 642124
rect 75992 642004 76468 642060
rect 76524 642004 76534 642060
rect 75936 641556 76188 641612
rect 76132 641164 76188 641556
rect 84634 641172 84644 641228
rect 84700 641172 85120 641228
rect 75936 641108 76188 641164
rect 75936 640212 76132 640268
rect 76188 640212 76198 640268
rect 77242 640052 77252 640108
rect 77308 640052 78820 640108
rect 78876 640052 78886 640108
rect 75936 639764 76356 639820
rect 76412 639764 76422 639820
rect 686308 633500 686364 634032
rect 704378 633556 704388 633612
rect 704444 633556 705236 633612
rect 705292 633556 705302 633612
rect 686298 633444 686308 633500
rect 686364 633444 686374 633500
rect 701866 633444 701876 633500
rect 701932 633444 704836 633500
rect 704892 633444 704902 633500
rect 704442 633332 704452 633388
rect 704508 633332 705284 633388
rect 705340 633332 705350 633388
rect 705674 633332 705684 633388
rect 705788 633332 705798 633388
rect 84186 626836 84196 626892
rect 84252 626836 85120 626892
rect 704378 626500 704388 626556
rect 704444 626500 704452 626556
rect 704508 626500 704518 626556
rect 705226 626276 705236 626332
rect 705340 626276 705350 626332
rect 705674 626276 705684 626332
rect 705788 626276 705798 626332
rect 704778 625380 704788 625436
rect 704892 625380 704902 625436
rect 72650 624596 72660 624652
rect 72716 624596 77588 624652
rect 77644 624596 77654 624652
rect 73546 624484 73556 624540
rect 73612 624484 77700 624540
rect 77756 624484 77766 624540
rect 73098 624372 73108 624428
rect 73164 624372 77924 624428
rect 77980 624372 77990 624428
rect 72202 624260 72212 624316
rect 72268 624260 78372 624316
rect 78428 624260 78438 624316
rect 686186 621348 686196 621404
rect 686252 621348 686262 621404
rect 686196 620816 686252 621348
rect 76346 618996 76356 619052
rect 76412 618996 84868 619052
rect 84924 618996 84934 619052
rect 72202 617652 72212 617708
rect 72268 617652 78596 617708
rect 78652 617652 78662 617708
rect 73546 617540 73556 617596
rect 73612 617540 77588 617596
rect 77644 617540 77654 617596
rect 84746 612612 84756 612668
rect 84812 612612 85120 612668
rect 701316 610180 702016 610236
rect 701316 609868 701372 610180
rect 689658 609812 689668 609868
rect 689724 609812 701372 609868
rect 701428 609756 702016 609788
rect 694474 609700 694484 609756
rect 694540 609732 702016 609756
rect 694540 609700 701484 609732
rect 701876 608836 702016 608892
rect 701876 608444 701932 608836
rect 701876 608388 702016 608444
rect 701316 607964 702016 607996
rect 695146 607908 695156 607964
rect 695212 607940 702016 607964
rect 695212 607908 701372 607940
rect 701316 607516 702016 607548
rect 694586 607460 694596 607516
rect 694652 607492 702016 607516
rect 694652 607460 701372 607492
rect 686532 606844 686588 607376
rect 701316 607044 702016 607100
rect 686522 606788 686532 606844
rect 686588 606788 686598 606844
rect 701316 606508 701372 607044
rect 686858 606452 686868 606508
rect 686924 606452 701372 606508
rect 76234 603092 76244 603148
rect 76300 603092 78148 603148
rect 78204 603092 78214 603148
rect 84410 601972 84420 602028
rect 84476 601972 84756 602028
rect 84812 601972 84822 602028
rect 75936 601900 76132 601956
rect 76188 601900 76198 601956
rect 75936 601452 76132 601508
rect 76188 601452 76198 601508
rect 75992 601004 76468 601060
rect 76524 601004 76534 601060
rect 80350 600628 80388 600684
rect 80444 600628 80454 600684
rect 75936 600556 76188 600612
rect 76132 600164 76188 600556
rect 75936 600108 76188 600164
rect 84942 599732 84980 599788
rect 85036 599732 85046 599788
rect 75936 599212 76132 599268
rect 76188 599212 76198 599268
rect 75936 598764 76356 598820
rect 76412 598764 76422 598820
rect 83738 598500 83748 598556
rect 83804 598500 83972 598556
rect 84028 598500 84038 598556
rect 85092 598108 85148 598304
rect 84970 598052 84980 598108
rect 85036 598052 85148 598108
rect 686644 593516 686700 594048
rect 686634 593460 686644 593516
rect 686700 593460 686710 593516
rect 701642 590436 701652 590492
rect 701708 590436 704836 590492
rect 704892 590436 704902 590492
rect 703994 590324 704004 590380
rect 704060 590324 705284 590380
rect 705340 590324 705350 590380
rect 704378 590212 704388 590268
rect 704444 590212 704452 590268
rect 704508 590212 704518 590268
rect 701866 589764 701876 589820
rect 701932 589764 705684 589820
rect 705740 589764 705750 589820
rect 83962 584052 83972 584108
rect 84028 584052 85120 584108
rect 701642 583268 701652 583324
rect 701708 583268 704836 583324
rect 704892 583268 704902 583324
rect 73434 582820 73444 582876
rect 73500 582820 76356 582876
rect 76412 582820 76422 582876
rect 703966 582820 704004 582876
rect 704060 582820 704070 582876
rect 704442 582820 704452 582876
rect 704508 582820 705284 582876
rect 705340 582820 705350 582876
rect 73770 582708 73780 582764
rect 73836 582708 77252 582764
rect 77308 582708 77318 582764
rect 72650 582596 72660 582652
rect 72716 582596 77476 582652
rect 77532 582596 77542 582652
rect 72202 582484 72212 582540
rect 72268 582484 78260 582540
rect 78316 582484 78326 582540
rect 705674 582372 705684 582428
rect 705788 582372 705798 582428
rect 686896 580692 688996 580748
rect 689052 580692 689062 580748
rect 76458 578676 76468 578732
rect 76524 578676 85204 578732
rect 85260 578676 85270 578732
rect 72202 576884 72212 576940
rect 72268 576884 78148 576940
rect 78204 576884 78214 576940
rect 73546 576772 73556 576828
rect 73612 576772 78484 576828
rect 78540 576772 78550 576828
rect 72650 576660 72660 576716
rect 72716 576660 77812 576716
rect 77868 576660 77878 576716
rect 73098 576548 73108 576604
rect 73164 576548 77924 576604
rect 77980 576548 77990 576604
rect 84298 569716 84308 569772
rect 84364 569716 85120 569772
rect 686868 566748 686924 567392
rect 701418 567180 701428 567236
rect 701484 567180 702016 567236
rect 694698 566804 694708 566860
rect 694764 566804 701484 566860
rect 701428 566788 701484 566804
rect 686868 566692 694932 566748
rect 694988 566692 694998 566748
rect 701428 566732 702016 566788
rect 690106 566132 690116 566188
rect 690172 566132 701428 566188
rect 701484 566132 701494 566188
rect 701876 565836 702016 565892
rect 701876 565444 701932 565836
rect 701876 565388 702016 565444
rect 694922 565012 694932 565068
rect 694988 565012 701372 565068
rect 701316 564996 701372 565012
rect 701316 564940 702016 564996
rect 701316 564508 702016 564548
rect 694698 564452 694708 564508
rect 694764 564492 702016 564508
rect 694764 564452 701372 564492
rect 701316 564044 702016 564100
rect 701316 562828 701372 564044
rect 686522 562772 686532 562828
rect 686588 562772 701372 562828
rect 76458 562660 76468 562716
rect 76524 562660 77700 562716
rect 77756 562660 77766 562716
rect 76794 562548 76804 562604
rect 76860 562548 78372 562604
rect 78428 562548 78438 562604
rect 76570 562436 76580 562492
rect 76636 562436 78596 562492
rect 78652 562436 78662 562492
rect 84522 561764 84532 561820
rect 84588 561764 84756 561820
rect 84812 561764 84822 561820
rect 75936 560900 76132 560956
rect 76188 560900 76198 560956
rect 75936 560476 76300 560508
rect 75936 560452 77140 560476
rect 76244 560420 77140 560452
rect 77196 560420 77206 560476
rect 75992 560004 76356 560060
rect 76412 560004 76422 560060
rect 75936 559556 76188 559612
rect 76132 559164 76188 559556
rect 84634 559412 84644 559468
rect 84700 559412 84756 559468
rect 84812 559412 84822 559468
rect 75936 559108 76188 559164
rect 75936 558212 76244 558268
rect 76300 558212 76310 558268
rect 83626 557844 83636 557900
rect 83692 557844 84084 557900
rect 84140 557844 84150 557900
rect 75936 557764 76132 557820
rect 76188 557764 76198 557820
rect 77242 557732 77252 557788
rect 77308 557732 78708 557788
rect 78764 557732 78774 557788
rect 83710 557732 83748 557788
rect 83804 557732 83814 557788
rect 84634 555492 84644 555548
rect 84700 555492 85120 555548
rect 686756 553532 686812 554064
rect 686746 553476 686756 553532
rect 686812 553476 686822 553532
rect 704974 547876 705012 547932
rect 705068 547876 705078 547932
rect 702090 547764 702100 547820
rect 702156 547764 704564 547820
rect 704620 547764 704630 547820
rect 704378 547652 704388 547708
rect 704444 547652 705124 547708
rect 705180 547652 705190 547708
rect 701866 543396 701876 543452
rect 701932 543396 705572 543452
rect 705628 543396 705638 543452
rect 73098 542500 73108 542556
rect 73164 542500 76356 542556
rect 76412 542500 76422 542556
rect 73546 542388 73556 542444
rect 73612 542388 76804 542444
rect 76860 542388 76870 542444
rect 72202 542276 72212 542332
rect 72268 542276 76580 542332
rect 76636 542276 76646 542332
rect 72650 542164 72660 542220
rect 72716 542164 77588 542220
rect 77644 542164 77654 542220
rect 84746 541156 84756 541212
rect 84812 541156 85120 541212
rect 686868 540204 686924 540736
rect 686858 540148 686868 540204
rect 686924 540148 686934 540204
rect 704554 540148 704564 540204
rect 704620 540148 705012 540204
rect 705068 540148 705078 540204
rect 702090 540036 702100 540092
rect 702156 540036 704676 540092
rect 704732 540036 704742 540092
rect 705086 540036 705124 540092
rect 705180 540036 705190 540092
rect 705674 539364 705684 539420
rect 705788 539364 705798 539420
rect 75348 536004 77252 536060
rect 77308 536004 77318 536060
rect 75348 535948 75404 536004
rect 73332 535892 75404 535948
rect 75460 535892 77364 535948
rect 77420 535892 77430 535948
rect 73332 535836 73388 535892
rect 75460 535836 75516 535892
rect 72202 535780 72212 535836
rect 72268 535780 73388 535836
rect 73546 535780 73556 535836
rect 73612 535780 75516 535836
rect 72650 535556 72660 535612
rect 72716 535556 77588 535612
rect 77644 535556 77654 535612
rect 84410 526932 84420 526988
rect 84476 526932 85120 526988
rect 686420 526876 686476 527408
rect 686410 526820 686420 526876
rect 686476 526820 686486 526876
rect 701316 524188 702016 524236
rect 690218 524132 690228 524188
rect 690284 524180 702016 524188
rect 690284 524132 701372 524180
rect 694810 523796 694820 523852
rect 694876 523796 701372 523852
rect 701316 523788 701372 523796
rect 701316 523732 702016 523788
rect 701876 522836 702016 522892
rect 701876 522444 701932 522836
rect 701876 522388 702016 522444
rect 695370 522004 695380 522060
rect 695436 522004 701372 522060
rect 701316 521996 701372 522004
rect 701316 521940 702016 521996
rect 701316 521500 702016 521548
rect 696266 521444 696276 521500
rect 696332 521492 702016 521500
rect 696332 521444 701372 521492
rect 686298 521108 686308 521164
rect 686364 521108 701372 521164
rect 701316 521100 701372 521108
rect 701316 521044 702016 521100
rect 75936 519900 76132 519956
rect 76188 519900 76198 519956
rect 75936 519452 76244 519508
rect 76300 519452 76310 519508
rect 84746 519092 84756 519148
rect 84812 519092 84868 519148
rect 84924 519092 84934 519148
rect 75992 519004 76468 519060
rect 76524 519004 76534 519060
rect 80238 518868 80276 518924
rect 80332 518868 80342 518924
rect 75936 518556 76188 518612
rect 76132 518164 76188 518556
rect 75936 518108 76188 518164
rect 84942 517860 84980 517916
rect 85036 517860 85046 517916
rect 75936 517212 76132 517268
rect 76188 517212 76198 517268
rect 75936 516764 76356 516820
rect 76412 516764 76422 516820
rect 83738 516404 83748 516460
rect 83804 516404 84196 516460
rect 84252 516404 84262 516460
rect 686868 513996 686924 514107
rect 686858 513940 686868 513996
rect 686924 513940 686934 513996
rect 84746 512596 84756 512652
rect 84812 512596 85120 512652
rect 704378 504532 704388 504588
rect 704444 504532 704452 504588
rect 704508 504532 704518 504588
rect 701642 504420 701652 504476
rect 701708 504420 704836 504476
rect 704892 504420 704902 504476
rect 703994 504308 704004 504364
rect 704060 504308 705284 504364
rect 705340 504308 705350 504364
rect 701866 504084 701876 504140
rect 701932 504084 705572 504140
rect 705628 504084 705638 504140
rect 73098 501620 73108 501676
rect 73164 501620 77924 501676
rect 77980 501620 77990 501676
rect 73546 501508 73556 501564
rect 73612 501508 77812 501564
rect 77868 501508 77878 501564
rect 72650 501396 72660 501452
rect 72716 501396 78484 501452
rect 78540 501396 78550 501452
rect 72202 501284 72212 501340
rect 72268 501284 78148 501340
rect 78204 501284 78214 501340
rect 686896 500724 693140 500780
rect 693196 500724 693206 500780
rect 84074 498372 84084 498428
rect 84140 498372 85120 498428
rect 686522 488180 686532 488236
rect 686588 488180 686598 488236
rect 686532 488012 686588 488180
rect 686532 487956 700532 488012
rect 700588 487956 700598 488012
rect 686308 487228 686364 487424
rect 686298 487172 686308 487228
rect 686364 487172 686374 487228
rect 84522 484036 84532 484092
rect 84588 484036 85120 484092
rect 686756 473788 686812 474096
rect 686746 473732 686756 473788
rect 686812 473732 686822 473788
rect 85092 469196 85148 469728
rect 84970 469140 84980 469196
rect 85036 469140 85148 469196
rect 686896 460740 693252 460796
rect 693308 460740 693318 460796
rect 84186 455476 84196 455532
rect 84252 455476 85120 455532
rect 686420 446908 686476 447440
rect 686410 446852 686420 446908
rect 686476 446852 686486 446908
rect 85092 440524 85148 441168
rect 85082 440468 85092 440524
rect 85148 440468 85158 440524
rect 686644 433468 686700 434112
rect 686634 433412 686644 433468
rect 686700 433412 686710 433468
rect 85092 426748 85148 426944
rect 85082 426692 85092 426748
rect 85148 426692 85158 426748
rect 686896 420756 693028 420812
rect 693084 420756 693094 420812
rect 76346 415716 76356 415772
rect 76412 415716 83412 415772
rect 83468 415716 83478 415772
rect 72202 412692 72212 412748
rect 72268 412692 78596 412748
rect 78652 412692 78662 412748
rect 73546 412580 73556 412636
rect 73612 412580 77700 412636
rect 77756 412580 77766 412636
rect 85092 412076 85148 412608
rect 84970 412020 84980 412076
rect 85036 412020 85148 412076
rect 686196 406812 686252 407456
rect 686186 406756 686196 406812
rect 686252 406756 686262 406812
rect 76570 399700 76580 399756
rect 76636 399700 77476 399756
rect 77532 399700 77542 399756
rect 76346 399588 76356 399644
rect 76412 399588 77588 399644
rect 77644 399588 77654 399644
rect 85204 398188 85260 398384
rect 85194 398132 85204 398188
rect 85260 398132 85270 398188
rect 75936 396900 76132 396956
rect 76188 396900 76198 396956
rect 83738 396900 83748 396956
rect 83804 396900 84308 396956
rect 84364 396900 84374 396956
rect 75936 396452 76132 396508
rect 76188 396452 76198 396508
rect 78922 396116 78932 396172
rect 78988 396116 80052 396172
rect 80108 396116 80118 396172
rect 75992 396004 77140 396060
rect 77196 396004 77206 396060
rect 75936 395556 76188 395612
rect 76132 395164 76188 395556
rect 75936 395108 76188 395164
rect 84634 394996 84644 395052
rect 84700 394996 84868 395052
rect 84924 394996 84934 395052
rect 75936 394212 76132 394268
rect 76188 394212 76198 394268
rect 686896 394100 689108 394156
rect 689164 394100 689174 394156
rect 75936 393764 76244 393820
rect 76300 393764 76310 393820
rect 83738 393652 83748 393708
rect 83804 393652 83972 393708
rect 84028 393652 84038 393708
rect 83598 393428 83636 393484
rect 83692 393428 83702 393484
rect 76122 387940 76132 387996
rect 76188 387940 77364 387996
rect 77420 387940 77430 387996
rect 84634 384020 84644 384076
rect 84700 384020 85120 384076
rect 686868 380156 686924 380800
rect 686868 380100 694820 380156
rect 694876 380100 694886 380156
rect 73770 377860 73780 377916
rect 73836 377860 76356 377916
rect 76412 377860 76422 377916
rect 72986 377748 72996 377804
rect 73052 377748 76132 377804
rect 76188 377748 76198 377804
rect 73098 377636 73108 377692
rect 73164 377636 76580 377692
rect 76636 377636 76646 377692
rect 72202 377524 72212 377580
rect 72268 377524 77252 377580
rect 77308 377524 77318 377580
rect 72202 371924 72212 371980
rect 72268 371924 77924 371980
rect 77980 371924 77990 371980
rect 73546 371812 73556 371868
rect 73612 371812 78148 371868
rect 78204 371812 78214 371868
rect 72650 371700 72660 371756
rect 72716 371700 77812 371756
rect 77868 371700 77878 371756
rect 73098 371588 73108 371644
rect 73164 371588 77588 371644
rect 77644 371588 77654 371644
rect 84858 369796 84868 369852
rect 84924 369796 85120 369852
rect 701642 368116 701652 368172
rect 701708 368116 704564 368172
rect 704620 368116 704630 368172
rect 703966 367780 704004 367836
rect 704060 367780 704070 367836
rect 704442 367780 704452 367836
rect 704508 367780 705284 367836
rect 705340 367780 705350 367836
rect 686308 366940 686364 367472
rect 705674 367332 705684 367388
rect 705788 367332 705798 367388
rect 686298 366884 686308 366940
rect 686364 366884 686374 366940
rect 84746 357140 84756 357196
rect 84812 357140 85428 357196
rect 85484 357140 85494 357196
rect 84410 356916 84420 356972
rect 84476 356916 84756 356972
rect 84812 356916 84822 356972
rect 76234 356356 76244 356412
rect 76300 356356 78260 356412
rect 78316 356356 78326 356412
rect 76794 356244 76804 356300
rect 76860 356244 78596 356300
rect 78652 356244 78662 356300
rect 76570 356132 76580 356188
rect 76636 356132 78372 356188
rect 78428 356132 78438 356188
rect 75936 355900 76132 355956
rect 76188 355900 76198 355956
rect 75936 355452 76132 355508
rect 76188 355452 76198 355508
rect 75992 355004 76468 355060
rect 76524 355004 76534 355060
rect 84718 355012 84756 355068
rect 84812 355012 84822 355068
rect 85316 354844 85372 355488
rect 85306 354788 85316 354844
rect 85372 354788 85382 354844
rect 75936 354556 76188 354612
rect 76132 354164 76188 354556
rect 75936 354108 76188 354164
rect 80126 354116 80164 354172
rect 80220 354116 80230 354172
rect 686532 353612 686588 354144
rect 686522 353556 686532 353612
rect 686588 353556 686598 353612
rect 75936 353212 76132 353268
rect 76188 353212 76198 353268
rect 75936 352764 76356 352820
rect 76412 352764 76422 352820
rect 694922 352212 694932 352268
rect 694988 352236 701372 352268
rect 694988 352212 702016 352236
rect 701316 352180 702016 352212
rect 695146 351764 695156 351820
rect 695212 351788 701372 351820
rect 695212 351764 702016 351788
rect 701316 351732 702016 351764
rect 701876 350836 702016 350892
rect 701876 350444 701932 350836
rect 701876 350388 702016 350444
rect 700522 349972 700532 350028
rect 700588 349996 701372 350028
rect 700588 349972 702016 349996
rect 701316 349940 702016 349972
rect 695034 349524 695044 349580
rect 695100 349548 701372 349580
rect 695100 349524 702016 349548
rect 701316 349492 702016 349524
rect 695370 349076 695380 349132
rect 695436 349100 701372 349132
rect 695436 349076 702016 349100
rect 701316 349044 702016 349076
rect 84298 341236 84308 341292
rect 84364 341236 85120 341292
rect 686532 340284 686588 340816
rect 686522 340228 686532 340284
rect 686588 340228 686598 340284
rect 73098 337540 73108 337596
rect 73164 337540 76580 337596
rect 76636 337540 76646 337596
rect 73546 337428 73556 337484
rect 73612 337428 76356 337484
rect 76412 337428 76422 337484
rect 72202 337316 72212 337372
rect 72268 337316 76804 337372
rect 76860 337316 76870 337372
rect 72650 337204 72660 337260
rect 72716 337204 77700 337260
rect 77756 337204 77766 337260
rect 686970 335972 686980 336028
rect 687036 335972 689108 336028
rect 689164 335972 689174 336028
rect 688986 334180 688996 334236
rect 689052 334180 695156 334236
rect 695212 334180 695222 334236
rect 686186 334068 686196 334124
rect 686252 334068 694820 334124
rect 694876 334068 694886 334124
rect 686634 333956 686644 334012
rect 686700 333956 695380 334012
rect 695436 333956 695446 334012
rect 222842 333732 222852 333788
rect 222908 333732 258916 333788
rect 258972 333732 258982 333788
rect 271002 333732 271012 333788
rect 271068 333732 388052 333788
rect 388108 333732 388118 333788
rect 393082 333732 393092 333788
rect 393148 333732 656740 333788
rect 656796 333732 656806 333788
rect 119130 333620 119140 333676
rect 119196 333620 171108 333676
rect 171164 333620 171174 333676
rect 209626 333620 209636 333676
rect 209692 333620 223412 333676
rect 223468 333620 223478 333676
rect 278282 333620 278292 333676
rect 278348 333620 406420 333676
rect 406476 333620 406486 333676
rect 160682 333508 160692 333564
rect 160748 333508 187124 333564
rect 187180 333508 187190 333564
rect 210634 333508 210644 333564
rect 210700 333508 221620 333564
rect 221676 333508 221686 333564
rect 320170 333508 320180 333564
rect 320236 333508 364532 333564
rect 364588 333508 364598 333564
rect 386026 333508 386036 333564
rect 386092 333508 460068 333564
rect 460124 333508 460134 333564
rect 127194 333396 127204 333452
rect 127260 333396 173460 333452
rect 173516 333396 173526 333452
rect 174570 333396 174580 333452
rect 174636 333396 191492 333452
rect 191548 333396 191558 333452
rect 216346 333396 216356 333452
rect 216412 333396 240996 333452
rect 241052 333396 241062 333452
rect 319946 333396 319956 333452
rect 320012 333396 370244 333452
rect 370300 333396 370310 333452
rect 370458 333396 370468 333452
rect 370524 333396 489412 333452
rect 489468 333396 489478 333452
rect 490531 333396 502347 333452
rect 490531 333340 490587 333396
rect 502291 333340 502347 333396
rect 525811 333396 549387 333452
rect 610922 333396 610932 333452
rect 610988 333396 688212 333452
rect 688268 333396 688278 333452
rect 525811 333340 525867 333396
rect 549331 333340 549387 333396
rect 162810 333284 162820 333340
rect 162876 333284 188636 333340
rect 217018 333284 217028 333340
rect 217084 333284 239092 333340
rect 239148 333284 239158 333340
rect 240538 333284 240548 333340
rect 240604 333284 304612 333340
rect 304668 333284 304678 333340
rect 353546 333284 353556 333340
rect 353612 333284 477540 333340
rect 477596 333284 477606 333340
rect 487946 333284 487956 333340
rect 488012 333284 490587 333340
rect 497326 333284 497364 333340
rect 497420 333284 497430 333340
rect 502291 333284 525867 333340
rect 533054 333284 533092 333340
rect 533148 333284 533158 333340
rect 549331 333284 626612 333340
rect 626668 333284 626678 333340
rect 188580 333228 188636 333284
rect 149034 333172 149044 333228
rect 149100 333172 173012 333228
rect 173068 333172 173078 333228
rect 173236 333172 181300 333228
rect 181356 333172 181366 333228
rect 184426 333172 184436 333228
rect 184492 333172 188356 333228
rect 188412 333172 188422 333228
rect 188570 333172 188580 333228
rect 188636 333172 188646 333228
rect 207498 333172 207508 333228
rect 207564 333172 217140 333228
rect 217196 333172 217206 333228
rect 218474 333172 218484 333228
rect 218540 333172 247044 333228
rect 247100 333172 247110 333228
rect 273130 333172 273140 333228
rect 273196 333172 393988 333228
rect 394044 333172 394054 333228
rect 421530 333172 421540 333228
rect 421596 333172 453684 333228
rect 453740 333172 453750 333228
rect 454906 333172 454916 333228
rect 454972 333172 603092 333228
rect 603148 333172 603158 333228
rect 173236 333116 173292 333172
rect 106698 333060 106708 333116
rect 106764 333060 135156 333116
rect 135212 333060 135222 333116
rect 146458 333060 146468 333116
rect 146524 333060 173292 333116
rect 173450 333060 173460 333116
rect 173516 333060 174020 333116
rect 174076 333060 174086 333116
rect 182186 333060 182196 333116
rect 182252 333060 194404 333116
rect 194460 333060 194470 333116
rect 211194 333060 211204 333116
rect 211260 333060 216132 333116
rect 216188 333060 216198 333116
rect 220154 333060 220164 333116
rect 220220 333060 253652 333116
rect 253708 333060 253718 333116
rect 290714 333060 290724 333116
rect 290780 333060 442372 333116
rect 442428 333060 442438 333116
rect 454682 333060 454692 333116
rect 454748 333060 609364 333116
rect 609420 333060 609430 333116
rect 701530 333060 701540 333116
rect 701596 333060 704836 333116
rect 704892 333060 704902 333116
rect 100650 332948 100660 333004
rect 100716 332948 133476 333004
rect 133532 332948 133542 333004
rect 140522 332948 140532 333004
rect 140588 332948 177212 333004
rect 178266 332948 178276 333004
rect 178332 332948 193732 333004
rect 193788 332948 193798 333004
rect 211754 332948 211764 333004
rect 211820 332948 227780 333004
rect 227836 332948 227846 333004
rect 286234 332948 286244 333004
rect 286300 332948 430500 333004
rect 430556 332948 430566 333004
rect 437658 332948 437668 333004
rect 437724 332948 591444 333004
rect 591500 332948 591510 333004
rect 177156 332892 177212 332948
rect 88778 332836 88788 332892
rect 88844 332836 133924 332892
rect 133980 332836 133990 332892
rect 134474 332836 134484 332892
rect 134540 332836 176932 332892
rect 176988 332836 176998 332892
rect 177156 332836 179172 332892
rect 179228 332836 179238 332892
rect 179396 332836 182756 332892
rect 182812 332836 182822 332892
rect 188346 332836 188356 332892
rect 188412 332836 194852 332892
rect 194908 332836 194918 332892
rect 203354 332836 203364 332892
rect 203420 332836 207956 332892
rect 208012 332836 208022 332892
rect 208954 332836 208964 332892
rect 209020 332836 219828 332892
rect 219884 332836 219894 332892
rect 225194 332836 225204 332892
rect 225260 332836 226044 332892
rect 229450 332836 229460 332892
rect 229516 332836 277508 332892
rect 277564 332836 277574 332892
rect 280634 332836 280644 332892
rect 280700 332836 418516 332892
rect 418572 332836 418582 332892
rect 421082 332836 421092 332892
rect 421148 332836 579460 332892
rect 579516 332836 579526 332892
rect 703994 332836 704004 332892
rect 704060 332836 705012 332892
rect 705068 332836 705078 332892
rect 179396 332780 179452 332836
rect 225988 332780 226044 332836
rect 98746 332724 98756 332780
rect 98812 332724 133700 332780
rect 133756 332724 133766 332780
rect 173002 332724 173012 332780
rect 173068 332724 179452 332780
rect 180170 332724 180180 332780
rect 180236 332724 195188 332780
rect 195244 332724 195254 332780
rect 196531 332724 198324 332780
rect 198380 332724 198390 332780
rect 205258 332724 205268 332780
rect 205324 332724 208124 332780
rect 208282 332724 208292 332780
rect 208348 332724 215908 332780
rect 215964 332724 215974 332780
rect 216122 332724 216132 332780
rect 216188 332724 225764 332780
rect 225820 332724 225830 332780
rect 225988 332724 265524 332780
rect 265580 332724 265590 332780
rect 277386 332724 277396 332780
rect 277452 332724 278292 332780
rect 278348 332724 278358 332780
rect 367882 332724 367892 332780
rect 367948 332724 567588 332780
rect 567644 332724 567654 332780
rect 701754 332724 701764 332780
rect 701820 332724 705572 332780
rect 705628 332724 705638 332780
rect 196531 332668 196587 332724
rect 208068 332668 208124 332724
rect 92810 332612 92820 332668
rect 92876 332612 118356 332668
rect 118412 332612 118422 332668
rect 176250 332612 176260 332668
rect 176316 332612 192276 332668
rect 192332 332612 192342 332668
rect 194170 332612 194180 332668
rect 194236 332612 196587 332668
rect 198090 332612 198100 332668
rect 198156 332612 201572 332668
rect 201628 332612 201638 332668
rect 208068 332612 209860 332668
rect 209916 332612 209926 332668
rect 210074 332612 210084 332668
rect 210140 332612 210644 332668
rect 210700 332612 210710 332668
rect 213322 332612 213332 332668
rect 213388 332612 231812 332668
rect 231868 332612 231878 332668
rect 233594 332612 233604 332668
rect 233660 332612 287364 332668
rect 287420 332612 287430 332668
rect 320394 332612 320404 332668
rect 320460 332612 358932 332668
rect 358988 332612 358998 332668
rect 418282 332612 418292 332668
rect 418348 332612 420532 332668
rect 420588 332612 420598 332668
rect 453674 332612 453684 332668
rect 453740 332612 454804 332668
rect 454860 332612 454870 332668
rect 551646 332612 551684 332668
rect 551740 332612 551750 332668
rect 623214 332612 623252 332668
rect 623308 332612 623318 332668
rect 673194 332612 673204 332668
rect 673260 332612 678916 332668
rect 678972 332612 678982 332668
rect 704378 332612 704388 332668
rect 704444 332612 704900 332668
rect 704956 332612 704966 332668
rect 324874 332500 324884 332556
rect 324940 332500 535780 332556
rect 535836 332500 535846 332556
rect 672270 332500 672308 332556
rect 672364 332500 672374 332556
rect 329242 332388 329252 332444
rect 329308 332388 547764 332444
rect 547820 332388 547830 332444
rect 359482 332276 359492 332332
rect 359548 332276 593460 332332
rect 593516 332276 593526 332332
rect 341786 332164 341796 332220
rect 341852 332164 575540 332220
rect 575596 332164 575606 332220
rect 144330 332052 144340 332108
rect 144396 332052 181636 332108
rect 181692 332052 181702 332108
rect 347722 332052 347732 332108
rect 347788 332052 362964 332108
rect 363020 332052 363030 332108
rect 366426 332052 366436 332108
rect 366492 332052 649012 332108
rect 649068 332052 649078 332108
rect 671290 332052 671300 332108
rect 671356 332052 687988 332108
rect 688044 332052 688054 332108
rect 76458 331940 76468 331996
rect 76524 331940 378756 331996
rect 378812 331940 378822 331996
rect 387146 331940 387156 331996
rect 387212 331940 658980 331996
rect 659036 331940 659046 331996
rect 671066 331940 671076 331996
rect 671132 331940 687876 331996
rect 687932 331940 687942 331996
rect 80490 331828 80500 331884
rect 80556 331828 672196 331884
rect 672252 331828 672262 331884
rect 80266 331716 80276 331772
rect 80332 331716 672084 331772
rect 672140 331716 672150 331772
rect 318266 331604 318276 331660
rect 318332 331604 517860 331660
rect 517916 331604 517926 331660
rect 267978 331492 267988 331548
rect 268044 331492 380772 331548
rect 380828 331492 380838 331548
rect 380986 331492 380996 331548
rect 381052 331492 565572 331548
rect 565628 331492 565638 331548
rect 274586 331380 274596 331436
rect 274652 331380 398692 331436
rect 398748 331380 398758 331436
rect 399690 331380 399700 331436
rect 399756 331380 434420 331436
rect 434476 331380 434486 331436
rect 272234 331268 272244 331324
rect 272300 331268 392756 331324
rect 392812 331268 392822 331324
rect 421754 331268 421764 331324
rect 421820 331268 440468 331324
rect 440524 331268 440534 331324
rect 270218 331156 270228 331212
rect 270284 331156 386820 331212
rect 386876 331156 386886 331212
rect 73882 331044 73892 331100
rect 73948 331044 78372 331100
rect 78428 331044 78438 331100
rect 367882 331044 367892 331100
rect 367948 331044 374836 331100
rect 374892 331044 374902 331100
rect 379642 331044 379652 331100
rect 379708 331044 428484 331100
rect 428540 331044 428550 331100
rect 75460 330932 77364 330988
rect 77420 330932 77430 330988
rect 75460 330876 75516 330932
rect 72202 330820 72212 330876
rect 72268 330820 75516 330876
rect 303034 330820 303044 330876
rect 303100 330820 476196 330876
rect 476252 330820 476262 330876
rect 216682 330708 216692 330764
rect 216748 330708 243684 330764
rect 243740 330708 243750 330764
rect 307514 330708 307524 330764
rect 307580 330708 488068 330764
rect 488124 330708 488134 330764
rect 72650 330596 72660 330652
rect 72716 330596 77476 330652
rect 77532 330596 77542 330652
rect 235274 330596 235284 330652
rect 235340 330596 291396 330652
rect 291452 330596 291462 330652
rect 311770 330596 311780 330652
rect 311836 330596 500052 330652
rect 500108 330596 500118 330652
rect 237402 330484 237412 330540
rect 237468 330484 297332 330540
rect 297388 330484 297398 330540
rect 316138 330484 316148 330540
rect 316204 330484 511924 330540
rect 511980 330484 511990 330540
rect 238522 330372 238532 330428
rect 238588 330372 301364 330428
rect 301420 330372 301430 330428
rect 353770 330372 353780 330428
rect 353836 330372 559636 330428
rect 559692 330372 559702 330428
rect 239642 330260 239652 330316
rect 239708 330260 303268 330316
rect 303324 330260 303334 330316
rect 336746 330260 336756 330316
rect 336812 330260 347060 330316
rect 347116 330260 347126 330316
rect 354106 330260 354116 330316
rect 354172 330260 581476 330316
rect 581532 330260 581542 330316
rect 245466 330148 245476 330204
rect 245532 330148 319172 330204
rect 319228 330148 319238 330204
rect 335962 330148 335972 330204
rect 336028 330148 356916 330204
rect 356972 330148 356982 330204
rect 359146 330148 359156 330204
rect 359212 330148 629188 330204
rect 629244 330148 629254 330204
rect 108714 330036 108724 330092
rect 108780 330036 168084 330092
rect 168140 330036 168150 330092
rect 215114 330036 215124 330092
rect 215180 330036 237748 330092
rect 237804 330036 237814 330092
rect 257114 330036 257124 330092
rect 257180 330036 350980 330092
rect 351036 330036 351046 330092
rect 359818 330036 359828 330092
rect 359884 330036 631204 330092
rect 631260 330036 631270 330092
rect 300794 329924 300804 329980
rect 300860 329924 470260 329980
rect 470316 329924 470326 329980
rect 296426 329812 296436 329868
rect 296492 329812 458276 329868
rect 458332 329812 458342 329868
rect 287242 329700 287252 329756
rect 287308 329700 399700 329756
rect 399756 329700 399766 329756
rect 285562 329588 285572 329644
rect 285628 329588 379652 329644
rect 379708 329588 379718 329644
rect 381434 329588 381444 329644
rect 381500 329588 411348 329644
rect 411404 329588 411414 329644
rect 346042 329476 346052 329532
rect 346108 329476 368900 329532
rect 368956 329476 368966 329532
rect 373594 329476 373604 329532
rect 373660 329476 380996 329532
rect 381052 329476 381062 329532
rect 346154 329364 346164 329420
rect 346220 329364 359492 329420
rect 359548 329364 359558 329420
rect 385466 329252 385476 329308
rect 385532 329252 387156 329308
rect 387212 329252 387222 329308
rect 156314 329140 156324 329196
rect 156380 329140 186452 329196
rect 186508 329140 186518 329196
rect 246250 329140 246260 329196
rect 246316 329140 321188 329196
rect 321244 329140 321254 329196
rect 342458 329140 342468 329196
rect 342524 329140 583492 329196
rect 583548 329140 583558 329196
rect 656730 329140 656740 329196
rect 656796 329140 666932 329196
rect 666988 329140 666998 329196
rect 150378 329028 150388 329084
rect 150444 329028 184212 329084
rect 184268 329028 184278 329084
rect 249946 329028 249956 329084
rect 250012 329028 331156 329084
rect 331212 329028 331222 329084
rect 344698 329028 344708 329084
rect 344764 329028 589428 329084
rect 589484 329028 589494 329084
rect 142426 328916 142436 328972
rect 142492 328916 180628 328972
rect 180684 328916 180694 328972
rect 214218 328916 214228 328972
rect 214284 328916 235732 328972
rect 235788 328916 235798 328972
rect 252074 328916 252084 328972
rect 252140 328916 337092 328972
rect 337148 328916 337158 328972
rect 349066 328916 349076 328972
rect 349132 328916 601412 328972
rect 601468 328916 601478 328972
rect 136490 328804 136500 328860
rect 136556 328804 178388 328860
rect 178444 328804 178454 328860
rect 225866 328804 225876 328860
rect 225932 328804 263620 328860
rect 263676 328804 263686 328860
rect 269546 328804 269556 328860
rect 269612 328804 384804 328860
rect 384860 328804 384870 328860
rect 388266 328804 388276 328860
rect 388332 328804 403396 328860
rect 403452 328804 403462 328860
rect 405738 328804 405748 328860
rect 405804 328804 660996 328860
rect 661052 328804 661062 328860
rect 130554 328692 130564 328748
rect 130620 328692 176260 328748
rect 176316 328692 176326 328748
rect 219370 328692 219380 328748
rect 219436 328692 245700 328748
rect 245756 328692 245766 328748
rect 254314 328692 254324 328748
rect 254380 328692 343028 328748
rect 343084 328692 343094 328748
rect 353434 328692 353444 328748
rect 353500 328692 613284 328748
rect 613340 328692 613350 328748
rect 116666 328580 116676 328636
rect 116732 328580 171892 328636
rect 171948 328580 171958 328636
rect 219930 328580 219940 328636
rect 219996 328580 249620 328636
rect 249676 328580 249686 328636
rect 254986 328580 254996 328636
rect 255052 328580 345044 328636
rect 345100 328580 345110 328636
rect 345258 328580 345268 328636
rect 345324 328580 352996 328636
rect 353052 328580 353062 328636
rect 365642 328580 365652 328636
rect 365708 328580 635124 328636
rect 635180 328580 635190 328636
rect 170314 328468 170324 328524
rect 170380 328468 190036 328524
rect 190092 328468 190102 328524
rect 222282 328468 222292 328524
rect 222348 328468 255668 328524
rect 255724 328468 255734 328524
rect 258570 328468 258580 328524
rect 258636 328468 355012 328524
rect 355068 328468 355078 328524
rect 364298 328468 364308 328524
rect 364364 328468 643076 328524
rect 643132 328468 643142 328524
rect 112634 328356 112644 328412
rect 112700 328356 169652 328412
rect 169708 328356 169718 328412
rect 172218 328356 172228 328412
rect 172284 328356 191492 328412
rect 191548 328356 191558 328412
rect 224410 328356 224420 328412
rect 224476 328356 261604 328412
rect 261660 328356 261670 328412
rect 265178 328356 265188 328412
rect 265244 328356 372820 328412
rect 372876 328356 372886 328412
rect 377850 328356 377860 328412
rect 377916 328356 672868 328412
rect 672924 328356 672934 328412
rect 166170 328244 166180 328300
rect 166236 328244 189364 328300
rect 189420 328244 189430 328300
rect 236730 328244 236740 328300
rect 236796 328244 293412 328300
rect 293468 328244 293478 328300
rect 334506 328244 334516 328300
rect 334572 328244 335972 328300
rect 336028 328244 336038 328300
rect 338090 328244 338100 328300
rect 338156 328244 571508 328300
rect 571564 328244 571574 328300
rect 168298 328132 168308 328188
rect 168364 328132 190820 328188
rect 190876 328132 190886 328188
rect 233146 328132 233156 328188
rect 233212 328132 285460 328188
rect 285516 328132 285526 328188
rect 297994 328132 298004 328188
rect 298060 328132 462308 328188
rect 462364 328132 462374 328188
rect 114650 328020 114660 328076
rect 114716 328020 170436 328076
rect 170492 328020 170502 328076
rect 232474 328020 232484 328076
rect 232540 328020 281428 328076
rect 281484 328020 281494 328076
rect 291498 328020 291508 328076
rect 291564 328020 444388 328076
rect 444444 328020 444454 328076
rect 230234 327908 230244 327964
rect 230300 327908 275492 327964
rect 275548 327908 275558 327964
rect 335178 327908 335188 327964
rect 335244 327908 343476 327964
rect 343532 327908 343542 327964
rect 343914 327908 343924 327964
rect 343980 327908 390740 327964
rect 390796 327908 390806 327964
rect 391178 327908 391188 327964
rect 391244 327908 421540 327964
rect 421596 327908 421606 327964
rect 335066 327796 335076 327852
rect 335132 327796 343476 327852
rect 343532 327796 343542 327852
rect 343690 327796 343700 327852
rect 343756 327796 367780 327852
rect 367836 327796 367846 327852
rect 381322 327796 381332 327852
rect 381388 327796 408660 327852
rect 408716 327796 408726 327852
rect 334394 327684 334404 327740
rect 334460 327684 347732 327740
rect 347788 327684 347798 327740
rect 358698 327684 358708 327740
rect 358764 327684 373604 327740
rect 373660 327684 373670 327740
rect 334282 327572 334292 327628
rect 334348 327572 346052 327628
rect 346108 327572 346118 327628
rect 367882 327572 367892 327628
rect 367948 327572 369684 327628
rect 369740 327572 369750 327628
rect 368666 327460 368676 327516
rect 368732 327460 369572 327516
rect 369628 327460 369638 327516
rect 376282 327460 376292 327516
rect 376348 327460 381444 327516
rect 381500 327460 381510 327516
rect 386362 327460 386372 327516
rect 386428 327460 391188 327516
rect 391244 327460 391254 327516
rect 453562 327460 453572 327516
rect 453628 327460 468244 327516
rect 468300 327460 468310 327516
rect 308970 327348 308980 327404
rect 309036 327348 492100 327404
rect 492156 327348 492166 327404
rect 317706 327236 317716 327292
rect 317772 327236 515956 327292
rect 516012 327236 516022 327292
rect 236058 327124 236068 327180
rect 236124 327124 295316 327180
rect 295372 327124 295382 327180
rect 319610 327124 319620 327180
rect 319676 327124 521892 327180
rect 521948 327124 521958 327180
rect 238298 327012 238308 327068
rect 238364 327012 299348 327068
rect 299404 327012 299414 327068
rect 335962 327012 335972 327068
rect 336028 327012 341012 327068
rect 341068 327012 341078 327068
rect 341786 327012 341796 327068
rect 341852 327012 354116 327068
rect 354172 327012 354182 327068
rect 354330 327012 354340 327068
rect 354396 327012 569604 327068
rect 569660 327012 569670 327068
rect 242666 326900 242676 326956
rect 242732 326900 311220 326956
rect 311276 326900 311286 326956
rect 328682 326900 328692 326956
rect 328748 326900 545748 326956
rect 545804 326900 545814 326956
rect 257898 326788 257908 326844
rect 257964 326788 345268 326844
rect 345324 326788 345334 326844
rect 350522 326788 350532 326844
rect 350588 326788 605332 326844
rect 605388 326788 605398 326844
rect 278394 326676 278404 326732
rect 278460 326676 381332 326732
rect 381388 326676 381398 326732
rect 382330 326676 382340 326732
rect 382396 326676 647108 326732
rect 647164 326676 647174 326732
rect 300206 326564 300244 326620
rect 300300 326564 300310 326620
rect 300458 326564 300468 326620
rect 300524 326564 456260 326620
rect 456316 326564 456326 326620
rect 293626 326452 293636 326508
rect 293692 326452 450324 326508
rect 450380 326452 450390 326508
rect 282762 326340 282772 326396
rect 282828 326340 418292 326396
rect 418348 326340 418358 326396
rect 295866 326228 295876 326284
rect 295932 326228 300468 326284
rect 300524 326228 300534 326284
rect 376730 326228 376740 326284
rect 376796 326228 379316 326284
rect 379372 326228 379382 326284
rect 470362 326116 470372 326172
rect 470428 326116 474180 326172
rect 474236 326116 474246 326172
rect 304602 326004 304612 326060
rect 304668 326004 480116 326060
rect 480172 326004 480182 326060
rect 381994 325780 382004 325836
rect 382060 325780 382340 325836
rect 382396 325780 382406 325836
rect 303818 325668 303828 325724
rect 303884 325668 353556 325724
rect 353612 325668 353622 325724
rect 360714 325668 360724 325724
rect 360780 325668 488404 325724
rect 488460 325668 488470 325724
rect 321290 325556 321300 325612
rect 321356 325556 525812 325612
rect 525868 325556 525878 325612
rect 292954 325444 292964 325500
rect 293020 325444 320068 325500
rect 320124 325444 320134 325500
rect 327898 325444 327908 325500
rect 327964 325444 542612 325500
rect 542668 325444 542678 325500
rect 244794 325332 244804 325388
rect 244860 325332 315812 325388
rect 315868 325332 315878 325388
rect 330138 325332 330148 325388
rect 330204 325332 549332 325388
rect 549388 325332 549398 325388
rect 247034 325220 247044 325276
rect 247100 325220 322532 325276
rect 322588 325220 322598 325276
rect 334506 325220 334516 325276
rect 334572 325220 561092 325276
rect 561148 325220 561158 325276
rect 162922 325108 162932 325164
rect 162988 325108 187908 325164
rect 187964 325108 187974 325164
rect 249162 325108 249172 325164
rect 249228 325108 327572 325164
rect 327628 325108 327638 325164
rect 340330 325108 340340 325164
rect 340396 325108 353892 325164
rect 353948 325108 353958 325164
rect 367210 325108 367220 325164
rect 367276 325108 650132 325164
rect 650188 325108 650198 325164
rect 703966 325108 704004 325164
rect 704060 325108 704070 325164
rect 704890 325108 704900 325164
rect 704956 325108 705124 325164
rect 705180 325108 705190 325164
rect 157882 324996 157892 325052
rect 157948 324996 185668 325052
rect 185724 324996 185734 325052
rect 251402 324996 251412 325052
rect 251468 324996 334292 325052
rect 334348 324996 334358 325052
rect 337418 324996 337428 325052
rect 337484 324996 354340 325052
rect 354396 324996 354406 325052
rect 367994 324996 368004 325052
rect 368060 324996 376292 325052
rect 376348 324996 376358 325052
rect 376506 324996 376516 325052
rect 376572 324996 673652 325052
rect 673708 324996 673718 325052
rect 701530 324996 701540 325052
rect 701596 324996 704564 325052
rect 704620 324996 704630 325052
rect 354106 324884 354116 324940
rect 354172 324884 471156 324940
rect 471212 324884 471222 324940
rect 505530 324884 505540 324940
rect 505596 324884 512372 324940
rect 512428 324884 512438 324940
rect 655498 324884 655508 324940
rect 655564 324884 661892 324940
rect 661948 324884 661958 324940
rect 349738 324772 349748 324828
rect 349804 324772 454916 324828
rect 454972 324772 454982 324828
rect 345370 324660 345380 324716
rect 345436 324660 437668 324716
rect 437724 324660 437734 324716
rect 295082 324548 295092 324604
rect 295148 324548 386372 324604
rect 386428 324548 386438 324604
rect 537562 324548 537572 324604
rect 537628 324548 537666 324604
rect 308186 324436 308196 324492
rect 308252 324436 370468 324492
rect 370524 324436 370534 324492
rect 554334 324436 554372 324492
rect 554428 324436 554438 324492
rect 161018 324324 161028 324380
rect 161084 324324 161700 324380
rect 161756 324324 161766 324380
rect 347722 324324 347732 324380
rect 347788 324324 353780 324380
rect 353836 324324 353846 324380
rect 375946 324324 375956 324380
rect 376012 324324 376516 324380
rect 376572 324324 376582 324380
rect 376730 324324 376740 324380
rect 376796 324324 376834 324380
rect 705674 324324 705684 324380
rect 705788 324324 705798 324380
rect 159898 324212 159908 324268
rect 159964 324212 161307 324268
rect 161251 324156 161307 324212
rect 161476 324212 161980 324268
rect 194842 324212 194852 324268
rect 194908 324212 195916 324268
rect 195972 324212 195982 324268
rect 199994 324212 200004 324268
rect 200060 324212 201068 324268
rect 201124 324212 201134 324268
rect 211754 324212 211764 324268
rect 211820 324212 212716 324268
rect 212772 324212 212782 324268
rect 216682 324212 216692 324268
rect 216748 324212 217868 324268
rect 217924 324212 217934 324268
rect 240202 324212 240212 324268
rect 240268 324212 241836 324268
rect 241892 324212 241902 324268
rect 274036 324212 396452 324268
rect 396508 324212 396518 324268
rect 161476 324156 161532 324212
rect 104094 324100 104132 324156
rect 104188 324100 104198 324156
rect 150164 324100 161028 324156
rect 161084 324100 161094 324156
rect 161251 324100 161532 324156
rect 161924 324156 161980 324212
rect 161924 324100 165340 324156
rect 165396 324100 165406 324156
rect 166282 324100 166292 324156
rect 166348 324100 166796 324156
rect 166852 324100 166862 324156
rect 169642 324100 169652 324156
rect 169764 324100 169774 324156
rect 186442 324100 186452 324156
rect 186564 324100 186574 324156
rect 191482 324100 191492 324156
rect 191548 324100 193004 324156
rect 193060 324100 193070 324156
rect 201562 324100 201572 324156
rect 201628 324100 201740 324156
rect 201796 324100 201806 324156
rect 203186 324100 203196 324156
rect 203252 324100 205044 324156
rect 205100 324100 205110 324156
rect 205258 324100 205268 324156
rect 205324 324100 206108 324156
rect 206164 324100 206174 324156
rect 208282 324100 208292 324156
rect 208404 324100 208414 324156
rect 213322 324100 213332 324156
rect 213444 324100 213454 324156
rect 214834 324100 214844 324156
rect 214900 324100 217476 324156
rect 217532 324100 217542 324156
rect 219314 324100 219324 324156
rect 219436 324100 219446 324156
rect 225810 324100 225820 324156
rect 225932 324100 225942 324156
rect 230178 324100 230188 324156
rect 230300 324100 230310 324156
rect 233594 324100 233604 324156
rect 233660 324100 234556 324156
rect 234612 324100 234622 324156
rect 236730 324100 236740 324156
rect 236852 324100 236862 324156
rect 253474 324100 253484 324156
rect 253596 324100 253606 324156
rect 255714 324100 255724 324156
rect 255836 324100 255846 324156
rect 258570 324100 258580 324156
rect 258692 324100 258702 324156
rect 259298 324100 259308 324156
rect 259364 324100 260932 324156
rect 260988 324100 260998 324156
rect 261538 324100 261548 324156
rect 261604 324100 262612 324156
rect 262668 324100 262678 324156
rect 263610 324100 263620 324156
rect 263732 324100 263742 324156
rect 269490 324100 269500 324156
rect 269612 324100 269622 324156
rect 273970 324100 273980 324156
rect 274036 324100 274092 324212
rect 291442 324100 291452 324156
rect 291564 324100 291574 324156
rect 295810 324100 295820 324156
rect 295932 324100 295942 324156
rect 299394 324100 299404 324156
rect 299516 324100 299526 324156
rect 302250 324100 302260 324156
rect 302372 324100 302382 324156
rect 306002 324100 306012 324156
rect 306124 324100 306134 324156
rect 308914 324100 308924 324156
rect 309036 324100 309046 324156
rect 311042 324100 311052 324156
rect 311164 324100 311174 324156
rect 317650 324100 317660 324156
rect 317772 324100 317782 324156
rect 330754 324100 330764 324156
rect 330820 324100 333172 324156
rect 333228 324100 333238 324156
rect 336578 324100 336588 324156
rect 336700 324100 336710 324156
rect 339490 324100 339500 324156
rect 339556 324100 341796 324156
rect 341852 324100 341862 324156
rect 347554 324100 347564 324156
rect 347676 324100 347686 324156
rect 356962 324100 356972 324156
rect 357084 324100 357094 324156
rect 358418 324100 358428 324156
rect 358540 324100 358550 324156
rect 361330 324100 361340 324156
rect 361396 324100 365652 324156
rect 365708 324100 365718 324156
rect 369394 324100 369404 324156
rect 369516 324100 369526 324156
rect 373762 324100 373772 324156
rect 373828 324100 377580 324156
rect 377822 324100 377860 324156
rect 377916 324100 377926 324156
rect 672410 324100 672420 324156
rect 672476 324100 683732 324156
rect 683788 324100 683798 324156
rect 135146 323988 135156 324044
rect 135212 323988 149492 324044
rect 149548 323988 149558 324044
rect 150164 323932 150220 324100
rect 151620 323988 161364 324044
rect 161420 323988 161430 324044
rect 161588 323988 166124 324044
rect 166180 323988 166190 324044
rect 260082 323988 260092 324044
rect 260204 323988 260214 324044
rect 325714 323988 325724 324044
rect 325836 323988 325846 324044
rect 330036 323988 334180 324044
rect 334236 323988 334246 324044
rect 335906 323988 335916 324044
rect 335972 323988 340452 324044
rect 340508 323988 340518 324044
rect 365698 323988 365708 324044
rect 365820 323988 365830 324044
rect 370850 323988 370860 324044
rect 370916 323988 374276 324044
rect 374332 323988 374342 324044
rect 374434 323988 374444 324044
rect 374500 323988 377188 324044
rect 377244 323988 377254 324044
rect 133466 323876 133476 323932
rect 133532 323876 150220 323932
rect 150602 323876 150612 323932
rect 150668 323876 151172 323932
rect 151228 323876 151238 323932
rect 151620 323820 151676 323988
rect 161588 323932 161644 323988
rect 330036 323932 330092 323988
rect 377524 323932 377580 324100
rect 377972 323988 384747 324044
rect 672634 323988 672644 324044
rect 672700 323988 682052 324044
rect 682108 323988 682118 324044
rect 377972 323932 378028 323988
rect 384691 323932 384747 323988
rect 159562 323876 159572 323932
rect 159628 323876 160972 323932
rect 161028 323876 161038 323932
rect 161130 323876 161140 323932
rect 161196 323876 161644 323932
rect 161802 323876 161812 323932
rect 161868 323876 162428 323932
rect 162484 323876 162494 323932
rect 162586 323876 162596 323932
rect 162652 323876 167580 323932
rect 167636 323876 167646 323932
rect 184874 323876 184884 323932
rect 184940 323876 197372 323932
rect 197428 323876 197438 323932
rect 241154 323876 241164 323932
rect 241220 323876 249396 323932
rect 249452 323876 249462 323932
rect 316866 323876 316876 323932
rect 316988 323876 316998 323932
rect 324146 323876 324156 323932
rect 324212 323876 330092 323932
rect 332210 323876 332220 323932
rect 332332 323876 332342 323932
rect 333666 323876 333676 323932
rect 333732 323876 347732 323932
rect 347788 323876 347798 323932
rect 371522 323876 371532 323932
rect 371644 323876 371654 323932
rect 372978 323876 372988 323932
rect 373044 323876 376852 323932
rect 376908 323876 376918 323932
rect 377290 323876 377300 323932
rect 377412 323876 377422 323932
rect 377524 323876 378028 323932
rect 378130 323876 378140 323932
rect 378196 323876 378644 323932
rect 378700 323876 378710 323932
rect 378802 323876 378812 323932
rect 378868 323876 379540 323932
rect 379596 323876 379606 323932
rect 384691 323876 485492 323932
rect 485548 323876 485558 323932
rect 149482 323764 149492 323820
rect 149548 323764 151676 323820
rect 151946 323764 151956 323820
rect 152012 323764 159908 323820
rect 159964 323764 159974 323820
rect 380286 323092 380324 323148
rect 380380 323092 380390 323148
rect 133914 322532 133924 322588
rect 133980 322532 159572 322588
rect 159628 322532 159638 322588
rect 672746 322532 672756 322588
rect 672812 322532 680372 322588
rect 680428 322532 680438 322588
rect 379764 322252 379820 322448
rect 379754 322196 379764 322252
rect 379820 322196 379830 322252
rect 159562 321188 159572 321244
rect 159628 321188 160048 321244
rect 379876 319564 379932 319984
rect 379866 319508 379876 319564
rect 379932 319508 379942 319564
rect 557694 319396 557732 319452
rect 557788 319396 557798 319452
rect 379764 317324 379820 317520
rect 379754 317268 379764 317324
rect 379820 317268 379830 317324
rect 159786 316260 159796 316316
rect 159852 316260 160048 316316
rect 75936 314900 76132 314956
rect 76188 314900 76198 314956
rect 379764 314860 379820 315056
rect 379754 314804 379764 314860
rect 379820 314804 379830 314860
rect 76468 314508 77252 314524
rect 75936 314468 77252 314508
rect 77308 314468 77318 314524
rect 75936 314452 76524 314468
rect 84494 314356 84532 314412
rect 84588 314356 84598 314412
rect 75992 314004 76356 314060
rect 76412 314004 76422 314060
rect 75936 313556 76188 313612
rect 76132 313164 76188 313556
rect 671514 313236 671524 313292
rect 671580 313236 687764 313292
rect 687820 313236 687830 313292
rect 75936 313108 76188 313164
rect 83962 312452 83972 312508
rect 84028 312452 84980 312508
rect 85036 312452 85046 312508
rect 379764 312396 379820 312592
rect 460254 312452 460292 312508
rect 460348 312452 460358 312508
rect 379754 312340 379764 312396
rect 379820 312340 379830 312396
rect 75936 312212 76132 312268
rect 76188 312212 76198 312268
rect 75936 311764 76356 311820
rect 76412 311764 76422 311820
rect 84046 311444 84084 311500
rect 84140 311444 84150 311500
rect 159674 311332 159684 311388
rect 159740 311332 160048 311388
rect 379764 309932 379820 310128
rect 379754 309876 379764 309932
rect 379820 309876 379830 309932
rect 458574 309204 458612 309260
rect 458668 309204 458678 309260
rect 695146 309204 695156 309260
rect 695212 309236 701372 309260
rect 695212 309204 702016 309236
rect 701316 309180 702016 309204
rect 164836 308756 173067 308812
rect 164836 308700 164892 308756
rect 173011 308700 173067 308756
rect 198660 308756 208347 308812
rect 198660 308700 198716 308756
rect 208291 308700 208347 308756
rect 309316 308756 321916 308812
rect 309316 308700 309372 308756
rect 164826 308644 164836 308700
rect 164892 308644 164902 308700
rect 173011 308644 195468 308700
rect 195524 308644 195534 308700
rect 198650 308644 198660 308700
rect 198716 308644 198726 308700
rect 199882 308644 199892 308700
rect 199948 308644 203644 308700
rect 208291 308644 211932 308700
rect 211988 308644 211998 308700
rect 220266 308644 220276 308700
rect 220332 308644 222348 308700
rect 222404 308644 222414 308700
rect 232082 308644 232092 308700
rect 232148 308644 240436 308700
rect 240492 308644 240502 308700
rect 247314 308644 247324 308700
rect 247380 308644 248500 308700
rect 248556 308644 248566 308700
rect 254034 308644 254044 308700
rect 254100 308644 254772 308700
rect 254828 308644 254838 308700
rect 257618 308644 257628 308700
rect 257684 308644 293972 308700
rect 294028 308644 294038 308700
rect 307010 308644 307020 308700
rect 307076 308644 309372 308700
rect 309474 308644 309484 308700
rect 309540 308644 321636 308700
rect 321692 308644 321702 308700
rect 203588 308588 203644 308644
rect 321860 308588 321916 308756
rect 384691 308756 670292 308812
rect 670348 308756 670358 308812
rect 384691 308700 384747 308756
rect 322074 308644 322084 308700
rect 322140 308644 337092 308700
rect 337148 308644 337158 308700
rect 341170 308644 341180 308700
rect 341236 308644 342580 308700
rect 342636 308644 342646 308700
rect 343634 308644 343644 308700
rect 343700 308644 344260 308700
rect 344316 308644 344326 308700
rect 356402 308644 356412 308700
rect 356468 308644 357700 308700
rect 357756 308644 357766 308700
rect 369842 308644 369852 308700
rect 369908 308644 370916 308700
rect 370972 308644 370982 308700
rect 377262 308644 377300 308700
rect 377356 308644 377366 308700
rect 377738 308644 377748 308700
rect 377804 308644 384747 308700
rect 701316 308732 702016 308788
rect 162922 308532 162932 308588
rect 162988 308532 164444 308588
rect 164500 308532 164510 308588
rect 164714 308532 164724 308588
rect 164780 308532 165564 308588
rect 165620 308532 165630 308588
rect 166170 308532 166180 308588
rect 166236 308532 188524 308588
rect 191482 308532 191492 308588
rect 191548 308532 192444 308588
rect 192500 308532 192510 308588
rect 193162 308532 193172 308588
rect 193228 308532 193676 308588
rect 193732 308532 193742 308588
rect 203242 308532 203252 308588
rect 203308 308532 203420 308588
rect 203476 308532 203486 308588
rect 203588 308532 212604 308588
rect 212660 308532 212670 308588
rect 213434 308532 213444 308588
rect 213500 308532 218652 308588
rect 218708 308532 218718 308588
rect 218810 308532 218820 308588
rect 218876 308532 221116 308588
rect 221172 308532 221182 308588
rect 231410 308532 231420 308588
rect 231476 308532 237356 308588
rect 237570 308532 237580 308588
rect 237636 308532 238420 308588
rect 238476 308532 238486 308588
rect 242386 308532 242396 308588
rect 242452 308532 262276 308588
rect 262332 308532 262342 308588
rect 262546 308532 262556 308588
rect 262612 308532 263620 308588
rect 263676 308532 263686 308588
rect 273802 308532 273812 308588
rect 273868 308532 274764 308588
rect 274820 308532 274830 308588
rect 279570 308532 279580 308588
rect 279636 308532 290667 308588
rect 296706 308532 296716 308588
rect 296772 308532 297220 308588
rect 297276 308532 297286 308588
rect 300682 308532 300692 308588
rect 300748 308532 302204 308588
rect 302260 308532 302270 308588
rect 307626 308532 307636 308588
rect 307692 308532 308924 308588
rect 308980 308532 308990 308588
rect 313170 308532 313180 308588
rect 313236 308532 313908 308588
rect 313964 308532 313974 308588
rect 316194 308532 316204 308588
rect 316260 308532 317380 308588
rect 317436 308532 317446 308588
rect 320450 308532 320460 308588
rect 320516 308532 320740 308588
rect 320796 308532 320806 308588
rect 320954 308532 320964 308588
rect 321020 308532 321692 308588
rect 321748 308532 321758 308588
rect 321850 308532 321860 308588
rect 321916 308532 321926 308588
rect 322868 308532 325947 308588
rect 188468 308476 188524 308532
rect 164602 308420 164612 308476
rect 164668 308420 166236 308476
rect 166292 308420 166302 308476
rect 168074 308420 168084 308476
rect 168140 308420 169260 308476
rect 169316 308420 169326 308476
rect 171322 308420 171332 308476
rect 171388 308420 172284 308476
rect 172340 308420 172350 308476
rect 173114 308420 173124 308476
rect 173180 308420 174188 308476
rect 174244 308420 174254 308476
rect 176362 308420 176372 308476
rect 176428 308420 177212 308476
rect 177268 308420 177278 308476
rect 179722 308420 179732 308476
rect 179788 308420 180908 308476
rect 180964 308420 180974 308476
rect 181402 308420 181412 308476
rect 181468 308420 182028 308476
rect 182084 308420 182094 308476
rect 183054 308420 183092 308476
rect 183148 308420 183158 308476
rect 184874 308420 184884 308476
rect 184940 308420 186396 308476
rect 186452 308420 186462 308476
rect 188468 308420 194908 308476
rect 194964 308420 194974 308476
rect 199994 308420 200004 308476
rect 200060 308420 200956 308476
rect 201012 308420 201022 308476
rect 201786 308420 201796 308476
rect 201852 308420 202860 308476
rect 202916 308420 202926 308476
rect 206602 308420 206612 308476
rect 206668 308420 207116 308476
rect 207172 308420 207182 308476
rect 209962 308420 209972 308476
rect 210028 308420 210700 308476
rect 210756 308420 210766 308476
rect 215114 308420 215124 308476
rect 215180 308420 219884 308476
rect 219940 308420 219950 308476
rect 225922 308420 225932 308476
rect 225988 308420 228452 308476
rect 228508 308420 228518 308476
rect 230178 308420 230188 308476
rect 230244 308420 237076 308476
rect 237132 308420 237142 308476
rect 237300 308364 237356 308532
rect 238522 308420 238532 308476
rect 238588 308420 240044 308476
rect 240100 308420 240110 308476
rect 241770 308420 241780 308476
rect 241892 308420 241902 308476
rect 243571 308420 258692 308476
rect 258748 308420 258758 308476
rect 260754 308420 260764 308476
rect 260820 308420 261940 308476
rect 261996 308420 262006 308476
rect 263778 308420 263788 308476
rect 263844 308420 265300 308476
rect 265356 308420 265366 308476
rect 265514 308420 265524 308476
rect 265580 308420 266812 308476
rect 266868 308420 266878 308476
rect 270442 308420 270452 308476
rect 270508 308420 271740 308476
rect 271796 308420 271806 308476
rect 280802 308420 280812 308476
rect 280868 308420 282100 308476
rect 282156 308420 282166 308476
rect 283882 308420 283892 308476
rect 283948 308420 285068 308476
rect 285124 308420 285134 308476
rect 285562 308420 285572 308476
rect 285628 308420 286972 308476
rect 287028 308420 287038 308476
rect 287354 308420 287364 308476
rect 287420 308420 288764 308476
rect 288820 308420 288830 308476
rect 243571 308364 243627 308420
rect 290611 308364 290667 308532
rect 322868 308476 322924 308532
rect 325891 308476 325947 308532
rect 329140 308532 376964 308588
rect 377020 308532 377030 308588
rect 329140 308476 329196 308532
rect 292282 308420 292292 308476
rect 292348 308420 293692 308476
rect 293748 308420 293758 308476
rect 294074 308420 294084 308476
rect 294140 308420 295484 308476
rect 295540 308420 295550 308476
rect 300794 308420 300804 308476
rect 300860 308420 301532 308476
rect 301588 308420 301598 308476
rect 302586 308420 302596 308476
rect 302652 308420 303996 308476
rect 304052 308420 304062 308476
rect 304154 308420 304164 308476
rect 304220 308420 305228 308476
rect 305284 308420 305294 308476
rect 307514 308420 307524 308476
rect 307580 308420 308252 308476
rect 308308 308420 308318 308476
rect 309194 308420 309204 308476
rect 309260 308420 310716 308476
rect 310772 308420 310782 308476
rect 310874 308420 310884 308476
rect 310940 308420 311948 308476
rect 312004 308420 312014 308476
rect 312498 308420 312508 308476
rect 312564 308420 313796 308476
rect 313852 308420 313862 308476
rect 314234 308420 314244 308476
rect 314300 308420 315644 308476
rect 315700 308420 315710 308476
rect 317482 308420 317492 308476
rect 317548 308420 318668 308476
rect 318724 308420 318734 308476
rect 319890 308420 319900 308476
rect 319956 308420 322924 308476
rect 324202 308420 324212 308476
rect 324268 308420 325388 308476
rect 325444 308420 325454 308476
rect 325891 308420 329196 308476
rect 329354 308420 329364 308476
rect 329420 308420 330876 308476
rect 330932 308420 330942 308476
rect 331034 308420 331044 308476
rect 331100 308420 331996 308476
rect 332052 308420 332062 308476
rect 332658 308420 332668 308476
rect 332724 308420 334180 308476
rect 334236 308420 334246 308476
rect 336186 308420 336196 308476
rect 336252 308420 336364 308476
rect 336420 308420 336430 308476
rect 337651 308420 361227 308476
rect 362562 308420 362572 308476
rect 362628 308420 362740 308476
rect 362796 308420 362806 308476
rect 363122 308420 363132 308476
rect 363188 308420 364420 308476
rect 364476 308420 364486 308476
rect 368610 308420 368620 308476
rect 368676 308420 369460 308476
rect 369516 308420 369526 308476
rect 377122 308420 377132 308476
rect 377188 308420 377860 308476
rect 377916 308420 377926 308476
rect 378074 308420 378084 308476
rect 378140 308420 379036 308476
rect 379092 308420 379102 308476
rect 337651 308364 337707 308420
rect 157882 308308 157892 308364
rect 157948 308308 189644 308364
rect 190558 308308 190596 308364
rect 190652 308308 190662 308364
rect 190810 308308 190820 308364
rect 190876 308308 206388 308364
rect 206444 308308 206454 308364
rect 216906 308308 216916 308364
rect 216972 308308 220388 308364
rect 220444 308308 220454 308364
rect 234574 308308 234612 308364
rect 234668 308308 234678 308364
rect 237300 308308 240324 308364
rect 240380 308308 240390 308364
rect 240650 308308 240660 308364
rect 240716 308308 243627 308364
rect 254762 308308 254772 308364
rect 254828 308308 287252 308364
rect 287308 308308 287318 308364
rect 290611 308308 308084 308364
rect 308140 308308 308150 308364
rect 310202 308308 310212 308364
rect 310268 308308 330036 308364
rect 330092 308308 330102 308364
rect 330250 308308 330260 308364
rect 330316 308308 337707 308364
rect 361171 308364 361227 308420
rect 361171 308308 377412 308364
rect 377468 308308 377478 308364
rect 189588 308252 189644 308308
rect 151162 308196 151172 308252
rect 151228 308196 189364 308252
rect 189420 308196 189430 308252
rect 189588 308196 191492 308252
rect 191548 308196 191558 308252
rect 196858 308196 196868 308252
rect 196924 308196 211316 308252
rect 211372 308196 211382 308252
rect 229674 308196 229684 308252
rect 229740 308196 235284 308252
rect 235340 308196 235350 308252
rect 243674 308196 243684 308252
rect 243740 308196 265412 308252
rect 265468 308196 265478 308252
rect 277274 308196 277284 308252
rect 277340 308196 336420 308252
rect 336476 308196 336486 308252
rect 378074 308196 378084 308252
rect 378140 308196 379428 308252
rect 379484 308196 379494 308252
rect 154634 308084 154644 308140
rect 154700 308084 191156 308140
rect 191212 308084 191222 308140
rect 193386 308084 193396 308140
rect 193452 308084 209412 308140
rect 209468 308084 209478 308140
rect 230906 308084 230916 308140
rect 230972 308084 238644 308140
rect 238700 308084 238710 308140
rect 241210 308084 241220 308140
rect 241276 308084 260596 308140
rect 260652 308084 260662 308140
rect 263610 308084 263620 308140
rect 263676 308084 305732 308140
rect 305788 308084 305798 308140
rect 313898 308084 313908 308140
rect 313964 308084 337428 308140
rect 337484 308084 337494 308140
rect 376618 308084 376628 308140
rect 376684 308084 548436 308140
rect 548492 308084 548502 308140
rect 92362 307972 92372 308028
rect 92428 307972 161252 308028
rect 161308 307972 161318 308028
rect 163034 307972 163044 308028
rect 163100 307972 166180 308028
rect 166236 307972 166246 308028
rect 173002 307972 173012 308028
rect 173068 307972 199668 308028
rect 199724 307972 199734 308028
rect 208394 307972 208404 308028
rect 208460 307972 216804 308028
rect 216860 307972 216870 308028
rect 237066 307972 237076 308028
rect 237132 307972 237412 308028
rect 237468 307972 237478 308028
rect 246698 307972 246708 308028
rect 246764 307972 272132 308028
rect 272188 307972 272198 308028
rect 281530 307972 281540 308028
rect 281596 307972 301700 308028
rect 301756 307972 301766 308028
rect 315018 307972 315028 308028
rect 315084 307972 414932 308028
rect 414988 307972 414998 308028
rect 106026 307860 106036 307916
rect 106092 307860 167412 307916
rect 167468 307860 167478 307916
rect 186554 307860 186564 307916
rect 186620 307860 190820 307916
rect 190876 307860 190886 307916
rect 194954 307860 194964 307916
rect 195020 307860 210084 307916
rect 210140 307860 210150 307916
rect 233370 307860 233380 307916
rect 233436 307860 243684 307916
rect 243740 307860 243750 307916
rect 251066 307860 251076 307916
rect 251132 307860 280644 307916
rect 280700 307860 280710 307916
rect 290611 307860 302372 307916
rect 302428 307860 302438 307916
rect 325994 307860 326004 307916
rect 326060 307860 438452 307916
rect 438508 307860 438518 307916
rect 290611 307804 290667 307860
rect 105802 307748 105812 307804
rect 105868 307748 167972 307804
rect 168028 307748 168038 307804
rect 191594 307748 191604 307804
rect 191660 307748 208292 307804
rect 208348 307748 208358 307804
rect 251934 307748 251972 307804
rect 252028 307748 252038 307804
rect 261370 307748 261380 307804
rect 261436 307748 290667 307804
rect 335738 307748 335748 307804
rect 335804 307748 462756 307804
rect 462812 307748 462822 307804
rect 532382 307748 532420 307804
rect 532476 307748 532486 307804
rect 104122 307636 104132 307692
rect 104188 307636 166740 307692
rect 166796 307636 166806 307692
rect 184762 307636 184772 307692
rect 184828 307636 205268 307692
rect 205324 307636 205334 307692
rect 210074 307636 210084 307692
rect 210140 307636 217364 307692
rect 217420 307636 217430 307692
rect 218586 307636 218596 307692
rect 218652 307636 221620 307692
rect 221676 307636 221686 307692
rect 233930 307636 233940 307692
rect 233996 307636 238700 307692
rect 238858 307636 238868 307692
rect 238924 307636 255332 307692
rect 255388 307636 255398 307692
rect 293066 307636 293076 307692
rect 293132 307636 336644 307692
rect 336700 307636 336710 307692
rect 344922 307636 344932 307692
rect 344988 307636 482916 307692
rect 482972 307636 482982 307692
rect 238644 307580 238700 307636
rect 100762 307524 100772 307580
rect 100828 307524 164948 307580
rect 165004 307524 165014 307580
rect 165386 307524 165396 307580
rect 165452 307524 182644 307580
rect 182700 307524 182710 307580
rect 183418 307524 183428 307580
rect 183484 307524 204596 307580
rect 204652 307524 204662 307580
rect 211866 307524 211876 307580
rect 211932 307524 218036 307580
rect 218092 307524 218102 307580
rect 229114 307524 229124 307580
rect 229180 307524 235172 307580
rect 235228 307524 235238 307580
rect 238644 307524 245252 307580
rect 245308 307524 245318 307580
rect 250394 307524 250404 307580
rect 250460 307524 278852 307580
rect 278908 307524 278918 307580
rect 282090 307524 282100 307580
rect 282156 307524 301476 307580
rect 301532 307524 301542 307580
rect 306506 307524 306516 307580
rect 306572 307524 319956 307580
rect 320012 307524 320022 307580
rect 322970 307524 322980 307580
rect 323036 307524 336756 307580
rect 336812 307524 336822 307580
rect 370906 307524 370916 307580
rect 370972 307524 534212 307580
rect 534268 307524 534278 307580
rect 701316 307468 701372 308732
rect 99054 307412 99092 307468
rect 99148 307412 99158 307468
rect 102442 307412 102452 307468
rect 102508 307412 102546 307468
rect 190026 307412 190036 307468
rect 190092 307412 207620 307468
rect 207676 307412 207686 307468
rect 213658 307412 213668 307468
rect 213724 307412 219156 307468
rect 219212 307412 219222 307468
rect 227210 307412 227220 307468
rect 227276 307412 230132 307468
rect 230188 307412 230198 307468
rect 232698 307412 232708 307468
rect 232764 307412 241892 307468
rect 241948 307412 241958 307468
rect 282762 307412 282772 307468
rect 282828 307412 289716 307468
rect 289772 307412 289782 307468
rect 303930 307412 303940 307468
rect 303996 307412 307860 307468
rect 307916 307412 307926 307468
rect 330026 307412 330036 307468
rect 330092 307412 337204 307468
rect 337260 307412 337270 307468
rect 377822 307412 377860 307468
rect 377916 307412 377926 307468
rect 426654 307412 426692 307468
rect 426748 307412 426758 307468
rect 550974 307412 551012 307468
rect 551068 307412 551078 307468
rect 686858 307412 686868 307468
rect 686924 307412 701372 307468
rect 701876 307836 702016 307892
rect 701876 307444 701932 307836
rect 701876 307388 702016 307444
rect 265066 307300 265076 307356
rect 265132 307300 310772 307356
rect 310828 307300 310838 307356
rect 358922 307300 358932 307356
rect 358988 307300 510692 307356
rect 510748 307300 510758 307356
rect 289370 307188 289380 307244
rect 289436 307188 361172 307244
rect 361228 307188 361238 307244
rect 371690 307188 371700 307244
rect 371756 307188 538580 307244
rect 538636 307188 538646 307244
rect 290042 307076 290052 307132
rect 290108 307076 362852 307132
rect 362908 307076 362918 307132
rect 372362 307076 372372 307132
rect 372428 307076 539252 307132
rect 539308 307076 539318 307132
rect 290490 306964 290500 307020
rect 290556 306964 364532 307020
rect 364588 306964 364598 307020
rect 371018 306964 371028 307020
rect 371084 306964 538356 307020
rect 538412 306964 538422 307020
rect 694922 306964 694932 307020
rect 694988 306996 701372 307020
rect 694988 306964 702016 306996
rect 701316 306940 702016 306964
rect 159674 306852 159684 306908
rect 159740 306852 337092 306908
rect 337148 306852 337158 306908
rect 374154 306852 374164 306908
rect 374220 306852 543396 306908
rect 543452 306852 543462 306908
rect 84858 306740 84868 306796
rect 84924 306740 657636 306796
rect 657692 306740 657702 306796
rect 85194 306628 85204 306684
rect 85260 306628 659316 306684
rect 659372 306628 659382 306684
rect 83402 306516 83412 306572
rect 83468 306516 670628 306572
rect 670684 306516 670694 306572
rect 695146 306516 695156 306572
rect 695212 306548 701372 306572
rect 695212 306516 702016 306548
rect 701316 306492 702016 306516
rect 264394 306404 264404 306460
rect 264460 306404 309092 306460
rect 309148 306404 309158 306460
rect 357130 306404 357140 306460
rect 357196 306404 508116 306460
rect 508172 306404 508182 306460
rect 344250 306292 344260 306348
rect 344316 306292 481236 306348
rect 481292 306292 481302 306348
rect 701316 306044 702016 306100
rect 701316 306012 701372 306044
rect 686746 305956 686756 306012
rect 686812 305956 701372 306012
rect 159898 305844 159908 305900
rect 159964 305844 160020 305900
rect 160076 305844 160086 305900
rect 84634 305732 84644 305788
rect 84700 305732 84756 305788
rect 84812 305732 84822 305788
rect 169754 305620 169764 305676
rect 169820 305620 170996 305676
rect 171052 305620 171062 305676
rect 174682 305620 174692 305676
rect 174748 305620 175924 305676
rect 175980 305620 175990 305676
rect 176474 305620 176484 305676
rect 176540 305620 177716 305676
rect 177772 305620 177782 305676
rect 252074 305620 252084 305676
rect 252140 305620 252756 305676
rect 252812 305620 252822 305676
rect 299226 305620 299236 305676
rect 299292 305620 300244 305676
rect 300300 305620 300310 305676
rect 302698 305620 302708 305676
rect 302764 305620 303380 305676
rect 303436 305620 303446 305676
rect 327674 305620 327684 305676
rect 327740 305620 328916 305676
rect 328972 305620 328982 305676
rect 349738 305620 349748 305676
rect 349804 305620 492996 305676
rect 493052 305620 493062 305676
rect 351642 305508 351652 305564
rect 351708 305508 496356 305564
rect 496412 305508 496422 305564
rect 352202 305396 352212 305452
rect 352268 305396 497252 305452
rect 497308 305396 497318 305452
rect 352874 305284 352884 305340
rect 352940 305284 498932 305340
rect 498988 305284 498998 305340
rect 364970 305172 364980 305228
rect 365036 305172 524916 305228
rect 524972 305172 524982 305228
rect 364410 305060 364420 305116
rect 364476 305060 523236 305116
rect 523292 305060 523302 305116
rect 367434 304948 367444 305004
rect 367500 304948 529956 305004
rect 530012 304948 530022 305004
rect 369338 304836 369348 304892
rect 369404 304836 532532 304892
rect 532588 304836 532598 304892
rect 347946 304724 347956 304780
rect 348012 304724 489636 304780
rect 489692 304724 489702 304780
rect 348506 304612 348516 304668
rect 348572 304612 488852 304668
rect 488908 304612 488918 304668
rect 372810 303940 372820 303996
rect 372876 303940 385924 303996
rect 385980 303940 385990 303996
rect 520510 303940 520548 303996
rect 520604 303940 520614 303996
rect 345482 303828 345492 303884
rect 345548 303828 482132 303884
rect 482188 303828 482198 303884
rect 285562 303716 285572 303772
rect 285628 303716 300692 303772
rect 300748 303716 300758 303772
rect 346714 303716 346724 303772
rect 346780 303716 485492 303772
rect 485548 303716 485558 303772
rect 522302 303716 522340 303772
rect 522396 303716 522406 303772
rect 258906 303604 258916 303660
rect 258972 303604 297332 303660
rect 297388 303604 297398 303660
rect 359370 303604 359380 303660
rect 359436 303604 513156 303660
rect 513212 303604 513222 303660
rect 253418 303492 253428 303548
rect 253484 303492 285908 303548
rect 285964 303492 285974 303548
rect 294298 303492 294308 303548
rect 294364 303492 341796 303548
rect 341852 303492 341862 303548
rect 374826 303492 374836 303548
rect 374892 303492 545076 303548
rect 545132 303492 545142 303548
rect 270554 303380 270564 303436
rect 270620 303380 320852 303436
rect 320908 303380 320918 303436
rect 373594 303380 373604 303436
rect 373660 303380 543508 303436
rect 543564 303380 543574 303436
rect 188122 303268 188132 303324
rect 188188 303268 201348 303324
rect 201404 303268 201414 303324
rect 279066 303268 279076 303324
rect 279132 303268 339332 303324
rect 339388 303268 339398 303324
rect 375386 303268 375396 303324
rect 375452 303268 546756 303324
rect 546812 303268 546822 303324
rect 171546 303156 171556 303212
rect 171612 303156 199108 303212
rect 199164 303156 199174 303212
rect 277834 303156 277844 303212
rect 277900 303156 337652 303212
rect 337708 303156 337718 303212
rect 375946 303156 375956 303212
rect 376012 303156 548548 303212
rect 548604 303156 548614 303212
rect 342458 303044 342468 303100
rect 342524 303044 477876 303100
rect 477932 303044 477942 303100
rect 83150 302372 83188 302428
rect 83244 302372 83254 302428
rect 335822 302260 335860 302316
rect 335916 302260 335926 302316
rect 285982 302148 286020 302204
rect 286076 302148 286086 302204
rect 285534 302036 285572 302092
rect 285628 302036 285638 302092
rect 282986 301924 282996 301980
rect 283052 301924 348516 301980
rect 348572 301924 348582 301980
rect 282314 301812 282324 301868
rect 282380 301812 349748 301868
rect 349804 301812 349814 301868
rect 354862 301812 354900 301868
rect 354956 301812 354966 301868
rect 283882 301700 283892 301756
rect 283948 301700 352772 301756
rect 352828 301700 352838 301756
rect 664346 301700 664356 301756
rect 664412 301700 670628 301756
rect 670684 301700 670694 301756
rect 248714 301588 248724 301644
rect 248780 301588 278964 301644
rect 279020 301588 279030 301644
rect 285758 301588 285796 301644
rect 285852 301588 285862 301644
rect 337082 301588 337092 301644
rect 337148 301588 560196 301644
rect 560252 301588 560262 301644
rect 662666 301588 662676 301644
rect 662732 301588 671188 301644
rect 671244 301588 671254 301644
rect 248938 301476 248948 301532
rect 249004 301476 277172 301532
rect 277228 301476 277238 301532
rect 278058 301476 278068 301532
rect 278124 301476 335748 301532
rect 335804 301476 335814 301532
rect 336858 301476 336868 301532
rect 336924 301476 566020 301532
rect 566076 301476 566086 301532
rect 657626 301476 657636 301532
rect 657692 301476 671188 301532
rect 671244 301476 671254 301532
rect 356094 301364 356132 301420
rect 356188 301364 356198 301420
rect 292254 300580 292292 300636
rect 292348 300580 292358 300636
rect 294494 300580 294532 300636
rect 294588 300580 294598 300636
rect 298974 300580 299012 300636
rect 299068 300580 299078 300636
rect 302558 300580 302596 300636
rect 302652 300580 302662 300636
rect 302782 300580 302820 300636
rect 302876 300580 302886 300636
rect 284218 300468 284228 300524
rect 284284 300468 335412 300524
rect 335468 300468 335478 300524
rect 337194 300468 337204 300524
rect 337260 300468 376628 300524
rect 376684 300468 376694 300524
rect 287914 300356 287924 300412
rect 287980 300356 359492 300412
rect 359548 300356 359558 300412
rect 287354 300244 287364 300300
rect 287420 300244 359940 300300
rect 359996 300244 360006 300300
rect 252298 300132 252308 300188
rect 252364 300132 283892 300188
rect 283948 300132 283958 300188
rect 300682 300132 300692 300188
rect 300748 300132 388164 300188
rect 388220 300132 388230 300188
rect 252074 300020 252084 300076
rect 252140 300020 284452 300076
rect 284508 300020 284518 300076
rect 302698 300020 302708 300076
rect 302764 300020 391524 300076
rect 391580 300020 391590 300076
rect 259018 299908 259028 299964
rect 259084 299908 299796 299964
rect 299852 299908 299862 299964
rect 304266 299908 304276 299964
rect 304332 299908 393316 299964
rect 393372 299908 393382 299964
rect 258794 299796 258804 299852
rect 258860 299796 299012 299852
rect 299068 299796 299078 299852
rect 307626 299796 307636 299852
rect 307692 299796 399812 299852
rect 399868 299796 399878 299852
rect 336634 299684 336644 299740
rect 336700 299684 369572 299740
rect 369628 299684 369638 299740
rect 381742 299684 381780 299740
rect 381836 299684 381846 299740
rect 389694 299684 389732 299740
rect 389788 299684 389798 299740
rect 295754 299572 295764 299628
rect 295820 299572 345156 299628
rect 345212 299572 345222 299628
rect 274250 298452 274260 298508
rect 274316 298452 318276 298508
rect 318332 298452 318342 298508
rect 265626 298340 265636 298396
rect 265692 298340 311332 298396
rect 311388 298340 311398 298396
rect 314234 298340 314244 298396
rect 314300 298340 335524 298396
rect 335580 298340 335590 298396
rect 294074 298228 294084 298284
rect 294140 298228 343700 298284
rect 343756 298228 343766 298284
rect 274026 298116 274036 298172
rect 274092 298116 329476 298172
rect 329532 298116 329542 298172
rect 272346 297780 272356 297836
rect 272412 297780 273028 297836
rect 273084 297780 273094 297836
rect 310958 297220 310996 297276
rect 311052 297220 311062 297276
rect 309194 296772 309204 296828
rect 309260 296772 335636 296828
rect 335692 296772 335702 296828
rect 305834 296660 305844 296716
rect 305900 296660 334628 296716
rect 334684 296660 334694 296716
rect 73098 296548 73108 296604
rect 73164 296548 77588 296604
rect 77644 296548 77654 296604
rect 270890 296548 270900 296604
rect 270956 296548 322868 296604
rect 322924 296548 322934 296604
rect 337418 296548 337428 296604
rect 337484 296548 397460 296604
rect 397516 296548 397526 296604
rect 73546 296436 73556 296492
rect 73612 296436 77812 296492
rect 77868 296436 77878 296492
rect 272458 296436 272468 296492
rect 272524 296436 326676 296492
rect 326732 296436 326742 296492
rect 336970 296436 336980 296492
rect 337036 296436 397236 296492
rect 397292 296436 397302 296492
rect 72202 296324 72212 296380
rect 72268 296324 77924 296380
rect 77980 296324 77990 296380
rect 72650 296212 72660 296268
rect 72716 296212 78148 296268
rect 78204 296212 78214 296268
rect 336970 294980 336980 295036
rect 337036 294980 403508 295036
rect 403564 294980 403574 295036
rect 337194 294868 337204 294924
rect 337260 294868 404852 294924
rect 404908 294868 404918 294924
rect 146122 294756 146132 294812
rect 146188 294756 186676 294812
rect 186732 294756 186742 294812
rect 275594 294756 275604 294812
rect 275660 294756 332724 294812
rect 332780 294756 332790 294812
rect 336186 294756 336196 294812
rect 336252 294756 463764 294812
rect 463820 294756 463830 294812
rect 502282 294308 502292 294364
rect 502348 294308 624708 294364
rect 624764 294308 624774 294364
rect 503962 294196 503972 294252
rect 504028 294196 625268 294252
rect 625324 294196 625334 294252
rect 483802 294084 483812 294140
rect 483868 294084 606116 294140
rect 606172 294084 606182 294140
rect 485482 293972 485492 294028
rect 485548 293972 618548 294028
rect 618604 293972 618614 294028
rect 490634 293860 490644 293916
rect 490700 293860 491316 293916
rect 491372 293860 491382 293916
rect 509002 293860 509012 293916
rect 509068 293860 509796 293916
rect 509852 293860 509862 293916
rect 514042 293860 514052 293916
rect 514108 293860 514836 293916
rect 514892 293860 514902 293916
rect 542602 293860 542612 293916
rect 542668 293860 543396 293916
rect 543452 293860 543462 293916
rect 544394 293860 544404 293916
rect 544460 293860 545076 293916
rect 545132 293860 545142 293916
rect 549546 293860 549556 293916
rect 549612 293860 550116 293916
rect 550172 293860 550182 293916
rect 494666 293636 494676 293692
rect 494732 293636 621908 293692
rect 621964 293636 621974 293692
rect 539214 293412 539252 293468
rect 539308 293412 539318 293468
rect 547642 293412 547652 293468
rect 547708 293412 548548 293468
rect 548604 293412 641508 293468
rect 641564 293412 641574 293468
rect 545962 293300 545972 293356
rect 546028 293300 546756 293356
rect 546812 293300 641060 293356
rect 641116 293300 641126 293356
rect 336746 293188 336756 293244
rect 336812 293188 418292 293244
rect 418348 293188 418358 293244
rect 544394 293188 544404 293244
rect 544460 293188 640612 293244
rect 640668 293188 640678 293244
rect 336074 293076 336084 293132
rect 336140 293076 465332 293132
rect 465388 293076 465398 293132
rect 542602 293076 542612 293132
rect 542668 293076 640052 293132
rect 640108 293076 640118 293132
rect 510654 292964 510692 293020
rect 510748 292964 510758 293020
rect 514042 292964 514052 293020
rect 514108 292964 629076 293020
rect 629132 292964 629142 293020
rect 488814 292852 488852 292908
rect 488908 292852 488918 292908
rect 490634 292852 490644 292908
rect 490700 292852 606116 292908
rect 606172 292852 606182 292908
rect 498894 292740 498932 292796
rect 498988 292740 498998 292796
rect 512362 292740 512372 292796
rect 512428 292740 513156 292796
rect 513212 292740 628628 292796
rect 628684 292740 628694 292796
rect 489066 292628 489076 292684
rect 489132 292628 489636 292684
rect 489692 292628 605780 292684
rect 605836 292628 605846 292684
rect 497214 292516 497252 292572
rect 497308 292516 497318 292572
rect 509002 292516 509012 292572
rect 509068 292516 627172 292572
rect 627228 292516 627238 292572
rect 502291 292404 623812 292460
rect 623868 292404 623878 292460
rect 502291 292348 502347 292404
rect 465294 292292 465332 292348
rect 465388 292292 465398 292348
rect 493882 292292 493892 292348
rect 493948 292292 494676 292348
rect 494732 292292 494742 292348
rect 499706 292292 499716 292348
rect 499772 292292 502347 292348
rect 609802 292292 609812 292348
rect 609868 292292 670292 292348
rect 670348 292292 670358 292348
rect 92362 292180 92372 292236
rect 92428 292180 92484 292236
rect 92540 292180 92550 292236
rect 320926 292180 320964 292236
rect 321020 292180 321030 292236
rect 321150 292180 321188 292236
rect 321244 292180 321254 292236
rect 321402 292180 321412 292236
rect 321468 292180 321506 292236
rect 507322 292180 507332 292236
rect 507388 292180 508116 292236
rect 508172 292180 508182 292236
rect 522666 292180 522676 292236
rect 522732 292180 523236 292236
rect 523292 292180 523302 292236
rect 540922 292180 540932 292236
rect 540988 292180 541716 292236
rect 541772 292180 541782 292236
rect 542714 292180 542724 292236
rect 542780 292180 543508 292236
rect 543564 292180 543574 292236
rect 613498 292068 613508 292124
rect 613564 292068 620900 292124
rect 620956 292068 620966 292124
rect 93146 291956 93156 292012
rect 93212 291956 669396 292012
rect 669452 291956 669462 292012
rect 173198 291844 173236 291900
rect 173292 291844 173302 291900
rect 316026 291844 316036 291900
rect 316092 291844 418964 291900
rect 419020 291844 419030 291900
rect 428782 291844 428820 291900
rect 428876 291844 428886 291900
rect 606218 291844 606228 291900
rect 606284 291844 621348 291900
rect 621404 291844 621414 291900
rect 152842 291732 152852 291788
rect 152908 291732 189924 291788
rect 189980 291732 189990 291788
rect 317706 291732 317716 291788
rect 317772 291732 421652 291788
rect 421708 291732 421718 291788
rect 428558 291732 428596 291788
rect 428652 291732 428662 291788
rect 508106 291732 508116 291788
rect 508172 291732 626612 291788
rect 626668 291732 626678 291788
rect 142986 291620 142996 291676
rect 143052 291620 184996 291676
rect 185052 291620 185062 291676
rect 315914 291620 315924 291676
rect 315980 291620 420196 291676
rect 420252 291620 420262 291676
rect 534174 291620 534212 291676
rect 534268 291620 534278 291676
rect 548426 291620 548436 291676
rect 548492 291620 642068 291676
rect 642124 291620 642134 291676
rect 648778 291620 648788 291676
rect 648844 291620 671524 291676
rect 671580 291620 671590 291676
rect 142762 291508 142772 291564
rect 142828 291508 185444 291564
rect 185500 291508 185510 291564
rect 317482 291508 317492 291564
rect 317548 291508 423444 291564
rect 423500 291508 423510 291564
rect 430350 291508 430388 291564
rect 430444 291508 430454 291564
rect 505978 291508 505988 291564
rect 506044 291508 506436 291564
rect 506492 291508 506502 291564
rect 525914 291508 525924 291564
rect 525980 291508 526596 291564
rect 526652 291508 536172 291564
rect 543498 291508 543508 291564
rect 543564 291508 639604 291564
rect 639660 291508 639670 291564
rect 647322 291508 647332 291564
rect 647388 291508 671076 291564
rect 671132 291508 671142 291564
rect 120922 291396 120932 291452
rect 120988 291396 174916 291452
rect 174972 291396 174982 291452
rect 369674 291396 369684 291452
rect 369740 291396 535892 291452
rect 535948 291396 535958 291452
rect 536116 291340 536172 291508
rect 537562 291396 537572 291452
rect 537628 291396 538356 291452
rect 538412 291396 637700 291452
rect 637756 291396 637766 291452
rect 645866 291396 645876 291452
rect 645932 291396 671300 291452
rect 671356 291396 671366 291452
rect 532494 291284 532532 291340
rect 532588 291284 532598 291340
rect 536116 291284 633332 291340
rect 633388 291284 633398 291340
rect 524122 291172 524132 291228
rect 524188 291172 524916 291228
rect 524972 291172 632884 291228
rect 632940 291172 632950 291228
rect 117870 291060 117908 291116
rect 117964 291060 117974 291116
rect 522666 291060 522676 291116
rect 522732 291060 632436 291116
rect 632492 291060 632502 291116
rect 521294 290948 521332 291004
rect 521388 290948 521398 291004
rect 609802 290948 609812 291004
rect 609868 290948 644868 291004
rect 644924 290948 644934 291004
rect 535854 290836 535892 290892
rect 535948 290836 535958 290892
rect 540922 290836 540932 290892
rect 540988 290836 639156 290892
rect 639212 290836 639222 290892
rect 463754 290724 463764 290780
rect 463820 290724 642964 290780
rect 643020 290724 643030 290780
rect 92558 290612 92596 290668
rect 92652 290612 92662 290668
rect 606330 290612 606340 290668
rect 606396 290612 614404 290668
rect 614460 290612 614470 290668
rect 614964 290612 615916 290668
rect 658858 290612 658868 290668
rect 658924 290612 670068 290668
rect 670124 290612 670134 290668
rect 614964 290556 615020 290612
rect 615860 290556 615916 290612
rect 475374 290500 475412 290556
rect 475468 290500 475478 290556
rect 482906 290500 482916 290556
rect 482972 290500 615020 290556
rect 615076 290500 615412 290556
rect 615468 290500 615478 290556
rect 615626 290500 615636 290556
rect 615692 290500 615730 290556
rect 615860 290500 617092 290556
rect 617148 290500 617158 290556
rect 637214 290500 637252 290556
rect 637308 290500 637318 290556
rect 643514 290500 643524 290556
rect 643580 290500 646548 290556
rect 646604 290500 646614 290556
rect 668378 290500 668388 290556
rect 668444 290500 669844 290556
rect 669900 290500 669910 290556
rect 689294 290500 689332 290556
rect 689388 290500 689398 290556
rect 615076 290444 615132 290500
rect 139178 290388 139188 290444
rect 139244 290388 165396 290444
rect 165452 290388 165462 290444
rect 481226 290388 481236 290444
rect 481292 290388 607796 290444
rect 607852 290388 607862 290444
rect 608020 290388 615132 290444
rect 615290 290388 615300 290444
rect 615356 290388 616084 290444
rect 616140 290388 616150 290444
rect 616410 290388 616420 290444
rect 616476 290388 619892 290444
rect 619948 290388 619958 290444
rect 666026 290388 666036 290444
rect 666092 290388 670292 290444
rect 670348 290388 670358 290444
rect 688174 290388 688212 290444
rect 688268 290388 688278 290444
rect 608020 290332 608076 290388
rect 79706 290276 79716 290332
rect 79772 290276 80276 290332
rect 80332 290276 80342 290332
rect 141754 290276 141764 290332
rect 141820 290276 168756 290332
rect 168812 290276 168822 290332
rect 472014 290276 472052 290332
rect 472108 290276 472118 290332
rect 477866 290276 477876 290332
rect 477932 290276 478660 290332
rect 478716 290276 608076 290332
rect 608906 290276 608916 290332
rect 608972 290276 614516 290332
rect 614572 290276 614582 290332
rect 614730 290276 614740 290332
rect 614796 290276 626667 290332
rect 666922 290276 666932 290332
rect 666988 290276 672420 290332
rect 672476 290276 672486 290332
rect 626611 290220 626667 290276
rect 160234 290164 160244 290220
rect 160300 290164 191716 290220
rect 191772 290164 191782 290220
rect 606302 290164 606340 290220
rect 606396 290164 606406 290220
rect 607786 290164 607796 290220
rect 607852 290164 614460 290220
rect 614730 290164 614740 290220
rect 614796 290164 614852 290220
rect 614908 290164 614918 290220
rect 615076 290164 616532 290220
rect 616588 290164 616598 290220
rect 617316 290164 620452 290220
rect 620508 290164 620518 290220
rect 626611 290164 648228 290220
rect 648284 290164 648294 290220
rect 662666 290164 662676 290220
rect 662732 290164 672084 290220
rect 672140 290164 672150 290220
rect 614404 290108 614460 290164
rect 615076 290108 615132 290164
rect 617316 290108 617372 290164
rect 72762 290052 72772 290108
rect 72828 290052 72838 290108
rect 78026 290052 78036 290108
rect 78092 290052 78820 290108
rect 78876 290052 78886 290108
rect 149482 290052 149492 290108
rect 149548 290052 188244 290108
rect 188300 290052 188310 290108
rect 606106 290052 606116 290108
rect 606172 290052 611044 290108
rect 611100 290052 611110 290108
rect 611492 290052 614180 290108
rect 614236 290052 614246 290108
rect 614404 290052 615132 290108
rect 615402 290052 615412 290108
rect 615468 290052 617372 290108
rect 617502 290052 617540 290108
rect 617596 290052 617606 290108
rect 619780 290052 629468 290108
rect 631754 290052 631764 290108
rect 631820 290052 642740 290108
rect 642796 290052 642806 290108
rect 643411 290052 646884 290108
rect 646940 290052 646950 290108
rect 664122 290052 664132 290108
rect 664188 290052 666932 290108
rect 666988 290052 666998 290108
rect 667146 290052 667156 290108
rect 667212 290052 671188 290108
rect 671244 290052 671254 290108
rect 72772 289996 72828 290052
rect 611492 289996 611548 290052
rect 619780 289996 619836 290052
rect 629412 289996 629468 290052
rect 643411 289996 643467 290052
rect 72772 289940 78092 289996
rect 150714 289940 150724 289996
rect 150780 289940 188356 289996
rect 188412 289940 188422 289996
rect 336746 289940 336756 289996
rect 336812 289940 432516 289996
rect 432572 289940 432582 289996
rect 610922 289940 610932 289996
rect 610988 289940 611268 289996
rect 611324 289940 611334 289996
rect 611482 289940 611492 289996
rect 611548 289940 611558 289996
rect 611930 289940 611940 289996
rect 611996 289940 619836 289996
rect 620666 289940 620676 289996
rect 620732 289940 629188 289996
rect 629244 289940 629254 289996
rect 629412 289940 643467 289996
rect 644186 289940 644196 289996
rect 644252 289940 656964 289996
rect 657020 289940 657030 289996
rect 667268 289940 671188 289996
rect 671244 289940 671254 289996
rect 78036 289884 78092 289940
rect 667268 289884 667324 289940
rect 72202 289828 72212 289884
rect 72268 289828 77700 289884
rect 77756 289828 77766 289884
rect 78026 289828 78036 289884
rect 78092 289828 78102 289884
rect 83066 289828 83076 289884
rect 83132 289828 651588 289884
rect 651644 289828 651654 289884
rect 652558 289828 652596 289884
rect 652652 289828 652662 289884
rect 657402 289828 657412 289884
rect 657468 289828 661948 289884
rect 663114 289828 663124 289884
rect 663180 289828 667324 289884
rect 670282 289828 670292 289884
rect 670348 289828 671300 289884
rect 671356 289828 671366 289884
rect 672270 289828 672308 289884
rect 672364 289828 672374 289884
rect 704638 289828 704676 289884
rect 704732 289828 704742 289884
rect 704974 289828 705012 289884
rect 705068 289828 705078 289884
rect 661892 289772 661948 289828
rect 73546 289716 73556 289772
rect 73612 289716 77924 289772
rect 77980 289716 77990 289772
rect 83850 289716 83860 289772
rect 83916 289716 596427 289772
rect 596371 289660 596427 289716
rect 603091 289716 620676 289772
rect 620732 289716 620742 289772
rect 622766 289716 622804 289772
rect 622860 289716 622870 289772
rect 623214 289716 623252 289772
rect 623308 289716 623318 289772
rect 626126 289716 626164 289772
rect 626220 289716 626230 289772
rect 628030 289716 628068 289772
rect 628124 289716 628134 289772
rect 629038 289716 629076 289772
rect 629132 289716 629142 289772
rect 629290 289716 629300 289772
rect 629356 289716 631764 289772
rect 631820 289716 631830 289772
rect 631950 289716 631988 289772
rect 632044 289716 632054 289772
rect 636206 289716 636244 289772
rect 636300 289716 636310 289772
rect 636654 289716 636692 289772
rect 636748 289716 636758 289772
rect 638110 289716 638148 289772
rect 638204 289716 638214 289772
rect 638670 289716 638708 289772
rect 638764 289716 638774 289772
rect 640014 289716 640052 289772
rect 640108 289716 640118 289772
rect 640574 289716 640612 289772
rect 640668 289716 640678 289772
rect 641022 289716 641060 289772
rect 641116 289716 641126 289772
rect 641470 289716 641508 289772
rect 641564 289716 641574 289772
rect 642478 289716 642516 289772
rect 642572 289716 642582 289772
rect 642730 289716 642740 289772
rect 642796 289716 644196 289772
rect 644252 289716 644262 289772
rect 644382 289716 644420 289772
rect 644476 289716 644486 289772
rect 652250 289716 652260 289772
rect 652316 289716 653044 289772
rect 653100 289716 653110 289772
rect 655470 289716 655508 289772
rect 655564 289716 655574 289772
rect 658270 289716 658308 289772
rect 658364 289716 658374 289772
rect 661630 289716 661668 289772
rect 661724 289716 661734 289772
rect 661892 289716 666932 289772
rect 666988 289716 666998 289772
rect 667230 289716 667268 289772
rect 667324 289716 667334 289772
rect 667454 289716 667492 289772
rect 667548 289716 667558 289772
rect 670842 289716 670852 289772
rect 670908 289716 671076 289772
rect 671132 289716 671142 289772
rect 671626 289716 671636 289772
rect 671692 289716 687652 289772
rect 687708 289716 687718 289772
rect 603091 289660 603147 289716
rect 73098 289604 73108 289660
rect 73164 289604 77812 289660
rect 77868 289604 77878 289660
rect 596371 289604 603147 289660
rect 609811 289604 611380 289660
rect 611436 289604 611446 289660
rect 609811 289548 609867 289604
rect 600506 289492 600516 289548
rect 600572 289492 609867 289548
rect 702090 289380 702100 289436
rect 702156 289380 704836 289436
rect 704892 289380 704902 289436
rect 479518 289268 479556 289324
rect 479612 289268 479622 289324
rect 337502 289156 337540 289212
rect 337596 289156 337606 289212
rect 600506 289156 600516 289212
rect 600572 289156 609812 289212
rect 609868 289156 609878 289212
rect 687502 289156 687540 289212
rect 687596 289156 687606 289212
rect 479546 289044 479556 289100
rect 479612 289044 608916 289100
rect 608972 289044 608982 289100
rect 701978 289044 701988 289100
rect 702044 289044 705572 289100
rect 705628 289044 705638 289100
rect 611342 288820 611380 288876
rect 611436 288820 611446 288876
rect 559178 288484 559188 288540
rect 559244 288484 603147 288540
rect 603091 288428 603147 288484
rect 468804 288372 470932 288428
rect 470988 288372 596427 288428
rect 603091 288372 611744 288428
rect 671552 288372 671860 288428
rect 671916 288372 671926 288428
rect 137946 288260 137956 288316
rect 138012 288260 165396 288316
rect 165452 288260 165462 288316
rect 337978 288260 337988 288316
rect 338044 288260 468580 288316
rect 468636 288260 468646 288316
rect 468804 288204 468860 288372
rect 596371 288316 596427 288372
rect 596371 288260 610708 288316
rect 610764 288260 610774 288316
rect 136602 288148 136612 288204
rect 136668 288148 165620 288204
rect 165676 288148 165686 288204
rect 339434 288148 339444 288204
rect 339500 288148 468860 288204
rect 474506 288148 474516 288204
rect 474572 288148 606340 288204
rect 606396 288148 606406 288204
rect 611006 288148 611044 288204
rect 611100 288148 611110 288204
rect 162250 288036 162260 288092
rect 162316 288036 193284 288092
rect 193340 288036 193350 288092
rect 337754 288036 337764 288092
rect 337820 288036 469140 288092
rect 469196 288036 469206 288092
rect 472826 288036 472836 288092
rect 472892 288036 606228 288092
rect 606284 288036 606294 288092
rect 468542 287252 468580 287308
rect 468636 287252 468646 287308
rect 469102 287252 469140 287308
rect 469196 287252 469206 287308
rect 474478 287252 474516 287308
rect 474572 287252 474582 287308
rect 114874 286580 114884 286636
rect 114940 286580 171668 286636
rect 171724 286580 171734 286636
rect 112298 286468 112308 286524
rect 112364 286468 169876 286524
rect 169932 286468 169942 286524
rect 90570 286356 90580 286412
rect 90636 286356 159684 286412
rect 159740 286356 159750 286412
rect 559066 286132 559076 286188
rect 559132 286132 611744 286188
rect 94042 285572 94052 285628
rect 94108 285572 94948 285628
rect 95004 285572 95014 285628
rect 142762 285572 142772 285628
rect 142828 285572 143668 285628
rect 143724 285572 143734 285628
rect 186554 285572 186564 285628
rect 186620 285572 187236 285628
rect 187292 285572 187302 285628
rect 208394 285572 208404 285628
rect 208460 285572 208964 285628
rect 209020 285572 209030 285628
rect 218586 285572 218596 285628
rect 218652 285572 219268 285628
rect 219324 285572 219334 285628
rect 230122 285572 230132 285628
rect 230188 285572 230692 285628
rect 230748 285572 230758 285628
rect 423322 285572 423332 285628
rect 423388 285572 424116 285628
rect 424172 285572 424182 285628
rect 428586 285572 428596 285628
rect 428652 285572 429268 285628
rect 429324 285572 429334 285628
rect 488842 285572 488852 285628
rect 488908 285572 489524 285628
rect 489580 285572 489590 285628
rect 493882 285572 493892 285628
rect 493948 285572 494564 285628
rect 494620 285572 494630 285628
rect 324426 285460 324436 285516
rect 324492 285460 332667 285516
rect 324202 285348 324212 285404
rect 324268 285348 330316 285404
rect 327870 285236 327908 285292
rect 327964 285236 327974 285292
rect 330260 285068 330316 285348
rect 332611 285180 332667 285460
rect 332611 285124 436324 285180
rect 436380 285124 436390 285180
rect 327786 285012 327796 285068
rect 327852 285012 329980 285068
rect 330260 285012 437668 285068
rect 437724 285012 437734 285068
rect 329924 284956 329980 285012
rect 117450 284900 117460 284956
rect 117516 284900 171444 284956
rect 171500 284900 171510 284956
rect 327646 284900 327684 284956
rect 327740 284900 327750 284956
rect 329550 284900 329588 284956
rect 329644 284900 329654 284956
rect 329924 284900 442708 284956
rect 442764 284900 442774 284956
rect 116106 284788 116116 284844
rect 116172 284788 171332 284844
rect 171388 284788 171398 284844
rect 325882 284788 325892 284844
rect 325948 284788 441476 284844
rect 441532 284788 441542 284844
rect 113530 284676 113540 284732
rect 113596 284676 169764 284732
rect 169820 284676 169830 284732
rect 377962 284676 377972 284732
rect 378028 284676 556724 284732
rect 556780 284676 556790 284732
rect 444014 284564 444052 284620
rect 444108 284564 444118 284620
rect 558842 283892 558852 283948
rect 558908 283892 611744 283948
rect 671552 283780 671860 283836
rect 671916 283780 671926 283836
rect 90346 283220 90356 283276
rect 90412 283220 609924 283276
rect 609980 283220 609990 283276
rect 78810 283108 78820 283164
rect 78876 283108 609924 283164
rect 609980 283108 609990 283164
rect 78474 282996 78484 283052
rect 78540 282996 609812 283052
rect 609868 282996 609878 283052
rect 334394 282212 334404 282268
rect 334460 282212 334470 282268
rect 334404 282156 334460 282212
rect 196522 282100 196532 282156
rect 196588 282100 196626 282156
rect 262014 282100 262052 282156
rect 262108 282100 262118 282156
rect 262378 282100 262388 282156
rect 262444 282100 263508 282156
rect 263564 282100 263574 282156
rect 334394 282100 334404 282156
rect 334460 282100 334470 282156
rect 334590 282100 334628 282156
rect 334684 282100 334694 282156
rect 391402 282100 391412 282156
rect 391468 282100 392756 282156
rect 392812 282100 392822 282156
rect 445246 282100 445284 282156
rect 445340 282100 445350 282156
rect 446590 282100 446628 282156
rect 446684 282100 446694 282156
rect 704666 282100 704676 282156
rect 704732 282100 705012 282156
rect 705068 282100 705078 282156
rect 168410 281988 168420 282044
rect 168476 281988 178164 282044
rect 178220 281988 178230 282044
rect 267530 281988 267540 282044
rect 267596 281988 274036 282044
rect 274092 281988 274102 282044
rect 314131 281988 320628 282044
rect 320684 281988 320694 282044
rect 320852 281988 329307 282044
rect 335402 281988 335412 282044
rect 335468 281988 351764 282044
rect 351820 281988 351830 282044
rect 704666 281988 704676 282044
rect 704732 281988 705012 282044
rect 705068 281988 705078 282044
rect 153738 281876 153748 281932
rect 153804 281876 159908 281932
rect 159964 281876 159974 281932
rect 173786 281876 173796 281932
rect 173852 281876 179732 281932
rect 179788 281876 179798 281932
rect 245354 281876 245364 281932
rect 245420 281876 269892 281932
rect 269948 281876 269958 281932
rect 140522 281764 140532 281820
rect 140588 281764 144844 281820
rect 145562 281764 145572 281820
rect 145628 281764 184884 281820
rect 184940 281764 184950 281820
rect 247034 281764 247044 281820
rect 247100 281764 276276 281820
rect 276332 281764 276342 281820
rect 144788 281708 144844 281764
rect 314131 281708 314187 281988
rect 320852 281932 320908 281988
rect 316810 281876 316820 281932
rect 316876 281876 320908 281932
rect 329251 281932 329307 281988
rect 329251 281876 344148 281932
rect 344204 281876 344214 281932
rect 702090 281876 702100 281932
rect 702156 281876 704836 281932
rect 704892 281876 704902 281932
rect 316586 281764 316596 281820
rect 316652 281764 318444 281820
rect 335850 281764 335860 281820
rect 335916 281764 381220 281820
rect 381276 281764 381286 281820
rect 397226 281764 397236 281820
rect 397292 281764 410676 281820
rect 410732 281764 410742 281820
rect 134026 281652 134036 281708
rect 134092 281652 143612 281708
rect 144788 281652 179787 281708
rect 253866 281652 253876 281708
rect 253932 281652 289044 281708
rect 289100 281652 289110 281708
rect 308186 281652 308196 281708
rect 308252 281652 314187 281708
rect 143556 281596 143612 281652
rect 179731 281596 179787 281652
rect 318388 281596 318444 281764
rect 320618 281652 320628 281708
rect 320684 281652 341572 281708
rect 341628 281652 341638 281708
rect 341786 281652 341796 281708
rect 341852 281652 342804 281708
rect 342860 281652 342870 281708
rect 352762 281652 352772 281708
rect 352828 281652 354340 281708
rect 354396 281652 354406 281708
rect 397450 281652 397460 281708
rect 397516 281652 412020 281708
rect 412076 281652 412086 281708
rect 143556 281540 173796 281596
rect 173852 281540 173862 281596
rect 179731 281540 183204 281596
rect 183260 281540 183270 281596
rect 196634 281540 196644 281596
rect 196700 281540 202020 281596
rect 202076 281540 202086 281596
rect 243786 281540 243796 281596
rect 243852 281540 267316 281596
rect 267372 281540 267382 281596
rect 267530 281540 267540 281596
rect 267596 281540 317268 281596
rect 317324 281540 317334 281596
rect 318388 281540 342804 281596
rect 342860 281540 342870 281596
rect 343466 281540 343476 281596
rect 343532 281540 373604 281596
rect 373660 281540 373670 281596
rect 377178 281540 377188 281596
rect 377244 281540 426132 281596
rect 426188 281540 426198 281596
rect 605546 281540 605556 281596
rect 605612 281540 611744 281596
rect 135370 281428 135380 281484
rect 135436 281428 181524 281484
rect 181580 281428 181590 281484
rect 182746 281428 182756 281484
rect 182812 281428 191547 281484
rect 191491 281372 191547 281428
rect 196531 281428 203812 281484
rect 203868 281428 203878 281484
rect 253642 281428 253652 281484
rect 253708 281428 290388 281484
rect 290444 281428 290454 281484
rect 301466 281428 301476 281484
rect 301532 281428 346724 281484
rect 346780 281428 346790 281484
rect 358474 281428 358484 281484
rect 358540 281428 362740 281484
rect 362796 281428 362806 281484
rect 377514 281428 377524 281484
rect 377580 281428 447860 281484
rect 447916 281428 447926 281484
rect 671552 281428 687316 281484
rect 687372 281428 687382 281484
rect 196531 281372 196587 281428
rect 126410 281316 126420 281372
rect 126476 281316 176148 281372
rect 176204 281316 176214 281372
rect 176362 281316 176372 281372
rect 176428 281316 185780 281372
rect 185836 281316 185846 281372
rect 191491 281316 196587 281372
rect 196746 281316 196756 281372
rect 196812 281316 201684 281372
rect 201740 281316 201750 281372
rect 267194 281316 267204 281372
rect 267260 281316 315924 281372
rect 315980 281316 315990 281372
rect 318266 281316 318276 281372
rect 318332 281316 332612 281372
rect 332668 281316 332678 281372
rect 335738 281316 335748 281372
rect 335804 281316 338996 281372
rect 339052 281316 339062 281372
rect 342580 281316 406868 281372
rect 406924 281316 406934 281372
rect 705674 281316 705684 281372
rect 705788 281316 705798 281372
rect 342580 281260 342636 281316
rect 128986 281204 128996 281260
rect 129052 281204 153972 281260
rect 154028 281204 154038 281260
rect 154196 281204 162316 281260
rect 162474 281204 162484 281260
rect 162540 281204 168420 281260
rect 168476 281204 168486 281260
rect 168644 281204 176596 281260
rect 176652 281204 176662 281260
rect 180170 281204 180180 281260
rect 180236 281204 201796 281260
rect 201852 281204 201862 281260
rect 270442 281204 270452 281260
rect 270508 281204 324884 281260
rect 324940 281204 324950 281260
rect 335626 281204 335636 281260
rect 335692 281204 342636 281260
rect 342794 281204 342804 281260
rect 342860 281204 372260 281260
rect 372316 281204 372326 281260
rect 377626 281204 377636 281260
rect 377692 281204 453012 281260
rect 453068 281204 453078 281260
rect 558730 281204 558740 281260
rect 558796 281204 570500 281260
rect 570556 281204 570566 281260
rect 154196 281148 154252 281204
rect 162260 281148 162316 281204
rect 168644 281148 168700 281204
rect 122490 281092 122500 281148
rect 122556 281092 122566 281148
rect 125066 281092 125076 281148
rect 125132 281092 154252 281148
rect 154308 281092 162204 281148
rect 162260 281092 168700 281148
rect 168756 281092 174804 281148
rect 174860 281092 174870 281148
rect 178938 281092 178948 281148
rect 179004 281092 185612 281148
rect 185770 281092 185780 281148
rect 185836 281092 200004 281148
rect 200060 281092 200070 281148
rect 237178 281092 237188 281148
rect 237244 281092 254436 281148
rect 254492 281092 254502 281148
rect 257114 281092 257124 281148
rect 257180 281092 294196 281148
rect 294252 281092 294262 281148
rect 314458 281092 314468 281148
rect 314524 281092 414596 281148
rect 414652 281092 414662 281148
rect 122500 281036 122556 281092
rect 154308 281036 154364 281092
rect 162148 281036 162204 281092
rect 168756 281036 168812 281092
rect 185556 281036 185612 281092
rect 122500 280980 154364 281036
rect 154420 280980 162092 281036
rect 162148 280980 168812 281036
rect 169642 280980 169652 281036
rect 169708 280980 169718 281036
rect 177930 280980 177940 281036
rect 177996 280980 185276 281036
rect 185556 280980 196644 281036
rect 196700 280980 196710 281036
rect 196970 280980 196980 281036
rect 197036 280980 197046 281036
rect 198314 280980 198324 281036
rect 198380 280980 198390 281036
rect 203578 280980 203588 281036
rect 203644 280980 213556 281036
rect 213612 280980 213622 281036
rect 238522 280980 238532 281036
rect 238588 280980 238598 281036
rect 243562 280980 243572 281036
rect 243628 280980 255387 281036
rect 273802 280980 273812 281036
rect 273868 280980 273878 281036
rect 274026 280980 274036 281036
rect 274092 280980 317828 281036
rect 317884 280980 317894 281036
rect 321626 280980 321636 281036
rect 321692 280980 398580 281036
rect 398636 280980 398646 281036
rect 558282 280980 558292 281036
rect 558348 280980 570388 281036
rect 570444 280980 570454 281036
rect 154420 280924 154476 280980
rect 162036 280924 162092 280980
rect 169652 280924 169708 280980
rect 185220 280924 185276 280980
rect 100762 280868 100772 280924
rect 100828 280868 101444 280924
rect 101500 280868 101510 280924
rect 111626 280868 111636 280924
rect 111692 280868 154476 280924
rect 154606 280868 154644 280924
rect 154700 280868 154710 280924
rect 159786 280868 159796 280924
rect 159852 280868 160580 280924
rect 160636 280868 160646 280924
rect 162036 280868 169708 280924
rect 175690 280868 175700 280924
rect 175756 280868 180740 280924
rect 180796 280868 180806 280924
rect 181598 280868 181636 280924
rect 181692 280868 181702 280924
rect 185220 280868 196756 280924
rect 196812 280868 196822 280924
rect 196980 280812 197036 280980
rect 109050 280756 109060 280812
rect 109116 280756 167972 280812
rect 168028 280756 168038 280812
rect 170538 280756 170548 280812
rect 170604 280756 197036 280812
rect 198324 280700 198380 280980
rect 92250 280644 92260 280700
rect 92316 280644 153748 280700
rect 153804 280644 153814 280700
rect 153962 280644 153972 280700
rect 154028 280644 162484 280700
rect 162540 280644 162550 280700
rect 171322 280644 171332 280700
rect 171388 280644 198380 280700
rect 238532 280700 238588 280980
rect 255331 280924 255387 280980
rect 273812 280924 273868 280980
rect 245242 280868 245252 280924
rect 245308 280868 246148 280924
rect 246204 280868 246214 280924
rect 255331 280868 267876 280924
rect 267932 280868 267942 280924
rect 272122 280868 272132 280924
rect 272188 280868 273252 280924
rect 273308 280868 273318 280924
rect 273812 280868 330932 280924
rect 330988 280868 330998 280924
rect 343690 280868 343700 280924
rect 343756 280868 374612 280924
rect 374668 280868 374678 280924
rect 378074 280868 378084 280924
rect 378140 280868 461748 280924
rect 461804 280868 461814 280924
rect 461962 280868 461972 280924
rect 462028 280868 462644 280924
rect 462700 280868 462710 280924
rect 477838 280868 477876 280924
rect 477932 280868 477942 280924
rect 482122 280868 482132 280924
rect 482188 280868 483028 280924
rect 483084 280868 483094 280924
rect 537562 280868 537572 280924
rect 537628 280868 538244 280924
rect 538300 280868 538310 280924
rect 557722 280868 557732 280924
rect 557788 280868 559076 280924
rect 559132 280868 559142 280924
rect 243571 280756 257684 280812
rect 257740 280756 257750 280812
rect 263498 280756 263508 280812
rect 263564 280756 306404 280812
rect 306460 280756 306470 280812
rect 307626 280756 307636 280812
rect 307692 280756 402388 280812
rect 402444 280756 402454 280812
rect 558618 280756 558628 280812
rect 558684 280756 570276 280812
rect 570332 280756 570342 280812
rect 243571 280700 243627 280756
rect 238532 280644 243627 280700
rect 245578 280644 245588 280700
rect 245644 280644 270452 280700
rect 270508 280644 270518 280700
rect 272570 280644 272580 280700
rect 272636 280644 328132 280700
rect 328188 280644 328198 280700
rect 338426 280644 338436 280700
rect 338492 280644 370468 280700
rect 370524 280644 370534 280700
rect 379754 280644 379764 280700
rect 379820 280644 554820 280700
rect 554876 280644 554886 280700
rect 559290 279636 559300 279692
rect 559356 279636 559366 279692
rect 559300 279104 559356 279636
rect 607226 279300 607236 279356
rect 607292 279300 611744 279356
rect 570378 277060 570388 277116
rect 570444 277060 611744 277116
rect 671552 276836 671748 276892
rect 671804 276836 671814 276892
rect 559290 276724 559300 276780
rect 559356 276724 559366 276780
rect 559300 276192 559356 276724
rect 603866 274708 603876 274764
rect 603932 274708 611744 274764
rect 671552 274484 687204 274540
rect 687260 274484 687270 274540
rect 76234 274036 76244 274092
rect 76300 274036 78708 274092
rect 78764 274036 78774 274092
rect 75936 273900 76132 273956
rect 76188 273900 76198 273956
rect 76346 273924 76356 273980
rect 76412 273924 78260 273980
rect 78316 273924 78326 273980
rect 76468 273812 78484 273868
rect 78540 273812 78550 273868
rect 76468 273508 76524 273812
rect 75936 273452 76524 273508
rect 559290 273476 559300 273532
rect 559356 273476 559366 273532
rect 559300 273280 559356 273476
rect 75992 273004 76468 273060
rect 76524 273004 76534 273060
rect 75936 272556 76244 272612
rect 76300 272556 76310 272612
rect 602298 272468 602308 272524
rect 602364 272468 611744 272524
rect 85054 272132 85092 272188
rect 85148 272132 85158 272188
rect 75936 271212 76132 271268
rect 76188 271212 76198 271268
rect 75936 270764 76244 270820
rect 76300 270764 76310 270820
rect 84158 270788 84196 270844
rect 84252 270788 84262 270844
rect 559290 270452 559300 270508
rect 559356 270452 559366 270508
rect 559300 270368 559356 270452
rect 570490 270340 570500 270396
rect 570556 270340 605556 270396
rect 605612 270340 605622 270396
rect 570266 270228 570276 270284
rect 570332 270228 611744 270284
rect 671552 269892 689220 269948
rect 689276 269892 689286 269948
rect 602186 267988 602196 268044
rect 602252 267988 611744 268044
rect 671552 267652 688436 267708
rect 688492 267652 688502 267708
rect 560308 267148 560364 267344
rect 560308 267092 607236 267148
rect 607292 267092 607302 267148
rect 694810 266196 694820 266252
rect 694876 266236 701372 266252
rect 694876 266196 702016 266236
rect 701316 266180 702016 266196
rect 693130 265748 693140 265804
rect 693196 265788 701372 265804
rect 693196 265748 702016 265788
rect 701316 265732 702016 265748
rect 600618 265636 600628 265692
rect 600684 265636 611744 265692
rect 559290 265076 559300 265132
rect 559356 265076 559366 265132
rect 559300 264432 559356 265076
rect 701876 264836 702016 264892
rect 701876 264444 701932 264836
rect 701876 264388 702016 264444
rect 701316 263940 702016 263996
rect 701316 263900 701372 263940
rect 686410 263844 686420 263900
rect 686476 263844 701372 263900
rect 697946 263508 697956 263564
rect 698012 263548 701372 263564
rect 698012 263508 702016 263548
rect 701316 263492 702016 263508
rect 559290 263396 559300 263452
rect 559356 263396 611744 263452
rect 701316 263044 702016 263100
rect 671552 262948 689220 263004
rect 689276 262948 689286 263004
rect 701316 262220 701372 263044
rect 686858 262164 686868 262220
rect 686924 262164 701372 262220
rect 560308 260764 560364 261520
rect 597146 261156 597156 261212
rect 597212 261156 611744 261212
rect 560308 260708 567867 260764
rect 671552 260708 688324 260764
rect 688380 260708 688390 260764
rect 567811 260428 567867 260708
rect 567811 260372 603876 260428
rect 603932 260372 603942 260428
rect 585386 258804 585396 258860
rect 585452 258804 611744 258860
rect 560308 257852 560364 258608
rect 560308 257796 567867 257852
rect 567811 257068 567867 257796
rect 567811 257012 602308 257068
rect 602364 257012 602374 257068
rect 560410 256564 560420 256620
rect 560476 256564 611744 256620
rect 559290 256116 559300 256172
rect 559356 256116 559366 256172
rect 671552 256116 689108 256172
rect 689164 256116 689174 256172
rect 559300 255584 559356 256116
rect 73098 255220 73108 255276
rect 73164 255220 76356 255276
rect 76412 255220 76422 255276
rect 73546 255108 73556 255164
rect 73612 255108 77476 255164
rect 77532 255108 77542 255164
rect 72538 254996 72548 255052
rect 72604 254996 77364 255052
rect 77420 254996 77430 255052
rect 72986 254884 72996 254940
rect 73052 254884 78372 254940
rect 78428 254884 78438 254940
rect 559626 254324 559636 254380
rect 559692 254324 611744 254380
rect 671552 253764 691236 253820
rect 691292 253764 691302 253820
rect 560308 252140 560364 252672
rect 560308 252084 602196 252140
rect 602252 252084 602262 252140
rect 608131 252084 611744 252140
rect 608131 252028 608187 252084
rect 560074 251972 560084 252028
rect 560140 251972 608187 252028
rect 560308 249116 560364 249760
rect 561091 249732 611744 249788
rect 561091 249676 561147 249732
rect 560858 249620 560868 249676
rect 560924 249620 561147 249676
rect 671552 249172 689556 249228
rect 689612 249172 689622 249228
rect 73210 249060 73220 249116
rect 73276 249060 78148 249116
rect 78204 249060 78214 249116
rect 560308 249060 561147 249116
rect 72202 248836 72212 248892
rect 72268 248836 77588 248892
rect 77644 248836 77654 248892
rect 561091 248780 561147 249060
rect 73546 248724 73556 248780
rect 73612 248724 77476 248780
rect 77532 248724 77542 248780
rect 561091 248724 600628 248780
rect 600684 248724 600694 248780
rect 72650 248612 72660 248668
rect 72716 248612 77364 248668
rect 77420 248612 77430 248668
rect 560634 247492 560644 247548
rect 560700 247492 611744 247548
rect 559300 246932 559524 246988
rect 559580 246932 559590 246988
rect 559300 246848 559356 246932
rect 671552 246820 689556 246876
rect 689612 246820 689622 246876
rect 704638 246820 704676 246876
rect 704732 246820 704742 246876
rect 704554 246260 704564 246316
rect 704620 246260 705284 246316
rect 705340 246260 705350 246316
rect 560970 245252 560980 245308
rect 561036 245252 611744 245308
rect 559300 243628 559356 243824
rect 559290 243572 559300 243628
rect 559356 243572 559366 243628
rect 583706 242900 583716 242956
rect 583772 242900 611744 242956
rect 671552 242228 689780 242284
rect 689836 242228 689846 242284
rect 560308 240380 560364 240912
rect 560522 240660 560532 240716
rect 560588 240660 611744 240716
rect 560308 240324 597156 240380
rect 597212 240324 597222 240380
rect 559738 240212 559748 240268
rect 559804 240212 560532 240268
rect 560588 240212 560598 240268
rect 671552 239876 692916 239932
rect 692972 239876 692982 239932
rect 704526 239092 704564 239148
rect 704620 239092 704630 239148
rect 560308 238420 560420 238476
rect 560476 238420 560486 238476
rect 561866 238420 561876 238476
rect 561932 238420 611744 238476
rect 704666 238420 704676 238476
rect 704732 238420 705284 238476
rect 705340 238420 705350 238476
rect 560308 238000 560364 238420
rect 560410 236180 560420 236236
rect 560476 236180 611744 236236
rect 671552 235284 689668 235340
rect 689724 235284 689734 235340
rect 559626 235172 559636 235228
rect 559692 235172 559702 235228
rect 559636 235088 559692 235172
rect 559962 233828 559972 233884
rect 560028 233828 611744 233884
rect 76346 233492 76356 233548
rect 76412 233492 78820 233548
rect 78876 233492 78886 233548
rect 671552 233044 694596 233100
rect 694652 233044 694662 233100
rect 75936 232900 76132 232956
rect 76188 232900 76198 232956
rect 560074 232708 560084 232764
rect 560140 232708 560150 232764
rect 75936 232452 76356 232508
rect 76412 232452 76422 232508
rect 75992 232004 76468 232060
rect 76524 232004 76534 232060
rect 84606 232036 84644 232092
rect 84700 232036 84710 232092
rect 560084 232064 560140 232708
rect 85166 231812 85204 231868
rect 85260 231812 85270 231868
rect 75936 231556 76244 231612
rect 76300 231556 76310 231612
rect 559850 231588 559860 231644
rect 559916 231588 611744 231644
rect 75936 230212 76132 230268
rect 76188 230212 76198 230268
rect 75936 229764 76356 229820
rect 76412 229764 76422 229820
rect 565226 229348 565236 229404
rect 565292 229348 611744 229404
rect 560336 229124 560868 229180
rect 560924 229124 560934 229180
rect 671552 228340 689892 228396
rect 689948 228340 689958 228396
rect 566906 226996 566916 227052
rect 566972 226996 611744 227052
rect 560336 226212 560644 226268
rect 560700 226212 560710 226268
rect 671552 226100 694708 226156
rect 694764 226100 694774 226156
rect 560858 224756 560868 224812
rect 560924 224756 611744 224812
rect 560336 223300 560980 223356
rect 561036 223300 561046 223356
rect 694922 223188 694932 223244
rect 694988 223236 701372 223244
rect 694988 223188 702016 223236
rect 701316 223180 702016 223188
rect 700522 222740 700532 222796
rect 700588 222788 701372 222796
rect 700588 222740 702016 222788
rect 701316 222732 702016 222740
rect 560634 222516 560644 222572
rect 560700 222516 611744 222572
rect 701876 221836 702016 221892
rect 671552 221508 690004 221564
rect 690060 221508 690070 221564
rect 701876 221444 701932 221836
rect 701876 221388 702016 221444
rect 701316 220940 702016 220996
rect 701316 220892 701372 220940
rect 690451 220836 701372 220892
rect 560074 220388 560084 220444
rect 560140 220388 561147 220444
rect 561091 220332 561147 220388
rect 560308 220220 560364 220304
rect 561091 220276 611744 220332
rect 560308 220164 583716 220220
rect 583772 220164 583782 220220
rect 690451 220108 690507 220836
rect 695034 220500 695044 220556
rect 695100 220548 701372 220556
rect 695100 220500 702016 220548
rect 701316 220492 702016 220500
rect 686298 220052 686308 220108
rect 686364 220052 690507 220108
rect 701418 220044 701428 220100
rect 701484 220044 702016 220100
rect 671552 219156 694596 219212
rect 694652 219156 694662 219212
rect 686746 218372 686756 218428
rect 686812 218372 701428 218428
rect 701484 218372 701494 218428
rect 559738 217924 559748 217980
rect 559804 217924 559814 217980
rect 578666 217924 578676 217980
rect 578732 217924 611744 217980
rect 559748 217392 559804 217924
rect 560970 215684 560980 215740
rect 561036 215684 611744 215740
rect 73098 214564 73108 214620
rect 73164 214564 77812 214620
rect 77868 214564 77878 214620
rect 671552 214564 689668 214620
rect 689724 214564 689734 214620
rect 73546 214452 73556 214508
rect 73612 214452 78036 214508
rect 78092 214452 78102 214508
rect 560336 214452 561876 214508
rect 561932 214452 561942 214508
rect 72202 214340 72212 214396
rect 72268 214340 77700 214396
rect 77756 214340 77766 214396
rect 72650 214228 72660 214284
rect 72716 214228 77924 214284
rect 77980 214228 77990 214284
rect 568586 213444 568596 213500
rect 568652 213444 611744 213500
rect 671552 212212 694708 212268
rect 694764 212212 694774 212268
rect 560336 211540 560532 211596
rect 560588 211540 560598 211596
rect 568698 211092 568708 211148
rect 568764 211092 611744 211148
rect 559290 209188 559300 209244
rect 559356 209188 561147 209244
rect 559962 209076 559972 209132
rect 560028 209076 560038 209132
rect 559972 208544 560028 209076
rect 561091 208908 561147 209188
rect 561091 208852 611744 208908
rect 72650 207844 72660 207900
rect 72716 207844 84644 207900
rect 84700 207844 84710 207900
rect 73546 207732 73556 207788
rect 73612 207732 78036 207788
rect 78092 207732 78102 207788
rect 72202 207620 72212 207676
rect 72268 207620 84756 207676
rect 84812 207620 84822 207676
rect 671552 207620 690116 207676
rect 690172 207620 690182 207676
rect 560410 206612 560420 206668
rect 560476 206612 611744 206668
rect 559850 206164 559860 206220
rect 559916 206164 559926 206220
rect 559860 205632 559916 206164
rect 671552 205268 696276 205324
rect 696332 205268 696342 205324
rect 570602 204372 570612 204428
rect 570668 204372 611744 204428
rect 701418 203588 701428 203644
rect 701484 203588 705732 203644
rect 705788 203588 705798 203644
rect 701642 203476 701652 203532
rect 701708 203476 704836 203532
rect 704892 203476 704902 203532
rect 703882 203364 703892 203420
rect 703948 203364 705284 203420
rect 705340 203364 705350 203420
rect 701866 203252 701876 203308
rect 701932 203252 704388 203308
rect 704444 203252 704454 203308
rect 560308 202076 560364 202720
rect 560308 202020 565236 202076
rect 565292 202020 565302 202076
rect 570490 202020 570500 202076
rect 570556 202020 611744 202076
rect 671552 200676 690228 200732
rect 690284 200676 690294 200732
rect 560308 199164 560364 199808
rect 570266 199780 570276 199836
rect 570332 199780 611744 199836
rect 560308 199108 566916 199164
rect 566972 199108 566982 199164
rect 671552 198436 695044 198492
rect 695100 198436 695110 198492
rect 570378 197540 570388 197596
rect 570444 197540 611744 197596
rect 560336 196756 560868 196812
rect 560924 196756 560934 196812
rect 701642 196196 701652 196252
rect 701708 196196 704564 196252
rect 704620 196196 704630 196252
rect 703854 196084 703892 196140
rect 703948 196084 703958 196140
rect 701866 195972 701876 196028
rect 701932 195972 705012 196028
rect 705068 195972 705078 196028
rect 705674 195412 705684 195468
rect 705788 195412 705798 195468
rect 560858 195188 560868 195244
rect 560924 195188 611744 195244
rect 560336 193844 560644 193900
rect 560700 193844 560710 193900
rect 671552 193732 694932 193788
rect 694988 193732 694998 193788
rect 560746 192948 560756 193004
rect 560812 192948 611744 193004
rect 75936 191900 76132 191956
rect 76188 191900 76198 191956
rect 75936 191452 76132 191508
rect 76188 191452 76198 191508
rect 671552 191492 695156 191548
rect 695212 191492 695222 191548
rect 560074 191380 560084 191436
rect 560140 191380 560150 191436
rect 90318 191268 90356 191324
rect 90412 191268 90422 191324
rect 75992 191004 76468 191060
rect 76524 191004 76534 191060
rect 84270 190932 84308 190988
rect 84364 190932 84374 190988
rect 560084 190960 560140 191380
rect 560634 190708 560644 190764
rect 560700 190708 611744 190764
rect 76356 190612 83860 190652
rect 75936 190596 83860 190612
rect 83916 190596 83926 190652
rect 75936 190556 76412 190596
rect 75936 189212 76132 189268
rect 76188 189212 76198 189268
rect 75936 188764 76244 188820
rect 76300 188764 76310 188820
rect 571946 188468 571956 188524
rect 572012 188468 611744 188524
rect 560308 187292 560364 188048
rect 560308 187236 561147 187292
rect 561091 186508 561147 187236
rect 671552 186900 695156 186956
rect 695212 186900 695222 186956
rect 561091 186452 578676 186508
rect 578732 186452 578742 186508
rect 559290 186116 559300 186172
rect 559356 186116 611744 186172
rect 559626 185668 559636 185724
rect 559692 185668 560308 185724
rect 560364 185668 560374 185724
rect 560336 184996 560980 185052
rect 561036 184996 561046 185052
rect 671552 184548 697956 184604
rect 698012 184548 698022 184604
rect 605546 183876 605556 183932
rect 605612 183876 611744 183932
rect 560298 182980 560308 183036
rect 560364 182980 560532 183036
rect 560588 182980 560598 183036
rect 560308 181468 560364 182112
rect 560522 181636 560532 181692
rect 560588 181636 611744 181692
rect 560308 181412 568596 181468
rect 568652 181412 568662 181468
rect 694586 180180 694596 180236
rect 694652 180180 702016 180236
rect 671552 179956 694820 180012
rect 694876 179956 694886 180012
rect 693018 179732 693028 179788
rect 693084 179732 702016 179788
rect 585610 179284 585620 179340
rect 585676 179284 611744 179340
rect 560308 178556 560364 179200
rect 701876 178836 702016 178892
rect 560308 178500 568708 178556
rect 568764 178500 568774 178556
rect 701876 178444 701932 178836
rect 701876 178388 702016 178444
rect 696154 177940 696164 177996
rect 696220 177940 702016 177996
rect 671552 177604 695044 177660
rect 695100 177604 695110 177660
rect 690451 177492 702016 177548
rect 603866 177044 603876 177100
rect 603932 177044 611744 177100
rect 690451 176652 690507 177492
rect 689546 176596 689556 176652
rect 689612 176596 690507 176652
rect 696276 177044 702016 177100
rect 696276 176540 696332 177044
rect 686634 176484 686644 176540
rect 686700 176484 696332 176540
rect 559290 176372 559300 176428
rect 559356 176372 559366 176428
rect 686410 176372 686420 176428
rect 686476 176372 696164 176428
rect 696220 176372 696230 176428
rect 559300 176288 559356 176372
rect 605658 174804 605668 174860
rect 605724 174804 611744 174860
rect 560308 173796 560420 173852
rect 560476 173796 560486 173852
rect 560308 173264 560364 173796
rect 671552 173012 694932 173068
rect 694988 173012 694998 173068
rect 73770 172900 73780 172956
rect 73836 172900 77364 172956
rect 77420 172900 77430 172956
rect 72986 172788 72996 172844
rect 73052 172788 77476 172844
rect 77532 172788 77542 172844
rect 73098 172676 73108 172732
rect 73164 172676 78148 172732
rect 78204 172676 78214 172732
rect 72202 172564 72212 172620
rect 72268 172564 77588 172620
rect 77644 172564 77654 172620
rect 561866 172564 561876 172620
rect 561932 172564 611744 172620
rect 671552 170660 689556 170716
rect 689612 170660 689622 170716
rect 560308 169708 560364 170352
rect 603978 170212 603988 170268
rect 604044 170212 611744 170268
rect 560308 169652 570612 169708
rect 570668 169652 570678 169708
rect 560410 167972 560420 168028
rect 560476 167972 611744 168028
rect 560308 166796 560364 167440
rect 560308 166740 570500 166796
rect 570556 166740 570566 166796
rect 671552 166068 694596 166124
rect 694652 166068 694662 166124
rect 585834 165732 585844 165788
rect 585900 165732 611744 165788
rect 560308 163884 560364 164528
rect 560308 163828 570276 163884
rect 570332 163828 570342 163884
rect 671552 163828 694708 163884
rect 694764 163828 694774 163884
rect 586058 163380 586068 163436
rect 586124 163380 611744 163436
rect 560308 161308 560364 161504
rect 671552 161476 671748 161532
rect 671804 161476 671814 161532
rect 560308 161252 570388 161308
rect 570444 161252 570454 161308
rect 600618 161140 600628 161196
rect 600684 161140 611744 161196
rect 704974 160804 705012 160860
rect 705068 160804 705078 160860
rect 702090 160356 702100 160412
rect 702156 160356 704836 160412
rect 704892 160356 704902 160412
rect 704378 160244 704388 160300
rect 704444 160244 705236 160300
rect 705292 160244 705302 160300
rect 701978 159684 701988 159740
rect 702044 159684 705572 159740
rect 705628 159684 705638 159740
rect 671552 159124 700532 159180
rect 700588 159124 700598 159180
rect 585386 158900 585396 158956
rect 585452 158900 611744 158956
rect 560336 158564 560868 158620
rect 560924 158564 560934 158620
rect 671552 156884 694596 156940
rect 694652 156884 694662 156940
rect 565226 156660 565236 156716
rect 565292 156660 611744 156716
rect 560336 155652 560756 155708
rect 560812 155652 560822 155708
rect 671552 154532 671748 154588
rect 671804 154532 671814 154588
rect 560298 154308 560308 154364
rect 560364 154308 611744 154364
rect 560336 152740 560644 152796
rect 560700 152740 560710 152796
rect 704378 152740 704388 152796
rect 704444 152740 705012 152796
rect 705068 152740 705078 152796
rect 705226 152740 705236 152796
rect 705340 152740 705350 152796
rect 702090 152516 702100 152572
rect 702156 152516 704836 152572
rect 704892 152516 704902 152572
rect 705674 152404 705684 152460
rect 705788 152404 705798 152460
rect 671552 152292 671748 152348
rect 671804 152292 671814 152348
rect 575306 152068 575316 152124
rect 575372 152068 611744 152124
rect 671552 149940 671860 149996
rect 671916 149940 671926 149996
rect 598826 149828 598836 149884
rect 598892 149828 611744 149884
rect 560308 149548 560364 149744
rect 560308 149492 571956 149548
rect 572012 149492 572022 149548
rect 671552 147588 672756 147644
rect 672812 147588 672822 147644
rect 585610 147476 585620 147532
rect 585676 147476 611744 147532
rect 559290 147364 559300 147420
rect 559356 147364 559366 147420
rect 559300 146832 559356 147364
rect 671552 145348 671860 145404
rect 671916 145348 671926 145404
rect 585834 145236 585844 145292
rect 585900 145236 611744 145292
rect 559412 143388 559468 143920
rect 559402 143332 559412 143388
rect 559468 143332 559478 143388
rect 585162 142996 585172 143052
rect 585228 142996 611744 143052
rect 671552 142996 672196 143052
rect 672252 142996 672262 143052
rect 671738 142660 671748 142716
rect 671804 142660 673540 142716
rect 673596 142660 673606 142716
rect 671822 142100 671860 142156
rect 671916 142100 671926 142156
rect 559374 141652 559412 141708
rect 559468 141652 559478 141708
rect 671934 141540 671972 141596
rect 672028 141540 672038 141596
rect 671710 141092 671748 141148
rect 671804 141092 671814 141148
rect 560308 140364 560364 141008
rect 611492 140756 611744 140812
rect 671552 140756 672084 140812
rect 672140 140756 672150 140812
rect 560308 140308 567867 140364
rect 567811 139468 567867 140308
rect 611492 140140 611548 140756
rect 611492 140084 611716 140140
rect 611772 140084 611782 140140
rect 619891 140084 624036 140140
rect 624092 140084 624102 140140
rect 619891 140028 619947 140084
rect 619098 139972 619108 140028
rect 619164 139972 619947 140028
rect 623326 139972 623364 140028
rect 623420 139972 623430 140028
rect 624670 139972 624708 140028
rect 624764 139972 624774 140028
rect 657038 139972 657076 140028
rect 657132 139972 657142 140028
rect 657710 139972 657748 140028
rect 657804 139972 657814 140028
rect 618874 139860 618884 139916
rect 618940 139860 630756 139916
rect 630812 139860 630822 139916
rect 631390 139860 631428 139916
rect 631484 139860 631494 139916
rect 655694 139860 655732 139916
rect 655788 139860 655798 139916
rect 665130 139860 665140 139916
rect 665196 139860 671188 139916
rect 671244 139860 671254 139916
rect 618202 139748 618212 139804
rect 618268 139748 622692 139804
rect 622748 139748 622758 139804
rect 659082 139748 659092 139804
rect 659148 139748 669956 139804
rect 670012 139748 670022 139804
rect 621982 139636 622020 139692
rect 622076 139636 622086 139692
rect 632734 139636 632772 139692
rect 632828 139636 632838 139692
rect 638782 139636 638820 139692
rect 638876 139636 638886 139692
rect 650654 139636 650692 139692
rect 650748 139636 650758 139692
rect 656366 139636 656404 139692
rect 656460 139636 656470 139692
rect 666446 139636 666484 139692
rect 666540 139636 666550 139692
rect 667818 139636 667828 139692
rect 667884 139636 670404 139692
rect 670460 139636 670470 139692
rect 618650 139524 618660 139580
rect 618716 139524 624932 139580
rect 624988 139524 624998 139580
rect 659978 139524 659988 139580
rect 660044 139524 670068 139580
rect 670124 139524 670134 139580
rect 567811 139412 605556 139468
rect 605612 139412 605622 139468
rect 618538 139412 618548 139468
rect 618604 139412 619108 139468
rect 619164 139412 619174 139468
rect 619882 139412 619892 139468
rect 619948 139412 621460 139468
rect 621516 139412 621526 139468
rect 648442 139412 648452 139468
rect 648508 139412 649012 139468
rect 649068 139412 649078 139468
rect 650794 139412 650804 139468
rect 650860 139412 658420 139468
rect 658476 139412 658486 139468
rect 669610 139412 669620 139468
rect 669676 139412 670852 139468
rect 670908 139412 670918 139468
rect 664458 138964 664468 139020
rect 664524 138964 670964 139020
rect 671020 138964 671030 139020
rect 663786 138740 663796 138796
rect 663852 138740 670740 138796
rect 670796 138740 670806 138796
rect 559290 138516 559300 138572
rect 559356 138516 559366 138572
rect 559300 137984 559356 138516
rect 660426 137956 660436 138012
rect 660492 137956 669620 138012
rect 669676 137956 669686 138012
rect 662442 137844 662452 137900
rect 662508 137844 669844 137900
rect 669900 137844 669910 137900
rect 661770 137732 661780 137788
rect 661836 137732 669732 137788
rect 669788 137732 669798 137788
rect 701316 137228 702016 137236
rect 700522 137172 700532 137228
rect 700588 137180 702016 137228
rect 700588 137172 701372 137180
rect 663450 136948 663460 137004
rect 663516 136948 670404 137004
rect 670460 136948 670470 137004
rect 661546 136836 661556 136892
rect 661612 136836 670292 136892
rect 670348 136836 670358 136892
rect 701316 136780 702016 136788
rect 694810 136724 694820 136780
rect 694876 136732 702016 136780
rect 694876 136724 701372 136732
rect 649422 136276 649460 136332
rect 649516 136276 649526 136332
rect 649786 136276 649796 136332
rect 649852 136276 653716 136332
rect 653772 136276 653782 136332
rect 649898 136164 649908 136220
rect 649964 136164 655060 136220
rect 655116 136164 655126 136220
rect 650010 136052 650020 136108
rect 650076 136052 654388 136108
rect 654444 136052 654454 136108
rect 560186 135604 560196 135660
rect 560252 135604 560262 135660
rect 622346 135604 622356 135660
rect 622412 135604 636132 135660
rect 636188 135604 636198 135660
rect 560196 135072 560252 135604
rect 622234 135492 622244 135548
rect 622300 135492 638148 135548
rect 638204 135492 638214 135548
rect 669946 135492 669956 135548
rect 670012 135492 670022 135548
rect 622794 135380 622804 135436
rect 622860 135380 635460 135436
rect 635516 135380 635526 135436
rect 622682 135268 622692 135324
rect 622748 135268 637476 135324
rect 637532 135268 637542 135324
rect 669956 135212 670012 135492
rect 701316 135436 702016 135444
rect 700522 135380 700532 135436
rect 700588 135388 702016 135436
rect 700588 135380 701372 135388
rect 622570 135156 622580 135212
rect 622636 135156 636804 135212
rect 636860 135156 636870 135212
rect 669610 135156 669620 135212
rect 669676 135156 669686 135212
rect 669946 135156 669956 135212
rect 670012 135156 670022 135212
rect 669620 135100 669676 135156
rect 669620 135044 669844 135100
rect 669900 135044 669910 135100
rect 669498 134932 669508 134988
rect 669564 134932 669620 134988
rect 669676 134932 669686 134988
rect 701316 134940 702016 134996
rect 701316 134876 701372 134940
rect 650010 134820 650020 134876
rect 650076 134820 650132 134876
rect 650188 134820 650198 134876
rect 690451 134820 701372 134876
rect 618314 134596 618324 134652
rect 618380 134596 621348 134652
rect 621404 134596 621414 134652
rect 620442 134484 620452 134540
rect 620508 134484 621460 134540
rect 621516 134484 621526 134540
rect 690451 134428 690507 134820
rect 701428 134540 702016 134548
rect 694698 134484 694708 134540
rect 694764 134492 702016 134540
rect 694764 134484 701484 134492
rect 618398 134372 618436 134428
rect 618492 134372 618502 134428
rect 621114 134372 621124 134428
rect 621180 134372 621348 134428
rect 621404 134372 621414 134428
rect 686186 134372 686196 134428
rect 686252 134372 690507 134428
rect 701418 134044 701428 134100
rect 701484 134044 702016 134100
rect 650122 133140 650132 133196
rect 650188 133140 650198 133196
rect 650131 133084 650187 133140
rect 650112 133028 650122 133084
rect 650178 133028 650188 133084
rect 649450 132692 649460 132748
rect 649516 132692 649572 132748
rect 649628 132692 649638 132748
rect 686970 132692 686980 132748
rect 687036 132692 701428 132748
rect 701484 132692 701494 132748
rect 650010 132580 650020 132636
rect 650076 132580 654378 132636
rect 654434 132580 654444 132636
rect 655171 132580 656394 132636
rect 656450 132580 656460 132636
rect 657934 132580 657972 132636
rect 658028 132580 658038 132636
rect 664542 132580 664580 132636
rect 664636 132580 664646 132636
rect 666810 132580 666820 132636
rect 666876 132580 666922 132636
rect 666978 132580 666988 132636
rect 667584 132580 667594 132636
rect 667650 132580 669620 132636
rect 669676 132580 669686 132636
rect 670170 132580 670180 132636
rect 670236 132580 670852 132636
rect 670908 132580 670918 132636
rect 649898 132468 649908 132524
rect 649964 132468 654836 132524
rect 654892 132468 654902 132524
rect 655171 132412 655227 132580
rect 659614 132468 659652 132524
rect 659708 132468 659718 132524
rect 661984 132468 661994 132524
rect 662050 132468 666987 132524
rect 668256 132468 668266 132524
rect 668322 132468 670516 132524
rect 670572 132468 670582 132524
rect 650654 132356 650692 132412
rect 650748 132356 650758 132412
rect 650906 132356 650916 132412
rect 650972 132356 655227 132412
rect 666931 132412 666987 132468
rect 666931 132356 669732 132412
rect 669788 132356 669798 132412
rect 649226 132244 649236 132300
rect 649292 132244 651578 132300
rect 651634 132244 651644 132300
rect 653716 132244 655722 132300
rect 655778 132244 655788 132300
rect 660640 132244 660650 132300
rect 660706 132244 669844 132300
rect 669900 132244 669910 132300
rect 560308 131516 560364 132160
rect 649114 132132 649124 132188
rect 649180 132132 652250 132188
rect 652306 132132 652316 132188
rect 653482 132132 653492 132188
rect 653548 132132 653594 132188
rect 653650 132132 653660 132188
rect 648890 132020 648900 132076
rect 648956 132020 652922 132076
rect 652978 132020 652988 132076
rect 653716 131964 653772 132244
rect 649674 131908 649684 131964
rect 649740 131908 653772 131964
rect 653828 132132 657178 132188
rect 657234 132132 657244 132188
rect 661312 132132 661322 132188
rect 661378 132132 670292 132188
rect 670348 132132 670358 132188
rect 653828 131852 653884 132132
rect 611482 131796 611492 131852
rect 611548 131796 612164 131852
rect 612220 131796 612230 131852
rect 649562 131796 649572 131852
rect 649628 131796 653884 131852
rect 655171 132020 657850 132076
rect 657906 132020 657916 132076
rect 668928 132020 668938 132076
rect 668994 132020 671524 132076
rect 671580 132020 671590 132076
rect 655171 131740 655227 132020
rect 665914 131908 665924 131964
rect 665980 131908 671188 131964
rect 671244 131908 671254 131964
rect 663450 131796 663460 131852
rect 663516 131796 670404 131852
rect 670460 131796 670470 131852
rect 649338 131684 649348 131740
rect 649404 131684 655227 131740
rect 666586 131684 666596 131740
rect 666652 131684 671636 131740
rect 671692 131684 671702 131740
rect 648330 131572 648340 131628
rect 648396 131572 654724 131628
rect 654780 131572 654790 131628
rect 560308 131460 561147 131516
rect 660090 131460 660100 131516
rect 660156 131460 670180 131516
rect 670236 131460 670246 131516
rect 561091 131068 561147 131460
rect 663226 131348 663236 131404
rect 663292 131348 670068 131404
rect 670124 131348 670134 131404
rect 561091 131012 605668 131068
rect 605724 131012 605734 131068
rect 665102 131012 665140 131068
rect 665196 131012 665206 131068
rect 560308 128604 560364 129248
rect 560308 128548 561147 128604
rect 561091 127708 561147 128548
rect 561091 127652 603876 127708
rect 603932 127652 603942 127708
rect 643626 127540 643636 127596
rect 643692 127540 654500 127596
rect 654556 127540 654566 127596
rect 646286 127428 646324 127484
rect 646380 127428 646390 127484
rect 645642 127204 645652 127260
rect 645708 127204 655396 127260
rect 655452 127204 655462 127260
rect 644970 126980 644980 127036
rect 645036 126980 655172 127036
rect 655228 126980 655238 127036
rect 644298 126868 644308 126924
rect 644364 126868 655284 126924
rect 655340 126868 655350 126924
rect 642282 126756 642292 126812
rect 642348 126756 654276 126812
rect 654332 126756 654342 126812
rect 655918 126644 655956 126700
rect 656012 126644 656022 126700
rect 559300 126028 559356 126224
rect 559290 125972 559300 126028
rect 559356 125972 559366 126028
rect 646958 125972 646996 126028
rect 647052 125972 647062 126028
rect 647658 125972 647668 126028
rect 647724 125972 655620 126028
rect 655676 125972 655686 126028
rect 626014 125860 626052 125916
rect 626108 125860 626118 125916
rect 628030 125860 628068 125916
rect 628124 125860 628134 125916
rect 628702 125860 628740 125916
rect 628796 125860 628806 125916
rect 641470 125860 641508 125916
rect 641564 125860 641574 125916
rect 642954 125748 642964 125804
rect 643020 125748 654612 125804
rect 654668 125748 654678 125804
rect 640826 125636 640836 125692
rect 640892 125636 655956 125692
rect 656012 125636 656022 125692
rect 640154 125524 640164 125580
rect 640220 125524 655844 125580
rect 655900 125524 655910 125580
rect 619098 125412 619108 125468
rect 619164 125412 630084 125468
rect 630140 125412 630150 125468
rect 639482 125412 639492 125468
rect 639548 125412 655732 125468
rect 655788 125412 655798 125468
rect 629402 125300 629412 125356
rect 629468 125300 655284 125356
rect 655340 125300 655350 125356
rect 627386 125188 627396 125244
rect 627452 125188 654948 125244
rect 655004 125188 655014 125244
rect 626714 125076 626724 125132
rect 626780 125076 655060 125132
rect 655116 125076 655126 125132
rect 670142 123508 670180 123564
rect 670236 123508 670246 123564
rect 620554 123396 620564 123452
rect 620620 123396 627284 123452
rect 627340 123396 627350 123452
rect 560308 122668 560364 123312
rect 620330 123284 620340 123340
rect 620396 123284 622132 123340
rect 622188 123284 622198 123340
rect 641162 123284 641172 123340
rect 641228 123284 642740 123340
rect 642796 123284 642806 123340
rect 647854 123284 647892 123340
rect 647948 123284 647958 123340
rect 654948 122892 655004 123088
rect 654938 122836 654948 122892
rect 655004 122836 655014 122892
rect 560308 122612 603988 122668
rect 604044 122612 604054 122668
rect 618650 122612 618660 122668
rect 618716 122612 618772 122668
rect 618828 122612 618838 122668
rect 655274 121492 655284 121548
rect 655340 121492 655350 121548
rect 655284 121296 655340 121492
rect 655274 120596 655284 120652
rect 655340 120596 655732 120652
rect 655788 120596 655798 120652
rect 560336 120372 561876 120428
rect 561932 120372 561942 120428
rect 655386 119812 655396 119868
rect 655452 119812 655462 119868
rect 655396 119616 655452 119812
rect 655386 118916 655396 118972
rect 655452 118916 655844 118972
rect 655900 118916 655910 118972
rect 655050 118356 655060 118412
rect 655116 118356 655126 118412
rect 655060 117824 655116 118356
rect 701642 118020 701652 118076
rect 701708 118020 704836 118076
rect 704892 118020 704902 118076
rect 704666 117796 704676 117852
rect 704732 117796 704900 117852
rect 704956 117796 704966 117852
rect 701866 117684 701876 117740
rect 701932 117684 705572 117740
rect 705628 117684 705638 117740
rect 703994 117572 704004 117628
rect 704060 117572 705012 117628
rect 705068 117572 705078 117628
rect 560336 117460 560532 117516
rect 560588 117460 560598 117516
rect 654938 116564 654948 116620
rect 655004 116564 655014 116620
rect 654948 116032 655004 116564
rect 655050 114996 655060 115052
rect 655116 114996 655126 115052
rect 559300 114268 559356 114464
rect 655060 114352 655116 114996
rect 559290 114212 559300 114268
rect 559356 114212 559366 114268
rect 654938 113204 654948 113260
rect 655004 113204 655014 113260
rect 654948 112560 655004 113204
rect 559300 110908 559356 111552
rect 655508 111076 655620 111132
rect 655676 111076 655686 111132
rect 559290 110852 559300 110908
rect 559356 110852 559366 110908
rect 655508 110880 655564 111076
rect 651914 110180 651924 110236
rect 651980 110180 655396 110236
rect 655452 110180 655462 110236
rect 703966 110068 704004 110124
rect 704060 110068 704070 110124
rect 704890 110068 704900 110124
rect 704956 110068 705012 110124
rect 705068 110068 705078 110124
rect 701642 109956 701652 110012
rect 701708 109956 704564 110012
rect 704620 109956 704630 110012
rect 652922 109620 652932 109676
rect 652988 109620 655284 109676
rect 655340 109620 655350 109676
rect 705674 109396 705684 109452
rect 705788 109396 705798 109452
rect 560308 107884 560364 108640
rect 560308 107828 561147 107884
rect 561091 107548 561147 107828
rect 561091 107492 600628 107548
rect 600684 107492 600694 107548
rect 559300 105196 559356 105728
rect 559290 105140 559300 105196
rect 559356 105140 559366 105196
rect 560308 102508 560364 102704
rect 560308 102452 575316 102508
rect 575372 102452 575382 102508
rect 619882 100660 619892 100716
rect 619948 100660 620564 100716
rect 620620 100660 620630 100716
rect 622346 100660 622356 100716
rect 622412 100660 625380 100716
rect 625436 100660 625446 100716
rect 647546 100660 647556 100716
rect 647612 100660 654724 100716
rect 654780 100660 654790 100716
rect 619770 100548 619780 100604
rect 619836 100548 619846 100604
rect 560298 100324 560308 100380
rect 560364 100324 560374 100380
rect 560308 99792 560364 100324
rect 619780 99904 619836 100548
rect 622794 100436 622804 100492
rect 622860 100436 623364 100492
rect 623420 100436 623430 100492
rect 628590 100436 628628 100492
rect 628684 100436 628694 100492
rect 631166 100436 631204 100492
rect 631260 100436 631270 100492
rect 649534 100436 649572 100492
rect 649628 100436 649638 100492
rect 652138 100436 652148 100492
rect 652204 100436 654612 100492
rect 654668 100436 654678 100492
rect 633742 99988 633780 100044
rect 633836 99988 633846 100044
rect 635758 99988 635796 100044
rect 635852 99988 635862 100044
rect 639006 99988 639044 100044
rect 639100 99988 639110 100044
rect 641694 99988 641732 100044
rect 641788 99988 641798 100044
rect 644942 99988 644980 100044
rect 645036 99988 645046 100044
rect 619546 98980 619556 99036
rect 619612 98980 619724 99036
rect 619668 98672 619724 98980
rect 653520 98868 654500 98924
rect 654556 98868 654566 98924
rect 619322 97412 619332 97468
rect 619388 97412 619696 97468
rect 560308 96236 560364 96880
rect 560308 96180 565236 96236
rect 565292 96180 565302 96236
rect 618986 96180 618996 96236
rect 619052 96180 619696 96236
rect 652922 95620 652932 95676
rect 652988 95620 652998 95676
rect 652932 95536 652988 95620
rect 619098 94948 619108 95004
rect 619164 94948 619696 95004
rect 701316 94180 702016 94236
rect 701316 94108 701372 94180
rect 673530 94052 673540 94108
rect 673596 94052 701372 94108
rect 560308 93324 560364 93968
rect 618874 93716 618884 93772
rect 618940 93716 619696 93772
rect 701418 93732 701428 93788
rect 701484 93732 702016 93788
rect 560308 93268 561147 93324
rect 561091 92428 561147 93268
rect 619098 92484 619108 92540
rect 619164 92484 619696 92540
rect 694586 92484 694596 92540
rect 694652 92484 701708 92540
rect 701652 92444 701708 92484
rect 561091 92372 598836 92428
rect 598892 92372 598902 92428
rect 686522 92372 686532 92428
rect 686588 92372 701428 92428
rect 701484 92372 701494 92428
rect 701652 92388 702016 92444
rect 653520 92260 655172 92316
rect 655228 92260 655238 92316
rect 701418 91940 701428 91996
rect 701484 91940 702016 91996
rect 701316 91532 702016 91548
rect 694586 91476 694596 91532
rect 694652 91492 702016 91532
rect 694652 91476 701372 91492
rect 618538 91252 618548 91308
rect 618604 91252 619696 91308
rect 701316 91044 702016 91100
rect 559300 90748 559356 90944
rect 701316 90860 701372 91044
rect 686522 90804 686532 90860
rect 686588 90804 701372 90860
rect 559290 90692 559300 90748
rect 559356 90692 559366 90748
rect 686298 90692 686308 90748
rect 686364 90692 701428 90748
rect 701484 90692 701494 90748
rect 618314 89908 618324 89964
rect 618380 89908 619696 89964
rect 652922 89012 652932 89068
rect 652988 89012 652998 89068
rect 652932 88928 652988 89012
rect 618650 88676 618660 88732
rect 618716 88676 619696 88732
rect 559300 87500 559356 88032
rect 559290 87444 559300 87500
rect 559356 87444 559366 87500
rect 618874 87444 618884 87500
rect 618940 87444 619696 87500
rect 618426 86212 618436 86268
rect 618492 86212 619696 86268
rect 653520 85540 655956 85596
rect 656012 85540 656022 85596
rect 559300 84476 559356 85120
rect 618314 84980 618324 85036
rect 618380 84980 619696 85036
rect 559290 84420 559300 84476
rect 559356 84420 559366 84476
rect 618202 83748 618212 83804
rect 618268 83748 619696 83804
rect 672186 83412 672196 83468
rect 672252 83412 672980 83468
rect 673036 83412 673046 83468
rect 652922 82964 652932 83020
rect 652988 82964 652998 83020
rect 618650 82516 618660 82572
rect 618716 82516 619696 82572
rect 652932 82320 652988 82964
rect 560308 81900 560364 82208
rect 560298 81844 560308 81900
rect 560364 81844 560374 81900
rect 559290 81732 559300 81788
rect 559356 81732 585172 81788
rect 585228 81732 585238 81788
rect 558506 81620 558516 81676
rect 558572 81620 559412 81676
rect 559468 81620 559478 81676
rect 561091 81620 585396 81676
rect 585452 81620 585462 81676
rect 561091 81564 561147 81620
rect 558282 81508 558292 81564
rect 558348 81508 561147 81564
rect 559066 81396 559076 81452
rect 559132 81396 586068 81452
rect 586124 81396 586134 81452
rect 558954 81284 558964 81340
rect 559020 81284 585844 81340
rect 585900 81284 585910 81340
rect 618538 81284 618548 81340
rect 618604 81284 619696 81340
rect 558730 81172 558740 81228
rect 558796 81172 585620 81228
rect 585676 81172 585686 81228
rect 92334 80836 92372 80892
rect 92428 80836 92438 80892
rect 335934 80724 335972 80780
rect 336028 80724 336038 80780
rect 628030 80612 628068 80668
rect 628124 80612 628134 80668
rect 645054 80612 645092 80668
rect 645148 80612 645158 80668
rect 93818 79044 93828 79100
rect 93884 79044 190596 79100
rect 190652 79044 560196 79100
rect 560252 79044 560262 79100
rect 123498 78932 123508 78988
rect 123564 78932 561876 78988
rect 561932 78932 561942 78988
rect 671962 74452 671972 74508
rect 672028 74452 705284 74508
rect 705340 74452 705350 74508
rect 672074 74228 672084 74284
rect 672140 74228 704836 74284
rect 704892 74228 704902 74284
rect 672746 74004 672756 74060
rect 672812 74004 704340 74060
rect 704396 74004 704406 74060
rect 672970 73892 672980 73948
rect 673036 73892 705684 73948
rect 705740 73892 705750 73948
rect 324846 72100 324884 72156
rect 324940 72100 324950 72156
rect 526362 72100 526372 72156
rect 526428 72100 560980 72156
rect 561036 72100 561046 72156
rect 459162 71988 459172 72044
rect 459228 71988 559412 72044
rect 559468 71988 559478 72044
rect 506762 71876 506772 71932
rect 506828 71876 617316 71932
rect 617372 71876 617382 71932
rect 392074 71764 392084 71820
rect 392140 71764 548548 71820
rect 548604 71764 548614 71820
rect 454570 71652 454580 71708
rect 454636 71652 614628 71708
rect 614684 71652 614694 71708
rect 396106 71540 396116 71596
rect 396172 71540 611492 71596
rect 611548 71540 611558 71596
rect 341674 71428 341684 71484
rect 341740 71428 613956 71484
rect 614012 71428 614022 71484
rect 231242 71316 231252 71372
rect 231308 71316 620564 71372
rect 620620 71316 620630 71372
rect 619294 71092 619332 71148
rect 619388 71092 619398 71148
rect 617950 70980 617988 71036
rect 618044 70980 618054 71036
rect 257758 70532 257796 70588
rect 257852 70532 257862 70588
rect 396026 70532 396036 70588
rect 396092 70532 396116 70588
rect 396172 70532 396182 70588
rect 559402 70532 559412 70588
rect 559468 70532 560890 70588
rect 560946 70532 560956 70588
rect 539130 70308 539140 70364
rect 539196 70308 549287 70364
rect 549343 70308 549353 70364
rect 176172 70084 176182 70140
rect 176238 70084 176260 70140
rect 176316 70084 176326 70140
rect 231172 70084 231182 70140
rect 231238 70084 231252 70140
rect 231308 70084 231318 70140
rect 451171 70084 451181 70140
rect 451237 70084 454580 70140
rect 454636 70084 454646 70140
rect 494277 70084 494287 70140
rect 494396 70084 494406 70140
rect 505866 70084 505876 70140
rect 505946 70084 505970 70140
rect 548422 70084 548432 70140
rect 548492 70084 548526 70140
rect 450880 69748 450890 69804
rect 450946 69748 469140 69804
rect 469196 69748 469206 69804
rect 506026 69748 506036 69804
rect 506092 69748 519652 69804
rect 519708 69748 519718 69804
<< via3 >>
rect 470260 949172 470316 949228
rect 106596 947732 106652 947788
rect 216580 947732 216636 947788
rect 271572 947732 271628 947788
rect 470260 947732 470316 947788
rect 525700 947732 525756 947788
rect 690340 947732 690396 947788
rect 251188 947604 251244 947660
rect 306068 947604 306124 947660
rect 361396 947492 361452 947548
rect 545860 947492 545916 947548
rect 581140 947492 581196 947548
rect 655844 947492 655900 947548
rect 697956 947492 698012 947548
rect 525588 947284 525644 947340
rect 690340 947284 690396 947340
rect 361284 947156 361340 947212
rect 581252 947156 581308 947212
rect 545860 947044 545916 947100
rect 655844 947044 655900 947100
rect 471268 946836 471324 946892
rect 545636 946836 545692 946892
rect 655620 946836 655676 946892
rect 692916 946820 692972 946876
rect 196084 946708 196140 946764
rect 251076 946708 251132 946764
rect 361172 946708 361228 946764
rect 526148 946708 526204 946764
rect 581028 946708 581084 946764
rect 75460 945924 75516 945980
rect 525700 946388 525756 946444
rect 545524 946388 545580 946444
rect 655508 946388 655564 946444
rect 581140 946260 581196 946316
rect 471268 945924 471324 945980
rect 704004 945812 704060 945868
rect 75460 945700 75516 945756
rect 121940 943348 121996 943404
rect 122388 943348 122444 943404
rect 289828 943348 289884 943404
rect 341236 943348 341292 943404
rect 342692 943348 342748 943404
rect 454244 943460 454300 943516
rect 561316 943348 561372 943404
rect 233492 943236 233548 943292
rect 564900 943348 564956 943404
rect 670292 943348 670348 943404
rect 565012 943236 565068 943292
rect 121940 942676 121996 942732
rect 85428 942564 85484 942620
rect 122388 942564 122444 942620
rect 106596 942340 106652 942396
rect 216580 942340 216636 942396
rect 306068 942340 306124 942396
rect 334292 942340 334348 942396
rect 361172 942340 361228 942396
rect 251188 942228 251244 942284
rect 271572 942228 271628 942284
rect 361396 942228 361452 942284
rect 251076 942116 251132 942172
rect 334292 942116 334348 942172
rect 361284 942116 361340 942172
rect 196084 942004 196140 942060
rect 282436 937412 282492 937468
rect 688212 937300 688268 937356
rect 687428 937188 687484 937244
rect 285684 937076 285740 937132
rect 141876 936964 141932 937020
rect 178724 936964 178780 937020
rect 688436 936964 688492 937020
rect 141652 936740 141708 936796
rect 141428 936628 141484 936684
rect 687988 936516 688044 936572
rect 688884 936404 688940 936460
rect 689332 936292 689388 936348
rect 84084 935732 84140 935788
rect 84308 935732 84364 935788
rect 84532 935732 84588 935788
rect 85428 935620 85484 935676
rect 587524 935620 587580 935676
rect 695380 935508 695436 935564
rect 694260 935284 694316 935340
rect 233492 935172 233548 935228
rect 694036 935060 694092 935116
rect 694932 934948 694988 935004
rect 341012 934836 341068 934892
rect 458500 934836 458556 934892
rect 686308 934836 686364 934892
rect 686980 934388 687036 934444
rect 686756 934276 686812 934332
rect 700532 934164 700588 934220
rect 76132 929900 76188 929956
rect 83748 929796 83804 929852
rect 76356 929452 76412 929508
rect 76132 929004 76188 929060
rect 78932 927332 78988 927388
rect 76244 927212 76300 927268
rect 704004 927220 704060 927276
rect 703892 927108 703948 927164
rect 84644 926884 84700 926940
rect 76356 926764 76412 926820
rect 704788 926324 704836 926380
rect 704836 926324 704844 926380
rect 705684 926324 705732 926380
rect 705732 926324 705740 926380
rect 697732 925092 697788 925148
rect 700532 908964 700588 909020
rect 76020 897092 76076 897148
rect 704788 840308 704836 840364
rect 704836 840308 704844 840364
rect 705124 840308 705180 840364
rect 705684 840308 705732 840364
rect 705732 840308 705740 840364
rect 700420 838292 700476 838348
rect 700644 838292 700700 838348
rect 686308 834820 686364 834876
rect 701316 821828 701372 821884
rect 686644 807716 686700 807772
rect 700532 806932 700588 806988
rect 703892 806260 703948 806316
rect 76356 783636 76412 783692
rect 83748 766052 83804 766108
rect 76132 765900 76188 765956
rect 76132 765452 76188 765508
rect 76244 765004 76300 765060
rect 84644 764484 84700 764540
rect 76244 763212 76300 763268
rect 80500 763140 80556 763196
rect 76132 762764 76188 762820
rect 82292 762804 82348 762860
rect 83748 762804 83804 762860
rect 84756 755412 84812 755468
rect 703892 755076 703948 755132
rect 704788 754404 704836 754460
rect 704836 754404 704844 754460
rect 705684 754404 705732 754460
rect 705732 754404 705740 754460
rect 699188 752500 699244 752556
rect 700420 752500 700476 752556
rect 75460 740964 75516 741020
rect 75460 740740 75516 740796
rect 700532 738724 700588 738780
rect 689556 735812 689612 735868
rect 686980 728084 687036 728140
rect 84644 725060 84700 725116
rect 76132 724900 76188 724956
rect 77140 724388 77196 724444
rect 76468 724004 76524 724060
rect 84644 722596 84700 722652
rect 77252 722372 77308 722428
rect 76132 722212 76188 722268
rect 76356 721764 76412 721820
rect 83748 720692 83804 720748
rect 686868 713972 686924 714028
rect 705684 711396 705732 711452
rect 705732 711396 705740 711452
rect 700420 710500 700476 710556
rect 686756 701428 686812 701484
rect 76356 701316 76412 701372
rect 694596 693924 694652 693980
rect 694596 693476 694652 693532
rect 84644 684292 84700 684348
rect 76132 683900 76188 683956
rect 76132 683452 76188 683508
rect 76468 683004 76524 683060
rect 84868 682276 84924 682332
rect 82292 682164 82348 682220
rect 76132 681212 76188 681268
rect 83748 681156 83804 681212
rect 76132 680764 76188 680820
rect 702100 676564 702156 676620
rect 705236 676452 705292 676508
rect 704452 676340 704508 676396
rect 701764 675444 701820 675500
rect 686532 673652 686588 673708
rect 702100 669060 702156 669116
rect 704452 668500 704508 668556
rect 705236 668500 705284 668556
rect 705284 668500 705292 668556
rect 705684 668388 705732 668444
rect 705732 668388 705740 668444
rect 701428 653180 701484 653236
rect 701428 651812 701484 651868
rect 694036 650916 694092 650972
rect 694708 650468 694764 650524
rect 694260 650020 694316 650076
rect 686420 648116 686476 648172
rect 76132 642900 76188 642956
rect 77140 642404 77196 642460
rect 83748 642292 83804 642348
rect 84756 642068 84812 642124
rect 76468 642004 76524 642060
rect 76132 640212 76188 640268
rect 77252 640052 77308 640108
rect 76356 639764 76412 639820
rect 705236 633556 705292 633612
rect 686308 633444 686364 633500
rect 701876 633444 701932 633500
rect 704452 633332 704508 633388
rect 705684 633332 705732 633388
rect 705732 633332 705740 633388
rect 704452 626500 704508 626556
rect 705236 626276 705284 626332
rect 705284 626276 705292 626332
rect 705684 626276 705732 626332
rect 705732 626276 705740 626332
rect 704788 625380 704836 625436
rect 704836 625380 704844 625436
rect 686196 621348 686252 621404
rect 76356 618996 76412 619052
rect 689668 609812 689724 609868
rect 686868 606452 686924 606508
rect 76244 603092 76300 603148
rect 84756 601972 84812 602028
rect 76132 601900 76188 601956
rect 76132 601452 76188 601508
rect 76468 601004 76524 601060
rect 80388 600628 80444 600684
rect 84980 599732 85036 599788
rect 76132 599212 76188 599268
rect 76356 598764 76412 598820
rect 83748 598500 83804 598556
rect 701652 590436 701708 590492
rect 704004 590324 704060 590380
rect 704452 590212 704508 590268
rect 701876 589764 701932 589820
rect 701652 583268 701708 583324
rect 76356 582820 76412 582876
rect 704004 582820 704060 582876
rect 704452 582820 704508 582876
rect 705684 582372 705732 582428
rect 705732 582372 705740 582428
rect 76468 578676 76524 578732
rect 85204 578676 85260 578732
rect 701428 567180 701484 567236
rect 701428 566132 701484 566188
rect 694932 565012 694988 565068
rect 686532 562772 686588 562828
rect 76468 562660 76524 562716
rect 76804 562548 76860 562604
rect 76580 562436 76636 562492
rect 84756 561764 84812 561820
rect 76132 560900 76188 560956
rect 77140 560420 77196 560476
rect 76356 560004 76412 560060
rect 84756 559412 84812 559468
rect 76244 558212 76300 558268
rect 83636 557844 83692 557900
rect 76132 557764 76188 557820
rect 77252 557732 77308 557788
rect 83748 557732 83804 557788
rect 686756 553476 686812 553532
rect 705012 547876 705068 547932
rect 702100 547764 702156 547820
rect 705124 547652 705180 547708
rect 701876 543396 701932 543452
rect 76356 542500 76412 542556
rect 76804 542388 76860 542444
rect 76580 542276 76636 542332
rect 84756 541156 84812 541212
rect 686868 540148 686924 540204
rect 705012 540148 705068 540204
rect 702100 540036 702156 540092
rect 705124 540036 705180 540092
rect 705684 539364 705732 539420
rect 705732 539364 705740 539420
rect 686420 526820 686476 526876
rect 694820 523796 694876 523852
rect 686308 521108 686364 521164
rect 76132 519900 76188 519956
rect 76244 519452 76300 519508
rect 84868 519092 84924 519148
rect 76468 519004 76524 519060
rect 80276 518868 80332 518924
rect 84980 517860 85036 517916
rect 76132 517212 76188 517268
rect 76356 516764 76412 516820
rect 83748 516404 83804 516460
rect 704452 504532 704508 504588
rect 701652 504420 701708 504476
rect 704004 504308 704060 504364
rect 701876 504084 701932 504140
rect 686308 487172 686364 487228
rect 85092 440468 85148 440524
rect 686644 433412 686700 433468
rect 76356 415716 76412 415772
rect 84980 412020 85036 412076
rect 686196 406756 686252 406812
rect 76580 399700 76636 399756
rect 76356 399588 76412 399644
rect 76132 396900 76188 396956
rect 83748 396900 83804 396956
rect 76132 396452 76188 396508
rect 78932 396116 78988 396172
rect 77140 396004 77196 396060
rect 84868 394996 84924 395052
rect 76132 394212 76188 394268
rect 76244 393764 76300 393820
rect 83748 393652 83804 393708
rect 83636 393428 83692 393484
rect 694820 380100 694876 380156
rect 76356 377860 76412 377916
rect 76580 377636 76636 377692
rect 84868 369796 84924 369852
rect 701652 368116 701708 368172
rect 704004 367780 704060 367836
rect 704452 367780 704508 367836
rect 705684 367332 705732 367388
rect 705732 367332 705740 367388
rect 84756 357140 84812 357196
rect 85428 357140 85484 357196
rect 84756 356916 84812 356972
rect 76244 356356 76300 356412
rect 76804 356244 76860 356300
rect 76580 356132 76636 356188
rect 76132 355900 76188 355956
rect 76132 355452 76188 355508
rect 76468 355004 76524 355060
rect 84756 355012 84812 355068
rect 85316 354788 85372 354844
rect 80164 354116 80220 354172
rect 76132 353212 76188 353268
rect 76356 352764 76412 352820
rect 694932 352212 694988 352268
rect 695044 349524 695100 349580
rect 686532 340228 686588 340284
rect 76580 337540 76636 337596
rect 76356 337428 76412 337484
rect 76804 337316 76860 337372
rect 393092 333732 393148 333788
rect 191492 333396 191548 333452
rect 370468 333396 370524 333452
rect 353556 333284 353612 333340
rect 487956 333284 488012 333340
rect 497364 333284 497420 333340
rect 533092 333284 533148 333340
rect 173012 333172 173068 333228
rect 188356 333172 188412 333228
rect 216132 333060 216188 333116
rect 701540 333060 701596 333116
rect 188356 332836 188412 332892
rect 704004 332836 704060 332892
rect 173012 332724 173068 332780
rect 205268 332724 205324 332780
rect 208292 332724 208348 332780
rect 216132 332724 216188 332780
rect 367892 332724 367948 332780
rect 701764 332724 701820 332780
rect 118356 332612 118412 332668
rect 201572 332612 201628 332668
rect 213332 332612 213388 332668
rect 320404 332612 320460 332668
rect 453684 332612 453740 332668
rect 551684 332612 551740 332668
rect 623252 332612 623308 332668
rect 704900 332612 704956 332668
rect 672308 332500 672364 332556
rect 341796 332164 341852 332220
rect 76468 331940 76524 331996
rect 378756 331940 378812 331996
rect 353780 330372 353836 330428
rect 336756 330260 336812 330316
rect 186452 329140 186508 329196
rect 656740 329140 656796 329196
rect 225876 328804 225932 328860
rect 269556 328804 269612 328860
rect 388276 328804 388332 328860
rect 405748 328804 405804 328860
rect 219380 328692 219436 328748
rect 365652 328580 365708 328636
rect 258580 328468 258636 328524
rect 169652 328356 169708 328412
rect 377860 328356 377916 328412
rect 236740 328244 236796 328300
rect 334516 328244 334572 328300
rect 291508 328020 291564 328076
rect 230244 327908 230300 327964
rect 343924 327908 343980 327964
rect 343476 327796 343532 327852
rect 334404 327684 334460 327740
rect 358708 327684 358764 327740
rect 334292 327572 334348 327628
rect 367892 327572 367948 327628
rect 453572 327460 453628 327516
rect 308980 327348 309036 327404
rect 317716 327236 317772 327292
rect 335972 327012 336028 327068
rect 300244 326564 300300 326620
rect 300468 326564 300524 326620
rect 295876 326228 295932 326284
rect 300468 326228 300524 326284
rect 376740 326228 376796 326284
rect 470372 326116 470428 326172
rect 382004 325780 382060 325836
rect 353556 325668 353612 325724
rect 704004 325108 704060 325164
rect 704900 325108 704956 325164
rect 376516 324996 376572 325052
rect 701540 324996 701596 325052
rect 505540 324884 505596 324940
rect 655508 324884 655564 324940
rect 537572 324548 537628 324604
rect 370468 324436 370524 324492
rect 554372 324436 554428 324492
rect 161028 324324 161084 324380
rect 347732 324324 347788 324380
rect 353780 324324 353836 324380
rect 376516 324324 376572 324380
rect 376740 324324 376796 324380
rect 705684 324324 705732 324380
rect 705732 324324 705740 324380
rect 104132 324100 104188 324156
rect 166292 324100 166348 324156
rect 169652 324100 169708 324156
rect 186452 324100 186508 324156
rect 191492 324100 191548 324156
rect 201572 324100 201628 324156
rect 205268 324100 205324 324156
rect 208292 324100 208348 324156
rect 213332 324100 213388 324156
rect 219380 324100 219436 324156
rect 225876 324100 225932 324156
rect 230244 324100 230300 324156
rect 236740 324100 236796 324156
rect 253540 324100 253596 324156
rect 255780 324100 255836 324156
rect 258580 324100 258636 324156
rect 260932 324100 260988 324156
rect 262612 324100 262668 324156
rect 263620 324100 263676 324156
rect 269556 324100 269612 324156
rect 291508 324100 291564 324156
rect 295876 324100 295932 324156
rect 299460 324100 299516 324156
rect 302260 324100 302316 324156
rect 306068 324100 306124 324156
rect 308980 324100 309036 324156
rect 311108 324100 311164 324156
rect 317716 324100 317772 324156
rect 333172 324100 333228 324156
rect 336644 324100 336700 324156
rect 341796 324100 341852 324156
rect 347620 324100 347676 324156
rect 357028 324100 357084 324156
rect 358484 324100 358540 324156
rect 365652 324100 365708 324156
rect 369460 324100 369516 324156
rect 377860 324100 377916 324156
rect 672420 324100 672476 324156
rect 260148 323988 260204 324044
rect 325780 323988 325836 324044
rect 334180 323988 334236 324044
rect 340452 323988 340508 324044
rect 365764 323988 365820 324044
rect 374276 323988 374332 324044
rect 377188 323988 377244 324044
rect 151172 323876 151228 323932
rect 672644 323988 672700 324044
rect 161812 323876 161868 323932
rect 316932 323876 316988 323932
rect 332276 323876 332332 323932
rect 347732 323876 347788 323932
rect 371588 323876 371644 323932
rect 376852 323876 376908 323932
rect 377300 323876 377356 323932
rect 378644 323876 378700 323932
rect 379540 323876 379596 323932
rect 380324 323092 380380 323148
rect 672756 322532 672812 322588
rect 379764 322196 379820 322252
rect 159572 321188 159628 321244
rect 379876 319508 379932 319564
rect 557732 319396 557788 319452
rect 379764 317268 379820 317324
rect 159796 316260 159852 316316
rect 76132 314900 76188 314956
rect 379764 314804 379820 314860
rect 84532 314356 84588 314412
rect 76356 314004 76412 314060
rect 83972 312452 84028 312508
rect 460292 312452 460348 312508
rect 379764 312340 379820 312396
rect 76132 312212 76188 312268
rect 76356 311764 76412 311820
rect 84084 311444 84140 311500
rect 159684 311332 159740 311388
rect 379764 309876 379820 309932
rect 458612 309204 458668 309260
rect 695156 309204 695212 309260
rect 248500 308644 248556 308700
rect 321636 308644 321692 308700
rect 322084 308644 322140 308700
rect 342580 308644 342636 308700
rect 344260 308644 344316 308700
rect 357700 308644 357756 308700
rect 377300 308644 377356 308700
rect 377748 308644 377804 308700
rect 162932 308532 162988 308588
rect 164724 308532 164780 308588
rect 166180 308532 166236 308588
rect 193172 308532 193228 308588
rect 203252 308532 203308 308588
rect 238420 308532 238476 308588
rect 297220 308532 297276 308588
rect 300692 308532 300748 308588
rect 307636 308532 307692 308588
rect 317380 308532 317436 308588
rect 320740 308532 320796 308588
rect 321860 308532 321916 308588
rect 164612 308420 164668 308476
rect 181412 308420 181468 308476
rect 183092 308420 183148 308476
rect 206612 308420 206668 308476
rect 209972 308420 210028 308476
rect 241780 308420 241836 308476
rect 261940 308420 261996 308476
rect 265300 308420 265356 308476
rect 282100 308420 282156 308476
rect 313796 308420 313852 308476
rect 334180 308420 334236 308476
rect 336196 308420 336252 308476
rect 362740 308420 362796 308476
rect 364420 308420 364476 308476
rect 369460 308420 369516 308476
rect 377860 308420 377916 308476
rect 190596 308308 190652 308364
rect 190820 308308 190876 308364
rect 234612 308308 234668 308364
rect 330036 308308 330092 308364
rect 378084 308196 378140 308252
rect 379428 308196 379484 308252
rect 337428 308084 337484 308140
rect 166180 307972 166236 308028
rect 190820 307860 190876 307916
rect 251972 307748 252028 307804
rect 462756 307748 462812 307804
rect 532420 307748 532476 307804
rect 99092 307412 99148 307468
rect 102452 307412 102508 307468
rect 303940 307412 303996 307468
rect 330036 307412 330092 307468
rect 377860 307412 377916 307468
rect 426692 307412 426748 307468
rect 551012 307412 551068 307468
rect 686868 307412 686924 307468
rect 538580 307188 538636 307244
rect 159684 306852 159740 306908
rect 85204 306628 85260 306684
rect 670628 306516 670684 306572
rect 686756 305956 686812 306012
rect 159908 305844 159964 305900
rect 84644 305732 84700 305788
rect 385924 303940 385980 303996
rect 520548 303940 520604 303996
rect 482132 303828 482188 303884
rect 285572 303716 285628 303772
rect 522340 303716 522396 303772
rect 201348 303268 201404 303324
rect 477876 303044 477932 303100
rect 83188 302372 83244 302428
rect 335860 302260 335916 302316
rect 286020 302148 286076 302204
rect 285572 302036 285628 302092
rect 354900 301812 354956 301868
rect 664356 301700 664412 301756
rect 285796 301588 285852 301644
rect 671188 301476 671244 301532
rect 356132 301364 356188 301420
rect 292292 300580 292348 300636
rect 294532 300580 294588 300636
rect 299012 300580 299068 300636
rect 302596 300580 302652 300636
rect 302820 300580 302876 300636
rect 337204 300468 337260 300524
rect 300692 300132 300748 300188
rect 381780 299684 381836 299740
rect 389732 299684 389788 299740
rect 343700 298228 343756 298284
rect 310996 297220 311052 297276
rect 335636 296772 335692 296828
rect 334628 296660 334684 296716
rect 337428 296548 337484 296604
rect 397460 296548 397516 296604
rect 336980 296436 337036 296492
rect 397236 296436 397292 296492
rect 336196 294756 336252 294812
rect 550116 293860 550172 293916
rect 539252 293412 539308 293468
rect 641508 293412 641564 293468
rect 641060 293300 641116 293356
rect 336756 293188 336812 293244
rect 640612 293188 640668 293244
rect 640052 293076 640108 293132
rect 510692 292964 510748 293020
rect 629076 292964 629132 293020
rect 488852 292852 488908 292908
rect 606116 292852 606172 292908
rect 498932 292740 498988 292796
rect 497252 292516 497308 292572
rect 465332 292292 465388 292348
rect 670292 292292 670348 292348
rect 92372 292180 92428 292236
rect 320964 292180 321020 292236
rect 321188 292180 321244 292236
rect 321412 292180 321468 292236
rect 541716 292180 541772 292236
rect 93156 291956 93212 292012
rect 173236 291844 173292 291900
rect 428820 291844 428876 291900
rect 428596 291732 428652 291788
rect 534212 291620 534268 291676
rect 430388 291508 430444 291564
rect 506436 291508 506492 291564
rect 532532 291284 532588 291340
rect 117908 291060 117964 291116
rect 521332 290948 521388 291004
rect 535892 290836 535948 290892
rect 92596 290612 92652 290668
rect 606340 290612 606396 290668
rect 475412 290500 475468 290556
rect 615636 290500 615692 290556
rect 637252 290500 637308 290556
rect 646548 290500 646604 290556
rect 669844 290500 669900 290556
rect 689332 290500 689388 290556
rect 165396 290388 165452 290444
rect 607796 290388 607852 290444
rect 616420 290388 616476 290444
rect 670292 290388 670348 290444
rect 688212 290388 688268 290444
rect 80276 290276 80332 290332
rect 472052 290276 472108 290332
rect 608916 290276 608972 290332
rect 614516 290276 614572 290332
rect 666932 290276 666988 290332
rect 606340 290164 606396 290220
rect 607796 290164 607852 290220
rect 614740 290164 614796 290220
rect 78820 290052 78876 290108
rect 606116 290052 606172 290108
rect 611044 290052 611100 290108
rect 615412 290052 615468 290108
rect 617540 290052 617596 290108
rect 631764 290052 631820 290108
rect 666932 290052 666988 290108
rect 671188 290052 671244 290108
rect 611268 289940 611324 289996
rect 611492 289940 611548 289996
rect 611940 289940 611996 289996
rect 620676 289940 620732 289996
rect 629188 289940 629244 289996
rect 644196 289940 644252 289996
rect 652596 289828 652652 289884
rect 671300 289828 671356 289884
rect 672308 289828 672364 289884
rect 704676 289828 704732 289884
rect 705012 289828 705068 289884
rect 620676 289716 620732 289772
rect 622804 289716 622860 289772
rect 623252 289716 623308 289772
rect 626164 289716 626220 289772
rect 628068 289716 628124 289772
rect 629076 289716 629132 289772
rect 629300 289716 629356 289772
rect 631764 289716 631820 289772
rect 631988 289716 632044 289772
rect 636244 289716 636300 289772
rect 636692 289716 636748 289772
rect 638148 289716 638204 289772
rect 638708 289716 638764 289772
rect 640052 289716 640108 289772
rect 640612 289716 640668 289772
rect 641060 289716 641116 289772
rect 641508 289716 641564 289772
rect 642516 289716 642572 289772
rect 644196 289716 644252 289772
rect 644420 289716 644476 289772
rect 652260 289716 652316 289772
rect 655508 289716 655564 289772
rect 658308 289716 658364 289772
rect 661668 289716 661724 289772
rect 667268 289716 667324 289772
rect 667492 289716 667548 289772
rect 671076 289716 671132 289772
rect 671636 289716 671692 289772
rect 600516 289492 600572 289548
rect 702100 289380 702156 289436
rect 479556 289268 479612 289324
rect 337540 289156 337596 289212
rect 687540 289156 687596 289212
rect 608916 289044 608972 289100
rect 701988 289044 702044 289100
rect 611380 288820 611436 288876
rect 559188 288484 559244 288540
rect 671860 288372 671916 288428
rect 468580 288260 468636 288316
rect 165620 288148 165676 288204
rect 474516 288148 474572 288204
rect 611044 288148 611100 288204
rect 469140 288036 469196 288092
rect 468580 287252 468636 287308
rect 469140 287252 469196 287308
rect 474516 287252 474572 287308
rect 559076 286132 559132 286188
rect 327908 285236 327964 285292
rect 327684 284900 327740 284956
rect 329588 284900 329644 284956
rect 377972 284676 378028 284732
rect 444052 284564 444108 284620
rect 558852 283892 558908 283948
rect 609924 283220 609980 283276
rect 609812 282996 609868 283052
rect 334404 282212 334460 282268
rect 196532 282100 196588 282156
rect 262052 282100 262108 282156
rect 334628 282100 334684 282156
rect 391412 282100 391468 282156
rect 445284 282100 445340 282156
rect 446628 282100 446684 282156
rect 705012 282100 705068 282156
rect 168420 281988 168476 282044
rect 274036 281988 274092 282044
rect 320628 281988 320684 282044
rect 704676 281988 704732 282044
rect 153748 281876 153804 281932
rect 173796 281876 173852 281932
rect 316820 281876 316876 281932
rect 702100 281876 702156 281932
rect 335860 281764 335916 281820
rect 397236 281764 397292 281820
rect 320628 281652 320684 281708
rect 342804 281652 342860 281708
rect 352772 281652 352828 281708
rect 397460 281652 397516 281708
rect 173796 281540 173852 281596
rect 196644 281540 196700 281596
rect 343476 281540 343532 281596
rect 185780 281316 185836 281372
rect 196756 281316 196812 281372
rect 705684 281316 705732 281372
rect 705732 281316 705740 281372
rect 153972 281204 154028 281260
rect 162484 281204 162540 281260
rect 168420 281204 168476 281260
rect 335636 281204 335692 281260
rect 342804 281204 342860 281260
rect 377636 281204 377692 281260
rect 558740 281204 558796 281260
rect 185780 281092 185836 281148
rect 196644 280980 196700 281036
rect 274036 280980 274092 281036
rect 321636 280980 321692 281036
rect 558292 280980 558348 281036
rect 100772 280868 100828 280924
rect 154644 280868 154700 280924
rect 159796 280868 159852 280924
rect 181636 280868 181692 280924
rect 196756 280868 196812 280924
rect 153748 280644 153804 280700
rect 153972 280644 154028 280700
rect 162484 280644 162540 280700
rect 245252 280868 245308 280924
rect 272132 280868 272188 280924
rect 343700 280868 343756 280924
rect 378084 280868 378140 280924
rect 461972 280868 462028 280924
rect 477876 280868 477932 280924
rect 482132 280868 482188 280924
rect 537572 280868 537628 280924
rect 557732 280868 557788 280924
rect 307636 280756 307692 280812
rect 558628 280756 558684 280812
rect 338436 280644 338492 280700
rect 559300 279636 559356 279692
rect 671748 276836 671804 276892
rect 559300 276724 559356 276780
rect 76244 274036 76300 274092
rect 76132 273900 76188 273956
rect 76356 273924 76412 273980
rect 559300 273476 559356 273532
rect 76468 273004 76524 273060
rect 76244 272556 76300 272612
rect 85092 272132 85148 272188
rect 76132 271212 76188 271268
rect 76244 270764 76300 270820
rect 84196 270788 84252 270844
rect 559300 270452 559356 270508
rect 559300 265076 559356 265132
rect 686420 263844 686476 263900
rect 559300 263396 559356 263452
rect 689220 262948 689276 263004
rect 559300 256116 559356 256172
rect 689108 256116 689164 256172
rect 76356 255220 76412 255276
rect 559524 246932 559580 246988
rect 689556 246820 689612 246876
rect 704676 246820 704732 246876
rect 704564 246260 704620 246316
rect 559300 243572 559356 243628
rect 704564 239092 704620 239148
rect 704676 238420 704732 238476
rect 76356 233492 76412 233548
rect 694596 233044 694652 233100
rect 76132 232900 76188 232956
rect 76356 232452 76412 232508
rect 76468 232004 76524 232060
rect 84644 232036 84700 232092
rect 85204 231812 85260 231868
rect 76244 231556 76300 231612
rect 76132 230212 76188 230268
rect 76356 229764 76412 229820
rect 694708 226100 694764 226156
rect 686308 220052 686364 220108
rect 701428 220044 701484 220100
rect 701428 218372 701484 218428
rect 689668 214564 689724 214620
rect 559300 209188 559356 209244
rect 84644 207844 84700 207900
rect 84756 207620 84812 207676
rect 701428 203588 701484 203644
rect 701652 203476 701708 203532
rect 703892 203364 703948 203420
rect 701876 203252 701932 203308
rect 695044 198436 695100 198492
rect 701652 196196 701708 196252
rect 703892 196084 703948 196140
rect 701876 195972 701932 196028
rect 705684 195412 705732 195468
rect 705732 195412 705740 195468
rect 694932 193732 694988 193788
rect 76132 191900 76188 191956
rect 76132 191452 76188 191508
rect 90356 191268 90412 191324
rect 76468 191004 76524 191060
rect 84308 190932 84364 190988
rect 83860 190596 83916 190652
rect 76132 189212 76188 189268
rect 76244 188764 76300 188820
rect 695156 186900 695212 186956
rect 559300 186116 559356 186172
rect 559636 185668 559692 185724
rect 696164 177940 696220 177996
rect 689556 176596 689612 176652
rect 686644 176484 686700 176540
rect 559300 176372 559356 176428
rect 696164 176372 696220 176428
rect 689556 170660 689612 170716
rect 671748 161476 671804 161532
rect 705012 160804 705068 160860
rect 702100 160356 702156 160412
rect 705236 160244 705292 160300
rect 701988 159684 702044 159740
rect 585396 158900 585452 158956
rect 705012 152740 705068 152796
rect 705236 152740 705284 152796
rect 705284 152740 705292 152796
rect 702100 152516 702156 152572
rect 705684 152404 705732 152460
rect 705732 152404 705740 152460
rect 671748 152292 671804 152348
rect 585620 147476 585676 147532
rect 559300 147364 559356 147420
rect 671860 145348 671916 145404
rect 585844 145236 585900 145292
rect 559412 143332 559468 143388
rect 585172 142996 585228 143052
rect 671748 142660 671804 142716
rect 671860 142100 671916 142156
rect 559412 141652 559468 141708
rect 671972 141540 672028 141596
rect 671748 141092 671804 141148
rect 623364 139972 623420 140028
rect 624708 139972 624764 140028
rect 657076 139972 657132 140028
rect 657748 139972 657804 140028
rect 631428 139860 631484 139916
rect 655732 139860 655788 139916
rect 671188 139860 671244 139916
rect 618212 139748 618268 139804
rect 669956 139748 670012 139804
rect 622020 139636 622076 139692
rect 632772 139636 632828 139692
rect 638820 139636 638876 139692
rect 650692 139636 650748 139692
rect 656404 139636 656460 139692
rect 666484 139636 666540 139692
rect 670404 139636 670460 139692
rect 618660 139524 618716 139580
rect 670068 139524 670124 139580
rect 619892 139412 619948 139468
rect 648452 139412 648508 139468
rect 650804 139412 650860 139468
rect 670852 139412 670908 139468
rect 670964 138964 671020 139020
rect 670740 138740 670796 138796
rect 559300 138516 559356 138572
rect 669620 137956 669676 138012
rect 669844 137844 669900 137900
rect 669732 137732 669788 137788
rect 670404 136948 670460 137004
rect 670292 136836 670348 136892
rect 694820 136724 694876 136780
rect 649460 136276 649516 136332
rect 649796 136276 649852 136332
rect 649908 136164 649964 136220
rect 650020 136052 650076 136108
rect 622356 135604 622412 135660
rect 622244 135492 622300 135548
rect 669956 135492 670012 135548
rect 622804 135380 622860 135436
rect 622692 135268 622748 135324
rect 700532 135380 700588 135436
rect 622580 135156 622636 135212
rect 669620 135156 669676 135212
rect 669956 135156 670012 135212
rect 669844 135044 669900 135100
rect 669620 134932 669676 134988
rect 650132 134820 650188 134876
rect 621460 134484 621516 134540
rect 618436 134372 618492 134428
rect 621348 134372 621404 134428
rect 686196 134372 686252 134428
rect 701428 134044 701484 134100
rect 650132 133140 650188 133196
rect 649460 132692 649516 132748
rect 701428 132692 701484 132748
rect 650020 132580 650076 132636
rect 657972 132580 658028 132636
rect 664580 132580 664636 132636
rect 666820 132580 666876 132636
rect 669620 132580 669676 132636
rect 670852 132580 670908 132636
rect 649908 132468 649964 132524
rect 659652 132468 659708 132524
rect 670516 132468 670572 132524
rect 650692 132356 650748 132412
rect 650916 132356 650972 132412
rect 669732 132356 669788 132412
rect 669844 132244 669900 132300
rect 653492 132132 653548 132188
rect 649684 131908 649740 131964
rect 670292 132132 670348 132188
rect 649572 131796 649628 131852
rect 671188 131908 671244 131964
rect 670404 131796 670460 131852
rect 649348 131684 649404 131740
rect 670180 131460 670236 131516
rect 670068 131348 670124 131404
rect 665140 131012 665196 131068
rect 654500 127540 654556 127596
rect 646324 127428 646380 127484
rect 654276 126756 654332 126812
rect 655956 126644 656012 126700
rect 559300 125972 559356 126028
rect 646996 125972 647052 126028
rect 655620 125972 655676 126028
rect 626052 125860 626108 125916
rect 628068 125860 628124 125916
rect 628740 125860 628796 125916
rect 641508 125860 641564 125916
rect 654612 125748 654668 125804
rect 655956 125636 656012 125692
rect 655844 125524 655900 125580
rect 655732 125412 655788 125468
rect 655284 125300 655340 125356
rect 670180 123508 670236 123564
rect 620564 123396 620620 123452
rect 620340 123284 620396 123340
rect 642740 123284 642796 123340
rect 647892 123284 647948 123340
rect 654948 122836 655004 122892
rect 618772 122612 618828 122668
rect 655284 121492 655340 121548
rect 655284 120596 655340 120652
rect 655732 120596 655788 120652
rect 655396 119812 655452 119868
rect 655396 118916 655452 118972
rect 655844 118916 655900 118972
rect 655060 118356 655116 118412
rect 701652 118020 701708 118076
rect 704900 117796 704956 117852
rect 701876 117684 701932 117740
rect 704004 117572 704060 117628
rect 559300 114212 559356 114268
rect 654948 113204 655004 113260
rect 655620 111076 655676 111132
rect 559300 110852 559356 110908
rect 651924 110180 651980 110236
rect 704004 110068 704060 110124
rect 704900 110068 704956 110124
rect 701652 109956 701708 110012
rect 652932 109620 652988 109676
rect 705684 109396 705732 109452
rect 705732 109396 705740 109452
rect 559300 105140 559356 105196
rect 619892 100660 619948 100716
rect 622356 100660 622412 100716
rect 654724 100660 654780 100716
rect 622804 100436 622860 100492
rect 628628 100436 628684 100492
rect 631204 100436 631260 100492
rect 649572 100436 649628 100492
rect 654612 100436 654668 100492
rect 633780 99988 633836 100044
rect 635796 99988 635852 100044
rect 639044 99988 639100 100044
rect 641732 99988 641788 100044
rect 644980 99988 645036 100044
rect 654500 98868 654556 98924
rect 619332 97412 619388 97468
rect 652932 95620 652988 95676
rect 619108 94948 619164 95004
rect 701428 93732 701484 93788
rect 694596 92484 694652 92540
rect 686532 92372 686588 92428
rect 701428 92372 701484 92428
rect 701428 91940 701484 91996
rect 618548 91252 618604 91308
rect 559300 90692 559356 90748
rect 701428 90692 701484 90748
rect 652932 89012 652988 89068
rect 618660 88676 618716 88732
rect 559300 87444 559356 87500
rect 618884 87444 618940 87500
rect 618324 84980 618380 85036
rect 559300 84420 559356 84476
rect 618212 83748 618268 83804
rect 652932 82964 652988 83020
rect 559300 81732 559356 81788
rect 585172 81732 585228 81788
rect 558516 81620 558572 81676
rect 558292 81508 558348 81564
rect 559076 81396 559132 81452
rect 558964 81284 559020 81340
rect 558740 81172 558796 81228
rect 92372 80836 92428 80892
rect 335972 80724 336028 80780
rect 628068 80612 628124 80668
rect 645092 80612 645148 80668
rect 93828 79044 93884 79100
rect 324884 72100 324940 72156
rect 559412 71988 559468 72044
rect 396116 71540 396172 71596
rect 231252 71316 231308 71372
rect 620564 71316 620620 71372
rect 619332 71092 619388 71148
rect 617988 70980 618044 71036
rect 257796 70532 257852 70588
rect 396116 70532 396172 70588
rect 559412 70532 559468 70588
rect 539140 70308 539196 70364
rect 176260 70084 176316 70140
rect 231252 70084 231308 70140
rect 494340 70084 494343 70140
rect 494343 70084 494396 70140
rect 505876 70084 505890 70140
rect 505890 70084 505932 70140
rect 548436 70084 548488 70140
rect 548488 70084 548492 70140
rect 519652 69748 519708 69804
<< metal4 >>
rect 470260 949228 470316 949238
rect 106596 947788 106652 947798
rect 75460 945980 75516 945990
rect 75460 945756 75516 945924
rect 75460 945690 75516 945700
rect 85428 942620 85484 942630
rect 84084 936928 84140 936938
rect 84084 935788 84140 936872
rect 84084 935722 84140 935732
rect 84308 936748 84364 936758
rect 84308 935788 84364 936692
rect 84308 935722 84364 935732
rect 84532 936568 84588 936578
rect 84532 935788 84588 936512
rect 84532 935722 84588 935732
rect 85428 935676 85484 942564
rect 106596 942396 106652 947732
rect 216580 947788 216636 947798
rect 196084 946764 196140 946774
rect 121940 943404 121996 943414
rect 121940 942732 121996 943348
rect 121940 942666 121996 942676
rect 122388 943404 122444 943414
rect 122388 942620 122444 943348
rect 122388 942554 122444 942564
rect 106596 942330 106652 942340
rect 196084 942060 196140 946708
rect 216580 942396 216636 947732
rect 271572 947788 271628 947798
rect 251188 947660 251244 947670
rect 251076 946764 251132 946774
rect 216580 942330 216636 942340
rect 233492 943292 233548 943302
rect 196084 941994 196140 942004
rect 141876 937020 141932 937030
rect 141876 936928 141932 936964
rect 141876 936862 141932 936872
rect 178724 937020 178780 937030
rect 141652 936796 141708 936806
rect 141428 936684 141484 936694
rect 141652 936682 141708 936692
rect 141428 936568 141484 936628
rect 141428 936502 141484 936512
rect 178724 936568 178780 936964
rect 178724 936502 178780 936512
rect 85428 935610 85484 935620
rect 233492 935228 233548 943236
rect 251076 942172 251132 946708
rect 251188 942284 251244 947604
rect 251188 942218 251244 942228
rect 271572 942284 271628 947732
rect 470260 947788 470316 949172
rect 470260 947722 470316 947732
rect 525700 947788 525756 947798
rect 306068 947660 306124 947670
rect 271572 942218 271628 942228
rect 289828 943404 289884 943414
rect 251076 942106 251132 942116
rect 282436 937468 282492 937506
rect 282436 937402 282492 937412
rect 289828 937468 289884 943348
rect 306068 942396 306124 947604
rect 361396 947548 361452 947558
rect 361284 947212 361340 947222
rect 361172 946764 361228 946774
rect 341236 943404 341292 943414
rect 306068 942330 306124 942340
rect 334292 942396 334348 942406
rect 334292 942172 334348 942340
rect 334292 942106 334348 942116
rect 289828 937402 289884 937412
rect 341012 937468 341068 937478
rect 285684 937132 285740 937142
rect 285684 936748 285740 937076
rect 285684 936682 285740 936692
rect 233492 935162 233548 935172
rect 341012 934892 341068 937412
rect 341236 937288 341292 943348
rect 342692 943404 342748 943414
rect 342692 937468 342748 943348
rect 361172 942396 361228 946708
rect 361172 942330 361228 942340
rect 361284 942172 361340 947156
rect 361396 942284 361452 947492
rect 525700 947548 525756 947732
rect 690340 947788 690396 947798
rect 525700 947482 525756 947492
rect 545860 947548 545916 947558
rect 545860 947454 545916 947492
rect 581140 947548 581196 947558
rect 581140 947454 581196 947492
rect 655844 947548 655900 947558
rect 655844 947454 655900 947492
rect 690340 947548 690396 947732
rect 690340 947482 690396 947492
rect 697956 947548 698012 947558
rect 697956 947454 698012 947492
rect 525588 947340 525644 947350
rect 471268 946892 471324 946902
rect 471268 945980 471324 946836
rect 525588 946288 525644 947284
rect 690340 947340 690396 947350
rect 581252 947212 581308 947222
rect 545860 947100 545916 947110
rect 545636 946892 545692 946902
rect 526148 946764 526204 946774
rect 525588 946222 525644 946232
rect 525700 946444 525756 946454
rect 525700 946108 525756 946388
rect 525700 946042 525756 946052
rect 471268 945914 471324 945924
rect 526148 945928 526204 946708
rect 545524 946444 545580 946454
rect 545524 946288 545580 946388
rect 545524 946222 545580 946232
rect 526148 945862 526204 945872
rect 545636 945928 545692 946836
rect 545860 946108 545916 947044
rect 545860 946042 545916 946052
rect 581028 946764 581084 946774
rect 581028 946108 581084 946708
rect 581140 946316 581196 946326
rect 581140 946222 581196 946232
rect 581028 946042 581084 946052
rect 545636 945862 545692 945872
rect 581252 945928 581308 947156
rect 655844 947100 655900 947110
rect 655620 946892 655676 946902
rect 581252 945862 581308 945872
rect 655508 946444 655564 946454
rect 655508 945928 655564 946388
rect 655620 946108 655676 946836
rect 655844 946288 655900 947044
rect 655844 946222 655900 946232
rect 655620 946042 655676 946052
rect 655508 945862 655564 945872
rect 690340 945928 690396 947284
rect 690340 945862 690396 945872
rect 692916 946876 692972 946886
rect 361396 942218 361452 942228
rect 454244 943516 454300 943526
rect 361284 942106 361340 942116
rect 454244 938188 454300 943460
rect 561316 943404 561372 943414
rect 454244 938122 454300 938132
rect 458500 938188 458556 938198
rect 342692 937402 342748 937412
rect 341236 937222 341292 937232
rect 341012 934826 341068 934836
rect 458500 934892 458556 938132
rect 561316 936928 561372 943348
rect 564900 943404 564956 943414
rect 564900 938368 564956 943348
rect 670292 943404 670348 943414
rect 564900 938302 564956 938312
rect 565012 943292 565068 943302
rect 565012 937108 565068 943236
rect 565012 937042 565068 937052
rect 587524 938368 587580 938378
rect 561316 936862 561372 936872
rect 587524 935676 587580 938312
rect 670292 936388 670348 943348
rect 688212 937356 688268 937366
rect 687428 937288 687484 937298
rect 687428 937178 687484 937188
rect 687988 936748 688044 936758
rect 687988 936572 688044 936692
rect 687988 936506 688044 936516
rect 670292 936322 670348 936332
rect 587524 935610 587580 935620
rect 686420 935668 686476 935678
rect 458500 934826 458556 934836
rect 686196 935488 686252 935498
rect 76132 929956 76188 929966
rect 76132 929842 76188 929852
rect 83748 929908 83804 929918
rect 83748 929786 83804 929796
rect 76356 929508 76412 929518
rect 76132 929060 76188 929070
rect 76132 902187 76188 929004
rect 76356 927388 76412 929452
rect 76356 927322 76412 927332
rect 78932 927388 78988 927398
rect 78932 927294 78988 927332
rect 76244 927268 76300 927278
rect 76244 926488 76300 927212
rect 84644 926940 84700 926950
rect 76244 926422 76300 926432
rect 76356 926820 76412 926830
rect 76020 902131 76188 902187
rect 76020 897148 76076 902131
rect 76020 897082 76076 897092
rect 76356 783692 76412 926764
rect 84644 926488 84700 926884
rect 84644 926422 84700 926432
rect 76356 783626 76412 783636
rect 76132 766108 76188 766118
rect 76132 765956 76188 766052
rect 83748 766108 83804 766118
rect 83748 766014 83804 766052
rect 76132 765890 76188 765900
rect 76132 765508 76188 765518
rect 76132 763228 76188 765452
rect 76244 765060 76300 765070
rect 76244 764488 76300 765004
rect 76244 764422 76300 764432
rect 84644 764540 84700 764550
rect 84644 764422 84700 764432
rect 76132 763162 76188 763172
rect 76244 763268 76300 763278
rect 76132 763048 76188 763058
rect 76132 762820 76188 762992
rect 76244 762868 76300 763212
rect 80500 763228 80556 763238
rect 80500 763130 80556 763140
rect 76244 762802 76300 762812
rect 82292 763048 82348 763058
rect 82292 762860 82348 762992
rect 82292 762794 82348 762804
rect 83748 762868 83804 762898
rect 83748 762794 83804 762804
rect 76132 762754 76188 762764
rect 84756 755468 84812 755478
rect 75460 741020 75516 741030
rect 75460 740796 75516 740964
rect 75460 740730 75516 740740
rect 84644 725116 84700 725126
rect 76132 725068 76188 725078
rect 76132 724956 76188 725012
rect 84644 725002 84700 725012
rect 76132 724890 76188 724900
rect 77140 724444 77196 724454
rect 76468 724060 76524 724070
rect 76468 722548 76524 724004
rect 77140 722548 77196 724388
rect 84644 722652 84700 722662
rect 84644 722548 84700 722596
rect 77140 722492 77308 722548
rect 76468 722482 76524 722492
rect 77252 722428 77308 722492
rect 84644 722482 84700 722492
rect 77252 722362 77308 722372
rect 76132 722268 76188 722278
rect 76132 720748 76188 722212
rect 76132 720682 76188 720692
rect 76356 721820 76412 721830
rect 76356 701372 76412 721764
rect 83748 720748 83804 720758
rect 83748 720654 83804 720692
rect 76356 701306 76412 701316
rect 84644 684348 84700 684358
rect 76132 684028 76188 684038
rect 76132 683956 76188 683972
rect 84644 684028 84700 684292
rect 84644 683962 84700 683972
rect 76132 683890 76188 683900
rect 76132 683508 76188 683518
rect 76132 682408 76188 683452
rect 76132 682342 76188 682352
rect 76468 683060 76524 683070
rect 76468 682228 76524 683004
rect 76468 682162 76524 682172
rect 82292 682408 82348 682418
rect 82292 682220 82348 682352
rect 82292 682154 82348 682164
rect 76132 681268 76188 681278
rect 76132 681148 76188 681212
rect 76132 681082 76188 681092
rect 83748 681212 83804 681222
rect 83748 681148 83804 681156
rect 83748 681082 83804 681092
rect 76132 680968 76188 680978
rect 76132 680820 76188 680912
rect 76132 680754 76188 680764
rect 84644 680968 84700 680978
rect 76132 642956 76188 642966
rect 76132 642268 76188 642900
rect 76132 642202 76188 642212
rect 77140 642460 77196 642470
rect 76468 642088 76524 642098
rect 76468 641994 76524 642004
rect 76132 640268 76188 640278
rect 76132 640108 76188 640212
rect 77140 640108 77196 642404
rect 83748 642348 83804 642358
rect 83748 642268 83804 642292
rect 83748 642202 83804 642212
rect 77252 640108 77308 640118
rect 77140 640052 77252 640108
rect 76132 640042 76188 640052
rect 77252 640042 77308 640052
rect 76356 639820 76412 639830
rect 76356 619052 76412 639764
rect 76356 618986 76412 618996
rect 76244 603148 76300 603158
rect 76132 601956 76188 601986
rect 76132 601882 76188 601892
rect 76132 601508 76188 601518
rect 76132 600688 76188 601452
rect 76132 600622 76188 600632
rect 76132 599268 76188 599278
rect 76132 598528 76188 599212
rect 76132 598462 76188 598472
rect 76244 596427 76300 603092
rect 76468 601060 76524 601070
rect 76468 599788 76524 601004
rect 80388 600688 80444 600722
rect 80388 600618 80444 600628
rect 76468 599722 76524 599732
rect 76356 598820 76412 598830
rect 76356 597628 76412 598764
rect 83748 598556 83804 598566
rect 83748 598462 83804 598472
rect 76356 597572 76524 597628
rect 76244 596371 76412 596427
rect 76356 582876 76412 596371
rect 76356 582810 76412 582820
rect 76468 578732 76524 597572
rect 76468 578666 76524 578676
rect 76468 562716 76524 562726
rect 76132 561808 76188 561818
rect 76132 560956 76188 561752
rect 76132 560890 76188 560900
rect 76356 560060 76412 560070
rect 76356 559468 76412 560004
rect 76356 559402 76412 559412
rect 76244 558268 76300 558278
rect 76132 558028 76188 558038
rect 76132 557820 76188 557972
rect 76244 557848 76300 558212
rect 76244 557782 76300 557792
rect 76132 557754 76188 557764
rect 76468 549387 76524 562660
rect 76804 562604 76860 562614
rect 76356 549331 76524 549387
rect 76580 562492 76636 562502
rect 76356 542556 76412 549331
rect 76356 542490 76412 542500
rect 76580 542332 76636 562436
rect 76804 542444 76860 562548
rect 77140 560476 77196 560486
rect 77140 557848 77196 560420
rect 83748 558028 83804 558038
rect 83636 557900 83692 557910
rect 77140 557792 77308 557848
rect 77252 557788 77308 557792
rect 83636 557782 83692 557792
rect 83748 557788 83804 557972
rect 77252 557722 77308 557732
rect 83748 557722 83804 557732
rect 76804 542378 76860 542388
rect 76580 542266 76636 542276
rect 76132 519956 76188 519966
rect 76132 519148 76188 519900
rect 76132 519082 76188 519092
rect 76244 519508 76300 519518
rect 76244 518968 76300 519452
rect 76244 518902 76300 518912
rect 76468 519060 76524 519070
rect 76468 517528 76524 519004
rect 80276 518968 80332 518978
rect 80276 518858 80332 518868
rect 76468 517462 76524 517472
rect 76132 517268 76188 517278
rect 76132 516448 76188 517212
rect 76132 516382 76188 516392
rect 76356 516820 76412 516830
rect 76356 415772 76412 516764
rect 83748 516460 83804 516470
rect 83748 516366 83804 516392
rect 76356 415706 76412 415716
rect 76580 399756 76636 399766
rect 76356 399644 76412 399654
rect 76132 396956 76188 396966
rect 76132 396862 76188 396872
rect 76132 396508 76188 396518
rect 76132 396208 76188 396452
rect 76132 396142 76188 396152
rect 76132 394268 76188 394278
rect 76132 393688 76188 394212
rect 76132 393622 76188 393632
rect 76244 393820 76300 393830
rect 76244 393508 76300 393764
rect 76244 393442 76300 393452
rect 76356 377916 76412 399588
rect 76356 377850 76412 377860
rect 76580 377692 76636 399700
rect 83748 396956 83804 396966
rect 83748 396862 83804 396872
rect 78932 396208 78988 396218
rect 78932 396106 78988 396116
rect 77140 396060 77196 396070
rect 77140 394948 77196 396004
rect 77140 394882 77196 394892
rect 83748 393708 83804 393718
rect 83748 393614 83804 393632
rect 83636 393508 83692 393522
rect 83636 393418 83692 393428
rect 76580 377626 76636 377636
rect 76132 356968 76188 356978
rect 76132 355956 76188 356912
rect 76132 355890 76188 355900
rect 76244 356412 76300 356422
rect 76132 355508 76188 355518
rect 76132 354268 76188 355452
rect 76132 354202 76188 354212
rect 76132 353268 76188 353278
rect 76132 352828 76188 353212
rect 76132 352762 76188 352772
rect 76244 349467 76300 356356
rect 76804 356300 76860 356310
rect 76580 356188 76636 356198
rect 76468 355060 76524 355070
rect 76468 354988 76524 355004
rect 76468 354922 76524 354932
rect 76356 352820 76412 352830
rect 76356 351208 76412 352764
rect 76356 351152 76524 351208
rect 76244 349411 76412 349467
rect 76356 337484 76412 349411
rect 76356 337418 76412 337428
rect 76468 331996 76524 351152
rect 76580 337596 76636 356132
rect 76580 337530 76636 337540
rect 76804 337372 76860 356244
rect 80164 354268 80220 354278
rect 80164 354172 80220 354212
rect 80164 354106 80220 354116
rect 76804 337306 76860 337316
rect 76468 331930 76524 331940
rect 76132 314956 76188 314966
rect 76132 314308 76188 314900
rect 76132 314242 76188 314252
rect 84532 314412 84588 314422
rect 84532 314308 84588 314356
rect 84532 314242 84588 314252
rect 76356 314060 76412 314070
rect 76356 312508 76412 314004
rect 76356 312442 76412 312452
rect 83972 312508 84028 312518
rect 83972 312414 84028 312452
rect 76132 312268 76188 312278
rect 76132 311428 76188 312212
rect 76132 311362 76188 311372
rect 76356 311820 76412 311830
rect 76356 301528 76412 311764
rect 84084 311500 84140 311510
rect 84084 311428 84140 311444
rect 84084 311362 84140 311372
rect 84644 305788 84700 680912
rect 84756 655227 84812 755412
rect 84868 682332 84924 682342
rect 84868 682228 84924 682276
rect 84868 682162 84924 682172
rect 84756 655171 84924 655227
rect 84756 642124 84812 642134
rect 84756 642022 84812 642032
rect 84868 640108 84924 655171
rect 84868 640042 84924 640052
rect 686196 621404 686252 935432
rect 686308 934892 686364 934902
rect 686308 834876 686364 934836
rect 686308 834810 686364 834820
rect 686420 648172 686476 935612
rect 686980 934444 687036 934454
rect 686644 934408 686700 934418
rect 686644 807772 686700 934352
rect 686644 807706 686700 807716
rect 686756 934332 686812 934342
rect 686756 701484 686812 934276
rect 686980 728140 687036 934388
rect 686980 728074 687036 728084
rect 686756 701418 686812 701428
rect 686868 714028 686924 714038
rect 686420 648106 686476 648116
rect 686532 673708 686588 673718
rect 686196 621338 686252 621348
rect 686308 633500 686364 633510
rect 84756 602028 84812 602038
rect 84756 601948 84812 601972
rect 84756 601882 84812 601892
rect 84980 599788 85036 599798
rect 84980 599694 85036 599732
rect 85204 578732 85260 578742
rect 84756 561820 84812 561830
rect 84756 561726 84812 561752
rect 84756 559468 84812 559478
rect 84756 559374 84812 559412
rect 84756 541212 84812 541222
rect 84756 357196 84812 541156
rect 84868 519148 84924 519158
rect 84868 519054 84924 519092
rect 84980 517916 85036 517926
rect 84980 517528 85036 517860
rect 84980 517462 85036 517472
rect 85092 440524 85148 440534
rect 84980 412076 85036 412086
rect 84868 395052 84924 395062
rect 84868 394948 84924 394996
rect 84868 394882 84924 394892
rect 84756 357130 84812 357140
rect 84868 369852 84924 369862
rect 84756 356972 84812 356982
rect 84756 356878 84812 356912
rect 84756 355068 84812 355078
rect 84756 354988 84812 355012
rect 84756 354922 84812 354932
rect 84644 305722 84700 305732
rect 83188 302428 83244 302466
rect 83188 302362 83244 302372
rect 76356 301462 76412 301472
rect 80276 290332 80332 290342
rect 78820 290108 78876 290118
rect 78820 289648 78876 290052
rect 80276 290008 80332 290276
rect 80276 289942 80332 289952
rect 78820 289582 78876 289592
rect 76132 274168 76188 274178
rect 76132 273956 76188 274112
rect 76132 273890 76188 273900
rect 76244 274092 76300 274102
rect 76244 272612 76300 274036
rect 76244 272546 76300 272556
rect 76356 273980 76412 273990
rect 76132 271268 76188 271278
rect 76132 270748 76188 271212
rect 76132 270682 76188 270692
rect 76244 270820 76300 270830
rect 76244 270568 76300 270764
rect 76244 270502 76300 270512
rect 76356 255276 76412 273924
rect 76468 273060 76524 273070
rect 76468 272188 76524 273004
rect 76468 272122 76524 272132
rect 84196 270844 84252 270854
rect 84196 270748 84252 270788
rect 84196 270682 84252 270692
rect 76356 255210 76412 255220
rect 76468 234388 76524 234398
rect 76356 233548 76412 233558
rect 76132 232956 76188 232966
rect 76132 231868 76188 232900
rect 76356 232508 76412 233492
rect 76356 232442 76412 232452
rect 76468 232228 76524 234332
rect 76132 231802 76188 231812
rect 76356 232172 76524 232228
rect 76244 231612 76300 231622
rect 76132 230428 76188 230438
rect 76132 230268 76188 230372
rect 76132 230202 76188 230212
rect 76244 230248 76300 231556
rect 76244 230182 76300 230192
rect 76356 229820 76412 232172
rect 84644 232092 84700 232102
rect 76468 232060 76524 232086
rect 76468 231982 76524 231992
rect 84644 231982 84700 231992
rect 76356 229754 76412 229764
rect 84644 207900 84700 207910
rect 84644 206668 84700 207844
rect 84756 207676 84812 207686
rect 84756 206848 84812 207620
rect 84756 206782 84812 206792
rect 84644 206602 84700 206612
rect 76132 191956 76188 191966
rect 76132 191842 76188 191852
rect 76132 191508 76188 191518
rect 76132 190828 76188 191452
rect 83860 191188 83916 191198
rect 76132 190762 76188 190772
rect 76468 191060 76524 191070
rect 76468 189928 76524 191004
rect 83860 190652 83916 191132
rect 83860 190586 83916 190596
rect 84308 190988 84364 190998
rect 76468 189862 76524 189872
rect 84308 189928 84364 190932
rect 84308 189862 84364 189872
rect 76132 189268 76188 189278
rect 76132 188668 76188 189212
rect 76132 188602 76188 188612
rect 76244 188820 76300 188830
rect 76244 188488 76300 188764
rect 84868 188668 84924 369796
rect 84980 230428 85036 412020
rect 85092 274168 85148 440468
rect 85204 306684 85260 578676
rect 686308 521164 686364 633444
rect 686532 562828 686588 673652
rect 686868 606508 686924 713972
rect 686868 606442 686924 606452
rect 686532 562762 686588 562772
rect 686756 553532 686812 553542
rect 686308 521098 686364 521108
rect 686420 526876 686476 526886
rect 686308 487228 686364 487238
rect 686196 406812 686252 406822
rect 85428 357196 85484 357206
rect 85204 306618 85260 306628
rect 85316 354844 85372 354854
rect 85092 274102 85148 274112
rect 85092 272188 85148 272198
rect 85092 272094 85148 272132
rect 85204 231868 85260 231906
rect 85204 231802 85260 231812
rect 84980 230362 85036 230372
rect 85316 191908 85372 354788
rect 85428 352828 85484 357140
rect 85428 352762 85484 352772
rect 393092 333788 393148 333798
rect 191492 333452 191548 333462
rect 173012 333228 173068 333238
rect 173012 332780 173068 333172
rect 188356 333228 188412 333238
rect 188356 332892 188412 333172
rect 188356 332826 188412 332836
rect 173012 332714 173068 332724
rect 118356 332668 118412 332678
rect 104132 324208 104188 324218
rect 104132 324090 104188 324100
rect 118356 324028 118412 332612
rect 186452 329196 186508 329206
rect 169652 328412 169708 328422
rect 118356 323962 118412 323972
rect 161028 324380 161084 324390
rect 151172 323932 151228 323942
rect 151172 323848 151228 323876
rect 151172 323782 151228 323792
rect 161028 323848 161084 324324
rect 166292 324208 166348 324218
rect 166292 324090 166348 324100
rect 169652 324156 169708 328356
rect 169652 324090 169708 324100
rect 186452 324156 186508 329140
rect 186452 324090 186508 324100
rect 191492 324156 191548 333396
rect 370468 333452 370524 333462
rect 353556 333340 353612 333350
rect 216132 333116 216188 333126
rect 205268 332780 205324 332790
rect 191492 324090 191548 324100
rect 201572 332668 201628 332678
rect 201572 324156 201628 332612
rect 201572 324090 201628 324100
rect 205268 324156 205324 332724
rect 205268 324090 205324 324100
rect 208292 332780 208348 332790
rect 208292 324156 208348 332724
rect 216132 332780 216188 333060
rect 216132 332714 216188 332724
rect 208292 324090 208348 324100
rect 213332 332668 213388 332678
rect 213332 324156 213388 332612
rect 320404 332668 320460 332678
rect 225876 328860 225932 328870
rect 213332 324090 213388 324100
rect 219380 328748 219436 328758
rect 219380 324156 219436 328692
rect 219380 324090 219436 324100
rect 225876 324156 225932 328804
rect 269556 328860 269612 328870
rect 258580 328524 258636 328534
rect 236740 328300 236796 328310
rect 225876 324090 225932 324100
rect 230244 327964 230300 327974
rect 230244 324156 230300 327908
rect 230244 324090 230300 324100
rect 236740 324156 236796 328244
rect 255780 325288 255836 325298
rect 236740 324090 236796 324100
rect 253540 325108 253596 325118
rect 253540 324156 253596 325052
rect 253540 324090 253596 324100
rect 255780 324156 255836 325232
rect 255780 324090 255836 324100
rect 258580 324156 258636 328468
rect 260932 326728 260988 326738
rect 258580 324090 258636 324100
rect 260148 325648 260204 325658
rect 260148 324044 260204 325592
rect 260932 324156 260988 326672
rect 263620 326368 263676 326378
rect 260932 324090 260988 324100
rect 262612 326188 262668 326198
rect 262612 324156 262668 326132
rect 262612 324090 262668 324100
rect 263620 324156 263676 326312
rect 263620 324090 263676 324100
rect 269556 324156 269612 328804
rect 269556 324090 269612 324100
rect 291508 328076 291564 328086
rect 291508 324156 291564 328020
rect 300244 327448 300300 327458
rect 300244 326620 300300 327392
rect 308980 327404 309036 327414
rect 299460 326548 299516 326558
rect 300244 326554 300300 326564
rect 300468 326620 300524 326630
rect 291508 324090 291564 324100
rect 295876 326284 295932 326294
rect 295876 324156 295932 326228
rect 295876 324090 295932 324100
rect 299460 324156 299516 326492
rect 300468 326284 300524 326564
rect 300468 326218 300524 326228
rect 299460 324090 299516 324100
rect 302260 326008 302316 326018
rect 302260 324156 302316 325952
rect 302260 324090 302316 324100
rect 306068 325468 306124 325478
rect 306068 324156 306124 325412
rect 306068 324090 306124 324100
rect 308980 324156 309036 327348
rect 317716 327292 317772 327302
rect 308980 324090 309036 324100
rect 311108 327268 311164 327278
rect 311108 324156 311164 327212
rect 311108 324090 311164 324100
rect 316932 324748 316988 324758
rect 161812 324028 161868 324038
rect 260148 323978 260204 323988
rect 161812 323932 161868 323972
rect 161812 323866 161868 323876
rect 316932 323932 316988 324692
rect 317716 324156 317772 327236
rect 320404 325648 320460 332612
rect 341796 332220 341852 332230
rect 336756 330316 336812 330326
rect 336644 328348 336700 328358
rect 334516 328300 334572 328310
rect 334404 327740 334460 327750
rect 334292 327628 334348 327638
rect 334180 327088 334236 327098
rect 320404 325582 320460 325592
rect 333172 326908 333228 326918
rect 317716 324090 317772 324100
rect 325780 324568 325836 324578
rect 325780 324044 325836 324512
rect 325780 323978 325836 323988
rect 332276 324388 332332 324398
rect 316932 323866 316988 323876
rect 332276 323932 332332 324332
rect 333172 324156 333228 326852
rect 333172 324090 333228 324100
rect 334180 324044 334236 327032
rect 334292 326368 334348 327572
rect 334292 326302 334348 326312
rect 334404 326188 334460 327684
rect 334516 326728 334572 328244
rect 334516 326662 334572 326672
rect 335972 327068 336028 327078
rect 334404 326122 334460 326132
rect 335972 325108 336028 327012
rect 335972 325042 336028 325052
rect 336644 324156 336700 328292
rect 336756 325288 336812 330260
rect 336756 325222 336812 325232
rect 340452 325648 340508 325658
rect 336644 324090 336700 324100
rect 334180 323978 334236 323988
rect 340452 324044 340508 325592
rect 341796 324156 341852 332164
rect 343476 327964 343980 327988
rect 343476 327932 343924 327964
rect 343476 327852 343532 327932
rect 343924 327898 343980 327908
rect 343476 327786 343532 327796
rect 353556 325724 353612 333284
rect 367892 332780 367948 332790
rect 353556 325658 353612 325668
rect 353780 330428 353836 330438
rect 341796 324090 341852 324100
rect 347620 325288 347676 325298
rect 347620 324156 347676 325232
rect 347620 324090 347676 324100
rect 347732 324380 347788 324390
rect 340452 323978 340508 323988
rect 332276 323866 332332 323876
rect 347732 323932 347788 324324
rect 353780 324380 353836 330372
rect 365652 328636 365708 328646
rect 358708 327740 358764 327750
rect 353780 324314 353836 324324
rect 357028 326728 357084 326738
rect 357028 324156 357084 326672
rect 358708 325648 358764 327684
rect 358708 325582 358764 325592
rect 357028 324090 357084 324100
rect 358484 325108 358540 325118
rect 358484 324156 358540 325052
rect 358484 324090 358540 324100
rect 365652 324156 365708 328580
rect 367892 328348 367948 332724
rect 367892 328282 367948 328292
rect 369460 328528 369516 328538
rect 367892 327628 367948 327638
rect 367892 325468 367948 327572
rect 367892 325402 367948 325412
rect 365652 324090 365708 324100
rect 365764 324928 365820 324938
rect 365764 324044 365820 324872
rect 369460 324156 369516 328472
rect 370468 324492 370524 333396
rect 378756 331996 378812 332006
rect 377860 328412 377916 328422
rect 376852 327628 376908 327638
rect 376740 326284 376796 326294
rect 370468 324426 370524 324436
rect 374276 325468 374332 325478
rect 369460 324090 369516 324100
rect 374276 324044 374332 325412
rect 376516 325052 376572 325062
rect 376516 324380 376572 324996
rect 376516 324314 376572 324324
rect 376740 324380 376796 326228
rect 376740 324314 376796 324324
rect 365764 323978 365820 323988
rect 371588 324028 371644 324038
rect 347732 323866 347788 323876
rect 374276 323978 374332 323988
rect 371588 323932 371644 323972
rect 371588 323866 371644 323876
rect 376852 323932 376908 327572
rect 377188 324152 377804 324208
rect 377188 324044 377244 324152
rect 377188 323978 377244 323988
rect 376852 323866 376908 323876
rect 377300 323932 377356 323942
rect 161028 323782 161084 323792
rect 159572 321244 159628 321254
rect 93828 320968 93884 320978
rect 92372 292236 92428 292246
rect 92372 270568 92428 292180
rect 93156 292012 93212 292022
rect 92372 270502 92428 270512
rect 92596 290668 92652 290678
rect 85316 191842 85372 191852
rect 92372 206668 92428 206678
rect 90356 191324 90412 191334
rect 90356 191188 90412 191268
rect 90356 191122 90412 191132
rect 84868 188602 84924 188612
rect 76244 188422 76300 188432
rect 92372 80892 92428 206612
rect 92596 191008 92652 290612
rect 93156 230248 93212 291956
rect 93380 291448 93436 291458
rect 93156 230182 93212 230192
rect 93268 289108 93324 289118
rect 92596 190942 92652 190952
rect 93156 206848 93212 206858
rect 93156 83008 93212 206792
rect 93268 188488 93324 289052
rect 93380 234388 93436 291392
rect 93380 234322 93436 234332
rect 93268 188422 93324 188432
rect 93156 82942 93212 82952
rect 92372 80826 92428 80836
rect 93828 79100 93884 320912
rect 159572 320968 159628 321188
rect 159572 320902 159628 320912
rect 159796 316316 159852 316326
rect 159796 314187 159852 316260
rect 159796 314131 159964 314187
rect 159684 311388 159740 311398
rect 99092 308188 99148 308198
rect 99092 307468 99148 308132
rect 154644 308008 154700 308018
rect 102452 307828 102508 307838
rect 99092 307402 99148 307412
rect 100772 307468 100828 307478
rect 100772 280924 100828 307412
rect 102452 307468 102508 307772
rect 102452 307402 102508 307412
rect 117908 291628 117964 291638
rect 117908 291116 117964 291572
rect 117908 291050 117964 291060
rect 100772 280858 100828 280868
rect 153748 281932 153804 281942
rect 153748 280700 153804 281876
rect 153748 280634 153804 280644
rect 153972 281260 154028 281270
rect 153972 280700 154028 281204
rect 154644 280924 154700 307952
rect 159684 306908 159740 311332
rect 159684 306842 159740 306852
rect 159796 307648 159852 307658
rect 154644 280858 154700 280868
rect 159796 280924 159852 307592
rect 159908 305900 159964 314131
rect 248500 308700 248556 308710
rect 162932 308588 162988 308598
rect 162932 308188 162988 308532
rect 164724 308588 164780 308598
rect 162932 308122 162988 308132
rect 164612 308476 164668 308486
rect 164612 307828 164668 308420
rect 164612 307762 164668 307772
rect 164724 307468 164780 308532
rect 166180 308588 166236 308598
rect 166180 308028 166236 308532
rect 193172 308588 193228 308598
rect 166180 307962 166236 307972
rect 181412 308476 181468 308486
rect 164724 307402 164780 307412
rect 165396 307828 165452 307838
rect 159908 305834 159964 305844
rect 165396 290444 165452 307772
rect 165396 290378 165452 290388
rect 165620 307468 165676 307478
rect 165620 288204 165676 307412
rect 181412 307468 181468 308420
rect 183092 308476 183148 308486
rect 181412 307402 181468 307412
rect 181636 308188 181692 308198
rect 173236 291900 173292 291910
rect 173236 291628 173292 291844
rect 173236 291562 173292 291572
rect 165620 288138 165676 288148
rect 168420 282044 168476 282054
rect 159796 280858 159852 280868
rect 162484 281260 162540 281270
rect 153972 280634 154028 280644
rect 162484 280700 162540 281204
rect 168420 281260 168476 281988
rect 173796 281932 173852 281942
rect 173796 281596 173852 281876
rect 173796 281530 173852 281540
rect 168420 281194 168476 281204
rect 181636 280924 181692 308132
rect 183092 307828 183148 308420
rect 190596 308364 190652 308374
rect 190596 308008 190652 308308
rect 190596 307942 190652 307952
rect 190820 308364 190876 308374
rect 190820 307916 190876 308308
rect 190820 307850 190876 307860
rect 183092 307762 183148 307772
rect 193172 307648 193228 308532
rect 203252 308588 203308 308598
rect 203252 308188 203308 308532
rect 238420 308588 238476 308598
rect 203252 308122 203308 308132
rect 206612 308476 206668 308486
rect 193172 307582 193228 307592
rect 196532 307648 196588 307658
rect 196532 282156 196588 307592
rect 201348 307468 201404 307478
rect 201348 303324 201404 307412
rect 206612 307468 206668 308420
rect 209972 308476 210028 308486
rect 209972 307648 210028 308420
rect 209972 307582 210028 307592
rect 234612 308364 234668 308374
rect 206612 307402 206668 307412
rect 234612 307468 234668 308308
rect 238420 308008 238476 308532
rect 238420 307942 238476 307952
rect 241780 308476 241836 308486
rect 241780 307648 241836 308420
rect 248500 307828 248556 308644
rect 321636 308700 322140 308728
rect 321692 308672 322084 308700
rect 321636 308634 321692 308644
rect 322084 308634 322140 308644
rect 342580 308700 342636 308710
rect 297220 308588 297276 308598
rect 261940 308476 261996 308486
rect 248500 307762 248556 307772
rect 251972 308008 252028 308018
rect 251972 307804 252028 307952
rect 251972 307738 252028 307748
rect 241780 307582 241836 307592
rect 234612 307402 234668 307412
rect 245252 307468 245308 307478
rect 201348 303258 201404 303268
rect 196532 282090 196588 282100
rect 196644 281596 196700 281606
rect 185780 281372 185836 281382
rect 185780 281148 185836 281316
rect 185780 281082 185836 281092
rect 196644 281036 196700 281540
rect 196644 280970 196700 280980
rect 196756 281372 196812 281382
rect 181636 280858 181692 280868
rect 196756 280924 196812 281316
rect 196756 280858 196812 280868
rect 245252 280924 245308 307412
rect 261940 307468 261996 308420
rect 265300 308476 265356 308486
rect 261940 307402 261996 307412
rect 262052 307648 262108 307658
rect 262052 282156 262108 307592
rect 265300 307648 265356 308420
rect 282100 308476 282156 308486
rect 282100 308008 282156 308420
rect 282100 307942 282156 307952
rect 265300 307582 265356 307592
rect 272132 307828 272188 307838
rect 262052 282090 262108 282100
rect 245252 280858 245308 280868
rect 272132 280924 272188 307772
rect 285572 307468 285628 307478
rect 285572 303772 285628 307412
rect 297220 307468 297276 308532
rect 297220 307402 297276 307412
rect 300692 308588 300748 308598
rect 285572 303706 285628 303716
rect 286020 302204 286076 302214
rect 285572 302092 285628 302102
rect 285572 301708 285628 302036
rect 286020 301888 286076 302148
rect 286020 301822 286076 301832
rect 285572 301642 285628 301652
rect 285796 301644 285852 301654
rect 285796 300808 285852 301588
rect 285796 300742 285852 300752
rect 292292 300636 292348 300646
rect 292292 299548 292348 300580
rect 292292 299482 292348 299492
rect 294532 300636 294588 300646
rect 294532 299368 294588 300580
rect 299012 300636 299068 300646
rect 299012 300088 299068 300580
rect 300692 300188 300748 308532
rect 307636 308588 307692 308598
rect 303940 307648 303996 307658
rect 303940 307468 303996 307592
rect 303940 307402 303996 307412
rect 300692 300122 300748 300132
rect 302596 300636 302652 300646
rect 299012 300022 299068 300032
rect 294532 299302 294588 299312
rect 302596 299188 302652 300580
rect 302820 300636 302876 300646
rect 302820 299908 302876 300580
rect 302820 299842 302876 299852
rect 302596 299122 302652 299132
rect 274036 282044 274092 282054
rect 274036 281036 274092 281988
rect 274036 280970 274092 280980
rect 272132 280858 272188 280868
rect 307636 280812 307692 308532
rect 317380 308588 317436 308598
rect 313796 308476 313852 308486
rect 313796 307648 313852 308420
rect 313796 307582 313852 307592
rect 316820 308008 316876 308018
rect 310996 297276 311052 297286
rect 310996 295768 311052 297220
rect 310996 295702 311052 295712
rect 316820 281932 316876 307952
rect 317380 307828 317436 308532
rect 320740 308588 320796 308598
rect 320740 308008 320796 308532
rect 320740 307942 320796 307952
rect 321860 308588 321916 308598
rect 317380 307762 317436 307772
rect 320964 292236 321020 292246
rect 320964 291808 321020 292180
rect 321188 292236 321244 292246
rect 321188 291988 321244 292180
rect 321188 291922 321244 291932
rect 321412 292236 321468 292246
rect 320964 291742 321020 291752
rect 321412 291628 321468 292180
rect 321412 291562 321468 291572
rect 321860 290667 321916 308532
rect 334180 308476 334236 308486
rect 330036 308364 330092 308374
rect 330036 307468 330092 308308
rect 334180 308188 334236 308420
rect 334180 308122 334236 308132
rect 336196 308476 336252 308486
rect 330036 307402 330092 307412
rect 335860 302316 335916 302326
rect 335636 296828 335692 296838
rect 334628 296716 334684 296726
rect 321636 290611 321916 290667
rect 334404 295768 334460 295778
rect 316820 281866 316876 281876
rect 320628 282044 320684 282054
rect 320628 281708 320684 281988
rect 320628 281642 320684 281652
rect 321636 281036 321692 290611
rect 327908 285292 327964 285302
rect 327684 284956 327740 284966
rect 327684 284068 327740 284900
rect 327908 284788 327964 285236
rect 327908 284722 327964 284732
rect 329588 284956 329644 284966
rect 329588 284248 329644 284900
rect 329588 284182 329644 284192
rect 327684 284002 327740 284012
rect 334404 282268 334460 295712
rect 334404 282202 334460 282212
rect 334628 282156 334684 296660
rect 334628 282090 334684 282100
rect 335636 281260 335692 296772
rect 335860 281820 335916 302260
rect 336196 294812 336252 308420
rect 337428 308140 337484 308150
rect 336196 294746 336252 294756
rect 336756 307828 336812 307838
rect 335972 294148 336028 294158
rect 335972 291448 336028 294092
rect 336756 293244 336812 307772
rect 336980 307648 337036 307658
rect 336980 296492 337036 307592
rect 337204 307468 337260 307478
rect 337204 300524 337260 307412
rect 337204 300458 337260 300468
rect 337428 296604 337484 308084
rect 342580 303508 342636 308644
rect 342580 303442 342636 303452
rect 344260 308700 344316 308710
rect 344260 303328 344316 308644
rect 344260 303262 344316 303272
rect 357700 308700 357756 308710
rect 357700 303148 357756 308644
rect 377300 308700 377356 323876
rect 377300 308634 377356 308644
rect 377748 308700 377804 324152
rect 377860 324156 377916 328356
rect 377860 324090 377916 324100
rect 378644 323932 378700 323942
rect 378644 322588 378700 323876
rect 378644 322522 378700 322532
rect 378196 322228 378252 322238
rect 377748 308634 377804 308644
rect 377972 317368 378028 317378
rect 362740 308476 362796 308486
rect 362740 304048 362796 308420
rect 362740 303982 362796 303992
rect 364420 308476 364476 308486
rect 364420 303868 364476 308420
rect 369460 308476 369516 308486
rect 369460 307828 369516 308420
rect 377860 308476 377916 308486
rect 369460 307762 369516 307772
rect 377636 308188 377692 308198
rect 364420 303802 364476 303812
rect 357700 303082 357756 303092
rect 354900 301888 354956 301906
rect 354900 301802 354956 301812
rect 356132 301708 356188 301718
rect 356132 301420 356188 301652
rect 356132 301354 356188 301364
rect 352772 300808 352828 300818
rect 337428 296538 337484 296548
rect 338436 299548 338492 299558
rect 336980 296426 337036 296436
rect 336756 293178 336812 293188
rect 335972 291382 336028 291392
rect 337540 289212 337596 289222
rect 337540 289108 337596 289156
rect 337540 289042 337596 289052
rect 335860 281754 335916 281764
rect 335636 281194 335692 281204
rect 321636 280970 321692 280980
rect 307636 280746 307692 280756
rect 162484 280634 162540 280644
rect 338436 280700 338492 299492
rect 343476 299368 343532 299378
rect 342804 281708 342860 281718
rect 342804 281260 342860 281652
rect 343476 281596 343532 299312
rect 343476 281530 343532 281540
rect 343700 298284 343756 298294
rect 342804 281194 342860 281204
rect 343700 280924 343756 298228
rect 352772 281708 352828 300752
rect 352772 281642 352828 281652
rect 377636 281260 377692 308132
rect 377860 307648 377916 308420
rect 377860 307582 377916 307592
rect 377860 307468 377916 307478
rect 377860 307374 377916 307412
rect 377972 284732 378028 317312
rect 377972 284666 378028 284676
rect 378084 308252 378140 308262
rect 377636 281194 377692 281204
rect 343700 280858 343756 280868
rect 378084 280924 378140 308196
rect 378196 294868 378252 322172
rect 378756 309988 378812 331940
rect 388276 328860 388332 328870
rect 388276 326548 388332 328804
rect 393092 328528 393148 333732
rect 487956 333340 488012 333350
rect 453684 332668 453740 332678
rect 393092 328462 393148 328472
rect 405748 328860 405804 328870
rect 388276 326482 388332 326492
rect 382004 325836 382060 325846
rect 382004 324928 382060 325780
rect 405748 325468 405804 328804
rect 453572 327516 453628 327526
rect 453572 327448 453628 327460
rect 453572 327382 453628 327392
rect 405748 325402 405804 325412
rect 453684 325288 453740 332612
rect 470372 326172 470428 326182
rect 470372 326008 470428 326116
rect 470372 325942 470428 325952
rect 453684 325222 453740 325232
rect 487956 325108 488012 333284
rect 497364 333340 497420 333350
rect 497364 327268 497420 333284
rect 497364 327202 497420 327212
rect 533092 333340 533148 333350
rect 533092 327088 533148 333284
rect 533092 327022 533148 327032
rect 551684 332668 551740 332678
rect 551684 326908 551740 332612
rect 551684 326842 551740 326852
rect 623252 332668 623308 332678
rect 623252 326728 623308 332612
rect 672308 332556 672364 332566
rect 656740 329196 656796 329206
rect 656740 327628 656796 329140
rect 656740 327562 656796 327572
rect 623252 326662 623308 326672
rect 487956 325042 488012 325052
rect 505540 324940 505596 324950
rect 382004 324862 382060 324872
rect 485492 324928 485548 324938
rect 485492 324028 485548 324872
rect 505540 324748 505596 324884
rect 655508 324940 655564 324950
rect 655508 324846 655564 324872
rect 505540 324682 505596 324692
rect 537572 324604 537628 324614
rect 537572 324502 537628 324512
rect 554372 324492 554428 324502
rect 554372 324388 554428 324436
rect 554372 324322 554428 324332
rect 485492 323962 485548 323972
rect 379540 323932 379596 323942
rect 379540 322768 379596 323876
rect 380324 323148 380380 323158
rect 380324 322948 380380 323092
rect 380324 322882 380380 322892
rect 379540 322702 379596 322712
rect 379764 322252 379820 322262
rect 379764 322158 379820 322172
rect 379876 319564 379932 319574
rect 379876 319462 379932 319472
rect 557732 319528 557788 319538
rect 557732 319452 557788 319472
rect 557732 319386 557788 319396
rect 379764 317368 379820 317378
rect 379764 317258 379820 317268
rect 379764 314860 379820 314870
rect 378756 309922 378812 309932
rect 379428 314804 379764 314848
rect 379428 314792 379820 314804
rect 379428 308252 379484 314792
rect 672308 314187 672364 332500
rect 672420 324156 672476 324166
rect 672420 322948 672476 324100
rect 672420 322882 672476 322892
rect 672644 324044 672700 324054
rect 672644 322768 672700 323988
rect 672644 322702 672700 322712
rect 672756 322588 672812 322598
rect 672756 322494 672812 322532
rect 672196 314131 672364 314187
rect 379764 312508 379820 312518
rect 379764 312396 379820 312452
rect 460292 312508 460348 312518
rect 460292 312414 460348 312452
rect 379764 312330 379820 312340
rect 664356 309988 664412 309998
rect 379764 309932 379820 309942
rect 379764 309808 379820 309876
rect 379540 309752 379820 309808
rect 379540 309268 379596 309752
rect 379540 309202 379596 309212
rect 458612 309268 458668 309298
rect 458612 309194 458668 309204
rect 379428 308186 379484 308196
rect 426692 308008 426748 308018
rect 426692 307468 426748 307952
rect 532420 307828 532476 307842
rect 426692 307402 426748 307412
rect 462756 307804 462812 307814
rect 385924 303996 385980 304006
rect 385924 302608 385980 303940
rect 385924 302542 385980 302552
rect 381780 300088 381836 300098
rect 381780 299740 381836 300032
rect 381780 299674 381836 299684
rect 389732 299908 389788 299918
rect 389732 299740 389788 299852
rect 389732 299674 389788 299684
rect 378196 294802 378252 294812
rect 391412 299188 391468 299198
rect 391412 282156 391468 299132
rect 397460 296604 397516 296614
rect 391412 282090 391468 282100
rect 397236 296492 397292 296502
rect 397236 281820 397292 296436
rect 397236 281754 397292 281764
rect 397460 281708 397516 296548
rect 461972 292168 462028 292178
rect 428820 291988 428876 291998
rect 428820 291900 428876 291932
rect 428820 291834 428876 291844
rect 428596 291808 428652 291826
rect 428596 291722 428652 291732
rect 430388 291628 430444 291638
rect 430388 291564 430444 291572
rect 430388 291498 430444 291508
rect 444052 284788 444108 284798
rect 444052 284620 444108 284732
rect 444052 284554 444108 284564
rect 446628 284248 446684 284258
rect 445284 284068 445340 284078
rect 445284 282156 445340 284012
rect 445284 282090 445340 282100
rect 446628 282156 446684 284192
rect 446628 282090 446684 282100
rect 397460 281642 397516 281652
rect 378084 280858 378140 280868
rect 461972 280924 462028 292112
rect 462756 292168 462812 307748
rect 532420 307738 532476 307748
rect 550116 307648 550172 307658
rect 538580 307244 538636 307254
rect 520548 304048 520604 304058
rect 520548 303930 520604 303940
rect 482132 303884 482188 303894
rect 474516 303508 474572 303518
rect 465332 292348 465388 292358
rect 465332 292254 465388 292292
rect 462756 292102 462812 292112
rect 472052 290368 472108 290378
rect 472052 290266 472108 290276
rect 468580 288316 468636 288326
rect 468580 287308 468636 288260
rect 474516 288204 474572 303452
rect 479556 303328 479612 303338
rect 477876 303100 477932 303110
rect 475412 290556 475468 290566
rect 475412 290462 475468 290492
rect 468580 287176 468636 287252
rect 469140 288092 469196 288102
rect 469140 287488 469196 288036
rect 469140 287308 469196 287432
rect 469140 287242 469196 287252
rect 474516 287308 474572 288148
rect 474516 287242 474572 287252
rect 477876 290188 477932 303044
rect 461972 280858 462028 280868
rect 477876 280924 477932 290132
rect 479556 289324 479612 303272
rect 479556 289258 479612 289268
rect 482132 294328 482188 303828
rect 522340 303868 522396 303878
rect 522340 303772 522396 303812
rect 522340 303706 522396 303716
rect 477876 280858 477932 280868
rect 482132 280924 482188 294272
rect 506436 303148 506492 303158
rect 488852 292908 488908 292918
rect 488852 292814 488908 292832
rect 498932 292796 498988 292806
rect 498932 292708 498988 292740
rect 498932 292642 498988 292652
rect 497252 292572 497308 292582
rect 497252 292462 497308 292472
rect 506436 291564 506492 303092
rect 537572 293968 537628 293978
rect 510692 293068 510748 293078
rect 510692 292954 510748 292964
rect 534212 291676 534268 291686
rect 534212 291562 534268 291572
rect 506436 291448 506492 291508
rect 506436 291382 506492 291392
rect 532532 291340 532588 291350
rect 532532 291268 532588 291284
rect 532532 291202 532588 291212
rect 521332 291088 521388 291098
rect 521332 291004 521388 291032
rect 521332 290938 521388 290948
rect 535892 290908 535948 290930
rect 535892 290826 535948 290836
rect 482132 280858 482188 280868
rect 537572 280924 537628 293912
rect 538580 293968 538636 307188
rect 538580 293248 538636 293912
rect 541716 302608 541772 302618
rect 539252 293468 539308 293478
rect 539252 293362 539308 293372
rect 538580 293182 538636 293192
rect 541716 292236 541772 302552
rect 550116 293916 550172 307592
rect 551012 307468 551068 307478
rect 551012 307374 551068 307412
rect 652260 302428 652316 302438
rect 550116 293608 550172 293860
rect 550116 293542 550172 293552
rect 557732 294868 557788 294878
rect 541716 292170 541772 292180
rect 537572 280858 537628 280868
rect 557732 280924 557788 294812
rect 611380 294328 611436 294338
rect 606116 292908 606172 292918
rect 606116 290108 606172 292852
rect 606228 292888 606284 292898
rect 606228 290728 606284 292832
rect 609924 292168 609980 292178
rect 609812 291988 609868 291998
rect 606228 290662 606284 290672
rect 606340 290668 606396 290678
rect 606340 290548 606396 290612
rect 606340 290482 606396 290492
rect 607796 290444 607852 290454
rect 606340 290368 606396 290378
rect 606340 290220 606396 290312
rect 606340 290154 606396 290164
rect 607796 290220 607852 290388
rect 607796 290154 607852 290164
rect 608916 290332 608972 290342
rect 606116 290042 606172 290052
rect 600516 289548 600572 289558
rect 559188 288540 559244 288550
rect 559076 286188 559132 286198
rect 558852 283948 558908 283958
rect 558740 281260 558796 281270
rect 557732 280858 557788 280868
rect 558292 281036 558348 281046
rect 338436 280634 338492 280644
rect 558292 270507 558348 280980
rect 558628 280812 558684 280822
rect 558628 270507 558684 280756
rect 558740 272188 558796 281204
rect 558852 276508 558908 283892
rect 559076 279208 559132 286132
rect 559188 285627 559244 288484
rect 600516 287308 600572 289492
rect 608916 289100 608972 290276
rect 608916 289034 608972 289044
rect 600516 287242 600572 287252
rect 559188 285571 559356 285627
rect 559300 279692 559356 285571
rect 609812 283052 609868 291932
rect 609924 283276 609980 292112
rect 611380 290728 611436 294272
rect 644420 293608 644476 293618
rect 641508 293468 641564 293478
rect 638708 293428 638764 293438
rect 638148 293248 638204 293258
rect 628068 293068 628124 293078
rect 623252 292708 623308 292718
rect 622804 292528 622860 292538
rect 620676 291988 620732 291998
rect 611380 290662 611436 290672
rect 614740 290728 614796 290738
rect 614740 290668 614796 290672
rect 614292 290612 614796 290668
rect 620676 290728 620732 291932
rect 620676 290662 620732 290672
rect 614292 290548 614348 290612
rect 615636 290556 615692 290566
rect 614292 290482 614348 290492
rect 614404 290492 615468 290548
rect 611044 290368 611100 290378
rect 611044 290108 611100 290312
rect 614292 290368 614348 290378
rect 614404 290368 614460 290492
rect 614348 290312 614460 290368
rect 614516 290332 614572 290342
rect 614292 290302 614348 290312
rect 614516 290188 614572 290276
rect 614740 290220 614796 290230
rect 611044 290042 611100 290052
rect 611268 290132 611660 290188
rect 614516 290164 614740 290188
rect 614516 290132 614796 290164
rect 611268 289996 611324 290132
rect 611492 289996 611548 290006
rect 611268 289930 611324 289940
rect 611380 289940 611492 289996
rect 611604 289996 611660 290132
rect 615412 290108 615468 290492
rect 615636 290188 615692 290500
rect 616420 290548 616476 290558
rect 616420 290444 616476 290492
rect 616420 290378 616476 290388
rect 615636 290122 615692 290132
rect 617540 290368 617596 290378
rect 615412 290042 615468 290052
rect 617540 290108 617596 290312
rect 617540 290042 617596 290052
rect 611940 289996 611996 290006
rect 611604 289940 611940 289996
rect 611380 288876 611436 289940
rect 611492 289930 611548 289940
rect 611940 289930 611996 289940
rect 620676 289996 620732 290006
rect 620676 289772 620732 289940
rect 620676 289706 620732 289716
rect 622804 289772 622860 292472
rect 622804 289706 622860 289716
rect 623252 289772 623308 292652
rect 623252 289706 623308 289716
rect 626164 291448 626220 291458
rect 626164 289772 626220 291392
rect 626164 289706 626220 289716
rect 628068 289772 628124 293012
rect 628068 289706 628124 289716
rect 629076 293020 629132 293030
rect 629076 289772 629132 292964
rect 636692 291628 636748 291638
rect 636244 291268 636300 291278
rect 631988 291088 632044 291098
rect 631764 290108 631820 290118
rect 629188 289996 629244 290006
rect 629188 289772 629244 289940
rect 629300 289772 629356 289782
rect 629188 289716 629300 289772
rect 629076 289706 629132 289716
rect 629300 289706 629356 289716
rect 631764 289772 631820 290052
rect 631764 289706 631820 289716
rect 631988 289772 632044 291032
rect 631988 289706 632044 289716
rect 636244 289772 636300 291212
rect 636244 289706 636300 289716
rect 636692 289772 636748 291572
rect 637252 290908 637308 290918
rect 637252 290556 637308 290852
rect 637252 290490 637308 290500
rect 636692 289706 636748 289716
rect 638148 289772 638204 293192
rect 638148 289706 638204 289716
rect 638708 289772 638764 293372
rect 641060 293356 641116 293366
rect 640612 293244 640668 293254
rect 638708 289706 638764 289716
rect 640052 293132 640108 293142
rect 640052 289772 640108 293076
rect 640052 289706 640108 289716
rect 640612 289772 640668 293188
rect 640612 289706 640668 289716
rect 641060 289772 641116 293300
rect 641060 289706 641116 289716
rect 641508 289772 641564 293412
rect 641508 289706 641564 289716
rect 642516 291808 642572 291818
rect 642516 289772 642572 291752
rect 642516 289706 642572 289716
rect 644196 289996 644252 290006
rect 644196 289772 644252 289940
rect 644196 289706 644252 289716
rect 644420 289772 644476 293552
rect 646548 292348 646604 292358
rect 646548 290556 646604 292292
rect 646548 290490 646604 290500
rect 644420 289706 644476 289716
rect 652260 289772 652316 302372
rect 664356 301756 664412 309932
rect 670628 306572 670684 306582
rect 670628 302427 670684 306516
rect 670628 302371 671020 302427
rect 664356 301690 664412 301700
rect 670404 301528 670460 301538
rect 670292 292348 670348 292358
rect 670292 290908 670348 292292
rect 670180 290852 670348 290908
rect 669844 290728 669900 290738
rect 667492 290548 667548 290558
rect 666932 290332 666988 290342
rect 666932 290108 666988 290276
rect 666932 290042 666988 290052
rect 667044 290188 667100 290198
rect 652596 290008 652652 290018
rect 652596 289884 652652 289952
rect 661668 290008 661724 290018
rect 652596 289818 652652 289828
rect 655508 289828 655564 289838
rect 652260 289706 652316 289716
rect 655508 289706 655564 289716
rect 658308 289828 658364 289838
rect 658308 289706 658364 289716
rect 661668 289772 661724 289952
rect 667044 289828 667100 290132
rect 667044 289762 667100 289772
rect 667268 289828 667324 289838
rect 661668 289706 661724 289716
rect 667268 289706 667324 289716
rect 667492 289772 667548 290492
rect 669844 290556 669900 290672
rect 669844 290490 669900 290500
rect 670180 290548 670236 290852
rect 670404 290667 670460 301472
rect 670180 290482 670236 290492
rect 670292 290611 670460 290667
rect 670292 290444 670348 290611
rect 670292 290378 670348 290388
rect 670964 290008 671020 302371
rect 671188 301532 671244 301542
rect 670964 289942 671020 289952
rect 671076 291988 671132 291998
rect 667492 289706 667548 289716
rect 671076 289772 671132 291932
rect 671188 290108 671244 301476
rect 671188 290042 671244 290052
rect 671300 294148 671356 294158
rect 671300 289884 671356 294092
rect 672196 290188 672252 314131
rect 672196 290122 672252 290132
rect 671300 289818 671356 289828
rect 672308 289884 672364 289894
rect 671076 289706 671132 289716
rect 671636 289772 671692 289782
rect 672308 289762 672364 289772
rect 611380 288810 611436 288820
rect 611044 288204 611100 288214
rect 611044 287488 611100 288148
rect 611044 287422 611100 287432
rect 609924 283210 609980 283220
rect 609812 282986 609868 282996
rect 559300 279626 559356 279636
rect 559076 279152 559356 279208
rect 559300 276780 559356 279152
rect 671636 278907 671692 289716
rect 671860 289108 671916 289118
rect 671860 288428 671916 289052
rect 671860 288362 671916 288372
rect 671636 278851 671804 278907
rect 671748 276892 671804 278851
rect 671748 276826 671804 276836
rect 559300 276714 559356 276724
rect 558852 276452 559356 276508
rect 559300 273532 559356 276452
rect 559300 273466 559356 273476
rect 558740 272132 559356 272188
rect 558292 270451 558460 270507
rect 558404 268768 558460 270451
rect 558404 268702 558460 268712
rect 558516 270451 558684 270507
rect 559300 270508 559356 272132
rect 558516 257248 558572 270451
rect 559300 270442 559356 270452
rect 559300 268768 559356 268778
rect 559300 265132 559356 268712
rect 559300 265066 559356 265076
rect 559300 263452 559356 263462
rect 559300 259048 559356 263396
rect 559300 258992 559468 259048
rect 559412 258747 559468 258992
rect 559412 258691 559580 258747
rect 558516 257182 558572 257192
rect 559300 257248 559356 257258
rect 559300 256172 559356 257192
rect 559300 256106 559356 256116
rect 559524 246988 559580 258691
rect 559524 246922 559580 246932
rect 559300 243628 559356 243638
rect 559300 220107 559356 243572
rect 558292 220051 559356 220107
rect 335972 83008 336028 83018
rect 335972 80780 336028 82952
rect 558292 81564 558348 220051
rect 559300 209244 559356 209254
rect 559300 196587 559356 209188
rect 558964 196531 559356 196587
rect 558404 185788 558460 185798
rect 558404 143668 558460 185732
rect 558964 185248 559020 196531
rect 559300 186172 559356 186182
rect 559300 185428 559356 186116
rect 559636 185788 559692 185798
rect 559636 185724 559692 185732
rect 559636 185658 559692 185668
rect 558852 185192 559020 185248
rect 559076 185372 559356 185428
rect 558628 184888 558684 184898
rect 558628 161307 558684 184832
rect 558852 176428 558908 185192
rect 559076 184888 559132 185372
rect 559076 184822 559132 184832
rect 559300 176428 559356 176438
rect 558852 176372 559300 176428
rect 559300 176362 559356 176372
rect 671748 161532 671804 161542
rect 671748 161307 671804 161476
rect 558628 161251 559356 161307
rect 559300 147420 559356 161251
rect 671636 161251 671804 161307
rect 559300 147354 559356 147364
rect 585396 158956 585452 158966
rect 558404 143602 558460 143612
rect 559300 143668 559356 143678
rect 558516 142588 558572 142598
rect 558404 96688 558460 96698
rect 558404 82288 558460 96632
rect 558404 82222 558460 82232
rect 558516 81676 558572 142532
rect 559300 138572 559356 143612
rect 559412 143388 559468 143398
rect 559412 142588 559468 143332
rect 559412 142522 559468 142532
rect 585172 143052 585228 143062
rect 559412 142048 559468 142058
rect 559412 141708 559468 141992
rect 559412 141642 559468 141652
rect 559300 138506 559356 138516
rect 559300 126028 559356 126038
rect 558740 125972 559300 126027
rect 558740 125971 559356 125972
rect 558628 90748 558684 90758
rect 558628 82108 558684 90692
rect 558628 82042 558684 82052
rect 558516 81610 558572 81620
rect 558292 81498 558348 81508
rect 558740 81228 558796 125971
rect 559300 125962 559356 125971
rect 559300 114268 559356 114278
rect 558964 114212 559300 114267
rect 558964 114211 559356 114212
rect 558964 81340 559020 114211
rect 559300 114202 559356 114211
rect 559300 110908 559356 110918
rect 559188 110852 559300 110908
rect 559188 90747 559244 110852
rect 559300 110842 559356 110852
rect 559300 105196 559356 105206
rect 559300 96688 559356 105140
rect 559300 96622 559356 96632
rect 559076 90691 559244 90747
rect 559300 90748 559356 90786
rect 559076 81452 559132 90691
rect 559300 90682 559356 90692
rect 559300 87500 559356 87510
rect 559300 84988 559356 87444
rect 559188 84932 559356 84988
rect 559188 81928 559244 84932
rect 559188 81862 559244 81872
rect 559300 84476 559356 84486
rect 559300 81788 559356 84420
rect 559300 81722 559356 81732
rect 585172 81788 585228 142996
rect 585396 82288 585452 158900
rect 585396 82222 585452 82232
rect 585620 147532 585676 147542
rect 585620 82108 585676 147476
rect 585620 82042 585676 82052
rect 585844 145292 585900 145302
rect 585844 81928 585900 145236
rect 671636 141868 671692 161251
rect 671748 152348 671804 152358
rect 671748 142716 671804 152292
rect 671748 142650 671804 142660
rect 671860 145404 671916 145414
rect 671860 142408 671916 145348
rect 671860 142352 672028 142408
rect 671860 142156 671916 142166
rect 671860 142048 671916 142100
rect 671860 141982 671916 141992
rect 671636 141802 671692 141812
rect 671972 141596 672028 142352
rect 671972 141530 672028 141540
rect 671748 141148 671804 141158
rect 671748 141054 671804 141092
rect 618884 140068 618940 140078
rect 619108 140068 619164 140078
rect 618212 139804 618268 139814
rect 618212 83804 618268 139748
rect 618324 139708 618380 139718
rect 618324 85036 618380 139652
rect 618660 139580 618716 139590
rect 618548 139528 618604 139538
rect 618324 84970 618380 84980
rect 618436 134428 618492 134438
rect 618212 83738 618268 83748
rect 585844 81862 585900 81872
rect 585172 81722 585228 81732
rect 559076 81386 559132 81396
rect 558964 81274 559020 81284
rect 558740 81162 558796 81172
rect 335972 80714 336028 80724
rect 93828 79034 93884 79044
rect 324884 72156 324940 72166
rect 231252 71372 231308 71382
rect 176260 71308 176316 71318
rect 176260 70140 176316 71252
rect 176260 70074 176316 70084
rect 231252 70140 231308 71316
rect 324884 70768 324940 72100
rect 559412 72044 559468 72054
rect 324884 70702 324940 70712
rect 396116 71596 396172 71606
rect 257796 70588 257852 70598
rect 257796 70494 257852 70532
rect 396116 70588 396172 71540
rect 396116 70522 396172 70532
rect 494340 71488 494396 71498
rect 231252 70074 231308 70084
rect 494340 70140 494396 71432
rect 519652 71128 519708 71138
rect 494340 70074 494396 70084
rect 505876 70948 505932 70958
rect 505876 70140 505932 70892
rect 505876 70074 505932 70084
rect 519652 69804 519708 71072
rect 548436 70768 548492 70778
rect 539140 70588 539196 70598
rect 539140 70364 539196 70532
rect 539140 70298 539196 70308
rect 548436 70140 548492 70712
rect 559412 70588 559468 71988
rect 618436 71488 618492 134372
rect 618548 91308 618604 139472
rect 618548 91242 618604 91252
rect 618660 88732 618716 139524
rect 618772 123148 618828 123158
rect 618772 122668 618828 123092
rect 618772 122602 618828 122612
rect 618660 88666 618716 88676
rect 618884 87500 618940 140012
rect 618996 140012 619108 140068
rect 618996 139708 619052 140012
rect 619108 140002 619164 140012
rect 623364 140068 623420 140078
rect 623364 139962 623420 139972
rect 624708 140068 624764 140078
rect 624708 139962 624764 139972
rect 649348 140068 649404 140078
rect 631428 139916 631484 139926
rect 618996 139642 619052 139652
rect 619108 139888 619164 139898
rect 619108 95004 619164 139832
rect 631428 139822 631484 139832
rect 619332 139708 619388 139718
rect 632772 139708 632828 139730
rect 619332 97468 619388 139652
rect 622020 139692 622076 139702
rect 622020 139528 622076 139636
rect 632772 139626 632828 139636
rect 638820 139692 638876 139702
rect 619892 139468 619948 139478
rect 622020 139462 622076 139472
rect 622468 139528 622524 139538
rect 619892 100716 619948 139412
rect 622356 135660 622412 135670
rect 622244 135548 622300 135558
rect 621460 134540 621516 134550
rect 621348 134428 621404 134438
rect 620564 123452 620620 123462
rect 619892 100650 619948 100660
rect 620340 123340 620396 123350
rect 619332 97402 619388 97412
rect 619108 94938 619164 94948
rect 618884 87434 618940 87444
rect 618436 71422 618492 71432
rect 620340 80668 620396 123284
rect 620340 71308 620396 80612
rect 620564 80848 620620 123396
rect 621348 122968 621404 134372
rect 621348 122902 621404 122912
rect 621460 122788 621516 134484
rect 621460 122722 621516 122732
rect 622244 99388 622300 135492
rect 622356 100716 622412 135604
rect 622356 100650 622412 100660
rect 622244 99322 622300 99332
rect 622468 99208 622524 139472
rect 638820 139528 638876 139636
rect 638820 139462 638876 139472
rect 648452 139468 648508 139478
rect 622804 135436 622860 135446
rect 622692 135324 622748 135334
rect 622580 135212 622636 135222
rect 622580 100648 622636 135156
rect 622580 100582 622636 100592
rect 622692 100468 622748 135268
rect 622804 100492 622860 135380
rect 646324 127484 646380 127494
rect 646324 126748 646380 127428
rect 646324 126682 646380 126692
rect 646996 126028 647052 126038
rect 646996 125934 647052 125972
rect 626052 125916 626108 125926
rect 626052 124408 626108 125860
rect 628068 125916 628124 125926
rect 628068 124588 628124 125860
rect 628740 125916 628796 125926
rect 628740 124768 628796 125860
rect 641508 125916 641564 125926
rect 641508 124948 641564 125860
rect 641508 124882 641564 124892
rect 628740 124702 628796 124712
rect 628068 124522 628124 124532
rect 626052 124342 626108 124352
rect 642740 124228 642796 124238
rect 642740 123340 642796 124172
rect 648452 124228 648508 139412
rect 649348 131740 649404 140012
rect 649572 140068 649628 140078
rect 649460 136332 649516 136342
rect 649460 132748 649516 136276
rect 649460 132682 649516 132692
rect 649572 131852 649628 140012
rect 657076 140068 657132 140078
rect 657076 139962 657132 139972
rect 657748 140068 657804 140078
rect 657748 139962 657804 139972
rect 655732 139916 655788 139926
rect 649684 139888 649740 139898
rect 649684 131964 649740 139832
rect 655732 139822 655788 139832
rect 671188 139916 671244 139926
rect 669956 139804 670012 139814
rect 650916 139708 650972 139718
rect 650692 139692 650748 139702
rect 649796 136332 649852 136342
rect 649796 132328 649852 136276
rect 649908 136220 649964 136230
rect 649908 132524 649964 136164
rect 650020 136108 650076 136118
rect 650020 132636 650076 136052
rect 650132 134876 650188 134886
rect 650132 133196 650188 134820
rect 650132 133130 650188 133140
rect 650020 132570 650076 132580
rect 649908 132458 649964 132468
rect 650692 132412 650748 139636
rect 650804 139468 650860 139478
rect 650804 132688 650860 139412
rect 650804 132622 650860 132632
rect 650692 132346 650748 132356
rect 650916 132412 650972 139652
rect 656404 139708 656460 139730
rect 656404 139626 656460 139636
rect 666484 139692 666540 139702
rect 666484 139528 666540 139636
rect 666484 139462 666540 139472
rect 669620 138012 669676 138022
rect 669620 135212 669676 137956
rect 669844 137900 669900 137910
rect 669620 135146 669676 135156
rect 669732 137788 669788 137798
rect 669620 134988 669676 134998
rect 657972 132688 658028 132698
rect 657972 132570 658028 132580
rect 664580 132688 664636 132698
rect 664580 132570 664636 132580
rect 666820 132636 666876 132646
rect 659652 132524 659708 132534
rect 659652 132430 659708 132452
rect 650916 132346 650972 132356
rect 649796 132262 649852 132272
rect 653492 132328 653548 132338
rect 653492 132188 653548 132272
rect 666820 132328 666876 132580
rect 669620 132636 669676 134932
rect 669620 132570 669676 132580
rect 669732 132412 669788 137732
rect 669844 135388 669900 137844
rect 669956 135548 670012 139748
rect 670404 139692 670460 139702
rect 670068 139580 670124 139590
rect 670068 137787 670124 139524
rect 670404 137787 670460 139636
rect 671076 139528 671132 139538
rect 670852 139468 670908 139478
rect 670740 138796 670796 138806
rect 670068 137731 670236 137787
rect 670404 137731 670572 137787
rect 669956 135482 670012 135492
rect 669844 135332 670124 135388
rect 669956 135212 670012 135222
rect 669732 132346 669788 132356
rect 669844 135100 669900 135110
rect 666820 132262 666876 132272
rect 669844 132300 669900 135044
rect 669956 132508 670012 135156
rect 669956 132442 670012 132452
rect 669844 132234 669900 132244
rect 653492 132122 653548 132132
rect 649684 131898 649740 131908
rect 649572 131786 649628 131796
rect 649348 131674 649404 131684
rect 670068 131404 670124 135332
rect 670180 131516 670236 137731
rect 670404 137004 670460 137014
rect 670292 136892 670348 136902
rect 670292 132188 670348 136836
rect 670292 132122 670348 132132
rect 670404 131852 670460 136948
rect 670516 132524 670572 137731
rect 670740 132688 670796 138740
rect 670740 132622 670796 132632
rect 670852 132636 670908 139412
rect 670852 132570 670908 132580
rect 670964 139020 671020 139030
rect 670516 132458 670572 132468
rect 670404 131786 670460 131796
rect 670180 131450 670236 131460
rect 670068 131338 670124 131348
rect 665140 131068 665196 131078
rect 665140 130974 665196 131012
rect 670964 131068 671020 138964
rect 671076 132328 671132 139472
rect 671076 132262 671132 132272
rect 671188 131964 671244 139860
rect 686196 134428 686252 406756
rect 686308 220108 686364 487172
rect 686420 263900 686476 526820
rect 686644 433468 686700 433478
rect 686420 263834 686476 263844
rect 686532 340284 686588 340294
rect 686308 220042 686364 220052
rect 686196 134362 686252 134372
rect 671188 131898 671244 131908
rect 670964 131002 671020 131012
rect 654500 127596 654556 127606
rect 648452 124162 648508 124172
rect 654276 126812 654332 126822
rect 642740 123274 642796 123284
rect 647892 123340 647948 123366
rect 647892 123262 647948 123272
rect 651812 110548 651868 110558
rect 622804 100426 622860 100436
rect 628628 100648 628684 100658
rect 628628 100492 628684 100592
rect 649572 100648 649628 100658
rect 628628 100426 628684 100436
rect 631204 100492 631260 100506
rect 622692 100402 622748 100412
rect 649572 100492 649628 100592
rect 649572 100426 649628 100436
rect 631204 100402 631260 100412
rect 633780 100044 633836 100054
rect 633780 99388 633836 99988
rect 633780 99322 633836 99332
rect 635796 100044 635852 100054
rect 622468 99142 622524 99152
rect 635796 99208 635852 99988
rect 635796 99142 635852 99152
rect 639044 100044 639100 100054
rect 639044 99208 639100 99988
rect 641732 100044 641788 100054
rect 641732 99388 641788 99988
rect 644980 100044 645036 100054
rect 644980 99568 645036 99988
rect 644980 99502 645036 99512
rect 641732 99322 641788 99332
rect 639044 99142 639100 99152
rect 651812 86608 651868 110492
rect 651924 110236 651980 110246
rect 651924 90747 651980 110180
rect 652932 109676 652988 109686
rect 652932 95676 652988 109620
rect 654276 100648 654332 126756
rect 654276 100582 654332 100592
rect 654500 98924 654556 127540
rect 655956 126748 656012 126758
rect 655956 126634 656012 126644
rect 655508 126028 655564 126038
rect 654612 125804 654668 125814
rect 654612 100492 654668 125748
rect 655284 125356 655340 125366
rect 654724 124948 654780 124958
rect 654724 100716 654780 124892
rect 655060 124588 655116 124598
rect 654948 122968 655004 122978
rect 654948 122892 655004 122912
rect 654948 122826 655004 122836
rect 654948 120808 655004 120818
rect 654948 113260 655004 120752
rect 655060 118412 655116 124532
rect 655172 124408 655228 124418
rect 655172 120808 655228 124352
rect 655284 121548 655340 125300
rect 655284 121482 655340 121492
rect 655396 124768 655452 124778
rect 655172 120742 655228 120752
rect 655060 118346 655116 118356
rect 655284 120652 655340 120662
rect 654948 113194 655004 113204
rect 654724 100650 654780 100660
rect 654612 100426 654668 100436
rect 655284 99208 655340 120596
rect 655396 119868 655452 124712
rect 655396 119802 655452 119812
rect 655396 118972 655452 118982
rect 655396 99388 655452 118916
rect 655508 110548 655564 125972
rect 655620 126028 655676 126038
rect 655620 111132 655676 125972
rect 655956 125692 656012 125702
rect 655844 125580 655900 125590
rect 655732 125468 655788 125478
rect 655732 120652 655788 125412
rect 655732 120586 655788 120596
rect 655844 118972 655900 125524
rect 655844 118906 655900 118916
rect 655620 111066 655676 111076
rect 655508 110482 655564 110492
rect 655956 102507 656012 125636
rect 670180 123564 670236 123574
rect 670180 122788 670236 123508
rect 670180 122722 670236 122732
rect 655732 102451 656012 102507
rect 655732 99568 655788 102451
rect 655732 99502 655788 99512
rect 655396 99322 655452 99332
rect 655284 99142 655340 99152
rect 654500 98858 654556 98868
rect 652932 95610 652988 95620
rect 686532 92428 686588 340228
rect 686644 176540 686700 433412
rect 686756 306012 686812 553476
rect 686868 540204 686924 540214
rect 686868 307468 686924 540148
rect 686868 307402 686924 307412
rect 686756 305946 686812 305956
rect 688212 290444 688268 937300
rect 688436 937108 688492 937118
rect 688436 937020 688492 937052
rect 688436 936954 688492 936964
rect 689220 936928 689276 936938
rect 688884 936568 688940 936578
rect 688884 936460 688940 936512
rect 688884 936394 688940 936404
rect 688212 290378 688268 290388
rect 689108 936388 689164 936398
rect 687540 289212 687596 289222
rect 687540 289108 687596 289156
rect 687540 289042 687596 289052
rect 689108 256172 689164 936332
rect 689220 263004 689276 936872
rect 689332 936348 689388 936358
rect 689332 290556 689388 936292
rect 692916 922888 692972 946820
rect 703892 945928 703948 945938
rect 695380 935668 695436 935678
rect 695380 935564 695436 935612
rect 695380 935498 695436 935508
rect 694820 935488 694876 935498
rect 694260 935340 694316 935350
rect 692916 922822 692972 922832
rect 694036 935116 694092 935126
rect 689332 290490 689388 290500
rect 689556 735868 689612 735878
rect 689220 262938 689276 262948
rect 689108 256106 689164 256116
rect 689556 246876 689612 735812
rect 694036 650972 694092 935060
rect 694036 650906 694092 650916
rect 694260 650076 694316 935284
rect 694596 934408 694652 934418
rect 694596 693980 694652 934352
rect 694596 693914 694652 693924
rect 694260 650010 694316 650020
rect 694596 693532 694652 693542
rect 689556 246810 689612 246820
rect 689668 609868 689724 609878
rect 689668 214620 689724 609812
rect 694596 233100 694652 693476
rect 694596 233034 694652 233044
rect 694708 650524 694764 650534
rect 694708 226156 694764 650468
rect 694820 523852 694876 935432
rect 694932 935004 694988 935014
rect 694932 565068 694988 934948
rect 700532 934220 700588 934230
rect 697732 925148 697788 925158
rect 697732 924688 697788 925092
rect 697732 924622 697788 924632
rect 700532 909020 700588 934164
rect 703892 927164 703948 945872
rect 704004 945868 704060 945878
rect 704004 927276 704060 945812
rect 704004 927210 704060 927220
rect 703892 927098 703948 927108
rect 704788 926380 704844 926390
rect 704788 924508 704844 926324
rect 705684 926380 705740 926390
rect 705684 924688 705740 926324
rect 705684 924622 705740 924632
rect 704788 924442 704844 924452
rect 700532 908954 700588 908964
rect 704788 840364 704844 840374
rect 700420 838828 700476 838838
rect 700420 838348 700476 838772
rect 700420 838282 700476 838292
rect 700644 838648 700700 838658
rect 700644 838348 700700 838592
rect 704788 838468 704844 840308
rect 705124 840364 705180 840374
rect 705124 838828 705180 840308
rect 705124 838762 705180 838772
rect 705684 840364 705740 840374
rect 705684 838648 705740 840308
rect 705684 838582 705740 838592
rect 704788 838402 704844 838412
rect 700644 838282 700700 838292
rect 701316 838288 701372 838298
rect 701316 821884 701372 838232
rect 701316 821818 701372 821828
rect 700532 806988 700588 806998
rect 699188 752608 699244 752618
rect 699188 752490 699244 752500
rect 700420 752556 700476 752566
rect 700420 752428 700476 752500
rect 700420 752362 700476 752372
rect 700532 738780 700588 806932
rect 703892 806316 703948 806326
rect 703892 755132 703948 806260
rect 703892 755066 703948 755076
rect 704788 754460 704844 754470
rect 704788 752608 704844 754404
rect 704788 752542 704844 752552
rect 705684 754460 705740 754470
rect 705684 752428 705740 754404
rect 705684 752362 705740 752372
rect 700532 738714 700588 738724
rect 705684 711452 705740 711462
rect 700420 710556 700476 710566
rect 700420 709408 700476 710500
rect 700420 709342 700476 709352
rect 705684 709408 705740 711396
rect 705684 709342 705740 709352
rect 702100 676620 702156 676630
rect 701764 675500 701820 675510
rect 701764 666388 701820 675444
rect 702100 669116 702156 676564
rect 705236 676508 705292 676518
rect 702100 669050 702156 669060
rect 704452 676396 704508 676406
rect 704452 668556 704508 676340
rect 704452 668490 704508 668500
rect 705236 668556 705292 676452
rect 705236 668490 705292 668500
rect 701764 666322 701820 666332
rect 705684 668444 705740 668454
rect 705684 666388 705740 668388
rect 705684 666322 705740 666332
rect 701428 653236 701484 653246
rect 701428 651868 701484 653180
rect 701428 651802 701484 651812
rect 705236 633612 705292 633622
rect 701876 633500 701932 633510
rect 701876 623188 701932 633444
rect 704452 633388 704508 633398
rect 704452 626556 704508 633332
rect 704452 626490 704508 626500
rect 705236 626332 705292 633556
rect 705236 626266 705292 626276
rect 705684 633388 705740 633398
rect 705684 626332 705740 633332
rect 705684 626266 705740 626276
rect 704788 625436 704844 625446
rect 704788 623368 704844 625380
rect 704788 623302 704844 623312
rect 701876 623122 701932 623132
rect 701652 590492 701708 590502
rect 701652 583324 701708 590436
rect 704004 590380 704060 590390
rect 701652 583258 701708 583268
rect 701876 589820 701932 589830
rect 701876 580528 701932 589764
rect 704004 582876 704060 590324
rect 704004 582810 704060 582820
rect 704452 590268 704508 590278
rect 704452 582876 704508 590212
rect 704452 582810 704508 582820
rect 701876 580462 701932 580472
rect 705684 582428 705740 582438
rect 705684 580528 705740 582372
rect 705684 580462 705740 580472
rect 701428 567236 701484 567246
rect 701428 566188 701484 567180
rect 701428 566122 701484 566132
rect 694932 565002 694988 565012
rect 705012 547932 705068 547942
rect 702100 547820 702156 547830
rect 701876 543452 701932 543462
rect 701876 537508 701932 543396
rect 702100 540092 702156 547764
rect 705012 540204 705068 547876
rect 705012 540138 705068 540148
rect 705124 547708 705180 547718
rect 702100 540026 702156 540036
rect 705124 540092 705180 547652
rect 705124 540026 705180 540036
rect 701876 537442 701932 537452
rect 705684 539420 705740 539430
rect 705684 537508 705740 539364
rect 705684 537442 705740 537452
rect 694820 523786 694876 523796
rect 704452 504588 704508 504598
rect 701652 504476 701708 504486
rect 694708 226090 694764 226100
rect 694820 380156 694876 380166
rect 689668 214554 689724 214564
rect 686644 176474 686700 176484
rect 689556 176652 689612 176662
rect 689556 170716 689612 176596
rect 689556 170650 689612 170660
rect 694596 141148 694652 141158
rect 694596 92540 694652 141092
rect 694820 136780 694876 380100
rect 701652 368172 701708 504420
rect 704004 504364 704060 504374
rect 701652 368106 701708 368116
rect 701876 504140 701932 504150
rect 701876 365428 701932 504084
rect 704004 367836 704060 504308
rect 704004 367770 704060 367780
rect 704452 367836 704508 504532
rect 704452 367770 704508 367780
rect 701876 365362 701932 365372
rect 705684 367388 705740 367398
rect 705684 365428 705740 367332
rect 705684 365362 705740 365372
rect 694932 352268 694988 352278
rect 694932 193788 694988 352212
rect 695044 349580 695100 349590
rect 695044 198492 695100 349524
rect 701540 333116 701596 333126
rect 701540 325052 701596 333060
rect 704004 332892 704060 332902
rect 701540 324986 701596 324996
rect 701764 332780 701820 332790
rect 701764 322408 701820 332724
rect 704004 325164 704060 332836
rect 704004 325098 704060 325108
rect 704900 332668 704956 332678
rect 704900 325164 704956 332612
rect 704900 325098 704956 325108
rect 701764 322342 701820 322352
rect 705684 324380 705740 324390
rect 705684 322408 705740 324324
rect 705684 322342 705740 322352
rect 695044 198426 695100 198436
rect 695156 309260 695212 309270
rect 694932 193722 694988 193732
rect 695156 186956 695212 309204
rect 704676 289884 704732 289894
rect 702100 289436 702156 289446
rect 701988 289100 702044 289110
rect 701988 279388 702044 289044
rect 702100 281932 702156 289380
rect 704676 282044 704732 289828
rect 705012 289884 705068 289894
rect 705012 282156 705068 289828
rect 705012 282090 705068 282100
rect 704676 281978 704732 281988
rect 702100 281866 702156 281876
rect 701988 279322 702044 279332
rect 705684 281372 705740 281382
rect 705684 279388 705740 281316
rect 705684 279322 705740 279332
rect 704676 246876 704732 246886
rect 704564 246316 704620 246326
rect 704564 239148 704620 246260
rect 704564 239082 704620 239092
rect 704676 238476 704732 246820
rect 704676 238410 704732 238420
rect 701428 220100 701484 220110
rect 701428 218428 701484 220044
rect 701428 218362 701484 218372
rect 701428 203644 701484 203654
rect 701428 193528 701484 203588
rect 701652 203532 701708 203542
rect 701652 196252 701708 203476
rect 703892 203420 703948 203430
rect 701652 196186 701708 196196
rect 701876 203308 701932 203318
rect 701876 196028 701932 203252
rect 703892 196140 703948 203364
rect 703892 196074 703948 196084
rect 701876 195962 701932 195972
rect 701428 193462 701484 193472
rect 705684 195468 705740 195478
rect 705684 193528 705740 195412
rect 705684 193462 705740 193472
rect 695156 186890 695212 186900
rect 696164 177996 696220 178006
rect 696164 176428 696220 177940
rect 696164 176362 696220 176372
rect 705012 160860 705068 160870
rect 702100 160412 702156 160422
rect 701988 159740 702044 159750
rect 701988 150508 702044 159684
rect 702100 152572 702156 160356
rect 705012 152796 705068 160804
rect 705012 152730 705068 152740
rect 705236 160300 705292 160310
rect 705236 152796 705292 160244
rect 705236 152730 705292 152740
rect 702100 152506 702156 152516
rect 701988 150442 702044 150452
rect 705684 152460 705740 152470
rect 705684 150508 705740 152404
rect 705684 150442 705740 150452
rect 694820 136714 694876 136724
rect 700532 141868 700588 141878
rect 700532 135436 700588 141812
rect 700532 135370 700588 135380
rect 701428 134100 701484 134110
rect 701428 132748 701484 134044
rect 701428 132682 701484 132692
rect 701652 118076 701708 118086
rect 701652 110012 701708 118020
rect 704900 117852 704956 117862
rect 701652 109946 701708 109956
rect 701876 117740 701932 117750
rect 701876 107488 701932 117684
rect 704004 117628 704060 117638
rect 704004 110124 704060 117572
rect 704004 110058 704060 110068
rect 704900 110124 704956 117796
rect 704900 110058 704956 110068
rect 701876 107422 701932 107432
rect 705684 109452 705740 109462
rect 705684 107488 705740 109396
rect 705684 107422 705740 107432
rect 694596 92474 694652 92484
rect 701428 93788 701484 93798
rect 686532 92362 686588 92372
rect 701428 92428 701484 93732
rect 701428 92362 701484 92372
rect 701428 91996 701484 92006
rect 701428 90748 701484 91940
rect 651924 90691 652988 90747
rect 652932 89068 652988 90691
rect 701428 90682 701484 90692
rect 652932 89002 652988 89012
rect 651812 86552 652988 86608
rect 652932 83020 652988 86552
rect 652932 82954 652988 82964
rect 620564 71372 620620 80792
rect 628068 80668 628124 80678
rect 628068 80574 628124 80612
rect 645092 80668 645148 80678
rect 645092 80574 645148 80612
rect 620564 71306 620620 71316
rect 620340 71242 620396 71252
rect 619332 71148 619388 71158
rect 619332 71054 619388 71072
rect 617988 71036 618044 71046
rect 617988 70948 618044 70980
rect 617988 70882 618044 70892
rect 559412 70522 559468 70532
rect 548436 70074 548492 70084
rect 519652 69738 519708 69748
<< via4 >>
rect 84084 936872 84140 936928
rect 84308 936692 84364 936748
rect 84532 936512 84588 936568
rect 141876 936872 141932 936928
rect 141652 936740 141708 936748
rect 141652 936692 141708 936740
rect 141428 936512 141484 936568
rect 178724 936512 178780 936568
rect 282436 937412 282492 937468
rect 289828 937412 289884 937468
rect 341012 937412 341068 937468
rect 285684 936692 285740 936748
rect 525700 947492 525756 947548
rect 545860 947492 545916 947548
rect 581140 947492 581196 947548
rect 655844 947492 655900 947548
rect 690340 947492 690396 947548
rect 697956 947492 698012 947548
rect 525588 946232 525644 946288
rect 525700 946052 525756 946108
rect 545524 946232 545580 946288
rect 526148 945872 526204 945928
rect 545860 946052 545916 946108
rect 581140 946260 581196 946288
rect 581140 946232 581196 946260
rect 581028 946052 581084 946108
rect 545636 945872 545692 945928
rect 581252 945872 581308 945928
rect 655844 946232 655900 946288
rect 655620 946052 655676 946108
rect 655508 945872 655564 945928
rect 690340 945872 690396 945928
rect 454244 938132 454300 938188
rect 458500 938132 458556 938188
rect 342692 937412 342748 937468
rect 341236 937232 341292 937288
rect 564900 938312 564956 938368
rect 565012 937052 565068 937108
rect 587524 938312 587580 938368
rect 561316 936872 561372 936928
rect 687428 937244 687484 937288
rect 687428 937232 687484 937244
rect 687988 936692 688044 936748
rect 670292 936332 670348 936388
rect 686420 935612 686476 935668
rect 686196 935432 686252 935488
rect 76132 929900 76188 929908
rect 76132 929852 76188 929900
rect 83748 929852 83804 929908
rect 76356 927332 76412 927388
rect 78932 927332 78988 927388
rect 76244 926432 76300 926488
rect 84644 926432 84700 926488
rect 76132 766052 76188 766108
rect 83748 766052 83804 766108
rect 76244 764432 76300 764488
rect 84644 764484 84700 764488
rect 84644 764432 84700 764484
rect 76132 763172 76188 763228
rect 76132 762992 76188 763048
rect 80500 763196 80556 763228
rect 80500 763172 80556 763196
rect 76244 762812 76300 762868
rect 82292 762992 82348 763048
rect 83748 762860 83804 762868
rect 83748 762812 83804 762860
rect 76132 725012 76188 725068
rect 84644 725060 84700 725068
rect 84644 725012 84700 725060
rect 76468 722492 76524 722548
rect 84644 722492 84700 722548
rect 76132 720692 76188 720748
rect 83748 720692 83804 720748
rect 76132 683972 76188 684028
rect 84644 683972 84700 684028
rect 76132 682352 76188 682408
rect 76468 682172 76524 682228
rect 82292 682352 82348 682408
rect 76132 681092 76188 681148
rect 83748 681092 83804 681148
rect 76132 680912 76188 680968
rect 84644 680912 84700 680968
rect 76132 642212 76188 642268
rect 76468 642060 76524 642088
rect 76468 642032 76524 642060
rect 76132 640052 76188 640108
rect 83748 642212 83804 642268
rect 76132 601900 76188 601948
rect 76132 601892 76188 601900
rect 76132 600632 76188 600688
rect 76132 598472 76188 598528
rect 80388 600684 80444 600688
rect 80388 600632 80444 600684
rect 76468 599732 76524 599788
rect 83748 598500 83804 598528
rect 83748 598472 83804 598500
rect 76132 561752 76188 561808
rect 76356 559412 76412 559468
rect 76132 557972 76188 558028
rect 76244 557792 76300 557848
rect 83748 557972 83804 558028
rect 83636 557844 83692 557848
rect 83636 557792 83692 557844
rect 76132 519092 76188 519148
rect 76244 518912 76300 518968
rect 80276 518924 80332 518968
rect 80276 518912 80332 518924
rect 76468 517472 76524 517528
rect 76132 516392 76188 516448
rect 83748 516404 83804 516448
rect 83748 516392 83804 516404
rect 76132 396900 76188 396928
rect 76132 396872 76188 396900
rect 76132 396152 76188 396208
rect 76132 393632 76188 393688
rect 76244 393452 76300 393508
rect 83748 396900 83804 396928
rect 83748 396872 83804 396900
rect 78932 396172 78988 396208
rect 78932 396152 78988 396172
rect 77140 394892 77196 394948
rect 83748 393652 83804 393688
rect 83748 393632 83804 393652
rect 83636 393484 83692 393508
rect 83636 393452 83692 393484
rect 76132 356912 76188 356968
rect 76132 354212 76188 354268
rect 76132 352772 76188 352828
rect 76468 354932 76524 354988
rect 80164 354212 80220 354268
rect 76132 314252 76188 314308
rect 84532 314252 84588 314308
rect 76356 312452 76412 312508
rect 83972 312452 84028 312508
rect 76132 311372 76188 311428
rect 84084 311372 84140 311428
rect 84868 682172 84924 682228
rect 84756 642068 84812 642088
rect 84756 642032 84812 642068
rect 84868 640052 84924 640108
rect 686644 934352 686700 934408
rect 84756 601892 84812 601948
rect 84980 599732 85036 599788
rect 84756 561764 84812 561808
rect 84756 561752 84812 561764
rect 84756 559412 84812 559468
rect 84868 519092 84924 519148
rect 84980 517472 85036 517528
rect 84868 394892 84924 394948
rect 84756 356916 84812 356968
rect 84756 356912 84812 356916
rect 84756 354932 84812 354988
rect 83188 302372 83244 302428
rect 76356 301472 76412 301528
rect 80276 289952 80332 290008
rect 78820 289592 78876 289648
rect 76132 274112 76188 274168
rect 76132 270692 76188 270748
rect 76244 270512 76300 270568
rect 76468 272132 76524 272188
rect 84196 270692 84252 270748
rect 76468 234332 76524 234388
rect 76132 231812 76188 231868
rect 76132 230372 76188 230428
rect 76244 230192 76300 230248
rect 76468 232004 76524 232048
rect 76468 231992 76524 232004
rect 84644 232036 84700 232048
rect 84644 231992 84700 232036
rect 84756 206792 84812 206848
rect 84644 206612 84700 206668
rect 76132 191900 76188 191908
rect 76132 191852 76188 191900
rect 83860 191132 83916 191188
rect 76132 190772 76188 190828
rect 76468 189872 76524 189928
rect 84308 189872 84364 189928
rect 76132 188612 76188 188668
rect 85092 274112 85148 274168
rect 85092 272132 85148 272188
rect 85204 231812 85260 231868
rect 84980 230372 85036 230428
rect 85428 352772 85484 352828
rect 104132 324156 104188 324208
rect 104132 324152 104188 324156
rect 118356 323972 118412 324028
rect 151172 323792 151228 323848
rect 166292 324156 166348 324208
rect 166292 324152 166348 324156
rect 255780 325232 255836 325288
rect 253540 325052 253596 325108
rect 260932 326672 260988 326728
rect 260148 325592 260204 325648
rect 263620 326312 263676 326368
rect 262612 326132 262668 326188
rect 300244 327392 300300 327448
rect 299460 326492 299516 326548
rect 302260 325952 302316 326008
rect 306068 325412 306124 325468
rect 311108 327212 311164 327268
rect 316932 324692 316988 324748
rect 161812 323972 161868 324028
rect 334180 327032 334236 327088
rect 320404 325592 320460 325648
rect 333172 326852 333228 326908
rect 325780 324512 325836 324568
rect 332276 324332 332332 324388
rect 334292 326312 334348 326368
rect 336644 328292 336700 328348
rect 334516 326672 334572 326728
rect 334404 326132 334460 326188
rect 335972 325052 336028 325108
rect 336756 325232 336812 325288
rect 340452 325592 340508 325648
rect 347620 325232 347676 325288
rect 357028 326672 357084 326728
rect 358708 325592 358764 325648
rect 358484 325052 358540 325108
rect 367892 328292 367948 328348
rect 369460 328472 369516 328528
rect 367892 325412 367948 325468
rect 365764 324872 365820 324928
rect 376852 327572 376908 327628
rect 374276 325412 374332 325468
rect 371588 323972 371644 324028
rect 161028 323792 161084 323848
rect 93828 320912 93884 320968
rect 92372 270512 92428 270568
rect 85316 191852 85372 191908
rect 92372 206612 92428 206668
rect 90356 191132 90412 191188
rect 84868 188612 84924 188668
rect 76244 188432 76300 188488
rect 93380 291392 93436 291448
rect 93156 230192 93212 230248
rect 93268 289052 93324 289108
rect 92596 190952 92652 191008
rect 93156 206792 93212 206848
rect 93380 234332 93436 234388
rect 93268 188432 93324 188488
rect 93156 82952 93212 83008
rect 159572 320912 159628 320968
rect 99092 308132 99148 308188
rect 154644 307952 154700 308008
rect 102452 307772 102508 307828
rect 100772 307412 100828 307468
rect 117908 291572 117964 291628
rect 159796 307592 159852 307648
rect 162932 308132 162988 308188
rect 164612 307772 164668 307828
rect 164724 307412 164780 307468
rect 165396 307772 165452 307828
rect 165620 307412 165676 307468
rect 181412 307412 181468 307468
rect 181636 308132 181692 308188
rect 173236 291572 173292 291628
rect 190596 307952 190652 308008
rect 183092 307772 183148 307828
rect 203252 308132 203308 308188
rect 193172 307592 193228 307648
rect 196532 307592 196588 307648
rect 201348 307412 201404 307468
rect 209972 307592 210028 307648
rect 206612 307412 206668 307468
rect 238420 307952 238476 308008
rect 248500 307772 248556 307828
rect 251972 307952 252028 308008
rect 241780 307592 241836 307648
rect 234612 307412 234668 307468
rect 245252 307412 245308 307468
rect 261940 307412 261996 307468
rect 262052 307592 262108 307648
rect 282100 307952 282156 308008
rect 265300 307592 265356 307648
rect 272132 307772 272188 307828
rect 285572 307412 285628 307468
rect 297220 307412 297276 307468
rect 286020 301832 286076 301888
rect 285572 301652 285628 301708
rect 285796 300752 285852 300808
rect 292292 299492 292348 299548
rect 303940 307592 303996 307648
rect 299012 300032 299068 300088
rect 294532 299312 294588 299368
rect 302820 299852 302876 299908
rect 302596 299132 302652 299188
rect 313796 307592 313852 307648
rect 316820 307952 316876 308008
rect 310996 295712 311052 295768
rect 320740 307952 320796 308008
rect 317380 307772 317436 307828
rect 321188 291932 321244 291988
rect 320964 291752 321020 291808
rect 321412 291572 321468 291628
rect 334180 308132 334236 308188
rect 334404 295712 334460 295768
rect 327908 284732 327964 284788
rect 329588 284192 329644 284248
rect 327684 284012 327740 284068
rect 336756 307772 336812 307828
rect 335972 294092 336028 294148
rect 336980 307592 337036 307648
rect 337204 307412 337260 307468
rect 342580 303452 342636 303508
rect 344260 303272 344316 303328
rect 378644 322532 378700 322588
rect 378196 322172 378252 322228
rect 377972 317312 378028 317368
rect 362740 303992 362796 304048
rect 369460 307772 369516 307828
rect 377636 308132 377692 308188
rect 364420 303812 364476 303868
rect 357700 303092 357756 303148
rect 354900 301868 354956 301888
rect 354900 301832 354956 301868
rect 356132 301652 356188 301708
rect 352772 300752 352828 300808
rect 338436 299492 338492 299548
rect 335972 291392 336028 291448
rect 337540 289052 337596 289108
rect 343476 299312 343532 299368
rect 377860 307592 377916 307648
rect 377860 307412 377916 307468
rect 393092 328472 393148 328528
rect 388276 326492 388332 326548
rect 453572 327392 453628 327448
rect 405748 325412 405804 325468
rect 470372 325952 470428 326008
rect 453684 325232 453740 325288
rect 497364 327212 497420 327268
rect 533092 327032 533148 327088
rect 551684 326852 551740 326908
rect 656740 327572 656796 327628
rect 623252 326672 623308 326728
rect 487956 325052 488012 325108
rect 382004 324872 382060 324928
rect 485492 324872 485548 324928
rect 655508 324884 655564 324928
rect 655508 324872 655564 324884
rect 505540 324692 505596 324748
rect 537572 324548 537628 324568
rect 537572 324512 537628 324548
rect 554372 324332 554428 324388
rect 485492 323972 485548 324028
rect 380324 322892 380380 322948
rect 379540 322712 379596 322768
rect 379764 322196 379820 322228
rect 379764 322172 379820 322196
rect 379876 319508 379932 319528
rect 379876 319472 379932 319508
rect 557732 319472 557788 319528
rect 379764 317324 379820 317368
rect 379764 317312 379820 317324
rect 378756 309932 378812 309988
rect 672420 322892 672476 322948
rect 672644 322712 672700 322768
rect 672756 322532 672812 322588
rect 379764 312452 379820 312508
rect 460292 312452 460348 312508
rect 664356 309932 664412 309988
rect 379540 309212 379596 309268
rect 458612 309260 458668 309268
rect 458612 309212 458668 309260
rect 426692 307952 426748 308008
rect 385924 302552 385980 302608
rect 381780 300032 381836 300088
rect 389732 299852 389788 299908
rect 378196 294812 378252 294868
rect 391412 299132 391468 299188
rect 461972 292112 462028 292168
rect 428820 291932 428876 291988
rect 428596 291788 428652 291808
rect 428596 291752 428652 291788
rect 430388 291572 430444 291628
rect 444052 284732 444108 284788
rect 446628 284192 446684 284248
rect 445284 284012 445340 284068
rect 532420 307804 532476 307828
rect 532420 307772 532476 307804
rect 550116 307592 550172 307648
rect 520548 303996 520604 304048
rect 520548 303992 520604 303996
rect 474516 303452 474572 303508
rect 465332 292292 465388 292348
rect 462756 292112 462812 292168
rect 472052 290332 472108 290368
rect 472052 290312 472108 290332
rect 479556 303272 479612 303328
rect 475412 290500 475468 290548
rect 475412 290492 475468 290500
rect 468580 287252 468636 287308
rect 469140 287432 469196 287488
rect 477876 290132 477932 290188
rect 522340 303812 522396 303868
rect 482132 294272 482188 294328
rect 506436 303092 506492 303148
rect 488852 292852 488908 292888
rect 488852 292832 488908 292852
rect 498932 292652 498988 292708
rect 497252 292516 497308 292528
rect 497252 292472 497308 292516
rect 537572 293912 537628 293968
rect 510692 293020 510748 293068
rect 510692 293012 510748 293020
rect 534212 291620 534268 291628
rect 534212 291572 534268 291620
rect 506436 291392 506492 291448
rect 532532 291212 532588 291268
rect 521332 291032 521388 291088
rect 535892 290892 535948 290908
rect 535892 290852 535948 290892
rect 538580 293912 538636 293968
rect 541716 302552 541772 302608
rect 539252 293412 539308 293428
rect 539252 293372 539308 293412
rect 538580 293192 538636 293248
rect 551012 307412 551068 307468
rect 652260 302372 652316 302428
rect 550116 293552 550172 293608
rect 557732 294812 557788 294868
rect 611380 294272 611436 294328
rect 606228 292832 606284 292888
rect 609924 292112 609980 292168
rect 606228 290672 606284 290728
rect 609812 291932 609868 291988
rect 606340 290492 606396 290548
rect 606340 290312 606396 290368
rect 600516 287252 600572 287308
rect 644420 293552 644476 293608
rect 638708 293372 638764 293428
rect 638148 293192 638204 293248
rect 628068 293012 628124 293068
rect 623252 292652 623308 292708
rect 622804 292472 622860 292528
rect 620676 291932 620732 291988
rect 611380 290672 611436 290728
rect 614740 290672 614796 290728
rect 620676 290672 620732 290728
rect 614292 290492 614348 290548
rect 611044 290312 611100 290368
rect 614292 290312 614348 290368
rect 616420 290492 616476 290548
rect 615636 290132 615692 290188
rect 617540 290312 617596 290368
rect 626164 291392 626220 291448
rect 636692 291572 636748 291628
rect 636244 291212 636300 291268
rect 631988 291032 632044 291088
rect 637252 290852 637308 290908
rect 642516 291752 642572 291808
rect 646548 292292 646604 292348
rect 670404 301472 670460 301528
rect 669844 290672 669900 290728
rect 667492 290492 667548 290548
rect 667044 290132 667100 290188
rect 652596 289952 652652 290008
rect 661668 289952 661724 290008
rect 655508 289772 655564 289828
rect 658308 289772 658364 289828
rect 667044 289772 667100 289828
rect 667268 289772 667324 289828
rect 670180 290492 670236 290548
rect 670964 289952 671020 290008
rect 671076 291932 671132 291988
rect 671300 294092 671356 294148
rect 672196 290132 672252 290188
rect 672308 289772 672364 289828
rect 611044 287432 611100 287488
rect 671860 289052 671916 289108
rect 558404 268712 558460 268768
rect 559300 268712 559356 268768
rect 558516 257192 558572 257248
rect 559300 257192 559356 257248
rect 335972 82952 336028 83008
rect 558404 185732 558460 185788
rect 559636 185732 559692 185788
rect 558628 184832 558684 184888
rect 559076 184832 559132 184888
rect 558404 143612 558460 143668
rect 559300 143612 559356 143668
rect 558516 142532 558572 142588
rect 558404 96632 558460 96688
rect 558404 82232 558460 82288
rect 559412 142532 559468 142588
rect 559412 141992 559468 142048
rect 558628 90692 558684 90748
rect 558628 82052 558684 82108
rect 559300 96632 559356 96688
rect 559300 90692 559356 90748
rect 559188 81872 559244 81928
rect 585396 82232 585452 82288
rect 585620 82052 585676 82108
rect 671860 141992 671916 142048
rect 671636 141812 671692 141868
rect 671748 141092 671804 141148
rect 618884 140012 618940 140068
rect 618324 139652 618380 139708
rect 618548 139472 618604 139528
rect 585844 81872 585900 81928
rect 176260 71252 176316 71308
rect 324884 70712 324940 70768
rect 257796 70532 257852 70588
rect 494340 71432 494396 71488
rect 519652 71072 519708 71128
rect 505876 70892 505932 70948
rect 548436 70712 548492 70768
rect 539140 70532 539196 70588
rect 618772 123092 618828 123148
rect 619108 140012 619164 140068
rect 623364 140028 623420 140068
rect 623364 140012 623420 140028
rect 624708 140028 624764 140068
rect 624708 140012 624764 140028
rect 649348 140012 649404 140068
rect 618996 139652 619052 139708
rect 619108 139832 619164 139888
rect 631428 139860 631484 139888
rect 631428 139832 631484 139860
rect 619332 139652 619388 139708
rect 632772 139692 632828 139708
rect 632772 139652 632828 139692
rect 622020 139472 622076 139528
rect 622468 139472 622524 139528
rect 618436 71432 618492 71488
rect 620340 80612 620396 80668
rect 620340 71252 620396 71308
rect 621348 122912 621404 122968
rect 621460 122732 621516 122788
rect 622244 99332 622300 99388
rect 638820 139472 638876 139528
rect 622580 100592 622636 100648
rect 622692 100412 622748 100468
rect 646324 126692 646380 126748
rect 646996 125972 647052 126028
rect 641508 124892 641564 124948
rect 628740 124712 628796 124768
rect 628068 124532 628124 124588
rect 626052 124352 626108 124408
rect 642740 124172 642796 124228
rect 649572 140012 649628 140068
rect 657076 140028 657132 140068
rect 657076 140012 657132 140028
rect 657748 140028 657804 140068
rect 657748 140012 657804 140028
rect 649684 139832 649740 139888
rect 655732 139860 655788 139888
rect 655732 139832 655788 139860
rect 650916 139652 650972 139708
rect 650804 132632 650860 132688
rect 656404 139692 656460 139708
rect 656404 139652 656460 139692
rect 666484 139472 666540 139528
rect 657972 132636 658028 132688
rect 657972 132632 658028 132636
rect 664580 132636 664636 132688
rect 664580 132632 664636 132636
rect 659652 132468 659708 132508
rect 659652 132452 659708 132468
rect 649796 132272 649852 132328
rect 653492 132272 653548 132328
rect 666820 132272 666876 132328
rect 669956 132452 670012 132508
rect 670740 132632 670796 132688
rect 671076 139472 671132 139528
rect 665140 131012 665196 131068
rect 671076 132272 671132 132328
rect 670964 131012 671020 131068
rect 648452 124172 648508 124228
rect 647892 123284 647948 123328
rect 647892 123272 647948 123284
rect 651812 110492 651868 110548
rect 628628 100592 628684 100648
rect 649572 100592 649628 100648
rect 631204 100436 631260 100468
rect 631204 100412 631260 100436
rect 633780 99332 633836 99388
rect 622468 99152 622524 99208
rect 635796 99152 635852 99208
rect 644980 99512 645036 99568
rect 641732 99332 641788 99388
rect 639044 99152 639100 99208
rect 654276 100592 654332 100648
rect 655956 126700 656012 126748
rect 655956 126692 656012 126700
rect 655508 125972 655564 126028
rect 654724 124892 654780 124948
rect 655060 124532 655116 124588
rect 654948 122912 655004 122968
rect 654948 120752 655004 120808
rect 655172 124352 655228 124408
rect 655396 124712 655452 124768
rect 655172 120752 655228 120808
rect 655508 110492 655564 110548
rect 670180 122732 670236 122788
rect 655732 99512 655788 99568
rect 655396 99332 655452 99388
rect 655284 99152 655340 99208
rect 688436 937052 688492 937108
rect 689220 936872 689276 936928
rect 688884 936512 688940 936568
rect 689108 936332 689164 936388
rect 687540 289052 687596 289108
rect 703892 945872 703948 945928
rect 695380 935612 695436 935668
rect 694820 935432 694876 935488
rect 692916 922832 692972 922888
rect 694596 934352 694652 934408
rect 697732 924632 697788 924688
rect 705684 924632 705740 924688
rect 704788 924452 704844 924508
rect 700420 838772 700476 838828
rect 700644 838592 700700 838648
rect 705124 838772 705180 838828
rect 705684 838592 705740 838648
rect 704788 838412 704844 838468
rect 701316 838232 701372 838288
rect 699188 752556 699244 752608
rect 699188 752552 699244 752556
rect 700420 752372 700476 752428
rect 704788 752552 704844 752608
rect 705684 752372 705740 752428
rect 700420 709352 700476 709408
rect 705684 709352 705740 709408
rect 701764 666332 701820 666388
rect 705684 666332 705740 666388
rect 704788 623312 704844 623368
rect 701876 623132 701932 623188
rect 701876 580472 701932 580528
rect 705684 580472 705740 580528
rect 701876 537452 701932 537508
rect 705684 537452 705740 537508
rect 694596 141092 694652 141148
rect 701876 365372 701932 365428
rect 705684 365372 705740 365428
rect 701764 322352 701820 322408
rect 705684 322352 705740 322408
rect 701988 279332 702044 279388
rect 705684 279332 705740 279388
rect 701428 193472 701484 193528
rect 705684 193472 705740 193528
rect 701988 150452 702044 150508
rect 705684 150452 705740 150508
rect 700532 141812 700588 141868
rect 701876 107432 701932 107488
rect 705684 107432 705740 107488
rect 620564 80792 620620 80848
rect 628068 80612 628124 80668
rect 645092 80612 645148 80668
rect 619332 71092 619388 71128
rect 619332 71072 619388 71092
rect 617988 70892 618044 70948
<< metal5 >>
rect 107500 1007600 119500 1019600
rect 162500 1007600 174500 1019600
rect 217500 1007600 229500 1019600
rect 272500 1007600 284500 1019600
rect 327500 1007600 339500 1019600
rect 382500 1007600 394500 1019600
rect 437500 1007600 449500 1019600
rect 492500 1007600 504500 1019600
rect 547500 1007600 559500 1019600
rect 602500 1007600 614500 1019600
rect 657500 1007600 669500 1019600
rect 525684 947548 545932 947564
rect 525684 947492 525700 947548
rect 525756 947492 545860 947548
rect 545916 947492 545932 947548
rect 525684 947476 545932 947492
rect 581124 947548 655916 947564
rect 581124 947492 581140 947548
rect 581196 947492 655844 947548
rect 655900 947492 655916 947548
rect 581124 947476 655916 947492
rect 690324 947548 698028 947564
rect 690324 947492 690340 947548
rect 690396 947492 697956 947548
rect 698012 947492 698028 947548
rect 690324 947476 698028 947492
rect 525572 946288 545596 946304
rect 525572 946232 525588 946288
rect 525644 946232 545524 946288
rect 545580 946232 545596 946288
rect 525572 946216 545596 946232
rect 581124 946288 655916 946304
rect 581124 946232 581140 946288
rect 581196 946232 655844 946288
rect 655900 946232 655916 946288
rect 581124 946216 655916 946232
rect 525684 946108 545932 946124
rect 525684 946052 525700 946108
rect 525756 946052 545860 946108
rect 545916 946052 545932 946108
rect 525684 946036 545932 946052
rect 581012 946108 655692 946124
rect 581012 946052 581028 946108
rect 581084 946052 655620 946108
rect 655676 946052 655692 946108
rect 581012 946036 655692 946052
rect 526132 945928 545708 945944
rect 526132 945872 526148 945928
rect 526204 945872 545636 945928
rect 545692 945872 545708 945928
rect 526132 945856 545708 945872
rect 581236 945928 655580 945944
rect 581236 945872 581252 945928
rect 581308 945872 655508 945928
rect 655564 945872 655580 945928
rect 581236 945856 655580 945872
rect 690324 945928 703964 945944
rect 690324 945872 690340 945928
rect 690396 945872 703892 945928
rect 703948 945872 703964 945928
rect 690324 945856 703964 945872
rect 564884 938368 587596 938384
rect 564884 938312 564900 938368
rect 564956 938312 587524 938368
rect 587580 938312 587596 938368
rect 564884 938296 587596 938312
rect 454228 938188 458572 938204
rect 454228 938132 454244 938188
rect 454300 938132 458500 938188
rect 458556 938132 458572 938188
rect 454228 938116 458572 938132
rect 282420 937468 289900 937484
rect 282420 937412 282436 937468
rect 282492 937412 289828 937468
rect 289884 937412 289900 937468
rect 282420 937396 289900 937412
rect 340996 937468 342764 937484
rect 340996 937412 341012 937468
rect 341068 937412 342692 937468
rect 342748 937412 342764 937468
rect 340996 937396 342764 937412
rect 341220 937288 687500 937304
rect 341220 937232 341236 937288
rect 341292 937232 687428 937288
rect 687484 937232 687500 937288
rect 341220 937216 687500 937232
rect 564996 937108 688508 937124
rect 564996 937052 565012 937108
rect 565068 937052 688436 937108
rect 688492 937052 688508 937108
rect 564996 937036 688508 937052
rect 84068 936928 141948 936944
rect 84068 936872 84084 936928
rect 84140 936872 141876 936928
rect 141932 936872 141948 936928
rect 84068 936856 141948 936872
rect 561300 936928 689292 936944
rect 561300 936872 561316 936928
rect 561372 936872 689220 936928
rect 689276 936872 689292 936928
rect 561300 936856 689292 936872
rect 84292 936748 141724 936764
rect 84292 936692 84308 936748
rect 84364 936692 141652 936748
rect 141708 936692 141724 936748
rect 84292 936676 141724 936692
rect 285668 936748 688060 936764
rect 285668 936692 285684 936748
rect 285740 936692 687988 936748
rect 688044 936692 688060 936748
rect 285668 936676 688060 936692
rect 84516 936568 141500 936584
rect 84516 936512 84532 936568
rect 84588 936512 141428 936568
rect 141484 936512 141500 936568
rect 84516 936496 141500 936512
rect 178708 936568 688956 936584
rect 178708 936512 178724 936568
rect 178780 936512 688884 936568
rect 688940 936512 688956 936568
rect 178708 936496 688956 936512
rect 670276 936388 689180 936404
rect 670276 936332 670292 936388
rect 670348 936332 689108 936388
rect 689164 936332 689180 936388
rect 670276 936316 689180 936332
rect 686404 935668 695452 935684
rect 686404 935612 686420 935668
rect 686476 935612 695380 935668
rect 695436 935612 695452 935668
rect 686404 935596 695452 935612
rect 686180 935488 694892 935504
rect 686180 935432 686196 935488
rect 686252 935432 694820 935488
rect 694876 935432 694892 935488
rect 686180 935416 694892 935432
rect 686628 934408 694668 934424
rect 686628 934352 686644 934408
rect 686700 934352 694596 934408
rect 694652 934352 694668 934408
rect 686628 934336 694668 934352
rect 76116 929908 83820 929924
rect 76116 929852 76132 929908
rect 76188 929852 83748 929908
rect 83804 929852 83820 929908
rect 76116 929836 83820 929852
rect 76340 927388 79004 927404
rect 76340 927332 76356 927388
rect 76412 927332 78932 927388
rect 78988 927332 79004 927388
rect 76340 927316 79004 927332
rect 76228 926488 84716 926504
rect 76228 926432 76244 926488
rect 76300 926432 84644 926488
rect 84700 926432 84716 926488
rect 76228 926416 84716 926432
rect 697716 924688 705756 924704
rect 697716 924632 697732 924688
rect 697788 924632 705684 924688
rect 705740 924632 705756 924688
rect 697716 924616 705756 924632
rect 704772 924508 704860 924524
rect 400 912500 12400 924500
rect 704772 924452 704788 924508
rect 704844 924452 704860 924508
rect 704772 922904 704860 924452
rect 692900 922888 704860 922904
rect 692900 922832 692916 922888
rect 692972 922832 704860 922888
rect 692900 922816 704860 922832
rect 765600 913500 777600 925500
rect 400 871500 12400 883500
rect 765600 870500 777600 882500
rect 400 830500 12400 842500
rect 700404 838828 705196 838844
rect 700404 838772 700420 838828
rect 700476 838772 705124 838828
rect 705180 838772 705196 838828
rect 700404 838756 705196 838772
rect 700628 838648 705756 838664
rect 700628 838592 700644 838648
rect 700700 838592 705684 838648
rect 705740 838592 705756 838648
rect 700628 838576 705756 838592
rect 704772 838468 704860 838484
rect 704772 838412 704788 838468
rect 704844 838412 704860 838468
rect 704772 838304 704860 838412
rect 701300 838288 704860 838304
rect 701300 838232 701316 838288
rect 701372 838232 704860 838288
rect 701300 838216 704860 838232
rect 765600 827500 777600 839500
rect 400 789500 12400 801500
rect 765600 784500 777600 796500
rect 76116 766108 83820 766124
rect 76116 766052 76132 766108
rect 76188 766052 83748 766108
rect 83804 766052 83820 766108
rect 76116 766036 83820 766052
rect 76228 764488 84716 764504
rect 76228 764432 76244 764488
rect 76300 764432 84644 764488
rect 84700 764432 84716 764488
rect 76228 764416 84716 764432
rect 76116 763228 80572 763244
rect 76116 763172 76132 763228
rect 76188 763172 80500 763228
rect 80556 763172 80572 763228
rect 76116 763156 80572 763172
rect 76116 763048 82364 763064
rect 76116 762992 76132 763048
rect 76188 762992 82292 763048
rect 82348 762992 82364 763048
rect 76116 762976 82364 762992
rect 76228 762868 83820 762884
rect 76228 762812 76244 762868
rect 76300 762812 83748 762868
rect 83804 762812 83820 762868
rect 76228 762796 83820 762812
rect 400 748500 12400 760500
rect 699172 752608 704860 752624
rect 699172 752552 699188 752608
rect 699244 752552 704788 752608
rect 704844 752552 704860 752608
rect 699172 752536 704860 752552
rect 700404 752428 705756 752444
rect 700404 752372 700420 752428
rect 700476 752372 705684 752428
rect 705740 752372 705756 752428
rect 700404 752356 705756 752372
rect 765600 741500 777600 753500
rect 76116 725068 84716 725084
rect 76116 725012 76132 725068
rect 76188 725012 84644 725068
rect 84700 725012 84716 725068
rect 76116 724996 84716 725012
rect 76452 722548 84716 722564
rect 76452 722492 76468 722548
rect 76524 722492 84644 722548
rect 84700 722492 84716 722548
rect 76452 722476 84716 722492
rect 76116 720748 83820 720764
rect 76116 720692 76132 720748
rect 76188 720692 83748 720748
rect 83804 720692 83820 720748
rect 76116 720676 83820 720692
rect 400 707500 12400 719500
rect 700404 709408 705756 709424
rect 700404 709352 700420 709408
rect 700476 709352 705684 709408
rect 705740 709352 705756 709408
rect 700404 709336 705756 709352
rect 765600 698500 777600 710500
rect 76116 684028 84716 684044
rect 76116 683972 76132 684028
rect 76188 683972 84644 684028
rect 84700 683972 84716 684028
rect 76116 683956 84716 683972
rect 76116 682408 82364 682424
rect 76116 682352 76132 682408
rect 76188 682352 82292 682408
rect 82348 682352 82364 682408
rect 76116 682336 82364 682352
rect 76452 682228 84940 682244
rect 76452 682172 76468 682228
rect 76524 682172 84868 682228
rect 84924 682172 84940 682228
rect 76452 682156 84940 682172
rect 76116 681148 83820 681164
rect 76116 681092 76132 681148
rect 76188 681092 83748 681148
rect 83804 681092 83820 681148
rect 76116 681076 83820 681092
rect 76116 680968 84716 680984
rect 76116 680912 76132 680968
rect 76188 680912 84644 680968
rect 84700 680912 84716 680968
rect 76116 680896 84716 680912
rect 400 666500 12400 678500
rect 701748 666388 705756 666404
rect 701748 666332 701764 666388
rect 701820 666332 705684 666388
rect 705740 666332 705756 666388
rect 701748 666316 705756 666332
rect 765600 655500 777600 667500
rect 76116 642268 83820 642284
rect 76116 642212 76132 642268
rect 76188 642212 83748 642268
rect 83804 642212 83820 642268
rect 76116 642196 83820 642212
rect 76452 642088 84828 642104
rect 76452 642032 76468 642088
rect 76524 642032 84756 642088
rect 84812 642032 84828 642088
rect 76452 642016 84828 642032
rect 76116 640108 84940 640124
rect 76116 640052 76132 640108
rect 76188 640052 84868 640108
rect 84924 640052 84940 640108
rect 76116 640036 84940 640052
rect 400 625500 12400 637500
rect 704772 623368 704860 623384
rect 704772 623312 704788 623368
rect 704844 623312 704860 623368
rect 704772 623204 704860 623312
rect 701860 623188 704860 623204
rect 701860 623132 701876 623188
rect 701932 623132 704860 623188
rect 701860 623116 704860 623132
rect 765600 612500 777600 624500
rect 76116 601948 84828 601964
rect 76116 601892 76132 601948
rect 76188 601892 84756 601948
rect 84812 601892 84828 601948
rect 76116 601876 84828 601892
rect 76116 600688 80460 600704
rect 76116 600632 76132 600688
rect 76188 600632 80388 600688
rect 80444 600632 80460 600688
rect 76116 600616 80460 600632
rect 76452 599788 85052 599804
rect 76452 599732 76468 599788
rect 76524 599732 84980 599788
rect 85036 599732 85052 599788
rect 76452 599716 85052 599732
rect 76116 598528 83820 598544
rect 76116 598472 76132 598528
rect 76188 598472 83748 598528
rect 83804 598472 83820 598528
rect 76116 598456 83820 598472
rect 400 584500 12400 596500
rect 701860 580528 705756 580544
rect 701860 580472 701876 580528
rect 701932 580472 705684 580528
rect 705740 580472 705756 580528
rect 701860 580456 705756 580472
rect 765600 569500 777600 581500
rect 76116 561808 84828 561824
rect 76116 561752 76132 561808
rect 76188 561752 84756 561808
rect 84812 561752 84828 561808
rect 76116 561736 84828 561752
rect 76340 559468 84828 559484
rect 76340 559412 76356 559468
rect 76412 559412 84756 559468
rect 84812 559412 84828 559468
rect 76340 559396 84828 559412
rect 76116 558028 83820 558044
rect 76116 557972 76132 558028
rect 76188 557972 83748 558028
rect 83804 557972 83820 558028
rect 76116 557956 83820 557972
rect 76228 557848 83708 557864
rect 76228 557792 76244 557848
rect 76300 557792 83636 557848
rect 83692 557792 83708 557848
rect 76228 557776 83708 557792
rect 400 543500 12400 555500
rect 701860 537508 705756 537524
rect 701860 537452 701876 537508
rect 701932 537452 705684 537508
rect 705740 537452 705756 537508
rect 701860 537436 705756 537452
rect 765600 526500 777600 538500
rect 76116 519148 84940 519164
rect 76116 519092 76132 519148
rect 76188 519092 84868 519148
rect 84924 519092 84940 519148
rect 76116 519076 84940 519092
rect 76228 518968 80348 518984
rect 76228 518912 76244 518968
rect 76300 518912 80276 518968
rect 80332 518912 80348 518968
rect 76228 518896 80348 518912
rect 76452 517528 85052 517544
rect 76452 517472 76468 517528
rect 76524 517472 84980 517528
rect 85036 517472 85052 517528
rect 76452 517456 85052 517472
rect 76116 516448 83820 516464
rect 76116 516392 76132 516448
rect 76188 516392 83748 516448
rect 83804 516392 83820 516448
rect 76116 516376 83820 516392
rect 400 502500 12400 514500
rect 765600 483500 777600 495500
rect 400 461500 12400 473500
rect 765600 440500 777600 452500
rect 400 420500 12400 432500
rect 765600 397500 777600 409500
rect 76116 396928 83820 396944
rect 76116 396872 76132 396928
rect 76188 396872 83748 396928
rect 83804 396872 83820 396928
rect 76116 396856 83820 396872
rect 76116 396208 79004 396224
rect 76116 396152 76132 396208
rect 76188 396152 78932 396208
rect 78988 396152 79004 396208
rect 76116 396136 79004 396152
rect 77124 394948 84940 394964
rect 77124 394892 77140 394948
rect 77196 394892 84868 394948
rect 84924 394892 84940 394948
rect 77124 394876 84940 394892
rect 76116 393688 83820 393704
rect 76116 393632 76132 393688
rect 76188 393632 83748 393688
rect 83804 393632 83820 393688
rect 76116 393616 83820 393632
rect 76228 393508 83708 393524
rect 76228 393452 76244 393508
rect 76300 393452 83636 393508
rect 83692 393452 83708 393508
rect 76228 393436 83708 393452
rect 400 379500 12400 391500
rect 701860 365428 705756 365444
rect 701860 365372 701876 365428
rect 701932 365372 705684 365428
rect 705740 365372 705756 365428
rect 701860 365356 705756 365372
rect 76116 356968 84828 356984
rect 76116 356912 76132 356968
rect 76188 356912 84756 356968
rect 84812 356912 84828 356968
rect 76116 356896 84828 356912
rect 76452 354988 84828 355004
rect 76452 354932 76468 354988
rect 76524 354932 84756 354988
rect 84812 354932 84828 354988
rect 76452 354916 84828 354932
rect 765600 354500 777600 366500
rect 76116 354268 80236 354284
rect 76116 354212 76132 354268
rect 76188 354212 80164 354268
rect 80220 354212 80236 354268
rect 76116 354196 80236 354212
rect 76116 352828 85500 352844
rect 76116 352772 76132 352828
rect 76188 352772 85428 352828
rect 85484 352772 85500 352828
rect 76116 352756 85500 352772
rect 400 338500 12400 350500
rect 369444 328528 393164 328544
rect 369444 328472 369460 328528
rect 369516 328472 393092 328528
rect 393148 328472 393164 328528
rect 369444 328456 393164 328472
rect 336628 328348 367964 328364
rect 336628 328292 336644 328348
rect 336700 328292 367892 328348
rect 367948 328292 367964 328348
rect 336628 328276 367964 328292
rect 376836 327628 656812 327644
rect 376836 327572 376852 327628
rect 376908 327572 656740 327628
rect 656796 327572 656812 327628
rect 376836 327556 656812 327572
rect 300228 327448 453644 327464
rect 300228 327392 300244 327448
rect 300300 327392 453572 327448
rect 453628 327392 453644 327448
rect 300228 327376 453644 327392
rect 311092 327268 497436 327284
rect 311092 327212 311108 327268
rect 311164 327212 497364 327268
rect 497420 327212 497436 327268
rect 311092 327196 497436 327212
rect 334164 327088 533164 327104
rect 334164 327032 334180 327088
rect 334236 327032 533092 327088
rect 533148 327032 533164 327088
rect 334164 327016 533164 327032
rect 333156 326908 551756 326924
rect 333156 326852 333172 326908
rect 333228 326852 551684 326908
rect 551740 326852 551756 326908
rect 333156 326836 551756 326852
rect 260916 326728 334588 326744
rect 260916 326672 260932 326728
rect 260988 326672 334516 326728
rect 334572 326672 334588 326728
rect 260916 326656 334588 326672
rect 357012 326728 623324 326744
rect 357012 326672 357028 326728
rect 357084 326672 623252 326728
rect 623308 326672 623324 326728
rect 357012 326656 623324 326672
rect 299444 326548 388348 326564
rect 299444 326492 299460 326548
rect 299516 326492 388276 326548
rect 388332 326492 388348 326548
rect 299444 326476 388348 326492
rect 263604 326368 334364 326384
rect 263604 326312 263620 326368
rect 263676 326312 334292 326368
rect 334348 326312 334364 326368
rect 263604 326296 334364 326312
rect 262596 326188 334476 326204
rect 262596 326132 262612 326188
rect 262668 326132 334404 326188
rect 334460 326132 334476 326188
rect 262596 326116 334476 326132
rect 302244 326008 470444 326024
rect 302244 325952 302260 326008
rect 302316 325952 470372 326008
rect 470428 325952 470444 326008
rect 302244 325936 470444 325952
rect 260132 325648 320476 325664
rect 260132 325592 260148 325648
rect 260204 325592 320404 325648
rect 320460 325592 320476 325648
rect 260132 325576 320476 325592
rect 340436 325648 358780 325664
rect 340436 325592 340452 325648
rect 340508 325592 358708 325648
rect 358764 325592 358780 325648
rect 340436 325576 358780 325592
rect 306052 325468 367964 325484
rect 306052 325412 306068 325468
rect 306124 325412 367892 325468
rect 367948 325412 367964 325468
rect 306052 325396 367964 325412
rect 374260 325468 405820 325484
rect 374260 325412 374276 325468
rect 374332 325412 405748 325468
rect 405804 325412 405820 325468
rect 374260 325396 405820 325412
rect 255764 325288 336828 325304
rect 255764 325232 255780 325288
rect 255836 325232 336756 325288
rect 336812 325232 336828 325288
rect 255764 325216 336828 325232
rect 347604 325288 453756 325304
rect 347604 325232 347620 325288
rect 347676 325232 453684 325288
rect 453740 325232 453756 325288
rect 347604 325216 453756 325232
rect 253524 325108 336044 325124
rect 253524 325052 253540 325108
rect 253596 325052 335972 325108
rect 336028 325052 336044 325108
rect 253524 325036 336044 325052
rect 358468 325108 488028 325124
rect 358468 325052 358484 325108
rect 358540 325052 487956 325108
rect 488012 325052 488028 325108
rect 358468 325036 488028 325052
rect 365748 324928 382076 324944
rect 365748 324872 365764 324928
rect 365820 324872 382004 324928
rect 382060 324872 382076 324928
rect 365748 324856 382076 324872
rect 485476 324928 655580 324944
rect 485476 324872 485492 324928
rect 485548 324872 655508 324928
rect 655564 324872 655580 324928
rect 485476 324856 655580 324872
rect 316916 324748 505612 324764
rect 316916 324692 316932 324748
rect 316988 324692 505540 324748
rect 505596 324692 505612 324748
rect 316916 324676 505612 324692
rect 325764 324568 537644 324584
rect 325764 324512 325780 324568
rect 325836 324512 537572 324568
rect 537628 324512 537644 324568
rect 325764 324496 537644 324512
rect 332260 324388 554444 324404
rect 332260 324332 332276 324388
rect 332332 324332 554372 324388
rect 554428 324332 554444 324388
rect 332260 324316 554444 324332
rect 104116 324208 166364 324224
rect 104116 324152 104132 324208
rect 104188 324152 166292 324208
rect 166348 324152 166364 324208
rect 104116 324136 166364 324152
rect 118340 324028 161884 324044
rect 118340 323972 118356 324028
rect 118412 323972 161812 324028
rect 161868 323972 161884 324028
rect 118340 323956 161884 323972
rect 371572 324028 485564 324044
rect 371572 323972 371588 324028
rect 371644 323972 485492 324028
rect 485548 323972 485564 324028
rect 371572 323956 485564 323972
rect 151156 323848 161100 323864
rect 151156 323792 151172 323848
rect 151228 323792 161028 323848
rect 161084 323792 161100 323848
rect 151156 323776 161100 323792
rect 380308 322948 672492 322964
rect 380308 322892 380324 322948
rect 380380 322892 672420 322948
rect 672476 322892 672492 322948
rect 380308 322876 672492 322892
rect 379524 322768 672716 322784
rect 379524 322712 379540 322768
rect 379596 322712 672644 322768
rect 672700 322712 672716 322768
rect 379524 322696 672716 322712
rect 378628 322588 672828 322604
rect 378628 322532 378644 322588
rect 378700 322532 672756 322588
rect 672812 322532 672828 322588
rect 378628 322516 672828 322532
rect 701748 322408 705756 322424
rect 701748 322352 701764 322408
rect 701820 322352 705684 322408
rect 705740 322352 705756 322408
rect 701748 322336 705756 322352
rect 378180 322228 379836 322244
rect 378180 322172 378196 322228
rect 378252 322172 379764 322228
rect 379820 322172 379836 322228
rect 378180 322156 379836 322172
rect 93812 320968 159644 320984
rect 93812 320912 93828 320968
rect 93884 320912 159572 320968
rect 159628 320912 159644 320968
rect 93812 320896 159644 320912
rect 379860 319528 557804 319544
rect 379860 319472 379876 319528
rect 379932 319472 557732 319528
rect 557788 319472 557804 319528
rect 379860 319456 557804 319472
rect 377956 317368 379836 317384
rect 377956 317312 377972 317368
rect 378028 317312 379764 317368
rect 379820 317312 379836 317368
rect 377956 317296 379836 317312
rect 76116 314308 84604 314324
rect 76116 314252 76132 314308
rect 76188 314252 84532 314308
rect 84588 314252 84604 314308
rect 76116 314236 84604 314252
rect 76340 312508 84044 312524
rect 76340 312452 76356 312508
rect 76412 312452 83972 312508
rect 84028 312452 84044 312508
rect 76340 312436 84044 312452
rect 379748 312508 460364 312524
rect 379748 312452 379764 312508
rect 379820 312452 460292 312508
rect 460348 312452 460364 312508
rect 379748 312436 460364 312452
rect 765600 311500 777600 323500
rect 76116 311428 84156 311444
rect 76116 311372 76132 311428
rect 76188 311372 84084 311428
rect 84140 311372 84156 311428
rect 76116 311356 84156 311372
rect 378740 309988 664428 310004
rect 378740 309932 378756 309988
rect 378812 309932 664356 309988
rect 664412 309932 664428 309988
rect 378740 309916 664428 309932
rect 400 297500 12400 309500
rect 379524 309268 458684 309284
rect 379524 309212 379540 309268
rect 379596 309212 458612 309268
rect 458668 309212 458684 309268
rect 379524 309196 458684 309212
rect 99076 308188 163004 308204
rect 99076 308132 99092 308188
rect 99148 308132 162932 308188
rect 162988 308132 163004 308188
rect 99076 308116 163004 308132
rect 181620 308188 203324 308204
rect 181620 308132 181636 308188
rect 181692 308132 203252 308188
rect 203308 308132 203324 308188
rect 181620 308116 203324 308132
rect 334164 308188 377708 308204
rect 334164 308132 334180 308188
rect 334236 308132 377636 308188
rect 377692 308132 377708 308188
rect 334164 308116 377708 308132
rect 154628 308008 190668 308024
rect 154628 307952 154644 308008
rect 154700 307952 190596 308008
rect 190652 307952 190668 308008
rect 154628 307936 190668 307952
rect 238404 308008 252044 308024
rect 238404 307952 238420 308008
rect 238476 307952 251972 308008
rect 252028 307952 252044 308008
rect 238404 307936 252044 307952
rect 282084 308008 316892 308024
rect 282084 307952 282100 308008
rect 282156 307952 316820 308008
rect 316876 307952 316892 308008
rect 282084 307936 316892 307952
rect 320724 308008 426764 308024
rect 320724 307952 320740 308008
rect 320796 307952 426692 308008
rect 426748 307952 426764 308008
rect 320724 307936 426764 307952
rect 102436 307828 164684 307844
rect 102436 307772 102452 307828
rect 102508 307772 164612 307828
rect 164668 307772 164684 307828
rect 102436 307756 164684 307772
rect 165380 307828 183164 307844
rect 165380 307772 165396 307828
rect 165452 307772 183092 307828
rect 183148 307772 183164 307828
rect 165380 307756 183164 307772
rect 248484 307828 272204 307844
rect 248484 307772 248500 307828
rect 248556 307772 272132 307828
rect 272188 307772 272204 307828
rect 248484 307756 272204 307772
rect 317364 307828 336828 307844
rect 317364 307772 317380 307828
rect 317436 307772 336756 307828
rect 336812 307772 336828 307828
rect 317364 307756 336828 307772
rect 369444 307828 532492 307844
rect 369444 307772 369460 307828
rect 369516 307772 532420 307828
rect 532476 307772 532492 307828
rect 369444 307756 532492 307772
rect 159780 307648 193244 307664
rect 159780 307592 159796 307648
rect 159852 307592 193172 307648
rect 193228 307592 193244 307648
rect 159780 307576 193244 307592
rect 196516 307648 210044 307664
rect 196516 307592 196532 307648
rect 196588 307592 209972 307648
rect 210028 307592 210044 307648
rect 196516 307576 210044 307592
rect 241764 307648 262124 307664
rect 241764 307592 241780 307648
rect 241836 307592 262052 307648
rect 262108 307592 262124 307648
rect 241764 307576 262124 307592
rect 265284 307648 304012 307664
rect 265284 307592 265300 307648
rect 265356 307592 303940 307648
rect 303996 307592 304012 307648
rect 265284 307576 304012 307592
rect 313780 307648 337052 307664
rect 313780 307592 313796 307648
rect 313852 307592 336980 307648
rect 337036 307592 337052 307648
rect 313780 307576 337052 307592
rect 377844 307648 550188 307664
rect 377844 307592 377860 307648
rect 377916 307592 550116 307648
rect 550172 307592 550188 307648
rect 377844 307576 550188 307592
rect 100756 307468 164796 307484
rect 100756 307412 100772 307468
rect 100828 307412 164724 307468
rect 164780 307412 164796 307468
rect 100756 307396 164796 307412
rect 165604 307468 181484 307484
rect 165604 307412 165620 307468
rect 165676 307412 181412 307468
rect 181468 307412 181484 307468
rect 165604 307396 181484 307412
rect 201332 307468 206684 307484
rect 201332 307412 201348 307468
rect 201404 307412 206612 307468
rect 206668 307412 206684 307468
rect 201332 307396 206684 307412
rect 234596 307468 245324 307484
rect 234596 307412 234612 307468
rect 234668 307412 245252 307468
rect 245308 307412 245324 307468
rect 234596 307396 245324 307412
rect 261924 307468 285644 307484
rect 261924 307412 261940 307468
rect 261996 307412 285572 307468
rect 285628 307412 285644 307468
rect 261924 307396 285644 307412
rect 297204 307468 337276 307484
rect 297204 307412 297220 307468
rect 297276 307412 337204 307468
rect 337260 307412 337276 307468
rect 297204 307396 337276 307412
rect 377844 307468 551084 307484
rect 377844 307412 377860 307468
rect 377916 307412 551012 307468
rect 551068 307412 551084 307468
rect 377844 307396 551084 307412
rect 362724 304048 520620 304064
rect 362724 303992 362740 304048
rect 362796 303992 520548 304048
rect 520604 303992 520620 304048
rect 362724 303976 520620 303992
rect 364404 303868 522412 303884
rect 364404 303812 364420 303868
rect 364476 303812 522340 303868
rect 522396 303812 522412 303868
rect 364404 303796 522412 303812
rect 342564 303508 474588 303524
rect 342564 303452 342580 303508
rect 342636 303452 474516 303508
rect 474572 303452 474588 303508
rect 342564 303436 474588 303452
rect 344244 303328 479628 303344
rect 344244 303272 344260 303328
rect 344316 303272 479556 303328
rect 479612 303272 479628 303328
rect 344244 303256 479628 303272
rect 357684 303148 506508 303164
rect 357684 303092 357700 303148
rect 357756 303092 506436 303148
rect 506492 303092 506508 303148
rect 357684 303076 506508 303092
rect 385908 302608 541788 302624
rect 385908 302552 385924 302608
rect 385980 302552 541716 302608
rect 541772 302552 541788 302608
rect 385908 302536 541788 302552
rect 83172 302428 652332 302444
rect 83172 302372 83188 302428
rect 83244 302372 652260 302428
rect 652316 302372 652332 302428
rect 83172 302356 652332 302372
rect 286004 301888 354972 301904
rect 286004 301832 286020 301888
rect 286076 301832 354900 301888
rect 354956 301832 354972 301888
rect 286004 301816 354972 301832
rect 285556 301708 356204 301724
rect 285556 301652 285572 301708
rect 285628 301652 356132 301708
rect 356188 301652 356204 301708
rect 285556 301636 356204 301652
rect 76340 301528 670476 301544
rect 76340 301472 76356 301528
rect 76412 301472 670404 301528
rect 670460 301472 670476 301528
rect 76340 301456 670476 301472
rect 285780 300808 352844 300824
rect 285780 300752 285796 300808
rect 285852 300752 352772 300808
rect 352828 300752 352844 300808
rect 285780 300736 352844 300752
rect 298996 300088 381852 300104
rect 298996 300032 299012 300088
rect 299068 300032 381780 300088
rect 381836 300032 381852 300088
rect 298996 300016 381852 300032
rect 302804 299908 389804 299924
rect 302804 299852 302820 299908
rect 302876 299852 389732 299908
rect 389788 299852 389804 299908
rect 302804 299836 389804 299852
rect 292276 299548 338508 299564
rect 292276 299492 292292 299548
rect 292348 299492 338436 299548
rect 338492 299492 338508 299548
rect 292276 299476 338508 299492
rect 294516 299368 343548 299384
rect 294516 299312 294532 299368
rect 294588 299312 343476 299368
rect 343532 299312 343548 299368
rect 294516 299296 343548 299312
rect 302580 299188 391484 299204
rect 302580 299132 302596 299188
rect 302652 299132 391412 299188
rect 391468 299132 391484 299188
rect 302580 299116 391484 299132
rect 310980 295768 334476 295784
rect 310980 295712 310996 295768
rect 311052 295712 334404 295768
rect 334460 295712 334476 295768
rect 310980 295696 334476 295712
rect 378180 294868 557804 294884
rect 378180 294812 378196 294868
rect 378252 294812 557732 294868
rect 557788 294812 557804 294868
rect 378180 294796 557804 294812
rect 482116 294328 611452 294344
rect 482116 294272 482132 294328
rect 482188 294272 611380 294328
rect 611436 294272 611452 294328
rect 482116 294256 611452 294272
rect 335956 294148 671372 294164
rect 335956 294092 335972 294148
rect 336028 294092 671300 294148
rect 671356 294092 671372 294148
rect 335956 294076 671372 294092
rect 537556 293968 538652 293984
rect 537556 293912 537572 293968
rect 537628 293912 538580 293968
rect 538636 293912 538652 293968
rect 537556 293896 538652 293912
rect 550100 293608 644492 293624
rect 550100 293552 550116 293608
rect 550172 293552 644420 293608
rect 644476 293552 644492 293608
rect 550100 293536 644492 293552
rect 539236 293428 638780 293444
rect 539236 293372 539252 293428
rect 539308 293372 638708 293428
rect 638764 293372 638780 293428
rect 539236 293356 638780 293372
rect 538564 293248 638220 293264
rect 538564 293192 538580 293248
rect 538636 293192 638148 293248
rect 638204 293192 638220 293248
rect 538564 293176 638220 293192
rect 510676 293068 628140 293084
rect 510676 293012 510692 293068
rect 510748 293012 628068 293068
rect 628124 293012 628140 293068
rect 510676 292996 628140 293012
rect 488836 292888 606300 292904
rect 488836 292832 488852 292888
rect 488908 292832 606228 292888
rect 606284 292832 606300 292888
rect 488836 292816 606300 292832
rect 498916 292708 623324 292724
rect 498916 292652 498932 292708
rect 498988 292652 623252 292708
rect 623308 292652 623324 292708
rect 498916 292636 623324 292652
rect 497236 292528 622876 292544
rect 497236 292472 497252 292528
rect 497308 292472 622804 292528
rect 622860 292472 622876 292528
rect 497236 292456 622876 292472
rect 465316 292348 646620 292364
rect 465316 292292 465332 292348
rect 465388 292292 646548 292348
rect 646604 292292 646620 292348
rect 465316 292276 646620 292292
rect 461956 292168 467083 292184
rect 461956 292112 461972 292168
rect 462028 292112 462756 292168
rect 462812 292112 467083 292168
rect 461956 292096 467083 292112
rect 609908 292168 626683 292184
rect 609908 292112 609924 292168
rect 609980 292112 626683 292168
rect 609908 292096 626683 292112
rect 321172 291988 428892 292004
rect 321172 291932 321188 291988
rect 321244 291932 428820 291988
rect 428876 291932 428892 291988
rect 321172 291916 428892 291932
rect 466995 291824 467083 292096
rect 626595 292004 626683 292096
rect 609796 291988 620748 292004
rect 609796 291932 609812 291988
rect 609868 291932 620676 291988
rect 620732 291932 620748 291988
rect 609796 291916 620748 291932
rect 626595 291988 671148 292004
rect 626595 291932 671076 291988
rect 671132 291932 671148 291988
rect 626595 291916 671148 291932
rect 320948 291808 428668 291824
rect 320948 291752 320964 291808
rect 321020 291752 428596 291808
rect 428652 291752 428668 291808
rect 320948 291736 428668 291752
rect 466995 291808 642588 291824
rect 466995 291752 642516 291808
rect 642572 291752 642588 291808
rect 466995 291736 642588 291752
rect 117892 291628 173308 291644
rect 117892 291572 117908 291628
rect 117964 291572 173236 291628
rect 173292 291572 173308 291628
rect 117892 291556 173308 291572
rect 321396 291628 430460 291644
rect 321396 291572 321412 291628
rect 321468 291572 430388 291628
rect 430444 291572 430460 291628
rect 321396 291556 430460 291572
rect 534196 291628 636764 291644
rect 534196 291572 534212 291628
rect 534268 291572 636692 291628
rect 636748 291572 636764 291628
rect 534196 291556 636764 291572
rect 93364 291448 336044 291464
rect 93364 291392 93380 291448
rect 93436 291392 335972 291448
rect 336028 291392 336044 291448
rect 93364 291376 336044 291392
rect 506420 291448 626236 291464
rect 506420 291392 506436 291448
rect 506492 291392 626164 291448
rect 626220 291392 626236 291448
rect 506420 291376 626236 291392
rect 532516 291268 636316 291284
rect 532516 291212 532532 291268
rect 532588 291212 636244 291268
rect 636300 291212 636316 291268
rect 532516 291196 636316 291212
rect 521316 291088 632060 291104
rect 521316 291032 521332 291088
rect 521388 291032 631988 291088
rect 632044 291032 632060 291088
rect 521316 291016 632060 291032
rect 535876 290908 637324 290924
rect 535876 290852 535892 290908
rect 535948 290852 637252 290908
rect 637308 290852 637324 290908
rect 535876 290836 637324 290852
rect 606212 290728 606636 290744
rect 606212 290672 606228 290728
rect 606284 290672 606636 290728
rect 606212 290656 606636 290672
rect 611364 290728 614588 290744
rect 611364 290672 611380 290728
rect 611436 290672 614588 290728
rect 611364 290656 614588 290672
rect 614724 290728 614923 290744
rect 614724 290672 614740 290728
rect 614796 290672 614923 290728
rect 614724 290656 614923 290672
rect 620660 290728 669916 290744
rect 620660 290672 620676 290728
rect 620732 290672 669844 290728
rect 669900 290672 669916 290728
rect 620660 290656 669916 290672
rect 606548 290564 606636 290656
rect 475396 290548 606412 290564
rect 475396 290492 475412 290548
rect 475468 290492 606340 290548
rect 606396 290492 606412 290548
rect 475396 290476 606412 290492
rect 606548 290548 614364 290564
rect 606548 290492 614292 290548
rect 614348 290492 614364 290548
rect 606548 290476 614364 290492
rect 614500 290384 614588 290656
rect 614835 290564 614923 290656
rect 614835 290548 616492 290564
rect 614835 290492 616420 290548
rect 616476 290492 616492 290548
rect 614835 290476 616492 290492
rect 667476 290548 670252 290564
rect 667476 290492 667492 290548
rect 667548 290492 670180 290548
rect 670236 290492 670252 290548
rect 667476 290476 670252 290492
rect 472036 290368 606412 290384
rect 472036 290312 472052 290368
rect 472108 290312 606340 290368
rect 606396 290312 606412 290368
rect 472036 290296 606412 290312
rect 611028 290368 614364 290384
rect 611028 290312 611044 290368
rect 611100 290312 614292 290368
rect 614348 290312 614364 290368
rect 611028 290296 614364 290312
rect 614500 290368 617612 290384
rect 614500 290312 617540 290368
rect 617596 290312 617612 290368
rect 614500 290296 617612 290312
rect 477860 290188 615708 290204
rect 477860 290132 477876 290188
rect 477932 290132 615636 290188
rect 615692 290132 615708 290188
rect 477860 290116 615708 290132
rect 667028 290188 672268 290204
rect 667028 290132 667044 290188
rect 667100 290132 672196 290188
rect 672252 290132 672268 290188
rect 667028 290116 672268 290132
rect 80260 290008 652668 290024
rect 80260 289952 80276 290008
rect 80332 289952 652596 290008
rect 652652 289952 652668 290008
rect 80260 289936 652668 289952
rect 661652 290008 671036 290024
rect 661652 289952 661668 290008
rect 661724 289952 670964 290008
rect 671020 289952 671036 290008
rect 661652 289936 671036 289952
rect 90675 289828 655580 289844
rect 90675 289772 655508 289828
rect 655564 289772 655580 289828
rect 90675 289756 655580 289772
rect 658292 289828 667116 289844
rect 658292 289772 658308 289828
rect 658364 289772 667044 289828
rect 667100 289772 667116 289828
rect 658292 289756 667116 289772
rect 667252 289828 672380 289844
rect 667252 289772 667268 289828
rect 667324 289772 672308 289828
rect 672364 289772 672380 289828
rect 667252 289756 672380 289772
rect 90675 289664 90763 289756
rect 78804 289648 90763 289664
rect 78804 289592 78820 289648
rect 78876 289592 90763 289648
rect 78804 289576 90763 289592
rect 93252 289108 337612 289124
rect 93252 289052 93268 289108
rect 93324 289052 337540 289108
rect 337596 289052 337612 289108
rect 93252 289036 337612 289052
rect 671844 289108 687612 289124
rect 671844 289052 671860 289108
rect 671916 289052 687540 289108
rect 687596 289052 687612 289108
rect 671844 289036 687612 289052
rect 469124 287488 611116 287504
rect 469124 287432 469140 287488
rect 469196 287432 611044 287488
rect 611100 287432 611116 287488
rect 469124 287416 611116 287432
rect 468564 287308 600588 287324
rect 468564 287252 468580 287308
rect 468636 287252 600516 287308
rect 600572 287252 600588 287308
rect 468564 287236 600588 287252
rect 327892 284788 444124 284804
rect 327892 284732 327908 284788
rect 327964 284732 444052 284788
rect 444108 284732 444124 284788
rect 327892 284716 444124 284732
rect 329572 284248 446700 284264
rect 329572 284192 329588 284248
rect 329644 284192 446628 284248
rect 446684 284192 446700 284248
rect 329572 284176 446700 284192
rect 327668 284068 445356 284084
rect 327668 284012 327684 284068
rect 327740 284012 445284 284068
rect 445340 284012 445356 284068
rect 327668 283996 445356 284012
rect 701972 279388 705756 279404
rect 701972 279332 701988 279388
rect 702044 279332 705684 279388
rect 705740 279332 705756 279388
rect 701972 279316 705756 279332
rect 76116 274168 85164 274184
rect 76116 274112 76132 274168
rect 76188 274112 85092 274168
rect 85148 274112 85164 274168
rect 76116 274096 85164 274112
rect 76452 272188 85164 272204
rect 76452 272132 76468 272188
rect 76524 272132 85092 272188
rect 85148 272132 85164 272188
rect 76452 272116 85164 272132
rect 76116 270748 84268 270764
rect 76116 270692 76132 270748
rect 76188 270692 84196 270748
rect 84252 270692 84268 270748
rect 76116 270676 84268 270692
rect 76228 270568 92444 270584
rect 76228 270512 76244 270568
rect 76300 270512 92372 270568
rect 92428 270512 92444 270568
rect 76228 270496 92444 270512
rect 558388 268768 559372 268784
rect 558388 268712 558404 268768
rect 558460 268712 559300 268768
rect 559356 268712 559372 268768
rect 558388 268696 559372 268712
rect 765600 268500 777600 280500
rect 400 256500 12400 268500
rect 558500 257248 559372 257264
rect 558500 257192 558516 257248
rect 558572 257192 559300 257248
rect 559356 257192 559372 257248
rect 558500 257176 559372 257192
rect 76452 234388 93452 234404
rect 76452 234332 76468 234388
rect 76524 234332 93380 234388
rect 93436 234332 93452 234388
rect 76452 234316 93452 234332
rect 76452 232048 84716 232064
rect 76452 231992 76468 232048
rect 76524 231992 84644 232048
rect 84700 231992 84716 232048
rect 76452 231976 84716 231992
rect 76116 231868 85276 231884
rect 76116 231812 76132 231868
rect 76188 231812 85204 231868
rect 85260 231812 85276 231868
rect 76116 231796 85276 231812
rect 76116 230428 85052 230444
rect 76116 230372 76132 230428
rect 76188 230372 84980 230428
rect 85036 230372 85052 230428
rect 76116 230356 85052 230372
rect 76228 230248 93228 230264
rect 76228 230192 76244 230248
rect 76300 230192 93156 230248
rect 93212 230192 93228 230248
rect 76228 230176 93228 230192
rect 400 215500 12400 227500
rect 765600 225500 777600 237500
rect 84740 206848 93228 206864
rect 84740 206792 84756 206848
rect 84812 206792 93156 206848
rect 93212 206792 93228 206848
rect 84740 206776 93228 206792
rect 84628 206668 92444 206684
rect 84628 206612 84644 206668
rect 84700 206612 92372 206668
rect 92428 206612 92444 206668
rect 84628 206596 92444 206612
rect 701412 193528 705756 193544
rect 701412 193472 701428 193528
rect 701484 193472 705684 193528
rect 705740 193472 705756 193528
rect 701412 193456 705756 193472
rect 76116 191908 85388 191924
rect 76116 191852 76132 191908
rect 76188 191852 85316 191908
rect 85372 191852 85388 191908
rect 76116 191836 85388 191852
rect 83844 191188 90428 191204
rect 83844 191132 83860 191188
rect 83916 191132 90356 191188
rect 90412 191132 90428 191188
rect 83844 191116 90428 191132
rect 78915 191008 92668 191024
rect 78915 190952 92596 191008
rect 92652 190952 92668 191008
rect 78915 190936 92668 190952
rect 78915 190844 79003 190936
rect 76116 190828 79003 190844
rect 76116 190772 76132 190828
rect 76188 190772 79003 190828
rect 76116 190756 79003 190772
rect 76452 189928 84380 189944
rect 76452 189872 76468 189928
rect 76524 189872 84308 189928
rect 84364 189872 84380 189928
rect 76452 189856 84380 189872
rect 76116 188668 84940 188684
rect 76116 188612 76132 188668
rect 76188 188612 84868 188668
rect 84924 188612 84940 188668
rect 76116 188596 84940 188612
rect 76228 188488 93340 188504
rect 76228 188432 76244 188488
rect 76300 188432 93268 188488
rect 93324 188432 93340 188488
rect 76228 188416 93340 188432
rect 400 174500 12400 186500
rect 558388 185788 559708 185804
rect 558388 185732 558404 185788
rect 558460 185732 559636 185788
rect 559692 185732 559708 185788
rect 558388 185716 559708 185732
rect 558612 184888 559148 184904
rect 558612 184832 558628 184888
rect 558684 184832 559076 184888
rect 559132 184832 559148 184888
rect 558612 184816 559148 184832
rect 765600 182500 777600 194500
rect 701972 150508 705756 150524
rect 701972 150452 701988 150508
rect 702044 150452 705684 150508
rect 705740 150452 705756 150508
rect 701972 150436 705756 150452
rect 400 133500 12400 145500
rect 558388 143668 559372 143684
rect 558388 143612 558404 143668
rect 558460 143612 559300 143668
rect 559356 143612 559372 143668
rect 558388 143596 559372 143612
rect 558500 142588 559484 142604
rect 558500 142532 558516 142588
rect 558572 142532 559412 142588
rect 559468 142532 559484 142588
rect 558500 142516 559484 142532
rect 559396 142048 671932 142064
rect 559396 141992 559412 142048
rect 559468 141992 671860 142048
rect 671916 141992 671932 142048
rect 559396 141976 671932 141992
rect 671620 141868 700604 141884
rect 671620 141812 671636 141868
rect 671692 141812 700532 141868
rect 700588 141812 700604 141868
rect 671620 141796 700604 141812
rect 671732 141148 694668 141164
rect 671732 141092 671748 141148
rect 671804 141092 694596 141148
rect 694652 141092 694668 141148
rect 671732 141076 694668 141092
rect 618868 140176 624780 140264
rect 618868 140068 618956 140176
rect 618868 140012 618884 140068
rect 618940 140012 618956 140068
rect 618868 139996 618956 140012
rect 619092 140068 623436 140084
rect 619092 140012 619108 140068
rect 619164 140012 623364 140068
rect 623420 140012 623436 140068
rect 619092 139996 623436 140012
rect 624692 140068 624780 140176
rect 624692 140012 624708 140068
rect 624764 140012 624780 140068
rect 624692 139996 624780 140012
rect 649332 140176 657820 140264
rect 649332 140068 649420 140176
rect 649332 140012 649348 140068
rect 649404 140012 649420 140068
rect 649332 139996 649420 140012
rect 649556 140068 657148 140084
rect 649556 140012 649572 140068
rect 649628 140012 657076 140068
rect 657132 140012 657148 140068
rect 649556 139996 657148 140012
rect 657732 140068 657820 140176
rect 657732 140012 657748 140068
rect 657804 140012 657820 140068
rect 657732 139996 657820 140012
rect 619092 139888 631500 139904
rect 619092 139832 619108 139888
rect 619164 139832 631428 139888
rect 631484 139832 631500 139888
rect 619092 139816 631500 139832
rect 649668 139888 655804 139904
rect 649668 139832 649684 139888
rect 649740 139832 655732 139888
rect 655788 139832 655804 139888
rect 649668 139816 655804 139832
rect 618308 139708 619068 139724
rect 618308 139652 618324 139708
rect 618380 139652 618996 139708
rect 619052 139652 619068 139708
rect 618308 139636 619068 139652
rect 619316 139708 632844 139724
rect 619316 139652 619332 139708
rect 619388 139652 632772 139708
rect 632828 139652 632844 139708
rect 619316 139636 632844 139652
rect 650900 139708 656476 139724
rect 650900 139652 650916 139708
rect 650972 139652 656404 139708
rect 656460 139652 656476 139708
rect 650900 139636 656476 139652
rect 618532 139528 622092 139544
rect 618532 139472 618548 139528
rect 618604 139472 622020 139528
rect 622076 139472 622092 139528
rect 618532 139456 622092 139472
rect 622452 139528 638892 139544
rect 622452 139472 622468 139528
rect 622524 139472 638820 139528
rect 638876 139472 638892 139528
rect 622452 139456 638892 139472
rect 666468 139528 671148 139544
rect 666468 139472 666484 139528
rect 666540 139472 671076 139528
rect 671132 139472 671148 139528
rect 765600 139500 777600 151500
rect 666468 139456 671148 139472
rect 650788 132688 658044 132704
rect 650788 132632 650804 132688
rect 650860 132632 657972 132688
rect 658028 132632 658044 132688
rect 650788 132616 658044 132632
rect 664564 132688 670812 132704
rect 664564 132632 664580 132688
rect 664636 132632 670740 132688
rect 670796 132632 670812 132688
rect 664564 132616 670812 132632
rect 659636 132508 670028 132524
rect 659636 132452 659652 132508
rect 659708 132452 669956 132508
rect 670012 132452 670028 132508
rect 659636 132436 670028 132452
rect 649780 132328 653564 132344
rect 649780 132272 649796 132328
rect 649852 132272 653492 132328
rect 653548 132272 653564 132328
rect 649780 132256 653564 132272
rect 666804 132328 671148 132344
rect 666804 132272 666820 132328
rect 666876 132272 671076 132328
rect 671132 132272 671148 132328
rect 666804 132256 671148 132272
rect 665124 131068 671036 131084
rect 665124 131012 665140 131068
rect 665196 131012 670964 131068
rect 671020 131012 671036 131068
rect 665124 130996 671036 131012
rect 646308 126748 656028 126764
rect 646308 126692 646324 126748
rect 646380 126692 655956 126748
rect 656012 126692 656028 126748
rect 646308 126676 656028 126692
rect 646980 126028 655580 126044
rect 646980 125972 646996 126028
rect 647052 125972 655508 126028
rect 655564 125972 655580 126028
rect 646980 125956 655580 125972
rect 641492 124948 654796 124964
rect 641492 124892 641508 124948
rect 641564 124892 654724 124948
rect 654780 124892 654796 124948
rect 641492 124876 654796 124892
rect 628724 124768 655468 124784
rect 628724 124712 628740 124768
rect 628796 124712 655396 124768
rect 655452 124712 655468 124768
rect 628724 124696 655468 124712
rect 628052 124588 655132 124604
rect 628052 124532 628068 124588
rect 628124 124532 655060 124588
rect 655116 124532 655132 124588
rect 628052 124516 655132 124532
rect 626036 124408 655244 124424
rect 626036 124352 626052 124408
rect 626108 124352 655172 124408
rect 655228 124352 655244 124408
rect 626036 124336 655244 124352
rect 642724 124228 648524 124244
rect 642724 124172 642740 124228
rect 642796 124172 648452 124228
rect 648508 124172 648524 124228
rect 642724 124156 648524 124172
rect 638355 123328 647964 123344
rect 638355 123272 647892 123328
rect 647948 123272 647964 123328
rect 638355 123256 647964 123272
rect 638355 123164 638443 123256
rect 618756 123148 638443 123164
rect 618756 123092 618772 123148
rect 618828 123092 638443 123148
rect 618756 123076 638443 123092
rect 621332 122968 655020 122984
rect 621332 122912 621348 122968
rect 621404 122912 654948 122968
rect 655004 122912 655020 122968
rect 621332 122896 655020 122912
rect 621444 122788 670252 122804
rect 621444 122732 621460 122788
rect 621516 122732 670180 122788
rect 670236 122732 670252 122788
rect 621444 122716 670252 122732
rect 654932 120808 655244 120824
rect 654932 120752 654948 120808
rect 655004 120752 655172 120808
rect 655228 120752 655244 120808
rect 654932 120736 655244 120752
rect 651796 110548 655580 110564
rect 651796 110492 651812 110548
rect 651868 110492 655508 110548
rect 655564 110492 655580 110548
rect 651796 110476 655580 110492
rect 701860 107488 705756 107504
rect 701860 107432 701876 107488
rect 701932 107432 705684 107488
rect 705740 107432 705756 107488
rect 701860 107416 705756 107432
rect 400 92500 12400 104500
rect 622564 100648 628700 100664
rect 622564 100592 622580 100648
rect 622636 100592 628628 100648
rect 628684 100592 628700 100648
rect 622564 100576 628700 100592
rect 649556 100648 654348 100664
rect 649556 100592 649572 100648
rect 649628 100592 654276 100648
rect 654332 100592 654348 100648
rect 649556 100576 654348 100592
rect 622676 100468 631276 100484
rect 622676 100412 622692 100468
rect 622748 100412 631204 100468
rect 631260 100412 631276 100468
rect 622676 100396 631276 100412
rect 644964 99568 655804 99584
rect 644964 99512 644980 99568
rect 645036 99512 655732 99568
rect 655788 99512 655804 99568
rect 644964 99496 655804 99512
rect 622228 99388 633852 99404
rect 622228 99332 622244 99388
rect 622300 99332 633780 99388
rect 633836 99332 633852 99388
rect 622228 99316 633852 99332
rect 641716 99388 655468 99404
rect 641716 99332 641732 99388
rect 641788 99332 655396 99388
rect 655452 99332 655468 99388
rect 641716 99316 655468 99332
rect 622452 99208 635868 99224
rect 622452 99152 622468 99208
rect 622524 99152 635796 99208
rect 635852 99152 635868 99208
rect 622452 99136 635868 99152
rect 639028 99208 655356 99224
rect 639028 99152 639044 99208
rect 639100 99152 655284 99208
rect 655340 99152 655356 99208
rect 639028 99136 655356 99152
rect 558388 96688 559372 96704
rect 558388 96632 558404 96688
rect 558460 96632 559300 96688
rect 559356 96632 559372 96688
rect 558388 96616 559372 96632
rect 765600 96500 777600 108500
rect 558612 90748 559372 90764
rect 558612 90692 558628 90748
rect 558684 90692 559300 90748
rect 559356 90692 559372 90748
rect 558612 90676 559372 90692
rect 93140 83008 336044 83024
rect 93140 82952 93156 83008
rect 93212 82952 335972 83008
rect 336028 82952 336044 83008
rect 93140 82936 336044 82952
rect 558388 82288 585468 82304
rect 558388 82232 558404 82288
rect 558460 82232 585396 82288
rect 585452 82232 585468 82288
rect 558388 82216 585468 82232
rect 558612 82108 585692 82124
rect 558612 82052 558628 82108
rect 558684 82052 585620 82108
rect 585676 82052 585692 82108
rect 558612 82036 585692 82052
rect 559172 81928 585916 81944
rect 559172 81872 559188 81928
rect 559244 81872 585844 81928
rect 585900 81872 585916 81928
rect 559172 81856 585916 81872
rect 620548 80848 631723 80864
rect 620548 80792 620564 80848
rect 620620 80792 631723 80848
rect 620548 80776 631723 80792
rect 631635 80684 631723 80776
rect 620324 80668 628140 80684
rect 620324 80612 620340 80668
rect 620396 80612 628068 80668
rect 628124 80612 628140 80668
rect 620324 80596 628140 80612
rect 631635 80668 645164 80684
rect 631635 80612 645092 80668
rect 645148 80612 645164 80668
rect 631635 80596 645164 80612
rect 494324 71488 618508 71504
rect 494324 71432 494340 71488
rect 494396 71432 618436 71488
rect 618492 71432 618508 71488
rect 494324 71416 618508 71432
rect 176244 71308 620412 71324
rect 176244 71252 176260 71308
rect 176316 71252 620340 71308
rect 620396 71252 620412 71308
rect 176244 71236 620412 71252
rect 519636 71128 619404 71144
rect 519636 71072 519652 71128
rect 519708 71072 619332 71128
rect 619388 71072 619404 71128
rect 519636 71056 619404 71072
rect 505860 70948 618060 70964
rect 505860 70892 505876 70948
rect 505932 70892 617988 70948
rect 618044 70892 618060 70948
rect 505860 70876 618060 70892
rect 324868 70768 548508 70784
rect 324868 70712 324884 70768
rect 324940 70712 548436 70768
rect 548492 70712 548508 70768
rect 324868 70696 548508 70712
rect 257780 70588 539212 70604
rect 257780 70532 257796 70588
rect 257852 70532 539140 70588
rect 539196 70532 539212 70588
rect 257780 70516 539212 70532
rect 108500 400 120500 12400
rect 163500 400 175500 12400
rect 218500 400 230500 12400
rect 273500 400 285500 12400
rect 328500 400 340500 12400
rect 383500 400 395500 12400
rect 438500 400 450500 12400
rect 493500 400 505500 12400
rect 548500 400 560500 12400
rect 603500 400 615500 12400
rect 658500 400 670500 12400
rect 0 0 1 1
use caravel_gf180_pdn  caravel_gf180_pdn_0
timestamp 1483923398
transform 1 0 0 0 1 0
box 69800 69800 708200 950200
use caravel_logo  caravel_logo_0
timestamp 1638586901
transform 1 0 192076 0 1 1481
box -1680 0 10000 10373
use caravel_motto  caravel_motto_0
timestamp 1668623937
transform 1 0 -1570920 0 1 -71280
box 1867050 75020 1886060 78420
use caravel_clocking  clock_ctrl
timestamp 1654631816
transform 1 0 619608 0 1 110000
box 4 410 36000 14000
use copyright_block  copyright_block_0
timestamp 1654652987
transform 1 0 132720 0 1 7725
box -429 -6331 18270 2667
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1655130296
transform -1 0 708000 0 -1 110000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1655130296
transform -1 0 708000 0 -1 153000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1655130296
transform 1 0 70000 0 1 255000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1655130296
transform 1 0 70000 0 1 214000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1655130296
transform 1 0 70000 0 1 173000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1655130296
transform -1 0 708000 0 -1 583000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1655130296
transform -1 0 708000 0 -1 626000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1655130296
transform -1 0 708000 0 -1 669000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1655130296
transform -1 0 708000 0 -1 712000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1655130296
transform -1 0 708000 0 -1 841000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1655130296
transform -1 0 708000 0 -1 755000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1655130296
transform -1 0 708000 0 -1 927000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1655130296
transform 0 1 656000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1655130296
transform 0 1 546000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1655130296
transform 0 1 491000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1655130296
transform 0 1 436000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1655130296
transform -1 0 708000 0 -1 196000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1655130296
transform -1 0 708000 0 -1 239000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1655130296
transform -1 0 708000 0 -1 282000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1655130296
transform -1 0 708000 0 -1 325000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1655130296
transform -1 0 708000 0 -1 368000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1655130296
transform -1 0 708000 0 -1 540000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1655130296
transform 0 1 326000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1655130296
transform 0 1 271000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1655130296
transform 0 1 216000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1655130296
transform 0 1 161000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1655130296
transform 0 1 106000 -1 0 950000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1655130296
transform 1 0 70000 0 1 911000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1655130296
transform 1 0 70000 0 1 747000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1655130296
transform 1 0 70000 0 1 706000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1655130296
transform 1 0 70000 0 1 665000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1655130296
transform 1 0 70000 0 1 624000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1655130296
transform 1 0 70000 0 1 583000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1655130296
transform 1 0 70000 0 1 542000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1655130296
transform 1 0 70000 0 1 501000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1655130296
transform 1 0 70000 0 1 378000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1655130296
transform 1 0 70000 0 1 337000
box -100 -200 6604 35200
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1655130296
transform 1 0 70000 0 1 296000
box -100 -200 6604 35200
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1654613330
transform -1 0 691000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1654613330
transform 0 -1 702000 1 0 892000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1654613330
transform -1 0 581000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1654613330
transform -1 0 526000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1654613330
transform -1 0 471000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1654613330
transform -1 0 306000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1654613330
transform -1 0 361000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1654613330
transform -1 0 251000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block_007  gpio_defaults_block_007_0
timestamp 1654613370
transform 0 -1 702000 1 0 247000
box 0 0 14271 1235
use gpio_defaults_block_007  gpio_defaults_block_007_1
timestamp 1654613370
transform 0 -1 702000 1 0 204000
box 0 0 14271 1235
use gpio_defaults_block_007  gpio_defaults_block_007_2
timestamp 1654613370
transform 0 -1 702000 1 0 161000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1654613330
transform -1 0 141000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1654613330
transform -1 0 196000 0 -1 944000
box 0 0 14271 1235
use gpio_defaults_block_009  gpio_defaults_block_009_0
timestamp 1654613388
transform 0 -1 702000 1 0 118000
box 0 0 14271 1235
use gpio_defaults_block_009  gpio_defaults_block_009_1
timestamp 1654613388
transform 0 -1 702000 1 0 75000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1654613330
transform 0 1 76000 -1 0 946000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1654613330
transform 0 -1 702000 1 0 806000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1654613330
transform 0 -1 702000 1 0 720000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1654613330
transform 0 1 76000 -1 0 741000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1654613330
transform 0 1 76000 -1 0 782000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1654613330
transform 0 -1 702000 1 0 677000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1654613330
transform 0 -1 702000 1 0 634000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1654613330
transform 0 1 76000 -1 0 618000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1654613330
transform 0 1 76000 -1 0 659000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1654613330
transform 0 1 76000 -1 0 700000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1654613330
transform 0 -1 702000 1 0 591000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1654613330
transform 0 -1 702000 1 0 548000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1654613330
transform 0 1 76000 -1 0 536000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1654613330
transform 0 1 76000 -1 0 577000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1654613330
transform 0 -1 702000 1 0 505000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1654613330
transform 0 1 76000 -1 0 413000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1654613330
transform 0 -1 702000 1 0 333000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1654613330
transform 0 1 76000 -1 0 372000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1654613330
transform 0 -1 702000 1 0 290000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1654613330
transform 0 1 76000 -1 0 331000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1654613330
transform 0 1 76000 -1 0 290000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1654613330
transform 0 1 76000 -1 0 249000
box 0 0 14271 1235
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1654613330
transform 0 1 76000 -1 0 208000
box 0 0 14271 1235
use housekeeping  housekeeping
timestamp 1654687298
transform 1 0 611608 0 1 139579
box -28 0 60000 150000
use mgmt_protect  mgmt_buffers
timestamp 1654981632
transform 1 0 160000 0 1 308800
box 0 0 220000 15000
use user_project_wrapper  mprj ../maglef
timestamp 1655473269
transform 1 0 85972 0 1 334184
box -3036 -1244 603020 601004
use open_source  open_source_0 hexdigits
timestamp 1638586442
transform 1 0 237080 0 1 -3420
box 660 4580 25800 14430
use chip_io  padframe
timestamp 1668016291
transform 1 0 0 0 1 0
box 0 0 776000 1014000
use digital_pll  pll
timestamp 1654786971
transform 1 0 619608 0 1 80600
box 0 0 34000 20000
use simple_por  simple_por_0 ../macros/simple_por/maglef
timestamp 1655473345
transform 0 -1 676702 1 0 98600
box 24 74 25112 8716
use mgmt_core_wrapper  soc ../maglef
timestamp 1655473382
transform 1 0 90000 0 1 80600
box -1060 -400 471012 200400
use spare_logic_block  spare_logic\[0\]
timestamp 1654780538
transform 1 0 630640 0 1 310218
box -56 -56 15000 14000
use spare_logic_block  spare_logic\[1\]
timestamp 1654780538
transform 1 0 486000 0 1 310728
box -56 -56 15000 14000
use spare_logic_block  spare_logic\[2\]
timestamp 1654780538
transform 1 0 386000 0 1 310728
box -56 -56 15000 14000
use spare_logic_block  spare_logic\[3\]
timestamp 1654780538
transform 1 0 112000 0 1 310728
box -56 -56 15000 14000
use user_id_textblock  user_id_textblock_0
timestamp 1668623287
transform 1 0 47200 0 1 580
box 0 0 50660 12090
use user_id_programming  user_id_value
timestamp 1655126753
transform 1 0 649450 0 1 132400
box 0 0 22053 2313
<< labels >>
flabel metal5 108500 400 120500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 163500 400 175500 12400 0 FreeSans 24000 0 0 0 resetb
port 446 nsew
flabel metal5 273500 400 285500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 328500 400 340500 12400 0 FreeSans 24000 0 0 0 flash_csb
port 5 nsew
flabel metal5 383500 400 395500 12400 0 FreeSans 24000 0 0 0 flash_clk
port 2 nsew
flabel metal5 438500 400 450500 12400 0 FreeSans 24000 0 0 0 flash_io0
port 8 nsew
flabel metal5 493500 400 505500 12400 0 FreeSans 24000 0 0 0 flash_io1
port 13 nsew
flabel metal5 548500 400 560500 12400 0 FreeSans 24000 0 0 0 gpio
port 18 nsew
flabel metal5 603500 400 615500 12400 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 658500 400 670500 12400 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 96500 777600 108500 0 FreeSans 24000 0 0 0 mprj_io[0]
port 29 nsew
flabel metal5 765600 139500 777600 151500 0 FreeSans 24000 0 0 0 mprj_io[1]
port 40 nsew
flabel metal5 765600 182500 777600 194500 0 FreeSans 24000 0 0 0 mprj_io[2]
port 51 nsew
flabel metal5 765600 225500 777600 237500 0 FreeSans 24000 0 0 0 mprj_io[3]
port 60 nsew
flabel metal5 765600 268500 777600 280500 0 FreeSans 24000 0 0 0 mprj_io[4]
port 61 nsew
flabel metal5 765600 311500 777600 323500 0 FreeSans 24000 0 0 0 mprj_io[5]
port 62 nsew
flabel metal5 765600 354500 777600 366500 0 FreeSans 24000 0 0 0 mprj_io[6]
port 63 nsew
flabel metal5 765600 397500 777600 409500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 765600 440500 777600 452500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 765600 483500 777600 495500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 526500 777600 538500 0 FreeSans 24000 0 0 0 mprj_io[7]
port 64 nsew
flabel metal5 765600 569500 777600 581500 0 FreeSans 24000 0 0 0 mprj_io[8]
port 65 nsew
flabel metal5 765600 612500 777600 624500 0 FreeSans 24000 0 0 0 mprj_io[9]
port 66 nsew
flabel metal5 765600 655500 777600 667500 0 FreeSans 24000 0 0 0 mprj_io[10]
port 30 nsew
flabel metal5 765600 698500 777600 710500 0 FreeSans 24000 0 0 0 mprj_io[11]
port 31 nsew
flabel metal5 765600 741500 777600 753500 0 FreeSans 24000 0 0 0 mprj_io[12]
port 32 nsew
flabel metal5 765600 784500 777600 796500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 827500 777600 839500 0 FreeSans 24000 0 0 0 mprj_io[13]
port 33 nsew
flabel metal5 765600 870500 777600 882500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 765600 913500 777600 925500 0 FreeSans 24000 0 0 0 mprj_io[14]
port 34 nsew
flabel metal5 657500 1007600 669500 1019600 0 FreeSans 24000 0 0 0 mprj_io[15]
port 35 nsew
flabel metal5 602500 1007600 614500 1019600 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 547500 1007600 559500 1019600 0 FreeSans 24000 0 0 0 mprj_io[16]
port 36 nsew
flabel metal5 492500 1007600 504500 1019600 0 FreeSans 24000 0 0 0 mprj_io[17]
port 37 nsew
flabel metal5 437500 1007600 449500 1019600 0 FreeSans 24000 0 0 0 mprj_io[18]
port 38 nsew
flabel metal5 382500 1007600 394500 1019600 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 327500 1007600 339500 1019600 0 FreeSans 24000 0 0 0 mprj_io[19]
port 39 nsew
flabel metal5 272500 1007600 284500 1019600 0 FreeSans 24000 0 0 0 mprj_io[20]
port 41 nsew
flabel metal5 217500 1007600 229500 1019600 0 FreeSans 24000 0 0 0 mprj_io[21]
port 42 nsew
flabel metal5 162500 1007600 174500 1019600 0 FreeSans 24000 0 0 0 mprj_io[22]
port 43 nsew
flabel metal5 107500 1007600 119500 1019600 0 FreeSans 24000 0 0 0 mprj_io[23]
port 44 nsew
flabel metal5 400 912500 12400 924500 0 FreeSans 24000 0 0 0 mprj_io[24]
port 45 nsew
flabel metal5 400 871500 12400 883500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 830500 12400 842500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 789500 12400 801500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 400 748500 12400 760500 0 FreeSans 24000 0 0 0 mprj_io[25]
port 46 nsew
flabel metal5 400 707500 12400 719500 0 FreeSans 24000 0 0 0 mprj_io[26]
port 47 nsew
flabel metal5 400 666500 12400 678500 0 FreeSans 24000 0 0 0 mprj_io[27]
port 48 nsew
flabel metal5 400 625500 12400 637500 0 FreeSans 24000 0 0 0 mprj_io[28]
port 49 nsew
flabel metal5 400 584500 12400 596500 0 FreeSans 24000 0 0 0 mprj_io[29]
port 50 nsew
flabel metal5 400 543500 12400 555500 0 FreeSans 24000 0 0 0 mprj_io[30]
port 52 nsew
flabel metal5 400 502500 12400 514500 0 FreeSans 24000 0 0 0 mprj_io[31]
port 53 nsew
flabel metal5 400 461500 12400 473500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 420500 12400 432500 0 FreeSans 24000 0 0 0 vss
port 449 nsew
flabel metal5 400 379500 12400 391500 0 FreeSans 24000 0 0 0 mprj_io[32]
port 54 nsew
flabel metal5 400 338500 12400 350500 0 FreeSans 24000 0 0 0 mprj_io[33]
port 55 nsew
flabel metal5 400 297500 12400 309500 0 FreeSans 24000 0 0 0 mprj_io[34]
port 56 nsew
flabel metal5 400 256500 12400 268500 0 FreeSans 24000 0 0 0 mprj_io[35]
port 57 nsew
flabel metal5 400 215500 12400 227500 0 FreeSans 24000 0 0 0 mprj_io[36]
port 58 nsew
flabel metal5 400 174500 12400 186500 0 FreeSans 24000 0 0 0 mprj_io[37]
port 59 nsew
flabel metal5 400 133500 12400 145500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 400 92500 12400 104500 0 FreeSans 24000 0 0 0 vdd
port 448 nsew
flabel metal5 218500 400 230500 12400 0 FreeSans 24000 0 0 0 clock
port 0 nsew
<< properties >>
string FIXED_BBOX 0 0 778000 1020000
<< end >>
