magic
tech minimum
timestamp 1670242872
<< properties >>
string FIXED_BBOX 0 0 388 507
<< end >>
