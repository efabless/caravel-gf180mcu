* NGSPICE file created from digital_pll.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_1 EN I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_2 EN I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

.subckt digital_pll VDD VSS clockp[0] clockp[1] dco div[0] div[1] div[2] div[3] div[4]
+ enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
XANTENNA__577__A1 _498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_501_ _501_/I _501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_432_ _411_/Z _432_/A2 _433_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_363_ _363_/I _367_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__568__A1 _495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayint0/I ringosc.dstage\[1\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_415_ _671_/Q _415_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_346_ _666_/Q _681_/Q _346_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__679__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[11\].id.delayen1 _603_/ZN ringosc.dstage\[11\].id.delayen1/I ringosc.dstage\[11\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_329_ _329_/I _478_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_680_ _680_/D _652_/Z _686_/I _680_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_594_ _565_/B _565_/C _580_/Z _594_/B1 _561_/Z _594_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.trim0bar/ZN ringosc.dstage\[10\].id.delayenb1/I
+ ringosc.dstage\[11\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_663_ _663_/D _612_/Z _686_/I _663_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.trim0bar/ZN ringosc.dstage\[9\].id.delayenb1/I
+ ringosc.dstage\[9\].id.delayen0/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_17_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_577_ _498_/Z _577_/A2 _578_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xringosc.dstage\[10\].id.trim0bar _534_/ZN ringosc.dstage\[10\].id.trim0bar/ZN VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_646_ _646_/I _646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_500_ _486_/Z _510_/A1 _500_/B _501_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_431_ _437_/A1 _423_/Z _431_/B _432_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_362_ _356_/Z _368_/A2 _362_/B _367_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_629_ _622_/Z _619_/Z _630_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_414_ _673_/Q _402_/I _414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_345_ input2/Z _396_/A2 _348_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input29_I ext_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_328_ _668_/Q _468_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__604__A1 _604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__669__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_662_ _662_/I _662_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.trim1bar/ZN ringosc.dstage\[9\].id.delayenb1/I
+ ringosc.dstage\[9\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_593_ _593_/I _594_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.trim1bar/ZN ringosc.dstage\[10\].id.delayenb1/I
+ ringosc.dstage\[10\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA_input11_I ext_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_576_ _576_/A1 _588_/A3 _582_/A4 _576_/A4 _578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_645_ _645_/I _645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_430_ _429_/Z _388_/Z _431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_361_ _669_/Q _684_/Q _362_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_559_ _420_/Z _588_/A3 _559_/B _559_/C _562_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_628_ _628_/I _628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_413_ _420_/I _412_/Z _604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_344_ _666_/Q _681_/Q _396_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xringosc.dstage\[4\].id.delayen0 _506_/ZN ringosc.dstage\[4\].id.delayen0/I ringosc.dstage\[5\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_14_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_327_ _327_/I _684_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_592_ _592_/I _592_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_661_ _486_/Z _609_/I _662_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xringosc.dstage\[4\].id.trim1bar _579_/Z ringosc.dstage\[4\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__513__A1 _604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_575_ _507_/Z _575_/A2 _575_/A3 _576_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_644_ _634_/Z _643_/Z _645_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[9\].id.delaybuf0/I ringosc.dstage\[9\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.trim0bar/ZN rebuffer2/I ringosc.ibufp10/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XTAP_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/ZN ringosc.dstage\[10\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_360_ _360_/A1 _360_/A2 _360_/B _360_/C _368_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_489_ _487_/Z _589_/A3 _570_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_558_ _507_/Z _428_/Z _429_/Z _420_/Z _559_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_627_ _622_/Z _619_/Z _628_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_412_ _674_/Q _673_/Q _412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_343_ _341_/Z _360_/A2 _343_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xringosc.dstage\[4\].id.delayen1 _579_/Z ringosc.dstage\[4\].id.delayen1/I ringosc.dstage\[4\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_9_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_326_ _684_/Q _324_/Z _473_/B _327_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_ringosc.dstage\[0\].id.trim1bar_I _546_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I osc VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_591_ _603_/A1 _591_/A2 _591_/B _592_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_660_ _660_/I _660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[3\].id.trim0bar _501_/Z ringosc.dstage\[3\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.trim1bar/ZN rebuffer1/Z ringosc.dstage\[5\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/I ringosc.dstage\[9\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/I ringosc.dstage\[10\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_574_ _340_/Z _428_/Z _576_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_643_ _643_/I _643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_488_ _428_/I _429_/Z _589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_557_ _487_/Z _575_/A3 _559_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_626_ _626_/I _626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__404__A1 _674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_411_ _504_/A2 _388_/Z _411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_342_ _666_/Q _681_/Q _360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_609_ _609_/I _609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_325_ _329_/I _473_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input27_I ext_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_ringosc.dstage\[0\].id.delaybuf1_I ringosc.dstage\[0\].id.delayenb1/I VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_590_ _498_/Z _590_/A2 _591_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__682__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_573_ _573_/A1 _604_/B _573_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_642_ _642_/I _642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_625_ _622_/Z _619_/Z _626_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__486__I _646_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[5\].id.delaybuf0/I rebuffer2/I VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_556_ _582_/A1 _556_/A2 _565_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_487_ _507_/I _487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input1_I dco VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.trim0bar/ZN ringosc.dstage\[1\].id.delayenb1/I
+ ringosc.dstage\[2\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_410_ _410_/A1 _563_/A2 _407_/I _425_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_341_ _667_/Q _682_/Q _341_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayint0/I ringosc.dstage\[8\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_539_ _539_/I _580_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_608_ _643_/I _609_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_324_ _669_/Q _324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_572_ _569_/Z _572_/A2 _582_/A4 _604_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_641_ _634_/Z _631_/Z _642_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput36 _686_/Z clockp[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_555_ _412_/Z _571_/A2 _556_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_624_ _624_/I _624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_486_ _646_/I _486_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__672__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[5\].id.delaybuf1 rebuffer2/Z ringosc.dstage\[5\].id.delayen1/I VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.trim1bar/ZN ringosc.dstage\[1\].id.delayenb1/I
+ ringosc.dstage\[1\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_538_ _538_/I _541_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_340_ _340_/I _340_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_607_ input7/Z _607_/A2 _643_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xringosc.dstage\[1\].id.delayen0 _493_/ZN ringosc.dstage\[1\].id.delayen0/I ringosc.dstage\[2\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_469_ _459_/Z _469_/A2 _469_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_323_ _323_/I _685_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_ringosc.dstage\[0\].id.delayen1_EN _546_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input32_I ext_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[1\].id.trim1bar _562_/ZN ringosc.dstage\[1\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_571_ _539_/I _571_/A2 _582_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_640_ _640_/I _640_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput37 output37/I clockp[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_554_ _554_/A1 _584_/A1 _565_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_485_ _510_/B _646_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_623_ _622_/Z _619_/Z _624_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xringosc.dstage\[1\].id.delayen1 _562_/ZN ringosc.dstage\[1\].id.delayen1/I ringosc.dstage\[1\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_537_ _537_/I _537_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_606_ _606_/I _606_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_468_ _332_/Z _335_/Z _468_/B _469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ _393_/Z _399_/A2 _457_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[1\].id.delaybuf0/I ringosc.dstage\[1\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_322_ _461_/A1 _464_/B _322_/B _323_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayint0/I ringosc.dstage\[4\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__685__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I ext_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[0\].id.trim0bar _484_/Z ringosc.dstage\[0\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xringosc.dstage\[9\].id.delayen0 _532_/ZN ringosc.dstage\[9\].id.delayen0/I ringosc.dstage\[9\].id.delayen0/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_570_ _570_/A1 _584_/A1 _572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_553_ _575_/A2 _522_/Z _588_/A3 _520_/Z _553_/C _584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_484_ _484_/I _484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_622_ _622_/I _622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[9\].id.trim1bar _598_/ZN ringosc.dstage\[9\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__564__A1 _604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_536_ _529_/Z _536_/A2 _505_/B _536_/B2 _537_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_605_ _529_/Z _605_/A2 _605_/B _606_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_467_ _670_/Q _324_/Z _459_/Z _475_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_398_ _398_/A1 _397_/Z _399_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/I ringosc.dstage\[1\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_321_ _685_/Q _464_/B _322_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_519_ _495_/Z _519_/A2 _563_/A2 _519_/B2 _519_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__519__A1 _495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input18_I ext_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__675__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[9\].id.delayen1 _598_/ZN ringosc.dstage\[9\].id.delayen1/I ringosc.dstage\[9\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_0_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_552_ _487_/Z _563_/A2 _588_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_483_ input8/Z _483_/I1 _561_/I _484_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_621_ _621_/I _621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_535_ _575_/A2 _570_/A1 _536_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_604_ _604_/A1 _563_/Z _604_/B _605_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_397_ _349_/B _397_/A2 _387_/B _397_/A4 _397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_466_ _466_/I _669_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[8\].id.trim0bar _528_/ZN ringosc.dstage\[8\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_320_ _329_/I _464_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_518_ _507_/Z _539_/I _622_/I _519_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_13_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_449_ _442_/Z _452_/B _450_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayint0/I ringosc.dstage\[0\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xringosc.iss.reseten0 _609_/Z ringosc.iss.reseten0/I ringosc.ibufp00/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_10_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input30_I ext_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_551_ _551_/A1 _569_/A2 _554_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_620_ _610_/Z _619_/Z _621_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__665__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_482_ _510_/B _561_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.trim0bar/ZN ringosc.dstage\[8\].id.delayenb1/I
+ ringosc.dstage\[9\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_603_ _603_/A1 _603_/A2 _603_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_534_ _534_/I _534_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_396_ input2/Z _396_/A2 _396_/B _396_/C _397_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_465_ _465_/A1 _465_/A2 _466_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_517_ _517_/I _519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_448_ _414_/Z _448_/A2 _448_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_379_ _324_/Z _684_/Q _380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__600__A2 _561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.iss.delayint0 ringosc.iss.delayint0/I ringosc.iss.delayen0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input23_I ext_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__594__B2 _561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__346__A1 _666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_550_ _340_/I _565_/A2 _550_/B _569_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_481_ _481_/I _663_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_679_ _679_/D _650_/Z _686_/I _680_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_533_ _529_/Z input9/Z _553_/C _534_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_602_ _498_/Z _602_/A2 _603_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_464_ _670_/Q _464_/A2 _464_/B _465_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.trim1bar/ZN ringosc.dstage\[8\].id.delayenb1/I
+ ringosc.dstage\[8\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_395_ _383_/I _395_/A2 _397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_516_ _516_/I _516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_447_ _447_/I _674_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__678__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_378_ _669_/Q _684_/Q _380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xringosc.dstage\[6\].id.delayen0 _519_/ZN ringosc.dstage\[6\].id.delayen0/I ringosc.dstage\[7\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA_input16_I ext_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__440__I _674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__346__A2 _681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I ext_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_480_ _663_/Q _473_/B _481_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[6\].id.trim1bar _587_/ZN ringosc.dstage\[6\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_678_ _678_/D _648_/Z _686_/I _679_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xringosc.iss.reseten0_38 ringosc.iss.reseten0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
X_601_ _601_/I _601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_532_ _532_/I _532_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_463_ _324_/Z _459_/Z _465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_394_ _664_/Q _665_/Q _663_/Q _329_/I _398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_515_ _538_/I _513_/Z _515_/B _516_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_446_ _441_/Z _446_/A2 _447_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_377_ _670_/Q _685_/Q _377_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[8\].id.delaybuf0/I ringosc.dstage\[8\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.trim0bar/ZN ringosc.dstage\[4\].id.delayenb1/I
+ ringosc.dstage\[5\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_429_ _429_/I _429_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[10\].id.delayen0 _534_/ZN ringosc.dstage\[10\].id.delayen0/I ringosc.dstage\[11\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xinput1 dco _510_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xringosc.dstage\[6\].id.delayen1 _587_/ZN ringosc.dstage\[6\].id.delayen1/I ringosc.dstage\[6\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__668__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xringosc.dstage\[10\].id.trim1bar _601_/Z ringosc.dstage\[10\].id.trim1bar/ZN VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__336__I0 _681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_677_ _677_/D _645_/Z _686_/I _677_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xringosc.dstage\[5\].id.trim0bar _516_/Z ringosc.dstage\[5\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_531_ _529_/Z _531_/A2 _505_/B _531_/B2 _532_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_600_ _340_/Z _561_/Z _600_/B _601_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_393_ _672_/Q _671_/Q _402_/I _483_/I1 _393_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_462_ _462_/I _670_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_514_ _498_/Z _514_/A2 _515_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/I ringosc.dstage\[8\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.trim1bar/ZN ringosc.dstage\[4\].id.delayenb1/I
+ ringosc.dstage\[4\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_445_ _442_/Z _388_/Z _450_/A1 _443_/Z _445_/B2 _446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_376_ _376_/A1 _376_/A2 _376_/B _387_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_428_ _428_/I _428_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_359_ _667_/Q _682_/Q _360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__634__I _646_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[10\].id.delayen1 _601_/Z ringosc.dstage\[10\].id.delayen1/I ringosc.dstage\[10\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XTAP_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 div[0] input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input21_I ext_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_676_ _676_/D _642_/Z _686_/I _676_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_19_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_530_ _420_/Z _570_/A1 _531_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_392_ _420_/I _510_/A1 _483_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_461_ _461_/A1 _464_/A2 _473_/B _462_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_659_ _486_/Z _609_/I _660_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_513_ _604_/A1 _571_/A2 _513_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_444_ _433_/S _443_/Z _450_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_375_ _374_/B _375_/A2 _375_/A3 _376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_427_ _427_/I _677_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_358_ _468_/B _683_/Q _360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[4\].id.delaybuf0/I ringosc.dstage\[4\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput3 div[1] input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayint0/I ringosc.dstage\[7\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.trim0bar/ZN ringosc.dstage\[0\].id.delayenb1/I
+ ringosc.dstage\[1\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_18_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input14_I ext_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__421__A1 _604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_675_ _675_/D _640_/Z _686_/I _675_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__412__A1 _674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_391_ _677_/Q _676_/Q _675_/Q _510_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_460_ _324_/Z _459_/Z _464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_589_ _340_/Z _441_/Z _589_/A3 _591_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_658_ _658_/I _658_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_512_ _507_/I _428_/I _429_/I _571_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_443_ _414_/Z _448_/A2 _443_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_374_ _375_/A2 _375_/A3 _374_/B _376_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xringosc.dstage\[3\].id.delayen0 _501_/Z ringosc.dstage\[3\].id.delayen0/I ringosc.dstage\[4\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_426_ _340_/Z _425_/Z _427_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 div[2] _363_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_357_ _332_/Z _682_/Q _360_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/I ringosc.dstage\[4\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.trim1bar/ZN ringosc.dstage\[0\].id.delayenb1/I
+ ringosc.dstage\[0\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_10_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_409_ _676_/Q _675_/Q _563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xringosc.iss.delayenb0 ringosc.iss.ctrlen0/ZN ringosc.iss.delayenb1/I ringosc.ibufp00/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_15_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__681__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[3\].id.trim1bar _573_/ZN ringosc.dstage\[3\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_674_ _674_/D _638_/Z _686_/I _674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_390_ _674_/Q _673_/Q _420_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_588_ _585_/B _522_/Z _588_/A3 _559_/B _603_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_657_ _486_/Z _609_/I _658_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_511_ _507_/Z _548_/I _553_/C _538_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_442_ _673_/Q _442_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_373_ _363_/I _370_/Z _376_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_425_ _445_/B2 _425_/I1 _425_/S _425_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_356_ _668_/Q _683_/Q _356_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xinput5 div[3] _374_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[3\].id.delayen1 _573_/ZN ringosc.dstage\[3\].id.delayen1/I ringosc.dstage\[3\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XTAP_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_408_ _388_/Z _433_/S _445_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_339_ _507_/I _340_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xringosc.iss.delayenb1 ringosc.iss.trim1bar/ZN ringosc.iss.delayenb1/I ringosc.iss.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/I ringosc.dstage\[0\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput30 ext_trim[6] _517_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayint0/I ringosc.dstage\[3\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_14_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[2\].id.trim0bar _497_/ZN ringosc.dstage\[2\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_673_ _673_/D _636_/Z _686_/I _673_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__671__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_587_ _587_/A1 _587_/A2 _587_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_656_ _656_/I _656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_441_ _539_/I _441_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_510_ _510_/A1 _575_/A2 _510_/B _553_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_372_ _372_/A1 _396_/B _396_/C _387_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_639_ _634_/Z _631_/Z _640_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_424_ _411_/Z _437_/A1 _423_/Z _425_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_355_ _380_/A1 _368_/B _380_/A3 _367_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput6 div[4] _383_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_338_ _677_/Q _507_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_407_ _407_/I _433_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/I ringosc.dstage\[0\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 ext_trim[20] _590_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 ext_trim[7] _525_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/I ringosc.iss.delayen1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_672_ _672_/D _633_/Z _686_/I _672_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input12_I ext_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_586_ _524_/Z _586_/A2 _587_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_655_ _646_/Z _609_/I _656_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input4_I div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_440_ _674_/Q _539_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_371_ _374_/B _375_/A2 _375_/A3 _363_/I _370_/Z _396_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_569_ _569_/A1 _569_/A2 _569_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_638_ _638_/I _638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_423_ _429_/I _402_/I _423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_354_ _668_/Q _683_/Q _341_/Z _346_/Z _364_/B _380_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__684__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 enable input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_406_ _457_/A2 _435_/A2 _407_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_337_ _337_/I _681_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__686__I _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 ext_trim[11] _536_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 ext_trim[8] _527_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 ext_trim[21] _593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__590__A1 _498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_671_ _671_/D _630_/Z _686_/I _671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_19_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__342__A1 _666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_ringosc.dstage\[0\].id.delayenb0_I ringosc.dstage\[0\].id.delayenb1/I VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_585_ _412_/Z _522_/Z _585_/B _587_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_654_ _654_/I _654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_637_ _634_/Z _631_/Z _638_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_370_ _370_/A1 _365_/Z _370_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_568_ _495_/Z _568_/A2 _573_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_499_ _498_/Z _499_/A2 _500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xringosc.dstage\[0\].id.delayen0 _484_/Z ringosc.dstage\[0\].id.delayen0/I ringosc.dstage\[1\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_422_ _675_/Q _429_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_10_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_353_ _667_/Q _682_/Q _364_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput8 ext_trim[0] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.trim0bar/ZN ringosc.dstage\[7\].id.delayenb1/I
+ ringosc.dstage\[8\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_405_ _504_/A2 _410_/A1 _405_/A3 _575_/A2 _435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_336_ _681_/Q _335_/Z _478_/S _337_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__674__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I resetb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[0\].id.trim1bar _546_/ZN ringosc.dstage\[0\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput11 ext_trim[12] _542_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 ext_trim[9] _531_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 ext_trim[22] _595_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_319_ _680_/D _680_/Q _329_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_670_ _670_/D _628_/Z _686_/I _670_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__342__A2 _681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_584_ _584_/A1 _580_/Z _584_/A3 _584_/B1 _561_/Z _584_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_16_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_653_ _646_/Z _643_/Z _654_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_567_ _567_/I _567_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_498_ _510_/B _498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_636_ _636_/I _636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _604_/A1 _414_/Z _448_/A2 _420_/Z _388_/Z _437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xringosc.dstage\[0\].id.delayen1 _546_/ZN ringosc.dstage\[0\].id.delayen1/I ringosc.dstage\[0\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xinput9 ext_trim[10] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_352_ _669_/Q _684_/Q _368_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_619_ _643_/I _619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.trim1bar/ZN ringosc.dstage\[7\].id.delayenb1/I
+ ringosc.dstage\[7\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_404_ _674_/Q _673_/Q _575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_335_ _666_/Q _335_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input28_I ext_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput12 ext_trim[13] _545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 ext_trim[23] _599_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput34 osc _678_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_318_ _670_/Q _461_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[8\].id.delayen0 _528_/ZN ringosc.dstage\[8\].id.delayen0/I ringosc.dstage\[9\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_19_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__664__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_583_ _583_/I _584_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_652_ _652_/I _652_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input10_I ext_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_566_ _529_/Z _566_/A2 _566_/B1 _566_/B2 _567_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_497_ _497_/A1 _497_/A2 _497_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_635_ _634_/Z _631_/Z _636_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xringosc.dstage\[8\].id.trim1bar _594_/ZN ringosc.dstage\[8\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input2_I div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _420_/I _420_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_351_ _468_/B _683_/Q _380_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_549_ _412_/Z _522_/I _550_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__390__A1 _674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_618_ _618_/I _618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_403_ _507_/I _675_/Q _672_/Q _671_/Q _405_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_334_ _334_/I _682_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput13 ext_trim[14] _560_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 ext_trim[24] _602_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 resetb _607_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[7\].id.delaybuf0/I ringosc.dstage\[7\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__584__B2 _561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.trim0bar/ZN ringosc.dstage\[3\].id.delayenb1/I
+ ringosc.dstage\[4\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayint0/I ringosc.dstage\[11\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[8\].id.delayen1 _594_/ZN ringosc.dstage\[8\].id.delayen1/I ringosc.dstage\[8\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_582_ _582_/A1 _597_/B _569_/Z _582_/A4 _584_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_16_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_651_ _646_/Z _643_/Z _652_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_565_ _507_/Z _565_/A2 _565_/B _565_/C _566_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_496_ _495_/Z _496_/A2 _497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_634_ _646_/I _634_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__677__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[7\].id.trim0bar _526_/ZN ringosc.dstage\[7\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_350_ _374_/B _367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_548_ _548_/I _565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_617_ _610_/Z _609_/Z _618_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_479_ _479_/I _664_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_402_ _402_/I _410_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_333_ _682_/Q _332_/Z _478_/S _334_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput14 ext_trim[15] _566_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput25 ext_trim[25] _605_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/I ringosc.dstage\[7\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.trim1bar/ZN ringosc.dstage\[3\].id.delayenb1/I
+ ringosc.dstage\[3\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_22_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input33_I ext_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__335__I _666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_650_ _650_/I _650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_581_ _539_/I _563_/Z _597_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_564_ _604_/A1 _563_/Z _566_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_495_ _622_/I _495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_633_ _633_/I _633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[11\].id.trim0bar _537_/ZN ringosc.dstage\[11\].id.trim0bar/ZN VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_547_ _604_/A1 _571_/A2 _551_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_616_ _616_/I _616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_478_ _664_/Q _663_/Q _478_/S _479_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__602__A1 _498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_401_ _428_/I _504_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_332_ _667_/Q _332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__667__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput15 ext_trim[16] _568_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 ext_trim[2] _496_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input26_I ext_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[3\].id.delaybuf0/I ringosc.dstage\[3\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayint0/I ringosc.dstage\[6\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_580_ _580_/A1 _442_/Z _563_/Z _580_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_21_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_563_ _487_/Z _563_/A2 _563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_632_ _622_/Z _631_/Z _633_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_494_ _510_/B _622_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_546_ _546_/A1 _546_/A2 _546_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xringosc.ibufp10 ringosc.ibufp10/I ringosc.ibufp11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_477_ _477_/I _665_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_615_ _610_/Z _609_/Z _616_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_400_ _676_/Q _428_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_331_ _331_/I _683_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__520__A1 _674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_529_ _646_/I _529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__529__I _646_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 ext_trim[17] _577_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__502__A1 _495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput27 ext_trim[3] _499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[5\].id.delayen0 _516_/Z ringosc.dstage\[5\].id.delayen0/I ringosc.ibufp10/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA_input19_I ext_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/I ringosc.dstage\[3\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[5\].id.trim1bar _584_/ZN ringosc.dstage\[5\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_562_ _565_/B _565_/C _562_/A3 _562_/B1 _561_/Z _562_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_493_ _493_/I _493_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_631_ _643_/I _631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_545_ _524_/Z _545_/A2 _546_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_476_ _665_/Q _664_/Q _478_/S _477_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xringosc.ibufp00 ringosc.ibufp00/I ringosc.ibufp01/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_614_ _614_/I _614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.ibufp11 ringosc.ibufp11/I output37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_330_ _683_/Q _468_/B _478_/S _331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_528_ _538_/I _528_/A2 _528_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_459_ _468_/B _332_/Z _335_/Z _459_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xinput17 ext_trim[18] _583_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 ext_trim[4] _502_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[5\].id.delayen1 _584_/ZN ringosc.dstage\[5\].id.delayen1/I ringosc.dstage\[5\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_22_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__496__A1 _495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input31_I ext_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_561_ _561_/I _561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_492_ _486_/Z _492_/A2 _585_/B _493_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_630_ _630_/I _630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[4\].id.trim0bar _506_/ZN ringosc.dstage\[4\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayint0/I ringosc.dstage\[2\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_14_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xringosc.ibufp01 ringosc.ibufp01/I _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XTAP_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_613_ _610_/Z _609_/Z _614_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_544_ _441_/Z _522_/Z _585_/B _546_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_475_ _335_/Z _464_/B _475_/A3 _666_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_527_ _524_/Z _527_/A2 _528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_389_ _389_/I _402_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_458_ _458_/I _671_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput18 ext_trim[19] _586_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput29 ext_trim[5] _514_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__646__I _646_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__680__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.trim0bar/ZN ringosc.dstage\[11\].id.delayenb1/I
+ ringosc.iss.delayenb1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_17_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input24_I ext_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_560_ _560_/I _562_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_491_ _570_/A1 _497_/A1 _585_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_12_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__605__A2 _605_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_543_ _578_/A1 _543_/A2 _543_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__599__A1 _561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_474_ _474_/I _667_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_612_ _612_/I _612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_526_ _526_/A1 _526_/A2 _526_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__514__A1 _498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_388_ _389_/I _388_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_457_ _415_/Z _457_/A2 _457_/B _458_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput19 ext_trim[1] _492_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_509_ _563_/A2 _412_/Z _575_/A3 _420_/Z _548_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.trim1bar/ZN ringosc.dstage\[11\].id.delayenb1/I
+ ringosc.dstage\[11\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_10_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input17_I ext_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__670__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I ext_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_490_ _487_/Z _428_/Z _561_/I _497_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_542_ _524_/Z _542_/A2 _543_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_473_ _475_/A3 _473_/A2 _473_/B _474_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_611_ _610_/Z _609_/Z _612_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_525_ _524_/Z _525_/A2 _526_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_456_ _415_/Z _452_/B _457_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_387_ _387_/A1 _387_/A2 _382_/Z _387_/B _389_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_11_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[2\].id.delayen0 _497_/ZN ringosc.dstage\[2\].id.delayen0/I ringosc.dstage\[3\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_508_ _428_/I _429_/I _575_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__499__A1 _498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_439_ _439_/I _675_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[2\].id.trim1bar _567_/ZN ringosc.dstage\[2\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.trim0bar/ZN ringosc.dstage\[6\].id.delayenb1/I
+ ringosc.dstage\[7\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[11\].id.delaybuf0/I ringosc.dstage\[11\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_541_ _541_/A1 _569_/A1 _578_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_472_ _332_/Z _335_/Z _473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_610_ _622_/I _610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__683__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_524_ _646_/I _524_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_386_ _670_/Q _685_/Q _386_/B1 _384_/Z _386_/C _387_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_455_ _455_/I _672_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[2\].id.delayen1 _567_/ZN ringosc.dstage\[2\].id.delayen1/I ringosc.dstage\[2\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xrebuffer1 rebuffer2/I rebuffer1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_507_ _507_/I _507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_438_ _429_/Z _433_/S _438_/B _439_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_369_ _380_/A1 _362_/B _380_/A3 _375_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.trim1bar/ZN ringosc.dstage\[6\].id.delayenb1/I
+ ringosc.dstage\[6\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA__562__B2 _561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/I ringosc.dstage\[11\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input22_I ext_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[1\].id.trim0bar _493_/ZN ringosc.dstage\[1\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_686_ _686_/I _686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_540_ _580_/A1 _442_/Z _571_/A2 _569_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_471_ _471_/I _668_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_669_ _669_/D _626_/Z _686_/I _669_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_523_ _520_/Z _522_/Z _585_/B _526_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xringosc.iss.delayen0 _543_/ZN ringosc.iss.delayen0/I ringosc.ibufp00/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
X_454_ _454_/A1 _433_/S _454_/B _455_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_385_ _377_/Z _385_/A2 _386_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__673__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer2 rebuffer2/I rebuffer2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_506_ _506_/A1 _506_/A2 _506_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_437_ _437_/A1 _423_/Z _437_/B _438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_368_ _356_/Z _368_/A2 _368_/B _375_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xringosc.iss.trim1bar _606_/ZN ringosc.iss.trim1bar/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I ext_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_685_ _685_/D _662_/Z _686_/I _685_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input7_I enable VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/I ringosc.dstage\[6\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.trim0bar/ZN ringosc.dstage\[2\].id.delayenb1/I
+ ringosc.dstage\[3\].id.delaybuf0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayint0/I ringosc.dstage\[9\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayint0/I ringosc.dstage\[10\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_599_ _561_/Z _599_/A2 _600_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_470_ _475_/A3 _469_/Z _473_/B _471_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_668_ _668_/D _624_/Z _686_/I _668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_522_ _522_/I _522_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xringosc.iss.delayen1 _606_/ZN ringosc.iss.delayen1/I ringosc.iss.delayint0/I VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
X_453_ _415_/Z _417_/Z _453_/B _454_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_384_ _377_/Z _385_/A2 _384_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_505_ _441_/Z _582_/A1 _505_/B _506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xringosc.dstage\[9\].id.trim0bar _532_/ZN ringosc.dstage\[9\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_436_ _437_/A1 _423_/Z _452_/B _437_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_367_ _367_/A1 _367_/A2 _367_/A3 _367_/B1 _367_/B2 _396_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_19_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_419_ _415_/Z _417_/Z _419_/B _448_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__663__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_684_ _684_/D _660_/Z _686_/I _684_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/I ringosc.dstage\[6\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.trim1bar/ZN ringosc.dstage\[2\].id.delayenb1/I
+ ringosc.dstage\[2\].id.delayint0/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_598_ _598_/A1 _598_/A2 _598_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_667_ _667_/D _621_/Z _686_/I _667_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_521_ _340_/I _676_/Q _675_/Q _522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_452_ _415_/Z _417_/Z _452_/B _453_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_383_ _383_/I _386_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_504_ _340_/Z _504_/A2 _622_/I _505_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_435_ _457_/A2 _435_/A2 _452_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_366_ _370_/A1 _365_/Z _367_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__344__A1 _666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_418_ _454_/A1 _402_/I _419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_349_ input3/Z _343_/Z _349_/B _372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__547__A1 _604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.iss.ctrlen0 _609_/Z _543_/ZN ringosc.iss.ctrlen0/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_683_ _683_/D _658_/Z _686_/I _683_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input20_I ext_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__676__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_597_ _441_/Z _559_/B _597_/B _597_/C _598_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_666_ _666_/D _618_/Z _686_/I _666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_520_ _674_/Q _442_/Z _520_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[2\].id.delaybuf0/I ringosc.dstage\[2\].id.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayint0/I ringosc.dstage\[5\].id.delayen0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_451_ _451_/I _673_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_649_ _646_/Z _643_/Z _650_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_382_ _383_/I _395_/A2 _382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_503_ _340_/I _428_/Z _429_/Z _582_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_434_ _434_/I _676_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_365_ _356_/Z _360_/B _365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__344__A2 _681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_417_ _454_/A1 _389_/I _417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_348_ _348_/A1 _347_/Z _349_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xringosc.dstage\[7\].id.delayen0 _526_/ZN ringosc.dstage\[7\].id.delayen0/I ringosc.dstage\[8\].id.delaybuf0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_20_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_682_ _682_/D _656_/Z _686_/I _682_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input13_I ext_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_596_ _565_/B _565_/C _580_/Z _597_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_665_ _665_/D _616_/Z _686_/I _665_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/I ringosc.dstage\[2\].id.delayen1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input5_I div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[7\].id.trim1bar _592_/Z ringosc.dstage\[7\].id.trim1bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_450_ _450_/A1 _448_/Z _450_/B _451_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_381_ _377_/Z _385_/A2 _395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_579_ _579_/I _579_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_648_ _648_/I _648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__666__CLK _686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_502_ _495_/Z _502_/A2 _506_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_433_ _428_/Z _433_/I1 _433_/S _434_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_364_ _341_/Z _346_/Z _364_/B _370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_416_ _672_/Q _454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_347_ input3/Z _341_/Z _346_/Z _347_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_5_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[11\].id.delayen0 _537_/ZN ringosc.dstage\[11\].id.delayen0/I ringosc.iss.delayenb1/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_2
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xringosc.dstage\[7\].id.delayen1 _592_/Z ringosc.dstage\[7\].id.delayen1/I ringosc.dstage\[7\].id.delayint0/I
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__invz_1
XFILLER_18_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_681_ _681_/D _654_/Z _686_/I _681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_ringosc.dstage\[0\].id.delayenb1_I ringosc.dstage\[0\].id.delayenb1/I VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_595_ _495_/Z _595_/A2 _598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_664_ _664_/D _614_/Z _686_/I _664_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__524__I _646_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xringosc.dstage\[11\].id.trim1bar _603_/ZN ringosc.dstage\[11\].id.trim1bar/ZN VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_380_ _380_/A1 _380_/A2 _380_/A3 _380_/B _385_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xringosc.dstage\[6\].id.trim0bar _519_/ZN ringosc.dstage\[6\].id.trim0bar/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_578_ _578_/A1 _578_/A2 _578_/B _579_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__595__A1 _495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_647_ _646_/Z _643_/Z _648_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
.ends

