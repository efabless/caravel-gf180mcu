* Simple Schmitt trigger inverter testbench (No. 3:  Running at 3.3V)
* (Layout-extracted netlist)

.include /usr/share/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /usr/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /usr/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.include ../mag/simple_por.spice

V0 VDD 0 3.3
V1 In 0 PWL(0 0 100u 3.3 200u 3.3 300u 0)

X0 VDD 0 In Out schmitt_inverter

.control
tran 500n 350u
plot V(In) V(Out)
.endc
